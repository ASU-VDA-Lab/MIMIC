module fake_ariane_1702_n_1666 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_136, n_28, n_80, n_97, n_14, n_88, n_141, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1666);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_136;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1666;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_143;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_699;
wire n_727;
wire n_590;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1649;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1635;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g142 ( 
.A(n_16),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_75),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g144 ( 
.A(n_140),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_3),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_128),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_89),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_47),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_29),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_4),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_62),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_44),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_108),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_47),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_52),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_101),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_74),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_80),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_57),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_117),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_36),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_127),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_85),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_106),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_77),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_48),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_17),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_133),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_110),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_60),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_93),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_124),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_81),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_119),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_120),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_32),
.Y(n_185)
);

BUFx5_ASAP7_75t_L g186 ( 
.A(n_10),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_92),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_12),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_76),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_9),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_66),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_53),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_107),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_83),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_28),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_16),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_27),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_20),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_114),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_41),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_104),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_91),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_123),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_19),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_17),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_103),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_27),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_9),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_90),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_26),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_1),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_70),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_125),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_73),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_48),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_30),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_39),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_15),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_102),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_136),
.Y(n_225)
);

INVx4_ASAP7_75t_R g226 ( 
.A(n_2),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_88),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_111),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_118),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_98),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_67),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_18),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_121),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_32),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_55),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_113),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_30),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_130),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_21),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_29),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_41),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_69),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_132),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_4),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_64),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_95),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_46),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_65),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_18),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_134),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_5),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_26),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_97),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_20),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_54),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_35),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_51),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_34),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_126),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_11),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_131),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_49),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_5),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_50),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_137),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_116),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_94),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_58),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_35),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_24),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_7),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_14),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_10),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_28),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_82),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_22),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_100),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_19),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_8),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_122),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_25),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_78),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_59),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_115),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_248),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_150),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_145),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_0),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_186),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_197),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_186),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_186),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_276),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_186),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_150),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_153),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_186),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_168),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_186),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_186),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_250),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_250),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_0),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_250),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_250),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_173),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_181),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_185),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_181),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_231),
.Y(n_318)
);

INVxp67_ASAP7_75t_SL g319 ( 
.A(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_253),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_253),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_192),
.Y(n_322)
);

NOR2xp67_ASAP7_75t_L g323 ( 
.A(n_245),
.B(n_1),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_196),
.Y(n_324)
);

INVxp67_ASAP7_75t_SL g325 ( 
.A(n_253),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_231),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_253),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_199),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_259),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_259),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_206),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_259),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_259),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_188),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_212),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_274),
.Y(n_339)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_188),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_261),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_274),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_261),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_215),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_3),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_277),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_201),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_220),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_277),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_284),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_201),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_284),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_149),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_208),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_222),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_149),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_208),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_154),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_230),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_271),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_154),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_189),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_210),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_210),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_240),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_146),
.B(n_6),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_189),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_227),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_155),
.B(n_7),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_161),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_294),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_291),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_297),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_302),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_217),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_315),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_359),
.B(n_227),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_308),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_297),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_299),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_299),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_317),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_308),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_318),
.Y(n_385)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_347),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_326),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_290),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_330),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_341),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_343),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_292),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_351),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_301),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_304),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_304),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_306),
.Y(n_403)
);

CKINVDCx8_ASAP7_75t_R g404 ( 
.A(n_303),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_354),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_307),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_335),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_335),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_307),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_R g412 ( 
.A(n_295),
.B(n_268),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_359),
.B(n_249),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_309),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_305),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_309),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_359),
.B(n_144),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_314),
.Y(n_418)
);

BUFx8_ASAP7_75t_L g419 ( 
.A(n_296),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_311),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_316),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g422 ( 
.A1(n_311),
.A2(n_160),
.B(n_157),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_312),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_322),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_312),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_342),
.B(n_162),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

NAND3xp33_ASAP7_75t_L g428 ( 
.A(n_369),
.B(n_151),
.C(n_142),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_320),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_345),
.B(n_262),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_321),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_357),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_321),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_296),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_329),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_329),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_331),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_363),
.B(n_364),
.Y(n_438)
);

NAND2x1_ASAP7_75t_L g439 ( 
.A(n_353),
.B(n_226),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_331),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_334),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_334),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_356),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_426),
.B(n_352),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_396),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_371),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_431),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_376),
.A2(n_293),
.B1(n_310),
.B2(n_324),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

AND2x2_ASAP7_75t_SL g454 ( 
.A(n_376),
.B(n_366),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_415),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_328),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_426),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_392),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_426),
.B(n_313),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_323),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_413),
.B(n_360),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_360),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

BUFx8_ASAP7_75t_SL g466 ( 
.A(n_387),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_434),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_392),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_392),
.Y(n_470)
);

BUFx8_ASAP7_75t_SL g471 ( 
.A(n_387),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_417),
.B(n_319),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_417),
.B(n_325),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_436),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_414),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_436),
.Y(n_477)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_434),
.B(n_313),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_404),
.B(n_332),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_327),
.Y(n_480)
);

NAND2xp33_ASAP7_75t_R g481 ( 
.A(n_390),
.B(n_338),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_437),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_414),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

BUFx8_ASAP7_75t_SL g485 ( 
.A(n_397),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_378),
.B(n_344),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_378),
.B(n_348),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_405),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_411),
.B(n_336),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_372),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_404),
.B(n_355),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_401),
.B(n_298),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_418),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_411),
.B(n_340),
.Y(n_495)
);

AND2x2_ASAP7_75t_SL g496 ( 
.A(n_390),
.B(n_262),
.Y(n_496)
);

BUFx8_ASAP7_75t_SL g497 ( 
.A(n_397),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_401),
.B(n_300),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_437),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_438),
.B(n_365),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_374),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_427),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_404),
.B(n_158),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_374),
.B(n_356),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_432),
.A2(n_263),
.B1(n_281),
.B2(n_240),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_380),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_373),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_427),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_380),
.B(n_381),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_386),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_382),
.Y(n_512)
);

AND2x2_ASAP7_75t_SL g513 ( 
.A(n_422),
.B(n_152),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_421),
.B(n_158),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_398),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_424),
.B(n_268),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_412),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_386),
.B(n_358),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_443),
.B(n_337),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_386),
.B(n_361),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_375),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_419),
.Y(n_524)
);

INVx5_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

BUFx3_ASAP7_75t_L g526 ( 
.A(n_399),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_428),
.B(n_164),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_377),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_399),
.B(n_361),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_430),
.B(n_337),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_400),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_400),
.B(n_362),
.Y(n_532)
);

INVx4_ASAP7_75t_L g533 ( 
.A(n_402),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_419),
.B(n_164),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_L g535 ( 
.A1(n_430),
.A2(n_422),
.B1(n_410),
.B2(n_443),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_402),
.Y(n_536)
);

NAND2xp33_ASAP7_75t_L g537 ( 
.A(n_402),
.B(n_163),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_443),
.B(n_339),
.Y(n_539)
);

BUFx2_ASAP7_75t_L g540 ( 
.A(n_419),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_419),
.B(n_263),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_410),
.Y(n_542)
);

INVx4_ASAP7_75t_L g543 ( 
.A(n_403),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_403),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_383),
.B(n_273),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_422),
.A2(n_214),
.B1(n_251),
.B2(n_234),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_414),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_419),
.B(n_165),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_406),
.B(n_367),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_406),
.B(n_367),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_414),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_406),
.B(n_165),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_438),
.B(n_281),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_422),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_406),
.B(n_368),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_416),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_416),
.B(n_368),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_429),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_429),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_422),
.A2(n_174),
.B1(n_265),
.B2(n_190),
.Y(n_560)
);

AO22x2_ASAP7_75t_L g561 ( 
.A1(n_412),
.A2(n_256),
.B1(n_205),
.B2(n_258),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_420),
.B(n_425),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_435),
.Y(n_563)
);

AND2x6_ASAP7_75t_L g564 ( 
.A(n_420),
.B(n_271),
.Y(n_564)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_414),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_440),
.B(n_166),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_440),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_385),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_435),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_388),
.B(n_273),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_394),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_441),
.A2(n_278),
.B1(n_241),
.B2(n_239),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_435),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_442),
.B(n_339),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_442),
.B(n_379),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_414),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_423),
.B(n_163),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_442),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_423),
.B(n_176),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g581 ( 
.A(n_433),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_379),
.B(n_207),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_379),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_384),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_526),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_454),
.B(n_166),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_526),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_458),
.B(n_167),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_489),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_490),
.B(n_395),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_459),
.B(n_171),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_517),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_459),
.B(n_246),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_445),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_454),
.B(n_235),
.Y(n_595)
);

O2A1O1Ixp33_ASAP7_75t_L g596 ( 
.A1(n_509),
.A2(n_198),
.B(n_221),
.C(n_223),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_447),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_533),
.B(n_235),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_533),
.B(n_272),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_505),
.A2(n_267),
.B1(n_242),
.B2(n_260),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_583),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_524),
.B(n_346),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_447),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_444),
.B(n_463),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_486),
.B(n_266),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_583),
.Y(n_606)
);

NOR3x1_ASAP7_75t_L g607 ( 
.A(n_516),
.B(n_159),
.C(n_156),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_524),
.B(n_346),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_455),
.Y(n_610)
);

A2O1A1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_549),
.A2(n_286),
.B(n_237),
.C(n_232),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_444),
.B(n_272),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_502),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_472),
.B(n_275),
.Y(n_614)
);

OR2x6_ASAP7_75t_L g615 ( 
.A(n_540),
.B(n_349),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_474),
.B(n_280),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_480),
.B(n_461),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_533),
.B(n_205),
.Y(n_618)
);

INVx2_ASAP7_75t_SL g619 ( 
.A(n_490),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_536),
.B(n_178),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_461),
.B(n_283),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_493),
.B(n_143),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_536),
.B(n_204),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_493),
.B(n_147),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_496),
.A2(n_180),
.B1(n_209),
.B2(n_211),
.Y(n_625)
);

A2O1A1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_496),
.A2(n_350),
.B(n_349),
.C(n_219),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_517),
.B(n_148),
.Y(n_627)
);

INVx3_ASAP7_75t_L g628 ( 
.A(n_538),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_536),
.B(n_233),
.Y(n_629)
);

AND3x1_ASAP7_75t_L g630 ( 
.A(n_450),
.B(n_350),
.C(n_216),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g631 ( 
.A(n_507),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_501),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_508),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_561),
.A2(n_230),
.B1(n_393),
.B2(n_409),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_538),
.B(n_169),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_538),
.B(n_170),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_487),
.B(n_216),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_495),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_527),
.B(n_216),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_540),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_543),
.B(n_244),
.Y(n_641)
);

A2O1A1Ixp33_ASAP7_75t_L g642 ( 
.A1(n_501),
.A2(n_257),
.B(n_264),
.C(n_269),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_530),
.B(n_172),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_543),
.B(n_270),
.Y(n_644)
);

OAI22x1_ASAP7_75t_SL g645 ( 
.A1(n_445),
.A2(n_282),
.B1(n_288),
.B2(n_285),
.Y(n_645)
);

AND2x4_ASAP7_75t_L g646 ( 
.A(n_464),
.B(n_384),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_530),
.B(n_464),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_508),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_511),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_530),
.B(n_177),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_530),
.B(n_179),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_515),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_515),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_531),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_531),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_464),
.B(n_384),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_511),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_561),
.A2(n_183),
.B1(n_279),
.B2(n_255),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_453),
.B(n_182),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_543),
.B(n_163),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_542),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_544),
.B(n_230),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_491),
.B(n_506),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_8),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_512),
.B(n_184),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_456),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_467),
.A2(n_542),
.B1(n_498),
.B2(n_544),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_503),
.B(n_11),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_519),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_562),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_519),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_495),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_561),
.A2(n_218),
.B1(n_187),
.B2(n_252),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_558),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_558),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_514),
.B(n_13),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_451),
.B(n_163),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_541),
.A2(n_433),
.B1(n_423),
.B2(n_229),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_520),
.B(n_522),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_559),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_521),
.B(n_539),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_539),
.B(n_191),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_451),
.B(n_163),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_498),
.B(n_193),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_456),
.B(n_194),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_575),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_566),
.B(n_13),
.Y(n_687)
);

AOI22x1_ASAP7_75t_L g688 ( 
.A1(n_446),
.A2(n_465),
.B1(n_448),
.B2(n_452),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_556),
.B(n_195),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_479),
.B(n_14),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_575),
.Y(n_691)
);

BUFx6f_ASAP7_75t_SL g692 ( 
.A(n_467),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_567),
.B(n_200),
.Y(n_693)
);

OAI22x1_ASAP7_75t_L g694 ( 
.A1(n_553),
.A2(n_228),
.B1(n_225),
.B2(n_213),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_451),
.B(n_163),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_559),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_573),
.B(n_243),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_557),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_561),
.A2(n_513),
.B1(n_546),
.B2(n_560),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_510),
.Y(n_700)
);

INVx8_ASAP7_75t_L g701 ( 
.A(n_564),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_446),
.B(n_448),
.Y(n_702)
);

NOR2xp67_ASAP7_75t_SL g703 ( 
.A(n_494),
.B(n_238),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_564),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_492),
.B(n_21),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_563),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_504),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_451),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_537),
.A2(n_423),
.B(n_433),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_470),
.B(n_175),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_481),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_552),
.B(n_22),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_534),
.B(n_23),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_494),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_563),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_548),
.B(n_23),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_569),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_462),
.A2(n_202),
.B1(n_203),
.B2(n_236),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_569),
.Y(n_719)
);

A2O1A1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_529),
.A2(n_393),
.B(n_389),
.C(n_409),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_466),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_475),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_470),
.B(n_476),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_532),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_477),
.B(n_407),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_482),
.Y(n_726)
);

INVxp67_ASAP7_75t_L g727 ( 
.A(n_466),
.Y(n_727)
);

BUFx3_ASAP7_75t_L g728 ( 
.A(n_581),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_513),
.A2(n_393),
.B1(n_389),
.B2(n_409),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_470),
.B(n_175),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_482),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_484),
.B(n_408),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_484),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_462),
.A2(n_433),
.B1(n_423),
.B2(n_175),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_545),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_588),
.B(n_478),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_597),
.Y(n_737)
);

AOI21xp5_ASAP7_75t_L g738 ( 
.A1(n_660),
.A2(n_537),
.B(n_449),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_660),
.A2(n_460),
.B(n_457),
.Y(n_739)
);

OAI21xp5_ASAP7_75t_L g740 ( 
.A1(n_720),
.A2(n_535),
.B(n_488),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_604),
.B(n_478),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_625),
.A2(n_528),
.B1(n_571),
.B2(n_462),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_702),
.A2(n_449),
.B(n_473),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_670),
.B(n_516),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_699),
.A2(n_553),
.B1(n_564),
.B2(n_545),
.Y(n_745)
);

BUFx3_ASAP7_75t_L g746 ( 
.A(n_594),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_723),
.A2(n_449),
.B(n_457),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_723),
.A2(n_623),
.B(n_620),
.Y(n_748)
);

OAI21xp33_ASAP7_75t_L g749 ( 
.A1(n_685),
.A2(n_570),
.B(n_568),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_603),
.Y(n_750)
);

INVx11_ASAP7_75t_L g751 ( 
.A(n_692),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_698),
.B(n_550),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_619),
.B(n_638),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_707),
.B(n_555),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_672),
.B(n_523),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_618),
.A2(n_468),
.B(n_473),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_724),
.B(n_488),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_618),
.A2(n_460),
.B(n_473),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_711),
.B(n_500),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_594),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_612),
.B(n_686),
.Y(n_761)
);

AND2x2_ASAP7_75t_SL g762 ( 
.A(n_630),
.B(n_500),
.Y(n_762)
);

BUFx8_ASAP7_75t_L g763 ( 
.A(n_692),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_598),
.A2(n_468),
.B(n_499),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_666),
.B(n_572),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_708),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_721),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_641),
.A2(n_469),
.B1(n_470),
.B2(n_554),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_610),
.A2(n_469),
.B1(n_554),
.B2(n_565),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_666),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_735),
.B(n_471),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_589),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_714),
.B(n_579),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_623),
.A2(n_577),
.B(n_565),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_629),
.A2(n_577),
.B(n_565),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_629),
.A2(n_577),
.B(n_578),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_691),
.B(n_564),
.Y(n_777)
);

OAI21xp33_ASAP7_75t_L g778 ( 
.A1(n_684),
.A2(n_580),
.B(n_574),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_681),
.B(n_564),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_644),
.A2(n_578),
.B(n_576),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_646),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_631),
.Y(n_782)
);

OAI21xp33_ASAP7_75t_L g783 ( 
.A1(n_622),
.A2(n_581),
.B(n_584),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_701),
.B(n_704),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_599),
.A2(n_476),
.B(n_551),
.Y(n_785)
);

AO22x1_ASAP7_75t_L g786 ( 
.A1(n_714),
.A2(n_471),
.B1(n_485),
.B2(n_497),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_668),
.A2(n_584),
.B(n_551),
.C(n_476),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_720),
.A2(n_547),
.B(n_525),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_644),
.A2(n_551),
.B(n_476),
.Y(n_789)
);

AOI21x1_ASAP7_75t_L g790 ( 
.A1(n_677),
.A2(n_408),
.B(n_391),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_668),
.A2(n_547),
.B(n_525),
.C(n_483),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_662),
.A2(n_547),
.B(n_525),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_663),
.A2(n_731),
.B(n_722),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_640),
.B(n_547),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_L g795 ( 
.A1(n_586),
.A2(n_389),
.B(n_391),
.C(n_407),
.Y(n_795)
);

INVx3_ASAP7_75t_L g796 ( 
.A(n_646),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_SL g797 ( 
.A(n_727),
.B(n_485),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_713),
.A2(n_525),
.B(n_483),
.C(n_433),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_627),
.A2(n_525),
.B(n_483),
.Y(n_799)
);

OAI22xp5_ASAP7_75t_L g800 ( 
.A1(n_632),
.A2(n_483),
.B1(n_433),
.B2(n_423),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_586),
.B(n_497),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_605),
.B(n_391),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_614),
.B(n_407),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_616),
.B(n_637),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_635),
.A2(n_224),
.B(n_207),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_602),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_637),
.B(n_408),
.Y(n_807)
);

AOI22x1_ASAP7_75t_L g808 ( 
.A1(n_652),
.A2(n_433),
.B1(n_423),
.B2(n_224),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_725),
.A2(n_732),
.B(n_654),
.Y(n_809)
);

BUFx8_ASAP7_75t_L g810 ( 
.A(n_587),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_653),
.A2(n_224),
.B(n_207),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_655),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_640),
.B(n_175),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_595),
.B(n_24),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_591),
.B(n_31),
.Y(n_815)
);

AO32x2_ASAP7_75t_L g816 ( 
.A1(n_600),
.A2(n_582),
.A3(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_593),
.B(n_31),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_661),
.A2(n_733),
.B(n_726),
.Y(n_818)
);

OAI21xp5_ASAP7_75t_L g819 ( 
.A1(n_709),
.A2(n_582),
.B(n_175),
.Y(n_819)
);

O2A1O1Ixp5_ASAP7_75t_L g820 ( 
.A1(n_664),
.A2(n_582),
.B(n_37),
.C(n_38),
.Y(n_820)
);

BUFx8_ASAP7_75t_L g821 ( 
.A(n_585),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_602),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_621),
.B(n_33),
.Y(n_823)
);

CKINVDCx8_ASAP7_75t_R g824 ( 
.A(n_602),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_624),
.B(n_38),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_677),
.A2(n_582),
.B(n_175),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_656),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_683),
.A2(n_582),
.B(n_175),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_639),
.B(n_40),
.Y(n_829)
);

NOR3xp33_ASAP7_75t_L g830 ( 
.A(n_676),
.B(n_40),
.C(n_42),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_656),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_683),
.A2(n_224),
.B(n_207),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_626),
.B(n_42),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_626),
.B(n_43),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_695),
.A2(n_43),
.B(n_45),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_639),
.B(n_46),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_690),
.B(n_49),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_695),
.A2(n_50),
.B(n_51),
.Y(n_838)
);

O2A1O1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_676),
.A2(n_52),
.B(n_53),
.C(n_56),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_L g840 ( 
.A1(n_710),
.A2(n_79),
.B(n_84),
.Y(n_840)
);

OAI22xp5_ASAP7_75t_L g841 ( 
.A1(n_699),
.A2(n_664),
.B1(n_592),
.B2(n_628),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_636),
.A2(n_86),
.B(n_96),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_728),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_601),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_609),
.B(n_129),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_609),
.B(n_615),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_690),
.B(n_705),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_682),
.B(n_634),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_716),
.A2(n_705),
.B1(n_712),
.B2(n_647),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_712),
.A2(n_687),
.B(n_643),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_634),
.B(n_592),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_628),
.A2(n_606),
.B1(n_697),
.B2(n_689),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_658),
.B(n_673),
.Y(n_853)
);

NOR2xp67_ASAP7_75t_L g854 ( 
.A(n_718),
.B(n_694),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_650),
.B(n_651),
.Y(n_855)
);

AOI21x1_ASAP7_75t_L g856 ( 
.A1(n_730),
.A2(n_675),
.B(n_696),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_608),
.Y(n_857)
);

AND2x6_ASAP7_75t_L g858 ( 
.A(n_701),
.B(n_704),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_728),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_701),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_609),
.B(n_615),
.Y(n_861)
);

CKINVDCx10_ASAP7_75t_R g862 ( 
.A(n_645),
.Y(n_862)
);

NAND2xp33_ASAP7_75t_L g863 ( 
.A(n_704),
.B(n_708),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_687),
.B(n_716),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_615),
.B(n_693),
.Y(n_865)
);

AOI21xp33_ASAP7_75t_L g866 ( 
.A1(n_678),
.A2(n_665),
.B(n_659),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_700),
.B(n_708),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_613),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_730),
.A2(n_688),
.B(n_706),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_611),
.A2(n_642),
.B(n_596),
.C(n_678),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_607),
.B(n_703),
.Y(n_871)
);

AOI21x1_ASAP7_75t_L g872 ( 
.A1(n_633),
.A2(n_674),
.B(n_717),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_648),
.A2(n_671),
.B(n_719),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_611),
.B(n_680),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_649),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_657),
.A2(n_669),
.B(n_715),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_729),
.A2(n_734),
.B(n_642),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_729),
.B(n_496),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_588),
.B(n_458),
.Y(n_879)
);

AOI21x1_ASAP7_75t_L g880 ( 
.A1(n_723),
.A2(n_660),
.B(n_677),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_588),
.B(n_518),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_723),
.A2(n_660),
.B(n_677),
.Y(n_882)
);

NOR3xp33_ASAP7_75t_L g883 ( 
.A(n_588),
.B(n_456),
.C(n_445),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_667),
.B(n_496),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_588),
.B(n_458),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_588),
.B(n_458),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_679),
.A2(n_660),
.B(n_723),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_588),
.A2(n_586),
.B(n_617),
.C(n_667),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_L g889 ( 
.A1(n_588),
.A2(n_670),
.B1(n_641),
.B2(n_458),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_597),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_720),
.A2(n_660),
.B(n_702),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_588),
.B(n_518),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_588),
.B(n_518),
.Y(n_893)
);

AOI22xp5_ASAP7_75t_L g894 ( 
.A1(n_588),
.A2(n_496),
.B1(n_518),
.B2(n_625),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_588),
.A2(n_586),
.B(n_617),
.C(n_667),
.Y(n_895)
);

A2O1A1Ixp33_ASAP7_75t_L g896 ( 
.A1(n_668),
.A2(n_713),
.B(n_716),
.C(n_712),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_588),
.B(n_458),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_597),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_L g899 ( 
.A(n_588),
.B(n_518),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_594),
.B(n_666),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_660),
.A2(n_679),
.B(n_702),
.Y(n_901)
);

OR2x2_ASAP7_75t_L g902 ( 
.A(n_590),
.B(n_490),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_781),
.B(n_796),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_786),
.B(n_900),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_889),
.A2(n_901),
.B(n_768),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_879),
.B(n_885),
.Y(n_906)
);

INVx5_ASAP7_75t_L g907 ( 
.A(n_858),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_886),
.B(n_897),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_766),
.Y(n_909)
);

OAI21x1_ASAP7_75t_L g910 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_910)
);

OAI21x1_ASAP7_75t_L g911 ( 
.A1(n_880),
.A2(n_882),
.B(n_740),
.Y(n_911)
);

OAI21x1_ASAP7_75t_L g912 ( 
.A1(n_788),
.A2(n_785),
.B(n_809),
.Y(n_912)
);

NAND3xp33_ASAP7_75t_L g913 ( 
.A(n_829),
.B(n_836),
.C(n_864),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_749),
.A2(n_847),
.B1(n_850),
.B2(n_736),
.C(n_744),
.Y(n_914)
);

AO21x1_ASAP7_75t_L g915 ( 
.A1(n_866),
.A2(n_884),
.B(n_804),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_SL g916 ( 
.A1(n_745),
.A2(n_830),
.B(n_894),
.Y(n_916)
);

AO31x2_ASAP7_75t_L g917 ( 
.A1(n_787),
.A2(n_841),
.A3(n_848),
.B(n_798),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_875),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_860),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_849),
.A2(n_895),
.B(n_888),
.C(n_881),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_743),
.A2(n_738),
.B(n_769),
.Y(n_921)
);

OAI21xp33_ASAP7_75t_L g922 ( 
.A1(n_837),
.A2(n_825),
.B(n_823),
.Y(n_922)
);

OR2x6_ASAP7_75t_SL g923 ( 
.A(n_767),
.B(n_902),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_741),
.B(n_892),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_753),
.B(n_861),
.Y(n_925)
);

OAI21xp33_ASAP7_75t_L g926 ( 
.A1(n_814),
.A2(n_761),
.B(n_834),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_743),
.A2(n_738),
.B(n_752),
.Y(n_927)
);

INVx2_ASAP7_75t_SL g928 ( 
.A(n_751),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_766),
.Y(n_929)
);

A2O1A1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_893),
.A2(n_899),
.B(n_870),
.C(n_877),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_755),
.B(n_759),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_737),
.Y(n_932)
);

AOI21xp33_ASAP7_75t_L g933 ( 
.A1(n_853),
.A2(n_878),
.B(n_839),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_754),
.A2(n_748),
.B(n_792),
.Y(n_934)
);

AO31x2_ASAP7_75t_L g935 ( 
.A1(n_791),
.A2(n_874),
.A3(n_805),
.B(n_802),
.Y(n_935)
);

AO21x2_ASAP7_75t_L g936 ( 
.A1(n_783),
.A2(n_872),
.B(n_818),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_748),
.A2(n_739),
.B(n_747),
.Y(n_937)
);

AOI21xp33_ASAP7_75t_L g938 ( 
.A1(n_833),
.A2(n_855),
.B(n_851),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_739),
.A2(n_852),
.B(n_799),
.Y(n_939)
);

NAND2x1p5_ASAP7_75t_L g940 ( 
.A(n_796),
.B(n_827),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_900),
.B(n_742),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_824),
.B(n_846),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_750),
.A2(n_898),
.B1(n_890),
.B2(n_812),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_765),
.A2(n_771),
.B1(n_822),
.B2(n_806),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_865),
.B(n_801),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_818),
.A2(n_764),
.B(n_873),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_784),
.A2(n_757),
.B(n_756),
.Y(n_947)
);

NOR2xp67_ASAP7_75t_L g948 ( 
.A(n_782),
.B(n_772),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_758),
.A2(n_780),
.B(n_789),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_815),
.A2(n_817),
.B(n_845),
.C(n_779),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_780),
.A2(n_776),
.B(n_793),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_773),
.B(n_746),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_873),
.A2(n_832),
.B(n_776),
.Y(n_953)
);

AO21x2_ASAP7_75t_L g954 ( 
.A1(n_832),
.A2(n_826),
.B(n_828),
.Y(n_954)
);

AO31x2_ASAP7_75t_L g955 ( 
.A1(n_811),
.A2(n_803),
.A3(n_777),
.B(n_807),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_760),
.B(n_770),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_810),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_774),
.A2(n_775),
.B(n_863),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_844),
.B(n_827),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_778),
.A2(n_854),
.B(n_838),
.C(n_835),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_774),
.A2(n_775),
.B(n_813),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_857),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_800),
.A2(n_842),
.B(n_794),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_835),
.A2(n_838),
.B(n_820),
.C(n_840),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_831),
.B(n_859),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_876),
.A2(n_819),
.B(n_795),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_843),
.A2(n_859),
.B(n_868),
.C(n_871),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_867),
.A2(n_766),
.B(n_843),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_858),
.B(n_810),
.Y(n_969)
);

OAI21x1_ASAP7_75t_L g970 ( 
.A1(n_808),
.A2(n_858),
.B(n_816),
.Y(n_970)
);

AOI21x1_ASAP7_75t_SL g971 ( 
.A1(n_816),
.A2(n_763),
.B(n_821),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_858),
.B(n_821),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_858),
.B(n_763),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_797),
.B(n_816),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_862),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_755),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_879),
.B(n_885),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_879),
.B(n_885),
.Y(n_978)
);

AND2x2_ASAP7_75t_L g979 ( 
.A(n_902),
.B(n_619),
.Y(n_979)
);

OAI21xp5_ASAP7_75t_L g980 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_980)
);

OAI22x1_ASAP7_75t_L g981 ( 
.A1(n_849),
.A2(n_553),
.B1(n_625),
.B2(n_500),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_767),
.Y(n_982)
);

BUFx4f_ASAP7_75t_L g983 ( 
.A(n_900),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_L g984 ( 
.A1(n_745),
.A2(n_496),
.B1(n_505),
.B2(n_762),
.Y(n_984)
);

A2O1A1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_864),
.A2(n_896),
.B(n_829),
.C(n_836),
.Y(n_985)
);

NOR2xp67_ASAP7_75t_L g986 ( 
.A(n_782),
.B(n_445),
.Y(n_986)
);

AO21x1_ASAP7_75t_L g987 ( 
.A1(n_864),
.A2(n_847),
.B(n_889),
.Y(n_987)
);

OAI21xp5_ASAP7_75t_L g988 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_875),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_772),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_875),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_889),
.A2(n_901),
.B(n_679),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_751),
.Y(n_993)
);

AOI21x1_ASAP7_75t_SL g994 ( 
.A1(n_879),
.A2(n_886),
.B(n_885),
.Y(n_994)
);

OAI22x1_ASAP7_75t_L g995 ( 
.A1(n_849),
.A2(n_553),
.B1(n_625),
.B2(n_500),
.Y(n_995)
);

OAI21x1_ASAP7_75t_L g996 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_996)
);

OAI21x1_ASAP7_75t_L g997 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_860),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_767),
.Y(n_999)
);

OAI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_755),
.Y(n_1001)
);

AND3x4_ASAP7_75t_L g1002 ( 
.A(n_883),
.B(n_666),
.C(n_594),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_879),
.B(n_885),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_1005)
);

OAI21x1_ASAP7_75t_L g1006 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_864),
.A2(n_896),
.B1(n_889),
.B2(n_879),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1008)
);

BUFx2_ASAP7_75t_L g1009 ( 
.A(n_755),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_879),
.B(n_885),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_879),
.B(n_885),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_902),
.B(n_619),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_737),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_902),
.B(n_619),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_879),
.B(n_885),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_879),
.B(n_885),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_879),
.B(n_885),
.Y(n_1021)
);

OAI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_1022)
);

INVx4_ASAP7_75t_L g1023 ( 
.A(n_751),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_751),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_SL g1025 ( 
.A(n_858),
.B(n_496),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_864),
.A2(n_896),
.B1(n_889),
.B2(n_879),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_766),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_864),
.A2(n_896),
.B(n_829),
.C(n_836),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_766),
.Y(n_1031)
);

OAI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_901),
.A2(n_891),
.B(n_887),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_790),
.A2(n_869),
.B(n_856),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_746),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_1034),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_979),
.B(n_1015),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_913),
.A2(n_985),
.B(n_1028),
.C(n_916),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_969),
.B(n_956),
.Y(n_1038)
);

AOI22xp33_ASAP7_75t_L g1039 ( 
.A1(n_981),
.A2(n_995),
.B1(n_984),
.B2(n_931),
.Y(n_1039)
);

BUFx12f_ASAP7_75t_L g1040 ( 
.A(n_982),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_SL g1041 ( 
.A1(n_1025),
.A2(n_974),
.B1(n_945),
.B2(n_924),
.Y(n_1041)
);

INVx5_ASAP7_75t_L g1042 ( 
.A(n_904),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1004),
.B(n_1014),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_989),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_991),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_906),
.B(n_908),
.Y(n_1046)
);

OAI21xp33_ASAP7_75t_L g1047 ( 
.A1(n_1007),
.A2(n_1026),
.B(n_920),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_906),
.B(n_908),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_916),
.A2(n_1007),
.B1(n_1026),
.B2(n_978),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_977),
.B(n_978),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_977),
.B(n_1019),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_930),
.A2(n_922),
.B(n_914),
.C(n_933),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1019),
.A2(n_1021),
.B1(n_1020),
.B2(n_1010),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_999),
.Y(n_1054)
);

OA21x2_ASAP7_75t_L g1055 ( 
.A1(n_980),
.A2(n_1005),
.B(n_1032),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_952),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1020),
.B(n_1021),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_932),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_1017),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_969),
.B(n_972),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_983),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_983),
.Y(n_1062)
);

NAND2x1p5_ASAP7_75t_L g1063 ( 
.A(n_907),
.B(n_941),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_925),
.B(n_976),
.Y(n_1064)
);

AOI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_987),
.A2(n_915),
.B(n_933),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_957),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_926),
.B(n_938),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_1001),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1016),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_1009),
.Y(n_1070)
);

BUFx2_ASAP7_75t_R g1071 ( 
.A(n_923),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_962),
.Y(n_1072)
);

CKINVDCx20_ASAP7_75t_R g1073 ( 
.A(n_1023),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_960),
.A2(n_950),
.B(n_938),
.C(n_964),
.Y(n_1074)
);

OR2x2_ASAP7_75t_L g1075 ( 
.A(n_990),
.B(n_942),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_943),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_959),
.Y(n_1077)
);

INVxp67_ASAP7_75t_L g1078 ( 
.A(n_948),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_928),
.B(n_993),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_905),
.A2(n_1025),
.B(n_974),
.C(n_967),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_965),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1023),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_965),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_986),
.B(n_944),
.Y(n_1084)
);

AND2x2_ASAP7_75t_SL g1085 ( 
.A(n_973),
.B(n_971),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_SL g1086 ( 
.A1(n_988),
.A2(n_1003),
.B(n_1032),
.C(n_1022),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_1024),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_903),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_940),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_1002),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_975),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_L g1092 ( 
.A(n_988),
.B(n_1005),
.C(n_1003),
.Y(n_1092)
);

OR2x2_ASAP7_75t_L g1093 ( 
.A(n_909),
.B(n_1031),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_1000),
.A2(n_1022),
.B(n_1011),
.C(n_951),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_909),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_917),
.B(n_1000),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_907),
.B(n_998),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_1011),
.A2(n_951),
.B(n_927),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_934),
.A2(n_937),
.B(n_911),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_947),
.A2(n_939),
.B(n_921),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_963),
.A2(n_949),
.B(n_958),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_910),
.A2(n_1033),
.B(n_1030),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_929),
.B(n_1031),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1031),
.B(n_929),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_929),
.B(n_1027),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_1027),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_919),
.B(n_1027),
.Y(n_1107)
);

INVx8_ASAP7_75t_L g1108 ( 
.A(n_968),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_SL g1109 ( 
.A1(n_994),
.A2(n_917),
.B1(n_970),
.B2(n_912),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_961),
.B(n_954),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_966),
.A2(n_953),
.B(n_946),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_936),
.A2(n_954),
.B1(n_1029),
.B2(n_1006),
.Y(n_1112)
);

NAND2xp33_ASAP7_75t_L g1113 ( 
.A(n_935),
.B(n_955),
.Y(n_1113)
);

BUFx6f_ASAP7_75t_L g1114 ( 
.A(n_996),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_955),
.Y(n_1115)
);

O2A1O1Ixp5_ASAP7_75t_SL g1116 ( 
.A1(n_997),
.A2(n_1008),
.B(n_1012),
.C(n_1013),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1018),
.B(n_1004),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_982),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1004),
.B(n_1014),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_983),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_916),
.A2(n_913),
.B1(n_829),
.B2(n_836),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_916),
.A2(n_913),
.B1(n_829),
.B2(n_836),
.Y(n_1122)
);

INVx3_ASAP7_75t_SL g1123 ( 
.A(n_982),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_1004),
.B(n_445),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_985),
.A2(n_1028),
.B1(n_913),
.B2(n_1026),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_907),
.Y(n_1126)
);

BUFx6f_ASAP7_75t_L g1127 ( 
.A(n_983),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_969),
.B(n_956),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_952),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_913),
.A2(n_864),
.B(n_896),
.C(n_985),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_983),
.Y(n_1131)
);

BUFx4_ASAP7_75t_SL g1132 ( 
.A(n_999),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1004),
.B(n_1014),
.Y(n_1133)
);

HB1xp67_ASAP7_75t_L g1134 ( 
.A(n_979),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_985),
.A2(n_1028),
.B1(n_913),
.B2(n_1026),
.Y(n_1135)
);

AND2x4_ASAP7_75t_L g1136 ( 
.A(n_969),
.B(n_956),
.Y(n_1136)
);

OAI22xp33_ASAP7_75t_L g1137 ( 
.A1(n_913),
.A2(n_541),
.B1(n_864),
.B2(n_879),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_976),
.B(n_902),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_1034),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_985),
.A2(n_1028),
.B(n_992),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_913),
.A2(n_302),
.B1(n_315),
.B2(n_291),
.Y(n_1141)
);

NAND3xp33_ASAP7_75t_L g1142 ( 
.A(n_913),
.B(n_1028),
.C(n_985),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_932),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_969),
.B(n_956),
.Y(n_1144)
);

INVx2_ASAP7_75t_SL g1145 ( 
.A(n_983),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_985),
.A2(n_1028),
.B(n_879),
.C(n_886),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_985),
.A2(n_1028),
.B(n_992),
.Y(n_1147)
);

BUFx2_ASAP7_75t_SL g1148 ( 
.A(n_999),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_969),
.B(n_956),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_985),
.A2(n_1028),
.B(n_992),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_932),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_983),
.Y(n_1152)
);

INVx5_ASAP7_75t_L g1153 ( 
.A(n_904),
.Y(n_1153)
);

INVxp67_ASAP7_75t_L g1154 ( 
.A(n_979),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_932),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_982),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_913),
.A2(n_864),
.B(n_896),
.C(n_985),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_918),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1004),
.B(n_1014),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_907),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_983),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_1004),
.B(n_445),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_907),
.Y(n_1163)
);

INVx8_ASAP7_75t_L g1164 ( 
.A(n_1042),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_1127),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1115),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_1070),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1072),
.Y(n_1168)
);

OAI22xp33_ASAP7_75t_L g1169 ( 
.A1(n_1121),
.A2(n_1122),
.B1(n_1049),
.B2(n_1133),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_1121),
.A2(n_1122),
.B1(n_1039),
.B2(n_1141),
.Y(n_1170)
);

OAI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1130),
.A2(n_1157),
.B(n_1124),
.Y(n_1171)
);

INVx1_ASAP7_75t_SL g1172 ( 
.A(n_1138),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1058),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1162),
.A2(n_1119),
.B1(n_1159),
.B2(n_1043),
.Y(n_1174)
);

BUFx2_ASAP7_75t_L g1175 ( 
.A(n_1055),
.Y(n_1175)
);

INVx3_ASAP7_75t_L g1176 ( 
.A(n_1126),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1049),
.B(n_1076),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_1047),
.A2(n_1137),
.B1(n_1041),
.B2(n_1142),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1069),
.Y(n_1179)
);

CKINVDCx10_ASAP7_75t_R g1180 ( 
.A(n_1132),
.Y(n_1180)
);

HB1xp67_ASAP7_75t_L g1181 ( 
.A(n_1056),
.Y(n_1181)
);

AOI22xp33_ASAP7_75t_L g1182 ( 
.A1(n_1047),
.A2(n_1142),
.B1(n_1053),
.B2(n_1129),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1143),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1035),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1052),
.A2(n_1146),
.B(n_1037),
.Y(n_1185)
);

BUFx2_ASAP7_75t_L g1186 ( 
.A(n_1055),
.Y(n_1186)
);

AND2x2_ASAP7_75t_SL g1187 ( 
.A(n_1113),
.B(n_1096),
.Y(n_1187)
);

BUFx2_ASAP7_75t_R g1188 ( 
.A(n_1054),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_1139),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1151),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1050),
.B(n_1051),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1053),
.A2(n_1129),
.B1(n_1153),
.B2(n_1042),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1155),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_SL g1194 ( 
.A1(n_1125),
.A2(n_1135),
.B1(n_1153),
.B2(n_1090),
.Y(n_1194)
);

NAND2x1p5_ASAP7_75t_L g1195 ( 
.A(n_1062),
.B(n_1120),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1126),
.Y(n_1196)
);

INVx2_ASAP7_75t_SL g1197 ( 
.A(n_1093),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_1073),
.Y(n_1198)
);

OR2x6_ASAP7_75t_L g1199 ( 
.A(n_1063),
.B(n_1108),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1044),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1045),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1095),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1125),
.A2(n_1135),
.B1(n_1057),
.B2(n_1048),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1158),
.Y(n_1204)
);

CKINVDCx20_ASAP7_75t_R g1205 ( 
.A(n_1156),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1084),
.A2(n_1051),
.B1(n_1050),
.B2(n_1046),
.Y(n_1206)
);

INVx1_ASAP7_75t_SL g1207 ( 
.A(n_1075),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1077),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1067),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1140),
.A2(n_1147),
.B(n_1150),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1160),
.Y(n_1211)
);

INVx8_ASAP7_75t_L g1212 ( 
.A(n_1127),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1117),
.Y(n_1213)
);

OR2x2_ASAP7_75t_L g1214 ( 
.A(n_1092),
.B(n_1086),
.Y(n_1214)
);

INVxp67_ASAP7_75t_L g1215 ( 
.A(n_1036),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_1114),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1116),
.A2(n_1111),
.B(n_1099),
.Y(n_1217)
);

INVx3_ASAP7_75t_L g1218 ( 
.A(n_1160),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_1099),
.A2(n_1111),
.B(n_1074),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1098),
.A2(n_1065),
.B(n_1094),
.Y(n_1220)
);

INVx3_ASAP7_75t_L g1221 ( 
.A(n_1163),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1059),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1134),
.Y(n_1223)
);

CKINVDCx6p67_ASAP7_75t_R g1224 ( 
.A(n_1123),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1106),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1068),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1068),
.A2(n_1064),
.B1(n_1063),
.B2(n_1071),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1060),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1102),
.A2(n_1112),
.B(n_1098),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_L g1230 ( 
.A(n_1154),
.B(n_1083),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_1040),
.Y(n_1231)
);

BUFx8_ASAP7_75t_SL g1232 ( 
.A(n_1118),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1103),
.B(n_1105),
.Y(n_1233)
);

OAI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1062),
.A2(n_1120),
.B1(n_1066),
.B2(n_1061),
.Y(n_1234)
);

AO21x1_ASAP7_75t_SL g1235 ( 
.A1(n_1088),
.A2(n_1089),
.B(n_1109),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1079),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1109),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1080),
.A2(n_1085),
.B1(n_1145),
.B2(n_1152),
.Y(n_1238)
);

CKINVDCx11_ASAP7_75t_R g1239 ( 
.A(n_1082),
.Y(n_1239)
);

AOI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1038),
.A2(n_1128),
.B1(n_1136),
.B2(n_1144),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1110),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1091),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1104),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1081),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1078),
.A2(n_1038),
.B1(n_1128),
.B2(n_1136),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1131),
.A2(n_1161),
.B1(n_1148),
.B2(n_1087),
.Y(n_1246)
);

BUFx4f_ASAP7_75t_L g1247 ( 
.A(n_1131),
.Y(n_1247)
);

BUFx12f_ASAP7_75t_SL g1248 ( 
.A(n_1131),
.Y(n_1248)
);

AO21x1_ASAP7_75t_SL g1249 ( 
.A1(n_1108),
.A2(n_1163),
.B(n_1097),
.Y(n_1249)
);

BUFx2_ASAP7_75t_L g1250 ( 
.A(n_1095),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1144),
.B(n_1149),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1149),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1161),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1107),
.B(n_1096),
.Y(n_1254)
);

HB1xp67_ASAP7_75t_L g1255 ( 
.A(n_1070),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1072),
.Y(n_1256)
);

BUFx12f_ASAP7_75t_L g1257 ( 
.A(n_1054),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1072),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1127),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1072),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1035),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1121),
.A2(n_995),
.B1(n_981),
.B2(n_984),
.Y(n_1262)
);

INVx6_ASAP7_75t_L g1263 ( 
.A(n_1062),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1116),
.A2(n_1100),
.B(n_1101),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1042),
.B(n_1153),
.Y(n_1265)
);

OAI22xp5_ASAP7_75t_L g1266 ( 
.A1(n_1121),
.A2(n_1122),
.B1(n_913),
.B2(n_1049),
.Y(n_1266)
);

CKINVDCx14_ASAP7_75t_R g1267 ( 
.A(n_1054),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1072),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_1095),
.Y(n_1270)
);

BUFx3_ASAP7_75t_L g1271 ( 
.A(n_1035),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1054),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1166),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1177),
.B(n_1241),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1177),
.B(n_1241),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1254),
.Y(n_1276)
);

BUFx2_ASAP7_75t_L g1277 ( 
.A(n_1175),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1171),
.A2(n_1266),
.B(n_1185),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1175),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1280)
);

INVx2_ASAP7_75t_SL g1281 ( 
.A(n_1254),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1174),
.B(n_1198),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1216),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1226),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1169),
.A2(n_1178),
.B(n_1210),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1167),
.Y(n_1286)
);

HB1xp67_ASAP7_75t_L g1287 ( 
.A(n_1255),
.Y(n_1287)
);

BUFx2_ASAP7_75t_L g1288 ( 
.A(n_1186),
.Y(n_1288)
);

OR2x2_ASAP7_75t_L g1289 ( 
.A(n_1214),
.B(n_1213),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1198),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1203),
.B(n_1172),
.Y(n_1291)
);

AND3x1_ASAP7_75t_L g1292 ( 
.A(n_1170),
.B(n_1262),
.C(n_1182),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1187),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1237),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1272),
.B(n_1205),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1237),
.B(n_1214),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1209),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1173),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1219),
.B(n_1179),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1199),
.A2(n_1238),
.B(n_1265),
.Y(n_1300)
);

BUFx8_ASAP7_75t_L g1301 ( 
.A(n_1257),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1219),
.B(n_1183),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1181),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1219),
.B(n_1190),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1193),
.Y(n_1305)
);

OR2x2_ASAP7_75t_L g1306 ( 
.A(n_1207),
.B(n_1222),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1233),
.B(n_1220),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1264),
.A2(n_1217),
.B(n_1229),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_R g1309 ( 
.A(n_1180),
.B(n_1236),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_L g1310 ( 
.A(n_1272),
.B(n_1205),
.Y(n_1310)
);

OR2x2_ASAP7_75t_L g1311 ( 
.A(n_1223),
.B(n_1220),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1164),
.A2(n_1251),
.B1(n_1194),
.B2(n_1252),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1233),
.B(n_1208),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1235),
.B(n_1228),
.Y(n_1314)
);

OR2x2_ASAP7_75t_L g1315 ( 
.A(n_1197),
.B(n_1243),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1168),
.Y(n_1316)
);

INVxp67_ASAP7_75t_L g1317 ( 
.A(n_1230),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1256),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1258),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1260),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_SL g1321 ( 
.A(n_1234),
.B(n_1227),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1176),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1225),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1235),
.B(n_1215),
.Y(n_1324)
);

AND2x4_ASAP7_75t_L g1325 ( 
.A(n_1252),
.B(n_1251),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1176),
.A2(n_1211),
.B(n_1269),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1268),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1197),
.B(n_1243),
.Y(n_1328)
);

OR2x2_ASAP7_75t_L g1329 ( 
.A(n_1250),
.B(n_1192),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1176),
.B(n_1221),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1196),
.A2(n_1211),
.B(n_1218),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1247),
.A2(n_1246),
.B(n_1195),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1200),
.A2(n_1204),
.B1(n_1201),
.B2(n_1244),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1196),
.B(n_1221),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1164),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1267),
.B(n_1188),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1196),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1211),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1218),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1307),
.B(n_1271),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1307),
.B(n_1249),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1277),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_1311),
.Y(n_1343)
);

HB1xp67_ASAP7_75t_L g1344 ( 
.A(n_1277),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1279),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1299),
.B(n_1218),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1299),
.B(n_1270),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1302),
.B(n_1202),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1279),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1296),
.B(n_1271),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1302),
.B(n_1240),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1304),
.B(n_1184),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1298),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1288),
.Y(n_1354)
);

OAI211xp5_ASAP7_75t_L g1355 ( 
.A1(n_1278),
.A2(n_1239),
.B(n_1267),
.C(n_1236),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1311),
.B(n_1189),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1313),
.B(n_1261),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1296),
.B(n_1261),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1289),
.B(n_1189),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1313),
.B(n_1274),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1309),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1289),
.B(n_1224),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1274),
.B(n_1224),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1286),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1275),
.B(n_1245),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1294),
.Y(n_1366)
);

OAI221xp5_ASAP7_75t_L g1367 ( 
.A1(n_1285),
.A2(n_1195),
.B1(n_1247),
.B2(n_1263),
.C(n_1231),
.Y(n_1367)
);

AOI21xp33_ASAP7_75t_L g1368 ( 
.A1(n_1291),
.A2(n_1282),
.B(n_1294),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1292),
.A2(n_1263),
.B1(n_1242),
.B2(n_1231),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1287),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1292),
.A2(n_1248),
.B1(n_1257),
.B2(n_1253),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1273),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1364),
.B(n_1303),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1360),
.B(n_1293),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1360),
.B(n_1293),
.Y(n_1375)
);

NAND3xp33_ASAP7_75t_L g1376 ( 
.A(n_1369),
.B(n_1323),
.C(n_1284),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1364),
.B(n_1306),
.Y(n_1377)
);

NAND3xp33_ASAP7_75t_L g1378 ( 
.A(n_1368),
.B(n_1297),
.C(n_1280),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1352),
.B(n_1276),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1372),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1352),
.B(n_1281),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1369),
.A2(n_1321),
.B1(n_1325),
.B2(n_1312),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1370),
.B(n_1306),
.Y(n_1383)
);

NOR3xp33_ASAP7_75t_L g1384 ( 
.A(n_1367),
.B(n_1332),
.C(n_1322),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1370),
.B(n_1317),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_L g1386 ( 
.A(n_1368),
.B(n_1371),
.C(n_1366),
.Y(n_1386)
);

NAND3xp33_ASAP7_75t_L g1387 ( 
.A(n_1371),
.B(n_1297),
.C(n_1305),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1352),
.B(n_1281),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1366),
.B(n_1305),
.Y(n_1389)
);

NAND3xp33_ASAP7_75t_L g1390 ( 
.A(n_1367),
.B(n_1338),
.C(n_1337),
.Y(n_1390)
);

NAND3xp33_ASAP7_75t_L g1391 ( 
.A(n_1359),
.B(n_1338),
.C(n_1337),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1341),
.B(n_1324),
.Y(n_1392)
);

AOI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1343),
.A2(n_1319),
.B1(n_1318),
.B2(n_1316),
.C(n_1327),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_SL g1394 ( 
.A1(n_1355),
.A2(n_1324),
.B(n_1336),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1372),
.Y(n_1395)
);

AOI221xp5_ASAP7_75t_L g1396 ( 
.A1(n_1343),
.A2(n_1327),
.B1(n_1320),
.B2(n_1318),
.C(n_1316),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1341),
.B(n_1339),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1359),
.B(n_1308),
.C(n_1339),
.Y(n_1398)
);

OAI221xp5_ASAP7_75t_SL g1399 ( 
.A1(n_1362),
.A2(n_1290),
.B1(n_1300),
.B2(n_1314),
.C(n_1329),
.Y(n_1399)
);

OAI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1355),
.A2(n_1326),
.B(n_1331),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_SL g1401 ( 
.A1(n_1341),
.A2(n_1310),
.B(n_1295),
.Y(n_1401)
);

NAND4xp25_ASAP7_75t_L g1402 ( 
.A(n_1342),
.B(n_1334),
.C(n_1330),
.D(n_1322),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_1356),
.B(n_1339),
.C(n_1328),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1340),
.B(n_1283),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_R g1405 ( 
.A(n_1361),
.B(n_1242),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1356),
.A2(n_1326),
.B(n_1331),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_SL g1407 ( 
.A(n_1362),
.B(n_1335),
.Y(n_1407)
);

NAND4xp25_ASAP7_75t_L g1408 ( 
.A(n_1342),
.B(n_1322),
.C(n_1315),
.D(n_1333),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1357),
.B(n_1350),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1357),
.B(n_1350),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1357),
.B(n_1315),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1358),
.B(n_1319),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1380),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1406),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1380),
.Y(n_1415)
);

NAND2xp5_ASAP7_75t_L g1416 ( 
.A(n_1395),
.B(n_1343),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1378),
.A2(n_1365),
.B1(n_1351),
.B2(n_1363),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1395),
.B(n_1353),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1389),
.Y(n_1419)
);

NOR2x1_ASAP7_75t_L g1420 ( 
.A(n_1376),
.B(n_1358),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_1405),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1374),
.B(n_1346),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1377),
.B(n_1342),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1397),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1383),
.B(n_1349),
.Y(n_1425)
);

NAND3xp33_ASAP7_75t_L g1426 ( 
.A(n_1386),
.B(n_1344),
.C(n_1345),
.Y(n_1426)
);

HB1xp67_ASAP7_75t_L g1427 ( 
.A(n_1391),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1373),
.B(n_1349),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1398),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1393),
.B(n_1353),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1412),
.B(n_1349),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1375),
.Y(n_1432)
);

INVx2_ASAP7_75t_SL g1433 ( 
.A(n_1397),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1391),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1403),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1398),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1385),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1400),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_1390),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1404),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1396),
.B(n_1353),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1379),
.B(n_1347),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1402),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1379),
.B(n_1347),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1381),
.B(n_1348),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1428),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1430),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1413),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1435),
.B(n_1408),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1430),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1441),
.Y(n_1451)
);

NAND2x1_ASAP7_75t_L g1452 ( 
.A(n_1420),
.B(n_1392),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1443),
.B(n_1392),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1439),
.B(n_1376),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1441),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1419),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1419),
.Y(n_1457)
);

INVxp33_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

NAND3xp33_ASAP7_75t_L g1459 ( 
.A(n_1439),
.B(n_1436),
.C(n_1438),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1437),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1437),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1418),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1418),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1435),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1443),
.B(n_1381),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1443),
.B(n_1388),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1413),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1439),
.B(n_1411),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1415),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1439),
.B(n_1409),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1415),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1415),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1434),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1434),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1434),
.B(n_1410),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1427),
.B(n_1344),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1428),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1423),
.B(n_1386),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_1427),
.B(n_1345),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1422),
.B(n_1388),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1422),
.B(n_1363),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1436),
.B(n_1354),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1428),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1431),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1436),
.B(n_1354),
.Y(n_1485)
);

NAND3xp33_ASAP7_75t_L g1486 ( 
.A(n_1459),
.B(n_1429),
.C(n_1438),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1454),
.B(n_1438),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1469),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1454),
.B(n_1453),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1454),
.B(n_1414),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1453),
.B(n_1414),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1447),
.B(n_1429),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1471),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1472),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1450),
.B(n_1414),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1451),
.A2(n_1426),
.B(n_1417),
.C(n_1394),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1465),
.B(n_1422),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1452),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1455),
.B(n_1426),
.Y(n_1499)
);

OR2x2_ASAP7_75t_L g1500 ( 
.A(n_1475),
.B(n_1423),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1475),
.B(n_1423),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1460),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1464),
.B(n_1425),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_SL g1504 ( 
.A(n_1458),
.B(n_1417),
.C(n_1401),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1461),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1473),
.B(n_1431),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1446),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1474),
.B(n_1413),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1477),
.B(n_1483),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1456),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1452),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1465),
.B(n_1442),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1478),
.B(n_1425),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1458),
.B(n_1478),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1484),
.B(n_1425),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1457),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1466),
.B(n_1442),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1446),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1448),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1448),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1467),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1466),
.B(n_1442),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1481),
.B(n_1444),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1481),
.B(n_1444),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1449),
.B(n_1421),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1462),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1463),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1467),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1525),
.B(n_1421),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1504),
.A2(n_1449),
.B1(n_1387),
.B2(n_1468),
.Y(n_1530)
);

INVx4_ASAP7_75t_L g1531 ( 
.A(n_1487),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1523),
.B(n_1524),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1490),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1489),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1523),
.B(n_1480),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1488),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1490),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1524),
.B(n_1480),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1486),
.A2(n_1387),
.B1(n_1468),
.B2(n_1470),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1512),
.B(n_1476),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1512),
.B(n_1479),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1489),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1517),
.B(n_1485),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1492),
.B(n_1502),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1517),
.B(n_1482),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1488),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1486),
.A2(n_1470),
.B1(n_1382),
.B2(n_1390),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1522),
.B(n_1444),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1493),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1492),
.B(n_1413),
.Y(n_1550)
);

OR2x2_ASAP7_75t_L g1551 ( 
.A(n_1499),
.B(n_1431),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1493),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1522),
.B(n_1445),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1494),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1494),
.Y(n_1555)
);

BUFx2_ASAP7_75t_L g1556 ( 
.A(n_1487),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1502),
.B(n_1432),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1499),
.B(n_1416),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1505),
.Y(n_1559)
);

NOR2x1_ASAP7_75t_L g1560 ( 
.A(n_1514),
.B(n_1496),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1498),
.B(n_1384),
.Y(n_1561)
);

INVxp67_ASAP7_75t_L g1562 ( 
.A(n_1507),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1507),
.Y(n_1563)
);

BUFx3_ASAP7_75t_L g1564 ( 
.A(n_1507),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1536),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1536),
.Y(n_1566)
);

O2A1O1Ixp33_ASAP7_75t_L g1567 ( 
.A1(n_1560),
.A2(n_1495),
.B(n_1491),
.C(n_1518),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1546),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1546),
.Y(n_1569)
);

OAI21xp5_ASAP7_75t_L g1570 ( 
.A1(n_1560),
.A2(n_1530),
.B(n_1539),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1534),
.B(n_1491),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1561),
.A2(n_1495),
.B1(n_1498),
.B2(n_1511),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.B(n_1497),
.Y(n_1573)
);

AOI221xp5_ASAP7_75t_L g1574 ( 
.A1(n_1530),
.A2(n_1528),
.B1(n_1519),
.B2(n_1520),
.C(n_1521),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1549),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_L g1576 ( 
.A1(n_1547),
.A2(n_1528),
.B1(n_1519),
.B2(n_1521),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1534),
.B(n_1513),
.Y(n_1577)
);

OAI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1531),
.A2(n_1513),
.B1(n_1511),
.B2(n_1501),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1542),
.Y(n_1579)
);

AOI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1539),
.A2(n_1508),
.B(n_1518),
.Y(n_1580)
);

OAI32xp33_ASAP7_75t_L g1581 ( 
.A1(n_1547),
.A2(n_1518),
.A3(n_1503),
.B1(n_1501),
.B2(n_1500),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1556),
.B(n_1497),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1532),
.A2(n_1508),
.B(n_1500),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1549),
.Y(n_1584)
);

OAI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1544),
.A2(n_1506),
.B1(n_1528),
.B2(n_1519),
.C(n_1521),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1552),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1556),
.B(n_1503),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1529),
.B(n_1361),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_SL g1589 ( 
.A1(n_1564),
.A2(n_1520),
.B1(n_1516),
.B2(n_1505),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1544),
.A2(n_1520),
.B1(n_1526),
.B2(n_1527),
.C(n_1516),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1577),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1565),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1566),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1568),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1570),
.A2(n_1537),
.B1(n_1531),
.B2(n_1533),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1567),
.B(n_1533),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1567),
.B(n_1564),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1571),
.B(n_1551),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1569),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1588),
.B(n_1531),
.Y(n_1601)
);

NOR2x2_ASAP7_75t_L g1602 ( 
.A(n_1579),
.B(n_1531),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1575),
.Y(n_1603)
);

OAI222xp33_ASAP7_75t_L g1604 ( 
.A1(n_1576),
.A2(n_1531),
.B1(n_1562),
.B2(n_1551),
.C1(n_1558),
.C2(n_1537),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1582),
.B(n_1537),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1572),
.B(n_1537),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1587),
.B(n_1564),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1537),
.Y(n_1608)
);

AOI22xp33_ASAP7_75t_L g1609 ( 
.A1(n_1574),
.A2(n_1563),
.B1(n_1562),
.B2(n_1559),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1583),
.A2(n_1589),
.B1(n_1580),
.B2(n_1585),
.Y(n_1610)
);

NAND3x1_ASAP7_75t_SL g1611 ( 
.A(n_1605),
.B(n_1590),
.C(n_1232),
.Y(n_1611)
);

AOI211xp5_ASAP7_75t_L g1612 ( 
.A1(n_1604),
.A2(n_1581),
.B(n_1578),
.C(n_1563),
.Y(n_1612)
);

NAND3xp33_ASAP7_75t_L g1613 ( 
.A(n_1610),
.B(n_1589),
.C(n_1586),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1603),
.Y(n_1614)
);

NOR3xp33_ASAP7_75t_L g1615 ( 
.A(n_1598),
.B(n_1584),
.C(n_1550),
.Y(n_1615)
);

OAI221xp5_ASAP7_75t_L g1616 ( 
.A1(n_1609),
.A2(n_1558),
.B1(n_1551),
.B2(n_1550),
.C(n_1559),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1599),
.B(n_1532),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1608),
.A2(n_1552),
.B1(n_1555),
.B2(n_1554),
.C(n_1558),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_SL g1619 ( 
.A(n_1601),
.B(n_1232),
.Y(n_1619)
);

AND3x1_ASAP7_75t_L g1620 ( 
.A(n_1606),
.B(n_1532),
.C(n_1535),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1596),
.B(n_1535),
.Y(n_1621)
);

AOI221xp5_ASAP7_75t_L g1622 ( 
.A1(n_1597),
.A2(n_1555),
.B1(n_1554),
.B2(n_1510),
.C(n_1527),
.Y(n_1622)
);

INVxp67_ASAP7_75t_SL g1623 ( 
.A(n_1612),
.Y(n_1623)
);

NOR3x1_ASAP7_75t_L g1624 ( 
.A(n_1613),
.B(n_1607),
.C(n_1595),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1619),
.B(n_1601),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1616),
.A2(n_1609),
.B(n_1591),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_SL g1627 ( 
.A(n_1615),
.B(n_1603),
.C(n_1593),
.Y(n_1627)
);

NOR3x1_ASAP7_75t_L g1628 ( 
.A(n_1621),
.B(n_1617),
.C(n_1614),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1620),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1618),
.B(n_1535),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_L g1631 ( 
.A(n_1611),
.B(n_1594),
.C(n_1592),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1622),
.B(n_1600),
.Y(n_1632)
);

AND4x1_ASAP7_75t_L g1633 ( 
.A(n_1628),
.B(n_1602),
.C(n_1301),
.D(n_1538),
.Y(n_1633)
);

NAND4xp25_ASAP7_75t_L g1634 ( 
.A(n_1624),
.B(n_1541),
.C(n_1540),
.D(n_1543),
.Y(n_1634)
);

OAI211xp5_ASAP7_75t_SL g1635 ( 
.A1(n_1623),
.A2(n_1239),
.B(n_1509),
.C(n_1557),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1632),
.Y(n_1636)
);

AOI211x1_ASAP7_75t_SL g1637 ( 
.A1(n_1626),
.A2(n_1557),
.B(n_1540),
.C(n_1541),
.Y(n_1637)
);

AOI211xp5_ASAP7_75t_SL g1638 ( 
.A1(n_1625),
.A2(n_1629),
.B(n_1627),
.C(n_1631),
.Y(n_1638)
);

AOI222xp33_ASAP7_75t_L g1639 ( 
.A1(n_1630),
.A2(n_1510),
.B1(n_1526),
.B2(n_1545),
.C1(n_1543),
.C2(n_1541),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1636),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1633),
.A2(n_1509),
.B1(n_1540),
.B2(n_1515),
.Y(n_1641)
);

NOR2x1_ASAP7_75t_L g1642 ( 
.A(n_1634),
.B(n_1543),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1639),
.Y(n_1643)
);

AOI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1635),
.A2(n_1545),
.B1(n_1538),
.B2(n_1553),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1637),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1638),
.B(n_1545),
.Y(n_1646)
);

NOR2x1_ASAP7_75t_L g1647 ( 
.A(n_1640),
.B(n_1301),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1642),
.B(n_1538),
.Y(n_1648)
);

NOR3xp33_ASAP7_75t_SL g1649 ( 
.A(n_1646),
.B(n_1643),
.C(n_1645),
.Y(n_1649)
);

AOI22xp33_ASAP7_75t_SL g1650 ( 
.A1(n_1641),
.A2(n_1301),
.B1(n_1553),
.B2(n_1548),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1644),
.B(n_1548),
.Y(n_1651)
);

XOR2x2_ASAP7_75t_L g1652 ( 
.A(n_1647),
.B(n_1301),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1648),
.Y(n_1653)
);

INVx2_ASAP7_75t_L g1654 ( 
.A(n_1651),
.Y(n_1654)
);

OA22x2_ASAP7_75t_L g1655 ( 
.A1(n_1654),
.A2(n_1649),
.B1(n_1650),
.B2(n_1553),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1655),
.B(n_1654),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1656),
.A2(n_1653),
.B1(n_1652),
.B2(n_1548),
.Y(n_1657)
);

OAI211xp5_ASAP7_75t_L g1658 ( 
.A1(n_1656),
.A2(n_1515),
.B(n_1363),
.C(n_1440),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_1657),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1658),
.A2(n_1416),
.B(n_1407),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1659),
.A2(n_1660),
.B(n_1247),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1659),
.B(n_1424),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_SL g1663 ( 
.A1(n_1661),
.A2(n_1433),
.B(n_1424),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1663),
.Y(n_1664)
);

OAI221xp5_ASAP7_75t_R g1665 ( 
.A1(n_1664),
.A2(n_1662),
.B1(n_1440),
.B2(n_1212),
.C(n_1433),
.Y(n_1665)
);

AOI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1399),
.B(n_1165),
.C(n_1259),
.Y(n_1666)
);


endmodule