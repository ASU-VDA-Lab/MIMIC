module real_jpeg_25978_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_1),
.A2(n_45),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_1),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_174),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_174),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_1),
.A2(n_67),
.B1(n_70),
.B2(n_174),
.Y(n_300)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_3),
.A2(n_46),
.B1(n_58),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_3),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_3),
.A2(n_33),
.B1(n_34),
.B2(n_80),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_80),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_3),
.A2(n_67),
.B1(n_70),
.B2(n_80),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_4),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_7),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_57),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_7),
.A2(n_57),
.B1(n_67),
.B2(n_70),
.Y(n_133)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_9),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_88),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_88),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_9),
.A2(n_67),
.B1(n_70),
.B2(n_88),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_10),
.A2(n_53),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_10),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_119),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_119),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_10),
.A2(n_67),
.B1(n_70),
.B2(n_119),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_11),
.B(n_175),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_11),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_11),
.B(n_55),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_11),
.B(n_28),
.C(n_30),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_228),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_11),
.B(n_37),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_228),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_11),
.B(n_67),
.C(n_69),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_11),
.A2(n_101),
.B(n_287),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_12),
.A2(n_44),
.B1(n_53),
.B2(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_12),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_145),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_145),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_12),
.A2(n_67),
.B1(n_70),
.B2(n_145),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_40),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_14),
.A2(n_40),
.B1(n_67),
.B2(n_70),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_15),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_15),
.A2(n_33),
.B1(n_34),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_48),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_15),
.A2(n_48),
.B1(n_67),
.B2(n_70),
.Y(n_183)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_16),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_95),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_94),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_21),
.B(n_81),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_41),
.B1(n_61),
.B2(n_62),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_23),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_37),
.B(n_38),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_37),
.B1(n_91),
.B2(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_24),
.B(n_179),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_24),
.A2(n_37),
.B1(n_193),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_25),
.A2(n_26),
.B1(n_39),
.B2(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_25),
.A2(n_26),
.B1(n_92),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_25),
.A2(n_26),
.B1(n_123),
.B2(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_25),
.A2(n_192),
.B(n_194),
.Y(n_191)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_25),
.A2(n_194),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_26),
.A2(n_141),
.B(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_26),
.A2(n_178),
.B(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_27),
.A2(n_28),
.B1(n_68),
.B2(n_69),
.Y(n_72)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_28),
.B(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_34),
.B1(n_51),
.B2(n_52),
.Y(n_55)
);

AOI32xp33_ASAP7_75t_L g196 ( 
.A1(n_33),
.A2(n_47),
.A3(n_52),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp33_ASAP7_75t_SL g198 ( 
.A(n_34),
.B(n_51),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_34),
.B(n_253),
.Y(n_252)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_37),
.B(n_179),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.B1(n_55),
.B2(n_56),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_54),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx8_ASAP7_75t_L g175 ( 
.A(n_47),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_47),
.A2(n_228),
.B(n_229),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_49),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_49),
.A2(n_55),
.B1(n_144),
.B2(n_173),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_49),
.A2(n_147),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_53),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_54),
.A2(n_78),
.B1(n_79),
.B2(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_54),
.A2(n_87),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_54),
.B(n_117),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_54),
.A2(n_115),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_75),
.C(n_77),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_75),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_86),
.C(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_64),
.A2(n_85),
.B1(n_90),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_71),
.B(n_73),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_65),
.A2(n_71),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_65),
.A2(n_71),
.B1(n_109),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_65),
.A2(n_71),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_65),
.B(n_225),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_66),
.A2(n_74),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_66),
.A2(n_125),
.B1(n_139),
.B2(n_185),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_66),
.A2(n_185),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_66),
.A2(n_224),
.B(n_260),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_66),
.B(n_228),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_66)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_67),
.B(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_70),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_71),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_143),
.B(n_146),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.C(n_89),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_82),
.A2(n_86),
.B1(n_157),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_86),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_86),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_89),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI31xp33_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_158),
.A3(n_164),
.B(n_343),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_148),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_97),
.B(n_148),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_120),
.C(n_128),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_98),
.A2(n_120),
.B1(n_121),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_98),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_111),
.Y(n_98)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_100),
.B(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_100),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_100),
.A2(n_107),
.B1(n_108),
.B2(n_112),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B(n_106),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_106),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_101),
.A2(n_103),
.B1(n_133),
.B2(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_101),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_101),
.A2(n_202),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_101),
.B(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_101),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_102),
.Y(n_288)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_105),
.B(n_228),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_110),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_124),
.B(n_127),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_122),
.B(n_124),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_125),
.A2(n_274),
.B(n_275),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_125),
.A2(n_275),
.B(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_128),
.A2(n_129),
.B1(n_338),
.B2(n_340),
.Y(n_337)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.C(n_142),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_130),
.A2(n_131),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_136),
.B1(n_137),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_135),
.A2(n_200),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_140),
.B(n_142),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_151),
.C(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_159),
.A2(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_160),
.B(n_163),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_336),
.B(n_342),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_213),
.B(n_335),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_206),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_167),
.B(n_206),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_186),
.C(n_188),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_168),
.A2(n_169),
.B1(n_186),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_176),
.B2(n_177),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_176),
.C(n_180),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_173),
.Y(n_190)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_181),
.B(n_184),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_199)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_186),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_188),
.B(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_195),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_189),
.B(n_191),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_195),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_196),
.B(n_199),
.Y(n_230)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_203),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_208),
.B(n_209),
.C(n_212),
.Y(n_341)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_245),
.B(n_329),
.C(n_334),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_239),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_239),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_230),
.C(n_231),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_216),
.A2(n_217),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_222),
.C(n_226),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_230),
.B(n_231),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.C(n_236),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_269),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_237),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_238),
.A2(n_300),
.B(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_240),
.B(n_243),
.C(n_244),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_323),
.B(n_328),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_276),
.B(n_322),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_265),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_250),
.B(n_265),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_258),
.C(n_262),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_251),
.B(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_256),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_257),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_258),
.A2(n_262),
.B1(n_263),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_258),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_261),
.Y(n_274)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_270),
.B2(n_271),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_272),
.C(n_273),
.Y(n_327)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_316),
.B(n_321),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_296),
.B(n_315),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_290),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_290),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_285),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_284),
.C(n_285),
.Y(n_320)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_291),
.A2(n_292),
.B1(n_294),
.B2(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_294),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_304),
.B(n_314),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_302),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_309),
.B(n_313),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_320),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_320),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_331),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_330),
.B(n_331),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_341),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_337),
.B(n_341),
.Y(n_342)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_338),
.Y(n_340)
);


endmodule