module fake_netlist_6_973_n_2168 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2168);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2168;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_541;
wire n_512;
wire n_2073;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_2083;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_2081;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_2112;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_570;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_33),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_122),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_108),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_124),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_142),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_208),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_31),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_30),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_118),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_185),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_109),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_153),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_4),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_9),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_7),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_138),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_166),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_128),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_180),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

CKINVDCx12_ASAP7_75t_R g239 ( 
.A(n_148),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_146),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_91),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_200),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_154),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_6),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_55),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_53),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_204),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_116),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_53),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_6),
.Y(n_250)
);

BUFx10_ASAP7_75t_L g251 ( 
.A(n_33),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_133),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_192),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_40),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_68),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_64),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_161),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_0),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_106),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_55),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_83),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_81),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_164),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_71),
.Y(n_267)
);

BUFx8_ASAP7_75t_SL g268 ( 
.A(n_64),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_127),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_28),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_25),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_156),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_63),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_51),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_58),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_78),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_193),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_169),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_201),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_8),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_76),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_140),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_190),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_178),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_69),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_45),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_159),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_15),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_15),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_9),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_2),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_104),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_94),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_63),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_96),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_211),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_26),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_175),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_147),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_205),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_32),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_34),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_176),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_141),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_198),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_110),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_143),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_173),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_144),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_194),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_89),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_135),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_69),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_93),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_132),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_39),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_77),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_98),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_112),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_111),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_10),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_36),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_196),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_172),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_38),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_26),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_71),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_67),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_126),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_38),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_137),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_11),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_188),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_199),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_187),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_48),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_22),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_101),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_125),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_50),
.Y(n_342)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_203),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_87),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_120),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_72),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_28),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_113),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_165),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_52),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_25),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_158),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_129),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_130),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_179),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_162),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_170),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_107),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_20),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_19),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_131),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_4),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_207),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_65),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_42),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_57),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_1),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_119),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_16),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_24),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_82),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_195),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_121),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_44),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_61),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_41),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_99),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_56),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_149),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_160),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_206),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_74),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_102),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_49),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_100),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_72),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_19),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_134),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_2),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_186),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_115),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_21),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_16),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_60),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_43),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_20),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_23),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_49),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_85),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_24),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_44),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_22),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_88),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_105),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_5),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_155),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_57),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_42),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_171),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_90),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_114),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g413 ( 
.A(n_136),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_56),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_27),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_47),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_46),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_12),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_48),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_65),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_117),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_79),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_1),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_151),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_21),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_270),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_254),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_270),
.Y(n_428)
);

INVxp33_ASAP7_75t_L g429 ( 
.A(n_395),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_270),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_270),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_270),
.Y(n_432)
);

INVx3_ASAP7_75t_L g433 ( 
.A(n_270),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_259),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_268),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_405),
.B(n_3),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_217),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_259),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_287),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_220),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_279),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_287),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_376),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

CKINVDCx14_ASAP7_75t_R g445 ( 
.A(n_405),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_218),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_413),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_224),
.B(n_3),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_224),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_221),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_266),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_288),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_228),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_230),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_254),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_332),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_245),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_307),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_245),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_234),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_378),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_378),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_246),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_394),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_304),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_415),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_235),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_380),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_246),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_292),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_292),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_292),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_295),
.Y(n_475)
);

INVxp67_ASAP7_75t_SL g476 ( 
.A(n_413),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_406),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_236),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_227),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_227),
.B(n_7),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_237),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_382),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_295),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_240),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_400),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_252),
.B(n_8),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_315),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_315),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_241),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_324),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_332),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_324),
.Y(n_492)
);

INVxp33_ASAP7_75t_L g493 ( 
.A(n_328),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_251),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_242),
.Y(n_495)
);

NOR2xp67_ASAP7_75t_L g496 ( 
.A(n_379),
.B(n_10),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_247),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_248),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_253),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_257),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_219),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_328),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_260),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_269),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_272),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_329),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_277),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_300),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g509 ( 
.A(n_223),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_329),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_280),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_252),
.B(n_12),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_334),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_282),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_283),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_339),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_262),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_284),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_262),
.B(n_13),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_285),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_339),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_346),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_346),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_R g524 ( 
.A(n_293),
.B(n_213),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_350),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_296),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_299),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_350),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_359),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_379),
.A2(n_297),
.B(n_263),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_379),
.B(n_13),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_301),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_359),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_306),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_310),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_508),
.B(n_311),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_431),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_431),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_433),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_433),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_530),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_426),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_426),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_530),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_428),
.Y(n_546)
);

OR2x6_ASAP7_75t_L g547 ( 
.A(n_496),
.B(n_300),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

BUFx8_ASAP7_75t_L g549 ( 
.A(n_448),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_472),
.B(n_300),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_430),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_430),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_432),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_432),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_472),
.B(n_309),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_436),
.B(n_229),
.Y(n_556)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_445),
.Y(n_557)
);

NAND2x1_ASAP7_75t_L g558 ( 
.A(n_531),
.B(n_379),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_455),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_475),
.Y(n_560)
);

AND3x2_ASAP7_75t_L g561 ( 
.A(n_448),
.B(n_297),
.C(n_263),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_475),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_483),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_479),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_479),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_517),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_437),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_434),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_476),
.B(n_312),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_473),
.A2(n_392),
.B(n_336),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_434),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_438),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_427),
.B(n_229),
.Y(n_575)
);

OA21x2_ASAP7_75t_L g576 ( 
.A1(n_438),
.A2(n_265),
.B(n_264),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_480),
.B(n_229),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_487),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_439),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_439),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g581 ( 
.A(n_440),
.Y(n_581)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_456),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_442),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_491),
.B(n_251),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_442),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_443),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_441),
.B(n_215),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_487),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_491),
.B(n_251),
.Y(n_589)
);

OAI21x1_ASAP7_75t_L g590 ( 
.A1(n_473),
.A2(n_392),
.B(n_336),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g591 ( 
.A(n_452),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_447),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_477),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_474),
.B(n_309),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_443),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_444),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_444),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_477),
.B(n_406),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_488),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_490),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_501),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_461),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_474),
.B(n_309),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_461),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_447),
.B(n_341),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_462),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_490),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_509),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_492),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_449),
.Y(n_611)
);

NOR3xp33_ASAP7_75t_L g612 ( 
.A(n_486),
.B(n_347),
.C(n_261),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_446),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_492),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_502),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_462),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_464),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_502),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_450),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_464),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_465),
.B(n_467),
.Y(n_621)
);

BUFx8_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

NAND2xp33_ASAP7_75t_L g623 ( 
.A(n_524),
.B(n_225),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_542),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_536),
.B(n_453),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_543),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_537),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_537),
.Y(n_628)
);

INVx1_ASAP7_75t_SL g629 ( 
.A(n_557),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_609),
.B(n_454),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_537),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_543),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_538),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_556),
.B(n_460),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_538),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_567),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_556),
.B(n_469),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_546),
.Y(n_638)
);

AND3x2_ASAP7_75t_L g639 ( 
.A(n_584),
.B(n_589),
.C(n_557),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_341),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_546),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_552),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_536),
.B(n_478),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_619),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_571),
.B(n_481),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_538),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_544),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_539),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_571),
.B(n_484),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_613),
.B(n_435),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_544),
.Y(n_652)
);

INVxp33_ASAP7_75t_L g653 ( 
.A(n_587),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_544),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_541),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_539),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_553),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_557),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_550),
.B(n_451),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_540),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_598),
.B(n_494),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_542),
.Y(n_662)
);

OAI21xp33_ASAP7_75t_SL g663 ( 
.A1(n_577),
.A2(n_519),
.B(n_512),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_594),
.B(n_489),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_609),
.B(n_497),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_577),
.B(n_499),
.Y(n_666)
);

BUFx3_ASAP7_75t_L g667 ( 
.A(n_606),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_550),
.B(n_458),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_540),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_542),
.B(n_500),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_594),
.B(n_592),
.Y(n_671)
);

AOI22xp33_ASAP7_75t_L g672 ( 
.A1(n_612),
.A2(n_429),
.B1(n_369),
.B2(n_398),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_547),
.B(n_341),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_593),
.Y(n_674)
);

INVxp33_ASAP7_75t_L g675 ( 
.A(n_587),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_560),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_553),
.Y(n_677)
);

BUFx4f_ASAP7_75t_L g678 ( 
.A(n_576),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_606),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_609),
.B(n_504),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_594),
.B(n_505),
.Y(n_681)
);

BUFx2_ASAP7_75t_L g682 ( 
.A(n_593),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_542),
.B(n_511),
.Y(n_683)
);

BUFx6f_ASAP7_75t_L g684 ( 
.A(n_542),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_598),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_553),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_598),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_554),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_554),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_554),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_541),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_541),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_564),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_612),
.A2(n_375),
.B1(n_398),
.B2(n_369),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_602),
.A2(n_498),
.B1(n_503),
.B2(n_495),
.Y(n_695)
);

INVx5_ASAP7_75t_L g696 ( 
.A(n_542),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_560),
.Y(n_697)
);

AND2x2_ASAP7_75t_SL g698 ( 
.A(n_623),
.B(n_225),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_564),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_550),
.B(n_465),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_564),
.Y(n_701)
);

INVx5_ASAP7_75t_L g702 ( 
.A(n_542),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_562),
.Y(n_703)
);

NAND3xp33_ASAP7_75t_L g704 ( 
.A(n_576),
.B(n_459),
.C(n_457),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_562),
.Y(n_705)
);

INVx1_ASAP7_75t_SL g706 ( 
.A(n_559),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_594),
.B(n_527),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_545),
.Y(n_708)
);

NOR3xp33_ASAP7_75t_L g709 ( 
.A(n_575),
.B(n_360),
.C(n_463),
.Y(n_709)
);

AND2x6_ASAP7_75t_L g710 ( 
.A(n_545),
.B(n_225),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_568),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_563),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_584),
.B(n_535),
.Y(n_713)
);

INVxp67_ASAP7_75t_SL g714 ( 
.A(n_545),
.Y(n_714)
);

BUFx3_ASAP7_75t_L g715 ( 
.A(n_606),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_611),
.B(n_559),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_563),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_589),
.B(n_507),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_606),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_555),
.B(n_467),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_594),
.B(n_222),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_602),
.A2(n_515),
.B1(n_518),
.B2(n_514),
.Y(n_722)
);

NOR2x1p5_ASAP7_75t_L g723 ( 
.A(n_613),
.B(n_375),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_555),
.B(n_468),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_568),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_611),
.B(n_493),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_622),
.B(n_520),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_569),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_548),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_613),
.B(n_526),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_569),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_578),
.Y(n_732)
);

INVx4_ASAP7_75t_L g733 ( 
.A(n_545),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_592),
.B(n_343),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_592),
.B(n_377),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_568),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_579),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_547),
.B(n_613),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_555),
.B(n_468),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_613),
.B(n_532),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_578),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_588),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_592),
.B(n_314),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_592),
.B(n_316),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_548),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_575),
.B(n_534),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_588),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_579),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_L g750 ( 
.A(n_545),
.B(n_225),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_548),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_579),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_579),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_579),
.Y(n_754)
);

BUFx10_ASAP7_75t_L g755 ( 
.A(n_561),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_604),
.B(n_506),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_606),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_599),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_559),
.B(n_521),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_622),
.B(n_229),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_582),
.B(n_471),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_549),
.A2(n_547),
.B1(n_545),
.B2(n_576),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_604),
.B(n_264),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_599),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_548),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_579),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_582),
.B(n_466),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_600),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_600),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_601),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_601),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_604),
.B(n_510),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_579),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_572),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_582),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_549),
.A2(n_408),
.B1(n_414),
.B2(n_417),
.Y(n_776)
);

CKINVDCx11_ASAP7_75t_R g777 ( 
.A(n_581),
.Y(n_777)
);

AND2x6_ASAP7_75t_L g778 ( 
.A(n_548),
.B(n_225),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_662),
.B(n_549),
.Y(n_779)
);

NOR2xp33_ASAP7_75t_L g780 ( 
.A(n_685),
.B(n_549),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_676),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_759),
.B(n_470),
.Y(n_782)
);

BUFx6f_ASAP7_75t_SL g783 ( 
.A(n_636),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_624),
.B(n_549),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_726),
.Y(n_785)
);

AOI22x1_ASAP7_75t_L g786 ( 
.A1(n_640),
.A2(n_278),
.B1(n_294),
.B2(n_265),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_714),
.B(n_622),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_666),
.A2(n_547),
.B1(n_485),
.B2(n_482),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_655),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_L g790 ( 
.A(n_624),
.B(n_319),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_634),
.A2(n_547),
.B1(n_623),
.B2(n_622),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_637),
.B(n_622),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_624),
.B(n_592),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_655),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_726),
.B(n_587),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_SL g796 ( 
.A(n_723),
.B(n_249),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_697),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_655),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_777),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_663),
.A2(n_547),
.B1(n_216),
.B2(n_326),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_685),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_624),
.B(n_592),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_R g803 ( 
.A(n_645),
.B(n_581),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_687),
.B(n_561),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_625),
.B(n_547),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_697),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_624),
.B(n_592),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_703),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_644),
.B(n_646),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_687),
.B(n_226),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_703),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_650),
.B(n_558),
.Y(n_812)
);

BUFx6f_ASAP7_75t_SL g813 ( 
.A(n_636),
.Y(n_813)
);

OR2x6_ASAP7_75t_L g814 ( 
.A(n_682),
.B(n_727),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_705),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_700),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_705),
.Y(n_817)
);

INVxp67_ASAP7_75t_L g818 ( 
.A(n_716),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_712),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_712),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_717),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_691),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_717),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_663),
.B(n_231),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_664),
.B(n_232),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_698),
.B(n_558),
.Y(n_826)
);

AND2x6_ASAP7_75t_SL g827 ( 
.A(n_747),
.B(n_408),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_691),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_716),
.B(n_516),
.Y(n_829)
);

OAI22xp33_ASAP7_75t_L g830 ( 
.A1(n_704),
.A2(n_417),
.B1(n_419),
.B2(n_414),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_698),
.B(n_728),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_684),
.B(n_708),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_698),
.B(n_558),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_761),
.B(n_608),
.Y(n_834)
);

BUFx6f_ASAP7_75t_SL g835 ( 
.A(n_636),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_728),
.B(n_573),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_684),
.B(n_225),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_645),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_684),
.B(n_361),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_750),
.A2(n_566),
.B(n_565),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_681),
.B(n_233),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_691),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_684),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_684),
.B(n_322),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_692),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_731),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_731),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_732),
.B(n_573),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_674),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_SL g850 ( 
.A1(n_653),
.A2(n_591),
.B1(n_290),
.B2(n_387),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_692),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_627),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_667),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_708),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_713),
.B(n_294),
.C(n_278),
.Y(n_855)
);

NOR3xp33_ASAP7_75t_L g856 ( 
.A(n_709),
.B(n_313),
.C(n_305),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_708),
.B(n_361),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_732),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_741),
.B(n_573),
.Y(n_859)
);

BUFx5_ASAP7_75t_L g860 ( 
.A(n_710),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_670),
.A2(n_608),
.B(n_614),
.C(n_610),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_678),
.A2(n_590),
.B(n_572),
.C(n_313),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_741),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_742),
.B(n_573),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_707),
.B(n_244),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_628),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_628),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_708),
.B(n_361),
.Y(n_868)
);

NAND2xp33_ASAP7_75t_L g869 ( 
.A(n_708),
.B(n_746),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_761),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_746),
.Y(n_871)
);

INVx2_ASAP7_75t_SL g872 ( 
.A(n_682),
.Y(n_872)
);

INVxp33_ASAP7_75t_L g873 ( 
.A(n_767),
.Y(n_873)
);

INVx3_ASAP7_75t_L g874 ( 
.A(n_667),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_742),
.B(n_573),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_659),
.B(n_621),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_631),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_661),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_668),
.B(n_250),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_668),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_706),
.B(n_621),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_631),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_746),
.B(n_361),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_748),
.B(n_586),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_700),
.B(n_621),
.Y(n_885)
);

A2O1A1Ixp33_ASAP7_75t_L g886 ( 
.A1(n_678),
.A2(n_572),
.B(n_590),
.C(n_383),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_748),
.B(n_586),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_704),
.B(n_267),
.C(n_258),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_630),
.B(n_271),
.Y(n_889)
);

BUFx5_ASAP7_75t_L g890 ( 
.A(n_710),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_758),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_758),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_706),
.B(n_610),
.Y(n_893)
);

INVx5_ASAP7_75t_L g894 ( 
.A(n_710),
.Y(n_894)
);

OR2x2_ASAP7_75t_L g895 ( 
.A(n_775),
.B(n_661),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_764),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_633),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_764),
.B(n_586),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_768),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_768),
.B(n_586),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_769),
.B(n_586),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_633),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_775),
.B(n_614),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_746),
.B(n_361),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_769),
.B(n_597),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_635),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_720),
.Y(n_907)
);

NOR2xp67_ASAP7_75t_L g908 ( 
.A(n_730),
.B(n_740),
.Y(n_908)
);

NAND3xp33_ASAP7_75t_L g909 ( 
.A(n_694),
.B(n_274),
.C(n_273),
.Y(n_909)
);

AO22x2_ASAP7_75t_L g910 ( 
.A1(n_760),
.A2(n_371),
.B1(n_388),
.B2(n_383),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_L g911 ( 
.A(n_718),
.B(n_317),
.C(n_305),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_665),
.B(n_275),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_746),
.B(n_361),
.Y(n_913)
);

OR2x6_ASAP7_75t_L g914 ( 
.A(n_695),
.B(n_419),
.Y(n_914)
);

AND2x2_ASAP7_75t_SL g915 ( 
.A(n_762),
.B(n_776),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_770),
.B(n_597),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_635),
.Y(n_917)
);

NOR3xp33_ASAP7_75t_L g918 ( 
.A(n_680),
.B(n_320),
.C(n_317),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_770),
.B(n_597),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_771),
.B(n_597),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_771),
.B(n_719),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_678),
.A2(n_576),
.B1(n_590),
.B2(n_363),
.Y(n_922)
);

NAND2x1_ASAP7_75t_L g923 ( 
.A(n_733),
.B(n_551),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_647),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_719),
.B(n_597),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_756),
.B(n_551),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_636),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_733),
.B(n_333),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_756),
.B(n_335),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_733),
.B(n_340),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_679),
.Y(n_931)
);

NAND3x1_ASAP7_75t_L g932 ( 
.A(n_721),
.B(n_321),
.C(n_320),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_715),
.B(n_276),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_772),
.B(n_551),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_715),
.B(n_281),
.Y(n_935)
);

NOR3xp33_ASAP7_75t_L g936 ( 
.A(n_722),
.B(n_331),
.C(n_321),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_679),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_772),
.B(n_615),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_SL g939 ( 
.A(n_733),
.B(n_344),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_757),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_626),
.B(n_551),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_757),
.B(n_286),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_647),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_629),
.B(n_615),
.Y(n_944)
);

OR2x2_ASAP7_75t_L g945 ( 
.A(n_629),
.B(n_618),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_843),
.B(n_809),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_873),
.B(n_658),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_843),
.A2(n_702),
.B(n_696),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_862),
.A2(n_640),
.B(n_710),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_854),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_872),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_869),
.A2(n_702),
.B(n_696),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_880),
.A2(n_683),
.B(n_632),
.C(n_638),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_880),
.B(n_658),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_885),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_908),
.B(n_696),
.Y(n_956)
);

NOR2xp67_ASAP7_75t_L g957 ( 
.A(n_927),
.B(n_720),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_885),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_781),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_876),
.B(n_696),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_812),
.A2(n_702),
.B(n_774),
.Y(n_961)
);

NOR2xp67_ASAP7_75t_L g962 ( 
.A(n_838),
.B(n_724),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_915),
.A2(n_723),
.B1(n_763),
.B2(n_738),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_852),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_854),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_797),
.Y(n_966)
);

CKINVDCx10_ASAP7_75t_R g967 ( 
.A(n_783),
.Y(n_967)
);

O2A1O1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_830),
.A2(n_632),
.B(n_638),
.C(n_626),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_832),
.A2(n_702),
.B(n_774),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_806),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_870),
.B(n_639),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_854),
.Y(n_972)
);

AOI21xp33_ASAP7_75t_L g973 ( 
.A1(n_824),
.A2(n_763),
.B(n_738),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_915),
.A2(n_763),
.B1(n_738),
.B2(n_739),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_938),
.B(n_763),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_808),
.B(n_724),
.Y(n_976)
);

AO21x1_ASAP7_75t_L g977 ( 
.A1(n_824),
.A2(n_792),
.B(n_830),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_922),
.A2(n_640),
.B1(n_672),
.B2(n_673),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_811),
.B(n_739),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_816),
.B(n_651),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_881),
.Y(n_981)
);

INVx11_ASAP7_75t_L g982 ( 
.A(n_803),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_815),
.B(n_641),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_817),
.B(n_641),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_799),
.Y(n_985)
);

OR2x6_ASAP7_75t_L g986 ( 
.A(n_849),
.B(n_673),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_819),
.B(n_642),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_832),
.A2(n_774),
.B(n_671),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_785),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_886),
.A2(n_710),
.B(n_643),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_805),
.A2(n_774),
.B(n_744),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_888),
.B(n_649),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_894),
.A2(n_774),
.B(n_743),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_894),
.A2(n_735),
.B(n_734),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_866),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_831),
.A2(n_643),
.B(n_642),
.C(n_649),
.Y(n_996)
);

INVx6_ASAP7_75t_L g997 ( 
.A(n_945),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_867),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_854),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_820),
.B(n_656),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_853),
.Y(n_1001)
);

OAI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_800),
.A2(n_895),
.B1(n_907),
.B2(n_870),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_894),
.A2(n_738),
.B(n_673),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_821),
.B(n_656),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_922),
.A2(n_673),
.B1(n_738),
.B2(n_403),
.Y(n_1005)
);

AND2x6_ASAP7_75t_L g1006 ( 
.A(n_791),
.B(n_729),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_879),
.A2(n_669),
.B(n_660),
.C(n_729),
.Y(n_1007)
);

OAI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_826),
.A2(n_710),
.B(n_729),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_894),
.A2(n_673),
.B(n_737),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_823),
.B(n_846),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_871),
.A2(n_749),
.B(n_737),
.Y(n_1011)
);

CKINVDCx6p67_ASAP7_75t_R g1012 ( 
.A(n_783),
.Y(n_1012)
);

O2A1O1Ixp5_ASAP7_75t_L g1013 ( 
.A1(n_928),
.A2(n_669),
.B(n_660),
.C(n_745),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_847),
.B(n_745),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_871),
.A2(n_752),
.B(n_749),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_877),
.Y(n_1016)
);

BUFx3_ASAP7_75t_L g1017 ( 
.A(n_801),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_871),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_858),
.B(n_863),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_891),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_871),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_882),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_921),
.A2(n_753),
.B(n_752),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_944),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_893),
.B(n_755),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_833),
.A2(n_844),
.B(n_790),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_SL g1027 ( 
.A(n_813),
.B(n_591),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_925),
.A2(n_754),
.B(n_753),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_829),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_926),
.A2(n_766),
.B(n_754),
.Y(n_1030)
);

AOI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_825),
.A2(n_651),
.B1(n_755),
.B2(n_765),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_903),
.B(n_675),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_892),
.B(n_745),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_896),
.B(n_751),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_899),
.B(n_751),
.Y(n_1035)
);

BUFx12f_ASAP7_75t_L g1036 ( 
.A(n_878),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_853),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_879),
.B(n_755),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_818),
.B(n_755),
.Y(n_1039)
);

OAI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_934),
.A2(n_765),
.B(n_751),
.Y(n_1040)
);

OAI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_836),
.A2(n_765),
.B(n_699),
.Y(n_1041)
);

A2O1A1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_825),
.A2(n_331),
.B(n_371),
.C(n_388),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_848),
.A2(n_699),
.B(n_693),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_841),
.B(n_693),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_841),
.B(n_701),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_923),
.A2(n_773),
.B(n_766),
.Y(n_1046)
);

BUFx2_ASAP7_75t_SL g1047 ( 
.A(n_813),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_928),
.A2(n_773),
.B(n_711),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_897),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_874),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_930),
.A2(n_711),
.B(n_701),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_780),
.B(n_348),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_930),
.A2(n_736),
.B(n_725),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_939),
.A2(n_802),
.B(n_793),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_818),
.A2(n_256),
.B1(n_337),
.B2(n_345),
.Y(n_1055)
);

AOI22xp5_ASAP7_75t_L g1056 ( 
.A1(n_865),
.A2(n_407),
.B1(n_349),
.B2(n_353),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_939),
.A2(n_736),
.B(n_725),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_859),
.A2(n_652),
.B(n_648),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_793),
.A2(n_652),
.B(n_648),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_874),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_802),
.A2(n_657),
.B(n_654),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_810),
.B(n_618),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_865),
.B(n_654),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_807),
.A2(n_677),
.B(n_657),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_889),
.A2(n_363),
.B(n_352),
.C(n_345),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_864),
.A2(n_884),
.B(n_875),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_807),
.A2(n_686),
.B(n_677),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_810),
.B(n_686),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_933),
.B(n_688),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_933),
.B(n_688),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_902),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_779),
.A2(n_690),
.B(n_689),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_935),
.B(n_689),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_787),
.A2(n_690),
.B(n_566),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_834),
.B(n_251),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_837),
.A2(n_566),
.B(n_565),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_837),
.A2(n_566),
.B(n_565),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_780),
.B(n_354),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_SL g1079 ( 
.A(n_835),
.B(n_238),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_839),
.A2(n_566),
.B(n_565),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_935),
.B(n_337),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_839),
.A2(n_565),
.B(n_551),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_795),
.B(n_289),
.Y(n_1083)
);

OAI21xp33_ASAP7_75t_L g1084 ( 
.A1(n_889),
.A2(n_912),
.B(n_936),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_857),
.A2(n_358),
.B(n_352),
.Y(n_1085)
);

NOR3xp33_ASAP7_75t_L g1086 ( 
.A(n_788),
.B(n_372),
.C(n_358),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_942),
.B(n_372),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_857),
.A2(n_883),
.B(n_868),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_929),
.A2(n_533),
.B(n_513),
.C(n_522),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_868),
.A2(n_580),
.B(n_574),
.Y(n_1090)
);

OAI21xp33_ASAP7_75t_L g1091 ( 
.A1(n_912),
.A2(n_298),
.B(n_291),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_782),
.B(n_255),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_883),
.A2(n_580),
.B(n_574),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_904),
.A2(n_580),
.B(n_574),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_904),
.A2(n_595),
.B(n_583),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_940),
.B(n_510),
.Y(n_1096)
);

INVx2_ASAP7_75t_SL g1097 ( 
.A(n_803),
.Y(n_1097)
);

BUFx4f_ASAP7_75t_L g1098 ( 
.A(n_814),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_L g1099 ( 
.A(n_850),
.B(n_303),
.C(n_302),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_906),
.Y(n_1100)
);

OAI21xp33_ASAP7_75t_L g1101 ( 
.A1(n_936),
.A2(n_318),
.B(n_308),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_804),
.B(n_323),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_R g1103 ( 
.A(n_796),
.B(n_355),
.Y(n_1103)
);

OAI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_887),
.A2(n_778),
.B(n_620),
.Y(n_1104)
);

INVx4_ASAP7_75t_L g1105 ( 
.A(n_835),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_911),
.B(n_356),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_913),
.A2(n_583),
.B(n_620),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_942),
.B(n_931),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_937),
.B(n_804),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_917),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_898),
.B(n_583),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_913),
.A2(n_595),
.B(n_620),
.Y(n_1112)
);

OAI321xp33_ASAP7_75t_L g1113 ( 
.A1(n_914),
.A2(n_522),
.A3(n_529),
.B1(n_533),
.B2(n_513),
.C(n_523),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_914),
.B(n_327),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_914),
.B(n_330),
.Y(n_1115)
);

HB1xp67_ASAP7_75t_L g1116 ( 
.A(n_814),
.Y(n_1116)
);

AOI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_911),
.A2(n_368),
.B1(n_412),
.B2(n_410),
.Y(n_1117)
);

INVx1_ASAP7_75t_SL g1118 ( 
.A(n_827),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_814),
.B(n_338),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_900),
.B(n_595),
.Y(n_1120)
);

NAND2x1p5_ASAP7_75t_L g1121 ( 
.A(n_784),
.B(n_570),
.Y(n_1121)
);

AOI21xp33_ASAP7_75t_L g1122 ( 
.A1(n_910),
.A2(n_399),
.B(n_384),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_856),
.B(n_255),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_901),
.A2(n_596),
.B(n_617),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_SL g1125 ( 
.A(n_909),
.B(n_238),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_905),
.B(n_596),
.Y(n_1126)
);

INVxp67_ASAP7_75t_L g1127 ( 
.A(n_918),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_910),
.A2(n_397),
.B1(n_390),
.B2(n_389),
.Y(n_1128)
);

AND2x2_ASAP7_75t_SL g1129 ( 
.A(n_856),
.B(n_523),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_784),
.B(n_342),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_916),
.B(n_570),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_919),
.A2(n_596),
.B(n_617),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_910),
.A2(n_402),
.B1(n_374),
.B2(n_418),
.Y(n_1133)
);

NAND3xp33_ASAP7_75t_SL g1134 ( 
.A(n_1084),
.B(n_918),
.C(n_855),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_959),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_966),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1038),
.B(n_962),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1130),
.A2(n_946),
.B(n_1102),
.C(n_973),
.Y(n_1138)
);

NAND2x1p5_ASAP7_75t_L g1139 ( 
.A(n_1018),
.B(n_789),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_970),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_SL g1141 ( 
.A(n_1005),
.B(n_860),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_1024),
.B(n_855),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_946),
.A2(n_961),
.B(n_1026),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_950),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1020),
.Y(n_1145)
);

CKINVDCx14_ASAP7_75t_R g1146 ( 
.A(n_1012),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_964),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_975),
.B(n_1044),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_947),
.B(n_920),
.Y(n_1149)
);

NOR2xp33_ASAP7_75t_L g1150 ( 
.A(n_997),
.B(n_941),
.Y(n_1150)
);

NOR2xp33_ASAP7_75t_L g1151 ( 
.A(n_997),
.B(n_794),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_991),
.A2(n_828),
.B(n_798),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1032),
.B(n_255),
.Y(n_1153)
);

NAND2x2_ASAP7_75t_L g1154 ( 
.A(n_985),
.B(n_255),
.Y(n_1154)
);

INVx5_ASAP7_75t_L g1155 ( 
.A(n_950),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1122),
.A2(n_861),
.B(n_924),
.C(n_943),
.Y(n_1156)
);

OR2x6_ASAP7_75t_L g1157 ( 
.A(n_1047),
.B(n_932),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_1062),
.B(n_860),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1096),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_952),
.A2(n_960),
.B(n_948),
.Y(n_1160)
);

OR2x6_ASAP7_75t_L g1161 ( 
.A(n_1036),
.B(n_997),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1002),
.B(n_362),
.C(n_425),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_982),
.Y(n_1163)
);

CKINVDCx14_ASAP7_75t_R g1164 ( 
.A(n_1105),
.Y(n_1164)
);

A2O1A1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_973),
.A2(n_851),
.B(n_845),
.C(n_822),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_981),
.B(n_1109),
.Y(n_1166)
);

HB1xp67_ASAP7_75t_L g1167 ( 
.A(n_951),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1086),
.B(n_786),
.C(n_840),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_995),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_998),
.Y(n_1170)
);

NAND2x1p5_ASAP7_75t_L g1171 ( 
.A(n_1018),
.B(n_842),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1029),
.B(n_351),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_976),
.B(n_860),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_978),
.A2(n_416),
.B1(n_364),
.B2(n_401),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1096),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_R g1176 ( 
.A(n_1027),
.B(n_860),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_R g1177 ( 
.A(n_1097),
.B(n_860),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_979),
.B(n_890),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1016),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1108),
.B(n_1010),
.Y(n_1180)
);

NOR2xp33_ASAP7_75t_R g1181 ( 
.A(n_967),
.B(n_890),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_978),
.A2(n_1005),
.B1(n_974),
.B2(n_963),
.Y(n_1182)
);

O2A1O1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1122),
.A2(n_529),
.B(n_528),
.C(n_525),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_950),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1081),
.A2(n_404),
.B(n_373),
.C(n_381),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_1019),
.B(n_890),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1087),
.B(n_890),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1022),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_983),
.B(n_890),
.Y(n_1189)
);

OR2x6_ASAP7_75t_SL g1190 ( 
.A(n_1055),
.B(n_1128),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1049),
.Y(n_1191)
);

INVx2_ASAP7_75t_SL g1192 ( 
.A(n_989),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1017),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_L g1194 ( 
.A(n_1105),
.B(n_357),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_965),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_984),
.B(n_987),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1000),
.B(n_1004),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1044),
.B(n_607),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_960),
.A2(n_391),
.B(n_385),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1083),
.B(n_365),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_949),
.A2(n_421),
.B(n_422),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1071),
.Y(n_1202)
);

NAND3xp33_ASAP7_75t_SL g1203 ( 
.A(n_1114),
.B(n_409),
.C(n_420),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1100),
.Y(n_1204)
);

NAND2x1p5_ASAP7_75t_L g1205 ( 
.A(n_965),
.B(n_607),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1045),
.B(n_607),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1110),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1127),
.A2(n_411),
.B(n_424),
.C(n_367),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_R g1209 ( 
.A(n_971),
.B(n_239),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_955),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1045),
.B(n_616),
.Y(n_1211)
);

NOR2xp67_ASAP7_75t_SL g1212 ( 
.A(n_1113),
.B(n_525),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_954),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_958),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1014),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1068),
.B(n_616),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1033),
.Y(n_1217)
);

O2A1O1Ixp33_ASAP7_75t_L g1218 ( 
.A1(n_1065),
.A2(n_528),
.B(n_616),
.C(n_617),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_1092),
.Y(n_1219)
);

BUFx2_ASAP7_75t_L g1220 ( 
.A(n_1116),
.Y(n_1220)
);

INVxp67_ASAP7_75t_SL g1221 ( 
.A(n_965),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_953),
.A2(n_393),
.B(n_423),
.C(n_396),
.Y(n_1222)
);

BUFx4f_ASAP7_75t_L g1223 ( 
.A(n_980),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_980),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1034),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1001),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1039),
.B(n_366),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_949),
.A2(n_605),
.B(n_603),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_993),
.A2(n_605),
.B(n_603),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1001),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1075),
.B(n_370),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1063),
.B(n_570),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1035),
.Y(n_1233)
);

O2A1O1Ixp5_ASAP7_75t_L g1234 ( 
.A1(n_977),
.A2(n_239),
.B(n_325),
.C(n_243),
.Y(n_1234)
);

NOR3xp33_ASAP7_75t_SL g1235 ( 
.A(n_1055),
.B(n_386),
.C(n_243),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1025),
.A2(n_238),
.B1(n_243),
.B2(n_325),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1069),
.B(n_570),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1129),
.B(n_238),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1070),
.B(n_570),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1073),
.B(n_570),
.Y(n_1240)
);

INVx4_ASAP7_75t_SL g1241 ( 
.A(n_972),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1123),
.B(n_243),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_968),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_957),
.B(n_75),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1098),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_996),
.Y(n_1246)
);

BUFx8_ASAP7_75t_L g1247 ( 
.A(n_972),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1037),
.B(n_570),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_986),
.A2(n_1098),
.B1(n_1031),
.B2(n_990),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_1119),
.B(n_570),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1037),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_972),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1050),
.Y(n_1253)
);

INVx3_ASAP7_75t_SL g1254 ( 
.A(n_1118),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_999),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1050),
.B(n_585),
.Y(n_1256)
);

AOI21x1_ASAP7_75t_L g1257 ( 
.A1(n_956),
.A2(n_778),
.B(n_605),
.Y(n_1257)
);

OAI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1091),
.A2(n_585),
.B(n_603),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_R g1259 ( 
.A(n_1079),
.B(n_80),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_SL g1260 ( 
.A(n_1060),
.B(n_325),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1060),
.B(n_605),
.Y(n_1261)
);

INVx2_ASAP7_75t_SL g1262 ( 
.A(n_1103),
.Y(n_1262)
);

BUFx3_ASAP7_75t_L g1263 ( 
.A(n_986),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_999),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1003),
.A2(n_212),
.B(n_210),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1089),
.Y(n_1266)
);

BUFx8_ASAP7_75t_L g1267 ( 
.A(n_999),
.Y(n_1267)
);

OAI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_990),
.A2(n_778),
.B(n_325),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1115),
.B(n_14),
.Y(n_1269)
);

BUFx6f_ASAP7_75t_L g1270 ( 
.A(n_1021),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1021),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_969),
.A2(n_605),
.B(n_603),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_L g1273 ( 
.A(n_1101),
.B(n_17),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_1021),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1066),
.B(n_605),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1056),
.B(n_17),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1125),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_986),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_L g1279 ( 
.A1(n_1042),
.A2(n_18),
.B(n_23),
.C(n_27),
.Y(n_1279)
);

AOI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_992),
.A2(n_778),
.B1(n_605),
.B2(n_603),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1111),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1106),
.Y(n_1282)
);

OAI22xp5_ASAP7_75t_L g1283 ( 
.A1(n_1008),
.A2(n_585),
.B1(n_603),
.B2(n_605),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1120),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1126),
.Y(n_1285)
);

O2A1O1Ixp33_ASAP7_75t_SL g1286 ( 
.A1(n_1007),
.A2(n_778),
.B(n_209),
.C(n_202),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1008),
.A2(n_603),
.B1(n_585),
.B2(n_30),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1117),
.B(n_1052),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1009),
.A2(n_603),
.B(n_585),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1078),
.B(n_585),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1066),
.B(n_1040),
.Y(n_1291)
);

HB1xp67_ASAP7_75t_L g1292 ( 
.A(n_1128),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1124),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_994),
.A2(n_585),
.B(n_778),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1121),
.A2(n_585),
.B1(n_29),
.B2(n_31),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_988),
.A2(n_778),
.B(n_197),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1180),
.B(n_1133),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1161),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1135),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1152),
.A2(n_1048),
.B(n_1072),
.Y(n_1300)
);

AND3x4_ASAP7_75t_L g1301 ( 
.A(n_1235),
.B(n_1099),
.C(n_1133),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1138),
.A2(n_1054),
.B(n_1013),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1143),
.A2(n_1040),
.B(n_1041),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1148),
.A2(n_1030),
.B(n_1023),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1136),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1287),
.A2(n_1121),
.B(n_1041),
.Y(n_1306)
);

BUFx10_ASAP7_75t_L g1307 ( 
.A(n_1269),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1275),
.A2(n_1074),
.B(n_1057),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1182),
.A2(n_1053),
.A3(n_1051),
.B(n_1088),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1148),
.A2(n_1131),
.B(n_1058),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1182),
.A2(n_1028),
.A3(n_1131),
.B(n_1132),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1140),
.Y(n_1312)
);

INVx1_ASAP7_75t_SL g1313 ( 
.A(n_1167),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1228),
.A2(n_1160),
.B(n_1290),
.Y(n_1314)
);

NAND3xp33_ASAP7_75t_L g1315 ( 
.A(n_1200),
.B(n_1085),
.C(n_1112),
.Y(n_1315)
);

AOI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1239),
.A2(n_1011),
.B(n_1015),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1145),
.Y(n_1317)
);

OR2x6_ASAP7_75t_L g1318 ( 
.A(n_1161),
.B(n_1059),
.Y(n_1318)
);

INVxp67_ASAP7_75t_L g1319 ( 
.A(n_1220),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1254),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1196),
.A2(n_1058),
.B(n_1043),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1149),
.B(n_1006),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1197),
.A2(n_1104),
.B1(n_1043),
.B2(n_1046),
.Y(n_1323)
);

INVx4_ASAP7_75t_L g1324 ( 
.A(n_1155),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1276),
.A2(n_1006),
.B1(n_1104),
.B2(n_1061),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1153),
.B(n_1076),
.Y(n_1326)
);

NOR2xp67_ASAP7_75t_L g1327 ( 
.A(n_1262),
.B(n_1064),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1243),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1163),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1227),
.A2(n_1067),
.B(n_1077),
.C(n_1080),
.Y(n_1330)
);

OA21x2_ASAP7_75t_L g1331 ( 
.A1(n_1165),
.A2(n_1107),
.B(n_1095),
.Y(n_1331)
);

BUFx6f_ASAP7_75t_L g1332 ( 
.A(n_1144),
.Y(n_1332)
);

OAI22x1_ASAP7_75t_L g1333 ( 
.A1(n_1292),
.A2(n_1006),
.B1(n_29),
.B2(n_32),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1229),
.A2(n_1094),
.B(n_1093),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_1172),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1272),
.A2(n_1090),
.B(n_1082),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1215),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1187),
.A2(n_1006),
.B(n_189),
.Y(n_1338)
);

AOI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1239),
.A2(n_184),
.B(n_183),
.Y(n_1339)
);

NAND3xp33_ASAP7_75t_L g1340 ( 
.A(n_1162),
.B(n_18),
.C(n_34),
.Y(n_1340)
);

NAND3xp33_ASAP7_75t_L g1341 ( 
.A(n_1273),
.B(n_35),
.C(n_36),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1291),
.A2(n_181),
.B(n_177),
.Y(n_1342)
);

AOI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1240),
.A2(n_168),
.B(n_167),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_SL g1344 ( 
.A1(n_1287),
.A2(n_163),
.B(n_157),
.Y(n_1344)
);

BUFx10_ASAP7_75t_L g1345 ( 
.A(n_1161),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1141),
.A2(n_152),
.B(n_150),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1166),
.B(n_35),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1141),
.A2(n_145),
.B(n_139),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1249),
.A2(n_37),
.A3(n_40),
.B(n_41),
.Y(n_1349)
);

OR2x6_ASAP7_75t_L g1350 ( 
.A(n_1245),
.B(n_1192),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1281),
.B(n_37),
.Y(n_1351)
);

BUFx2_ASAP7_75t_SL g1352 ( 
.A(n_1193),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1268),
.A2(n_103),
.B(n_97),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1258),
.A2(n_95),
.B(n_92),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1231),
.B(n_43),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1219),
.B(n_46),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1247),
.Y(n_1357)
);

INVx3_ASAP7_75t_L g1358 ( 
.A(n_1144),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1240),
.A2(n_86),
.B(n_84),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_SL g1360 ( 
.A(n_1223),
.B(n_1277),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1268),
.A2(n_73),
.B(n_50),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_SL g1362 ( 
.A1(n_1282),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_1362)
);

AND2x4_ASAP7_75t_L g1363 ( 
.A(n_1263),
.B(n_54),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1224),
.B(n_54),
.Y(n_1364)
);

O2A1O1Ixp33_ASAP7_75t_SL g1365 ( 
.A1(n_1288),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_1365)
);

AO32x2_ASAP7_75t_L g1366 ( 
.A1(n_1249),
.A2(n_59),
.A3(n_61),
.B1(n_62),
.B2(n_66),
.Y(n_1366)
);

AOI31xp67_ASAP7_75t_L g1367 ( 
.A1(n_1232),
.A2(n_62),
.A3(n_66),
.B(n_67),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_1213),
.B(n_68),
.Y(n_1368)
);

NOR2xp67_ASAP7_75t_L g1369 ( 
.A(n_1203),
.B(n_1147),
.Y(n_1369)
);

AOI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1246),
.A2(n_70),
.B(n_73),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1150),
.A2(n_70),
.B1(n_1190),
.B2(n_1137),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1217),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1201),
.A2(n_1178),
.B(n_1173),
.Y(n_1373)
);

OAI22x1_ASAP7_75t_L g1374 ( 
.A1(n_1236),
.A2(n_1238),
.B1(n_1213),
.B2(n_1242),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1159),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1134),
.A2(n_1234),
.B(n_1222),
.C(n_1156),
.Y(n_1376)
);

AOI21xp33_ASAP7_75t_L g1377 ( 
.A1(n_1174),
.A2(n_1175),
.B(n_1250),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1284),
.B(n_1285),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1225),
.B(n_1233),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1151),
.B(n_1142),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1223),
.B(n_1210),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1198),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1247),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1214),
.B(n_1206),
.Y(n_1384)
);

OAI221xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1279),
.A2(n_1183),
.B1(n_1208),
.B2(n_1164),
.C(n_1157),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1267),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1174),
.A2(n_1209),
.B1(n_1278),
.B2(n_1260),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1237),
.A2(n_1211),
.B(n_1189),
.Y(n_1388)
);

NOR2xp67_ASAP7_75t_L g1389 ( 
.A(n_1169),
.B(n_1191),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1294),
.A2(n_1289),
.B(n_1257),
.Y(n_1390)
);

OAI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1186),
.A2(n_1168),
.B(n_1199),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1202),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1204),
.Y(n_1393)
);

AO32x2_ASAP7_75t_L g1394 ( 
.A1(n_1295),
.A2(n_1283),
.A3(n_1212),
.B1(n_1286),
.B2(n_1265),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1293),
.A2(n_1216),
.B(n_1168),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1267),
.Y(n_1396)
);

AND2x6_ASAP7_75t_L g1397 ( 
.A(n_1244),
.B(n_1195),
.Y(n_1397)
);

INVx6_ASAP7_75t_L g1398 ( 
.A(n_1278),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1207),
.B(n_1188),
.Y(n_1399)
);

AO31x2_ASAP7_75t_L g1400 ( 
.A1(n_1283),
.A2(n_1295),
.A3(n_1266),
.B(n_1296),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1158),
.A2(n_1261),
.B(n_1256),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1278),
.Y(n_1402)
);

O2A1O1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1185),
.A2(n_1157),
.B(n_1218),
.C(n_1170),
.Y(n_1403)
);

NAND2x1p5_ASAP7_75t_L g1404 ( 
.A(n_1155),
.B(n_1184),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1248),
.A2(n_1221),
.B(n_1139),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1146),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1139),
.A2(n_1171),
.B(n_1244),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_SL g1408 ( 
.A(n_1176),
.B(n_1259),
.Y(n_1408)
);

AOI21x1_ASAP7_75t_SL g1409 ( 
.A1(n_1157),
.A2(n_1154),
.B(n_1177),
.Y(n_1409)
);

AO31x2_ASAP7_75t_L g1410 ( 
.A1(n_1251),
.A2(n_1230),
.A3(n_1253),
.B(n_1226),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1179),
.B(n_1271),
.Y(n_1411)
);

AO21x1_ASAP7_75t_L g1412 ( 
.A1(n_1205),
.A2(n_1171),
.B(n_1280),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1264),
.B(n_1255),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1205),
.A2(n_1255),
.B(n_1252),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1252),
.A2(n_1194),
.B(n_1241),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1241),
.A2(n_1144),
.B(n_1184),
.Y(n_1416)
);

O2A1O1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1181),
.A2(n_1241),
.B(n_1195),
.C(n_1184),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1195),
.A2(n_1084),
.B1(n_1276),
.B2(n_1269),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1270),
.A2(n_1084),
.B(n_1269),
.C(n_1200),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1270),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1270),
.Y(n_1421)
);

AOI221x1_ASAP7_75t_L g1422 ( 
.A1(n_1274),
.A2(n_1084),
.B1(n_1086),
.B2(n_1138),
.C(n_1287),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1274),
.B(n_1180),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1274),
.B(n_1155),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1180),
.B(n_946),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1138),
.A2(n_1084),
.B(n_809),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1152),
.A2(n_1160),
.B(n_1143),
.Y(n_1427)
);

AOI211x1_ASAP7_75t_L g1428 ( 
.A1(n_1134),
.A2(n_1084),
.B(n_977),
.C(n_1122),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1167),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1269),
.A2(n_1084),
.B(n_1138),
.C(n_1200),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1143),
.A2(n_684),
.B(n_624),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1269),
.A2(n_1084),
.B(n_1200),
.C(n_556),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1143),
.A2(n_684),
.B(n_624),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1200),
.B(n_873),
.Y(n_1434)
);

AO31x2_ASAP7_75t_L g1435 ( 
.A1(n_1182),
.A2(n_977),
.A3(n_1138),
.B(n_1287),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1153),
.B(n_1032),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1144),
.Y(n_1437)
);

AO31x2_ASAP7_75t_L g1438 ( 
.A1(n_1182),
.A2(n_977),
.A3(n_1138),
.B(n_1287),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1135),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1152),
.A2(n_1160),
.B(n_1143),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_SL g1441 ( 
.A1(n_1138),
.A2(n_1288),
.B(n_1084),
.C(n_792),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1200),
.A2(n_1084),
.B1(n_747),
.B2(n_782),
.Y(n_1442)
);

INVx5_ASAP7_75t_L g1443 ( 
.A(n_1144),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1143),
.A2(n_684),
.B(n_624),
.Y(n_1444)
);

A2O1A1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1269),
.A2(n_1084),
.B(n_1138),
.C(n_1200),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1135),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1167),
.Y(n_1447)
);

NOR4xp25_ASAP7_75t_L g1448 ( 
.A(n_1269),
.B(n_1084),
.C(n_663),
.D(n_1134),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1152),
.A2(n_1160),
.B(n_1143),
.Y(n_1449)
);

AOI31xp67_ASAP7_75t_L g1450 ( 
.A1(n_1288),
.A2(n_792),
.A3(n_1290),
.B(n_1275),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1161),
.B(n_1047),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1200),
.B(n_873),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1152),
.A2(n_1160),
.B(n_1143),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1269),
.A2(n_1084),
.B(n_1200),
.C(n_556),
.Y(n_1454)
);

O2A1O1Ixp5_ASAP7_75t_L g1455 ( 
.A1(n_1200),
.A2(n_977),
.B(n_792),
.C(n_1234),
.Y(n_1455)
);

A2O1A1Ixp33_ASAP7_75t_L g1456 ( 
.A1(n_1269),
.A2(n_1084),
.B(n_1138),
.C(n_1200),
.Y(n_1456)
);

A2O1A1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1269),
.A2(n_1084),
.B(n_1138),
.C(n_1200),
.Y(n_1457)
);

AO31x2_ASAP7_75t_L g1458 ( 
.A1(n_1182),
.A2(n_977),
.A3(n_1138),
.B(n_1287),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1180),
.B(n_946),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1152),
.A2(n_1160),
.B(n_1143),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1143),
.A2(n_684),
.B(n_624),
.Y(n_1461)
);

BUFx3_ASAP7_75t_L g1462 ( 
.A(n_1161),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1180),
.B(n_946),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1180),
.A2(n_946),
.B1(n_1138),
.B2(n_1084),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1143),
.A2(n_684),
.B(n_624),
.Y(n_1465)
);

AOI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1143),
.A2(n_684),
.B(n_624),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_L g1467 ( 
.A1(n_1143),
.A2(n_684),
.B(n_624),
.Y(n_1467)
);

AOI221x1_ASAP7_75t_L g1468 ( 
.A1(n_1138),
.A2(n_1084),
.B1(n_1086),
.B2(n_1287),
.C(n_1269),
.Y(n_1468)
);

BUFx4f_ASAP7_75t_L g1469 ( 
.A(n_1329),
.Y(n_1469)
);

NAND2x1p5_ASAP7_75t_L g1470 ( 
.A(n_1324),
.B(n_1437),
.Y(n_1470)
);

OAI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1442),
.A2(n_1361),
.B1(n_1341),
.B2(n_1425),
.Y(n_1471)
);

BUFx12f_ASAP7_75t_L g1472 ( 
.A(n_1406),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1437),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1320),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1418),
.A2(n_1456),
.B1(n_1457),
.B2(n_1430),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1301),
.A2(n_1362),
.B1(n_1426),
.B2(n_1371),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1312),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1437),
.Y(n_1478)
);

BUFx4_ASAP7_75t_R g1479 ( 
.A(n_1357),
.Y(n_1479)
);

INVx8_ASAP7_75t_L g1480 ( 
.A(n_1443),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1340),
.A2(n_1297),
.B1(n_1353),
.B2(n_1333),
.Y(n_1481)
);

NAND2x1p5_ASAP7_75t_L g1482 ( 
.A(n_1443),
.B(n_1408),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1317),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1352),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1464),
.A2(n_1307),
.B1(n_1374),
.B2(n_1452),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1317),
.Y(n_1486)
);

BUFx8_ASAP7_75t_SL g1487 ( 
.A(n_1451),
.Y(n_1487)
);

INVx3_ASAP7_75t_L g1488 ( 
.A(n_1397),
.Y(n_1488)
);

OAI22x1_ASAP7_75t_L g1489 ( 
.A1(n_1328),
.A2(n_1434),
.B1(n_1337),
.B2(n_1372),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1445),
.A2(n_1463),
.B1(n_1459),
.B2(n_1454),
.Y(n_1490)
);

BUFx4_ASAP7_75t_SL g1491 ( 
.A(n_1451),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1436),
.B(n_1355),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1307),
.A2(n_1368),
.B1(n_1380),
.B2(n_1347),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1342),
.A2(n_1351),
.B1(n_1335),
.B2(n_1328),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1439),
.Y(n_1495)
);

BUFx12f_ASAP7_75t_L g1496 ( 
.A(n_1345),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1439),
.Y(n_1497)
);

INVx4_ASAP7_75t_L g1498 ( 
.A(n_1404),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1446),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1398),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_SL g1501 ( 
.A1(n_1364),
.A2(n_1335),
.B1(n_1356),
.B2(n_1366),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1337),
.A2(n_1372),
.B1(n_1378),
.B2(n_1364),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1350),
.Y(n_1503)
);

BUFx3_ASAP7_75t_L g1504 ( 
.A(n_1398),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1397),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1432),
.A2(n_1387),
.B1(n_1419),
.B2(n_1379),
.Y(n_1506)
);

BUFx3_ASAP7_75t_L g1507 ( 
.A(n_1298),
.Y(n_1507)
);

CKINVDCx11_ASAP7_75t_R g1508 ( 
.A(n_1345),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1397),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1322),
.A2(n_1325),
.B1(n_1348),
.B2(n_1346),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1305),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_L g1512 ( 
.A1(n_1377),
.A2(n_1382),
.B1(n_1369),
.B2(n_1326),
.Y(n_1512)
);

INVx6_ASAP7_75t_L g1513 ( 
.A(n_1350),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1428),
.A2(n_1385),
.B1(n_1319),
.B2(n_1423),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1462),
.Y(n_1515)
);

INVx4_ASAP7_75t_L g1516 ( 
.A(n_1424),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1447),
.Y(n_1517)
);

CKINVDCx11_ASAP7_75t_R g1518 ( 
.A(n_1313),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1448),
.A2(n_1383),
.B1(n_1386),
.B2(n_1396),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_SL g1520 ( 
.A1(n_1366),
.A2(n_1360),
.B1(n_1363),
.B2(n_1468),
.Y(n_1520)
);

CKINVDCx11_ASAP7_75t_R g1521 ( 
.A(n_1429),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1381),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1376),
.A2(n_1389),
.B1(n_1375),
.B2(n_1402),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1332),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1366),
.A2(n_1354),
.B1(n_1302),
.B2(n_1344),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1392),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1318),
.A2(n_1382),
.B1(n_1327),
.B2(n_1315),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1411),
.B(n_1393),
.Y(n_1528)
);

BUFx12f_ASAP7_75t_L g1529 ( 
.A(n_1332),
.Y(n_1529)
);

BUFx12f_ASAP7_75t_L g1530 ( 
.A(n_1332),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1399),
.Y(n_1531)
);

INVxp67_ASAP7_75t_SL g1532 ( 
.A(n_1395),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1397),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1358),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1420),
.Y(n_1535)
);

CKINVDCx11_ASAP7_75t_R g1536 ( 
.A(n_1318),
.Y(n_1536)
);

CKINVDCx11_ASAP7_75t_R g1537 ( 
.A(n_1409),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1410),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1391),
.A2(n_1384),
.B1(n_1338),
.B2(n_1373),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_SL g1540 ( 
.A1(n_1323),
.A2(n_1435),
.B1(n_1458),
.B2(n_1438),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1413),
.Y(n_1541)
);

BUFx10_ASAP7_75t_L g1542 ( 
.A(n_1417),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1321),
.A2(n_1395),
.B1(n_1303),
.B2(n_1310),
.Y(n_1543)
);

BUFx4f_ASAP7_75t_SL g1544 ( 
.A(n_1416),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1415),
.Y(n_1545)
);

CKINVDCx11_ASAP7_75t_R g1546 ( 
.A(n_1367),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1388),
.A2(n_1304),
.B1(n_1359),
.B2(n_1412),
.Y(n_1547)
);

INVx4_ASAP7_75t_L g1548 ( 
.A(n_1359),
.Y(n_1548)
);

INVx5_ASAP7_75t_L g1549 ( 
.A(n_1422),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1349),
.Y(n_1550)
);

OAI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1370),
.A2(n_1407),
.B1(n_1441),
.B2(n_1339),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1435),
.A2(n_1438),
.B1(n_1458),
.B2(n_1401),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1349),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1349),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1435),
.A2(n_1458),
.B1(n_1438),
.B2(n_1331),
.Y(n_1555)
);

BUFx4f_ASAP7_75t_SL g1556 ( 
.A(n_1365),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1394),
.Y(n_1557)
);

AOI22xp33_ASAP7_75t_L g1558 ( 
.A1(n_1331),
.A2(n_1405),
.B1(n_1414),
.B2(n_1455),
.Y(n_1558)
);

OAI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1306),
.A2(n_1461),
.B1(n_1431),
.B2(n_1466),
.Y(n_1559)
);

INVx11_ASAP7_75t_L g1560 ( 
.A(n_1403),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1343),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1309),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1309),
.Y(n_1563)
);

INVxp67_ASAP7_75t_SL g1564 ( 
.A(n_1433),
.Y(n_1564)
);

BUFx2_ASAP7_75t_SL g1565 ( 
.A(n_1444),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1465),
.A2(n_1467),
.B1(n_1330),
.B2(n_1314),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1394),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1309),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1394),
.A2(n_1400),
.B1(n_1450),
.B2(n_1460),
.Y(n_1569)
);

CKINVDCx11_ASAP7_75t_R g1570 ( 
.A(n_1400),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1400),
.Y(n_1571)
);

BUFx3_ASAP7_75t_L g1572 ( 
.A(n_1390),
.Y(n_1572)
);

INVx6_ASAP7_75t_L g1573 ( 
.A(n_1316),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1311),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_SL g1575 ( 
.A1(n_1427),
.A2(n_1453),
.B1(n_1449),
.B2(n_1440),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1308),
.A2(n_1311),
.B1(n_1300),
.B2(n_1336),
.Y(n_1576)
);

BUFx4f_ASAP7_75t_SL g1577 ( 
.A(n_1311),
.Y(n_1577)
);

INVx5_ASAP7_75t_L g1578 ( 
.A(n_1334),
.Y(n_1578)
);

BUFx2_ASAP7_75t_L g1579 ( 
.A(n_1421),
.Y(n_1579)
);

CKINVDCx5p33_ASAP7_75t_R g1580 ( 
.A(n_1329),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1299),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1299),
.Y(n_1582)
);

BUFx10_ASAP7_75t_L g1583 ( 
.A(n_1406),
.Y(n_1583)
);

OAI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1442),
.A2(n_1190),
.B1(n_1361),
.B2(n_1141),
.Y(n_1584)
);

BUFx10_ASAP7_75t_L g1585 ( 
.A(n_1406),
.Y(n_1585)
);

INVx2_ASAP7_75t_SL g1586 ( 
.A(n_1398),
.Y(n_1586)
);

OAI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1442),
.A2(n_1190),
.B1(n_1361),
.B2(n_1141),
.Y(n_1587)
);

OAI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1418),
.A2(n_1442),
.B1(n_1445),
.B2(n_1430),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1442),
.A2(n_1190),
.B1(n_1361),
.B2(n_1141),
.Y(n_1589)
);

BUFx3_ASAP7_75t_L g1590 ( 
.A(n_1421),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_1437),
.Y(n_1591)
);

BUFx12f_ASAP7_75t_L g1592 ( 
.A(n_1406),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1328),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1301),
.A2(n_1084),
.B1(n_1269),
.B2(n_1276),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1328),
.Y(n_1595)
);

CKINVDCx20_ASAP7_75t_R g1596 ( 
.A(n_1421),
.Y(n_1596)
);

CKINVDCx6p67_ASAP7_75t_R g1597 ( 
.A(n_1357),
.Y(n_1597)
);

BUFx8_ASAP7_75t_L g1598 ( 
.A(n_1329),
.Y(n_1598)
);

AOI22xp5_ASAP7_75t_SL g1599 ( 
.A1(n_1333),
.A2(n_1269),
.B1(n_1276),
.B2(n_747),
.Y(n_1599)
);

INVx6_ASAP7_75t_L g1600 ( 
.A(n_1437),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1442),
.A2(n_1200),
.B1(n_747),
.B2(n_1434),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1301),
.A2(n_1084),
.B1(n_1269),
.B2(n_1276),
.Y(n_1602)
);

CKINVDCx9p33_ASAP7_75t_R g1603 ( 
.A(n_1434),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1361),
.A2(n_1269),
.B1(n_1084),
.B2(n_1276),
.Y(n_1604)
);

CKINVDCx20_ASAP7_75t_R g1605 ( 
.A(n_1421),
.Y(n_1605)
);

CKINVDCx11_ASAP7_75t_R g1606 ( 
.A(n_1329),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1431),
.A2(n_946),
.B(n_1433),
.Y(n_1607)
);

INVx2_ASAP7_75t_SL g1608 ( 
.A(n_1398),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1442),
.A2(n_1200),
.B1(n_747),
.B2(n_1434),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1299),
.Y(n_1610)
);

OAI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1442),
.A2(n_1190),
.B1(n_1361),
.B2(n_1141),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1432),
.A2(n_1454),
.B(n_1445),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1299),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1421),
.Y(n_1614)
);

INVx6_ASAP7_75t_L g1615 ( 
.A(n_1437),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1398),
.Y(n_1616)
);

AOI21xp33_ASAP7_75t_L g1617 ( 
.A1(n_1432),
.A2(n_1454),
.B(n_1084),
.Y(n_1617)
);

AOI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1442),
.A2(n_1200),
.B1(n_747),
.B2(n_1434),
.Y(n_1618)
);

OAI21xp5_ASAP7_75t_SL g1619 ( 
.A1(n_1442),
.A2(n_747),
.B(n_639),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1299),
.Y(n_1620)
);

BUFx4f_ASAP7_75t_SL g1621 ( 
.A(n_1421),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1381),
.B(n_1298),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1361),
.A2(n_1269),
.B1(n_1084),
.B2(n_1276),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1538),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1572),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1593),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1536),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1553),
.B(n_1562),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1594),
.A2(n_1602),
.B1(n_1623),
.B2(n_1604),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1593),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1540),
.B(n_1557),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1545),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1595),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1604),
.A2(n_1623),
.B1(n_1601),
.B2(n_1618),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1477),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1483),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1528),
.Y(n_1637)
);

BUFx2_ASAP7_75t_L g1638 ( 
.A(n_1595),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1588),
.A2(n_1476),
.B1(n_1475),
.B2(n_1609),
.Y(n_1639)
);

INVxp33_ASAP7_75t_SL g1640 ( 
.A(n_1474),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1486),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1540),
.B(n_1612),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1497),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_R g1644 ( 
.A(n_1596),
.B(n_1605),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1499),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1581),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1563),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1574),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1532),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1582),
.Y(n_1650)
);

OAI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1607),
.A2(n_1576),
.B(n_1566),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1513),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1517),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1607),
.A2(n_1558),
.B(n_1547),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1532),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1550),
.Y(n_1656)
);

O2A1O1Ixp33_ASAP7_75t_SL g1657 ( 
.A1(n_1584),
.A2(n_1611),
.B(n_1587),
.C(n_1589),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1495),
.Y(n_1658)
);

OAI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1619),
.A2(n_1549),
.B1(n_1589),
.B2(n_1611),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1571),
.B(n_1555),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1544),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1513),
.Y(n_1662)
);

BUFx12f_ASAP7_75t_L g1663 ( 
.A(n_1606),
.Y(n_1663)
);

HB1xp67_ASAP7_75t_SL g1664 ( 
.A(n_1598),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1493),
.B(n_1531),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1567),
.Y(n_1666)
);

OAI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1558),
.A2(n_1547),
.B(n_1543),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1565),
.B(n_1554),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1567),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1490),
.A2(n_1617),
.B(n_1564),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1476),
.A2(n_1584),
.B1(n_1587),
.B2(n_1506),
.Y(n_1671)
);

AOI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1471),
.A2(n_1481),
.B1(n_1549),
.B2(n_1556),
.Y(n_1672)
);

BUFx2_ASAP7_75t_L g1673 ( 
.A(n_1489),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1555),
.B(n_1552),
.Y(n_1674)
);

HB1xp67_ASAP7_75t_L g1675 ( 
.A(n_1511),
.Y(n_1675)
);

BUFx3_ASAP7_75t_L g1676 ( 
.A(n_1544),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1610),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1613),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1620),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1526),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1573),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1493),
.B(n_1541),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1568),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1568),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1548),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1599),
.A2(n_1485),
.B1(n_1502),
.B2(n_1481),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1577),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1577),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1561),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1552),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1564),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1569),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1471),
.A2(n_1549),
.B1(n_1556),
.B2(n_1501),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1569),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1548),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1570),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1543),
.Y(n_1697)
);

BUFx2_ASAP7_75t_SL g1698 ( 
.A(n_1542),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1549),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1539),
.A2(n_1527),
.B(n_1510),
.Y(n_1700)
);

AND2x4_ASAP7_75t_L g1701 ( 
.A(n_1488),
.B(n_1505),
.Y(n_1701)
);

INVx6_ASAP7_75t_L g1702 ( 
.A(n_1533),
.Y(n_1702)
);

NAND2x1_ASAP7_75t_L g1703 ( 
.A(n_1510),
.B(n_1512),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1578),
.Y(n_1704)
);

CKINVDCx12_ASAP7_75t_R g1705 ( 
.A(n_1519),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1578),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1578),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1578),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1514),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_1488),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1512),
.A2(n_1494),
.B(n_1523),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1513),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1551),
.Y(n_1713)
);

AO31x2_ASAP7_75t_L g1714 ( 
.A1(n_1525),
.A2(n_1546),
.A3(n_1559),
.B(n_1575),
.Y(n_1714)
);

INVx3_ASAP7_75t_L g1715 ( 
.A(n_1560),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1575),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1559),
.Y(n_1717)
);

INVx3_ASAP7_75t_L g1718 ( 
.A(n_1505),
.Y(n_1718)
);

BUFx2_ASAP7_75t_L g1719 ( 
.A(n_1482),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1482),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1520),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1485),
.B(n_1502),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1520),
.B(n_1501),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1525),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1494),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1542),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1509),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1492),
.B(n_1622),
.Y(n_1728)
);

OAI21x1_ASAP7_75t_L g1729 ( 
.A1(n_1470),
.A2(n_1491),
.B(n_1537),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1470),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1491),
.Y(n_1731)
);

HB1xp67_ASAP7_75t_L g1732 ( 
.A(n_1534),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1473),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1473),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1507),
.B(n_1478),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1579),
.B(n_1590),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1600),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1518),
.A2(n_1521),
.B1(n_1496),
.B2(n_1508),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1600),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1500),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1524),
.B(n_1522),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1615),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1503),
.A2(n_1484),
.B1(n_1535),
.B2(n_1515),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1487),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1478),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1675),
.B(n_1608),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1680),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1638),
.B(n_1586),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1728),
.B(n_1616),
.Y(n_1749)
);

A2O1A1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1639),
.A2(n_1469),
.B(n_1603),
.C(n_1480),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1661),
.B(n_1676),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1638),
.B(n_1597),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1661),
.B(n_1676),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1670),
.B(n_1498),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1634),
.A2(n_1504),
.B1(n_1603),
.B2(n_1469),
.C(n_1614),
.Y(n_1755)
);

NOR2xp33_ASAP7_75t_L g1756 ( 
.A(n_1640),
.B(n_1621),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1741),
.B(n_1516),
.Y(n_1757)
);

AND2x4_ASAP7_75t_L g1758 ( 
.A(n_1676),
.B(n_1591),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1741),
.B(n_1529),
.Y(n_1759)
);

OAI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1629),
.A2(n_1580),
.B(n_1479),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1696),
.B(n_1530),
.Y(n_1761)
);

AOI221xp5_ASAP7_75t_L g1762 ( 
.A1(n_1657),
.A2(n_1480),
.B1(n_1591),
.B2(n_1621),
.C(n_1585),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1642),
.B(n_1583),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1686),
.A2(n_1472),
.B1(n_1592),
.B2(n_1598),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1687),
.B(n_1583),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1734),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1696),
.B(n_1585),
.Y(n_1767)
);

OR2x6_ASAP7_75t_L g1768 ( 
.A(n_1711),
.B(n_1668),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1642),
.B(n_1725),
.Y(n_1769)
);

OAI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1671),
.A2(n_1672),
.B(n_1693),
.C(n_1709),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1667),
.A2(n_1654),
.B(n_1711),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1637),
.B(n_1673),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1649),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1673),
.B(n_1626),
.Y(n_1774)
);

NOR2x1_ASAP7_75t_SL g1775 ( 
.A(n_1668),
.B(n_1698),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1721),
.A2(n_1659),
.B1(n_1722),
.B2(n_1723),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1626),
.B(n_1630),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1682),
.B(n_1665),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1703),
.A2(n_1725),
.B(n_1726),
.C(n_1722),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1687),
.B(n_1688),
.Y(n_1780)
);

NAND2x1_ASAP7_75t_L g1781 ( 
.A(n_1691),
.B(n_1689),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1736),
.B(n_1658),
.Y(n_1782)
);

NOR2x1_ASAP7_75t_SL g1783 ( 
.A(n_1668),
.B(n_1698),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1703),
.A2(n_1700),
.B(n_1724),
.C(n_1726),
.Y(n_1784)
);

OAI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1721),
.A2(n_1724),
.B1(n_1715),
.B2(n_1627),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1689),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1715),
.B(n_1740),
.Y(n_1787)
);

AOI221xp5_ASAP7_75t_L g1788 ( 
.A1(n_1717),
.A2(n_1690),
.B1(n_1697),
.B2(n_1713),
.C(n_1694),
.Y(n_1788)
);

INVx5_ASAP7_75t_L g1789 ( 
.A(n_1668),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1653),
.B(n_1712),
.Y(n_1790)
);

OR2x2_ASAP7_75t_SL g1791 ( 
.A(n_1702),
.B(n_1731),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_SL g1792 ( 
.A(n_1691),
.B(n_1699),
.Y(n_1792)
);

AO21x2_ASAP7_75t_L g1793 ( 
.A1(n_1651),
.A2(n_1713),
.B(n_1706),
.Y(n_1793)
);

BUFx5_ASAP7_75t_L g1794 ( 
.A(n_1706),
.Y(n_1794)
);

AO32x2_ASAP7_75t_L g1795 ( 
.A1(n_1652),
.A2(n_1662),
.A3(n_1631),
.B1(n_1692),
.B2(n_1694),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_L g1796 ( 
.A1(n_1717),
.A2(n_1715),
.B(n_1700),
.C(n_1697),
.Y(n_1796)
);

CKINVDCx5p33_ASAP7_75t_R g1797 ( 
.A(n_1644),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1633),
.B(n_1660),
.Y(n_1798)
);

BUFx8_ASAP7_75t_L g1799 ( 
.A(n_1663),
.Y(n_1799)
);

CKINVDCx6p67_ASAP7_75t_R g1800 ( 
.A(n_1663),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1628),
.Y(n_1801)
);

A2O1A1Ixp33_ASAP7_75t_L g1802 ( 
.A1(n_1715),
.A2(n_1729),
.B(n_1627),
.C(n_1652),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1649),
.Y(n_1803)
);

A2O1A1Ixp33_ASAP7_75t_L g1804 ( 
.A1(n_1729),
.A2(n_1627),
.B(n_1662),
.C(n_1699),
.Y(n_1804)
);

OA21x2_ASAP7_75t_L g1805 ( 
.A1(n_1716),
.A2(n_1695),
.B(n_1692),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1635),
.B(n_1636),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1635),
.B(n_1636),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1641),
.B(n_1643),
.Y(n_1808)
);

OA21x2_ASAP7_75t_L g1809 ( 
.A1(n_1716),
.A2(n_1695),
.B(n_1685),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_SL g1810 ( 
.A(n_1744),
.B(n_1702),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1643),
.B(n_1645),
.Y(n_1811)
);

OR2x6_ASAP7_75t_L g1812 ( 
.A(n_1656),
.B(n_1681),
.Y(n_1812)
);

NAND4xp25_ASAP7_75t_L g1813 ( 
.A(n_1738),
.B(n_1690),
.C(n_1744),
.D(n_1720),
.Y(n_1813)
);

O2A1O1Ixp33_ASAP7_75t_SL g1814 ( 
.A1(n_1743),
.A2(n_1727),
.B(n_1732),
.C(n_1705),
.Y(n_1814)
);

AO32x2_ASAP7_75t_L g1815 ( 
.A1(n_1631),
.A2(n_1714),
.A3(n_1669),
.B1(n_1666),
.B2(n_1628),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1645),
.B(n_1646),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1646),
.B(n_1650),
.Y(n_1817)
);

A2O1A1Ixp33_ASAP7_75t_L g1818 ( 
.A1(n_1719),
.A2(n_1720),
.B(n_1705),
.C(n_1674),
.Y(n_1818)
);

AO21x2_ASAP7_75t_L g1819 ( 
.A1(n_1707),
.A2(n_1708),
.B(n_1704),
.Y(n_1819)
);

AO21x2_ASAP7_75t_L g1820 ( 
.A1(n_1707),
.A2(n_1708),
.B(n_1704),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1674),
.A2(n_1744),
.B1(n_1656),
.B2(n_1702),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1702),
.A2(n_1735),
.B1(n_1701),
.B2(n_1730),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1655),
.Y(n_1823)
);

INVx3_ASAP7_75t_L g1824 ( 
.A(n_1819),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1815),
.B(n_1714),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1773),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1815),
.B(n_1714),
.Y(n_1827)
);

INVxp67_ASAP7_75t_SL g1828 ( 
.A(n_1781),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1815),
.B(n_1714),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1786),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1778),
.B(n_1679),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1778),
.B(n_1801),
.Y(n_1832)
);

AND2x4_ASAP7_75t_SL g1833 ( 
.A(n_1751),
.B(n_1753),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1791),
.Y(n_1834)
);

AND2x4_ASAP7_75t_L g1835 ( 
.A(n_1789),
.B(n_1625),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1773),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1803),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1801),
.B(n_1769),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1795),
.B(n_1669),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1769),
.B(n_1677),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1747),
.B(n_1823),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1795),
.B(n_1768),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1768),
.B(n_1683),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1768),
.B(n_1805),
.Y(n_1844)
);

AND2x4_ASAP7_75t_L g1845 ( 
.A(n_1819),
.B(n_1625),
.Y(n_1845)
);

AND2x2_ASAP7_75t_L g1846 ( 
.A(n_1805),
.B(n_1798),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1782),
.B(n_1774),
.Y(n_1847)
);

CKINVDCx16_ASAP7_75t_R g1848 ( 
.A(n_1810),
.Y(n_1848)
);

BUFx2_ASAP7_75t_L g1849 ( 
.A(n_1812),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1807),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1807),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1808),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1786),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_SL g1854 ( 
.A1(n_1770),
.A2(n_1710),
.B1(n_1701),
.B2(n_1718),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1806),
.B(n_1816),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1808),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1811),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1809),
.B(n_1817),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1809),
.B(n_1684),
.Y(n_1859)
);

INVxp67_ASAP7_75t_SL g1860 ( 
.A(n_1754),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1777),
.Y(n_1861)
);

NOR2x1_ASAP7_75t_L g1862 ( 
.A(n_1804),
.B(n_1632),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1788),
.B(n_1678),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1820),
.B(n_1647),
.Y(n_1864)
);

OAI222xp33_ASAP7_75t_L g1865 ( 
.A1(n_1776),
.A2(n_1730),
.B1(n_1664),
.B2(n_1742),
.C1(n_1739),
.C2(n_1733),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1820),
.B(n_1624),
.Y(n_1866)
);

NAND2xp33_ASAP7_75t_SL g1867 ( 
.A(n_1831),
.B(n_1797),
.Y(n_1867)
);

AOI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1863),
.A2(n_1776),
.B1(n_1779),
.B2(n_1755),
.C(n_1760),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1826),
.Y(n_1869)
);

BUFx2_ASAP7_75t_L g1870 ( 
.A(n_1834),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1860),
.B(n_1788),
.Y(n_1871)
);

OAI33xp33_ASAP7_75t_L g1872 ( 
.A1(n_1863),
.A2(n_1785),
.A3(n_1763),
.B1(n_1779),
.B2(n_1772),
.B3(n_1746),
.Y(n_1872)
);

OA211x2_ASAP7_75t_L g1873 ( 
.A1(n_1831),
.A2(n_1810),
.B(n_1755),
.C(n_1762),
.Y(n_1873)
);

NAND2xp33_ASAP7_75t_L g1874 ( 
.A(n_1862),
.B(n_1802),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1842),
.B(n_1847),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1842),
.B(n_1793),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1847),
.B(n_1790),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1826),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1859),
.Y(n_1879)
);

AOI211xp5_ASAP7_75t_SL g1880 ( 
.A1(n_1865),
.A2(n_1770),
.B(n_1814),
.C(n_1762),
.Y(n_1880)
);

OR2x6_ASAP7_75t_L g1881 ( 
.A(n_1834),
.B(n_1796),
.Y(n_1881)
);

INVxp67_ASAP7_75t_SL g1882 ( 
.A(n_1830),
.Y(n_1882)
);

INVx4_ASAP7_75t_L g1883 ( 
.A(n_1848),
.Y(n_1883)
);

INVx5_ASAP7_75t_SL g1884 ( 
.A(n_1835),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1845),
.B(n_1775),
.Y(n_1885)
);

OAI33xp33_ASAP7_75t_L g1886 ( 
.A1(n_1841),
.A2(n_1785),
.A3(n_1763),
.B1(n_1748),
.B2(n_1754),
.B3(n_1813),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1836),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1846),
.B(n_1771),
.Y(n_1888)
);

INVxp67_ASAP7_75t_L g1889 ( 
.A(n_1832),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1859),
.Y(n_1890)
);

AND2x4_ASAP7_75t_L g1891 ( 
.A(n_1845),
.B(n_1783),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1845),
.Y(n_1892)
);

OAI31xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1854),
.A2(n_1760),
.A3(n_1813),
.B(n_1796),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1858),
.Y(n_1894)
);

AND2x2_ASAP7_75t_L g1895 ( 
.A(n_1844),
.B(n_1794),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1845),
.Y(n_1896)
);

INVxp67_ASAP7_75t_L g1897 ( 
.A(n_1832),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1836),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1844),
.B(n_1794),
.Y(n_1899)
);

OR2x2_ASAP7_75t_L g1900 ( 
.A(n_1838),
.B(n_1784),
.Y(n_1900)
);

OA21x2_ASAP7_75t_L g1901 ( 
.A1(n_1825),
.A2(n_1818),
.B(n_1648),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1834),
.Y(n_1902)
);

BUFx3_ASAP7_75t_L g1903 ( 
.A(n_1849),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1837),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1837),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1827),
.B(n_1821),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1827),
.B(n_1821),
.Y(n_1907)
);

HB1xp67_ASAP7_75t_L g1908 ( 
.A(n_1853),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1838),
.B(n_1766),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1841),
.B(n_1766),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1864),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1850),
.B(n_1792),
.Y(n_1912)
);

INVx3_ASAP7_75t_L g1913 ( 
.A(n_1824),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1870),
.B(n_1902),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1870),
.B(n_1829),
.Y(n_1915)
);

INVx1_ASAP7_75t_SL g1916 ( 
.A(n_1902),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1875),
.B(n_1833),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1869),
.Y(n_1918)
);

AND2x4_ASAP7_75t_L g1919 ( 
.A(n_1885),
.B(n_1862),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1879),
.Y(n_1920)
);

INVxp67_ASAP7_75t_SL g1921 ( 
.A(n_1874),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1908),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1869),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1889),
.B(n_1861),
.Y(n_1924)
);

INVx1_ASAP7_75t_SL g1925 ( 
.A(n_1900),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1897),
.B(n_1861),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1867),
.B(n_1800),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1871),
.B(n_1840),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1900),
.B(n_1840),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1878),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1895),
.B(n_1849),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1878),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1887),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1871),
.B(n_1850),
.Y(n_1934)
);

OR2x2_ASAP7_75t_L g1935 ( 
.A(n_1894),
.B(n_1855),
.Y(n_1935)
);

AND2x4_ASAP7_75t_L g1936 ( 
.A(n_1885),
.B(n_1843),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1912),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1895),
.B(n_1839),
.Y(n_1938)
);

AND2x4_ASAP7_75t_L g1939 ( 
.A(n_1885),
.B(n_1843),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1887),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1898),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1898),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1912),
.Y(n_1943)
);

NAND2x1_ASAP7_75t_L g1944 ( 
.A(n_1881),
.B(n_1824),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1879),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1904),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1879),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1904),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1905),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1890),
.Y(n_1950)
);

AOI22xp33_ASAP7_75t_L g1951 ( 
.A1(n_1873),
.A2(n_1764),
.B1(n_1780),
.B2(n_1767),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1905),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1885),
.B(n_1864),
.Y(n_1953)
);

AOI221xp5_ASAP7_75t_L g1954 ( 
.A1(n_1872),
.A2(n_1857),
.B1(n_1851),
.B2(n_1856),
.C(n_1852),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1910),
.Y(n_1955)
);

AND2x4_ASAP7_75t_L g1956 ( 
.A(n_1891),
.B(n_1866),
.Y(n_1956)
);

INVx1_ASAP7_75t_SL g1957 ( 
.A(n_1903),
.Y(n_1957)
);

BUFx2_ASAP7_75t_L g1958 ( 
.A(n_1883),
.Y(n_1958)
);

INVx1_ASAP7_75t_SL g1959 ( 
.A(n_1903),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1925),
.B(n_1909),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1921),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1918),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1919),
.B(n_1891),
.Y(n_1963)
);

NOR2xp33_ASAP7_75t_L g1964 ( 
.A(n_1925),
.B(n_1886),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1920),
.Y(n_1965)
);

NOR2xp33_ASAP7_75t_L g1966 ( 
.A(n_1928),
.B(n_1886),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1929),
.B(n_1935),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1918),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1919),
.B(n_1899),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1923),
.Y(n_1970)
);

INVxp67_ASAP7_75t_L g1971 ( 
.A(n_1958),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1923),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1920),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1929),
.B(n_1909),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1919),
.B(n_1891),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1930),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1930),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1935),
.B(n_1882),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1922),
.B(n_1877),
.Y(n_1979)
);

AND2x4_ASAP7_75t_L g1980 ( 
.A(n_1919),
.B(n_1891),
.Y(n_1980)
);

INVx2_ASAP7_75t_L g1981 ( 
.A(n_1920),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1958),
.B(n_1884),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1914),
.B(n_1884),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1937),
.B(n_1877),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1945),
.Y(n_1985)
);

OR2x6_ASAP7_75t_L g1986 ( 
.A(n_1944),
.B(n_1883),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1932),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1943),
.B(n_1934),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1914),
.B(n_1884),
.Y(n_1989)
);

INVxp67_ASAP7_75t_L g1990 ( 
.A(n_1934),
.Y(n_1990)
);

NAND2x1p5_ASAP7_75t_L g1991 ( 
.A(n_1916),
.B(n_1883),
.Y(n_1991)
);

INVxp67_ASAP7_75t_L g1992 ( 
.A(n_1916),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1945),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1955),
.B(n_1883),
.Y(n_1994)
);

AND2x4_ASAP7_75t_L g1995 ( 
.A(n_1936),
.B(n_1892),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1954),
.B(n_1906),
.Y(n_1996)
);

INVx1_ASAP7_75t_SL g1997 ( 
.A(n_1957),
.Y(n_1997)
);

NAND4xp75_ASAP7_75t_L g1998 ( 
.A(n_1927),
.B(n_1873),
.C(n_1868),
.D(n_1901),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_SL g1999 ( 
.A(n_1951),
.B(n_1893),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1924),
.B(n_1906),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1924),
.B(n_1907),
.Y(n_2001)
);

NOR3xp33_ASAP7_75t_L g2002 ( 
.A(n_1944),
.B(n_1872),
.C(n_1868),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1926),
.B(n_1911),
.Y(n_2003)
);

INVx2_ASAP7_75t_SL g2004 ( 
.A(n_1957),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1932),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1945),
.Y(n_2006)
);

AND2x4_ASAP7_75t_L g2007 ( 
.A(n_2004),
.B(n_1936),
.Y(n_2007)
);

AND2x2_ASAP7_75t_SL g2008 ( 
.A(n_2002),
.B(n_1893),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1991),
.B(n_1936),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1991),
.B(n_1936),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1983),
.B(n_1939),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1966),
.B(n_1959),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1962),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1968),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1970),
.Y(n_2015)
);

OAI21xp33_ASAP7_75t_L g2016 ( 
.A1(n_1999),
.A2(n_1880),
.B(n_1926),
.Y(n_2016)
);

AOI211x1_ASAP7_75t_L g2017 ( 
.A1(n_1999),
.A2(n_1915),
.B(n_1907),
.C(n_1876),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_1966),
.B(n_1964),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1972),
.Y(n_2019)
);

HB1xp67_ASAP7_75t_L g2020 ( 
.A(n_2004),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1976),
.Y(n_2021)
);

OA21x2_ASAP7_75t_L g2022 ( 
.A1(n_1998),
.A2(n_1950),
.B(n_1947),
.Y(n_2022)
);

NAND2x1p5_ASAP7_75t_L g2023 ( 
.A(n_1982),
.B(n_1959),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1967),
.B(n_1888),
.Y(n_2024)
);

INVx2_ASAP7_75t_SL g2025 ( 
.A(n_1983),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1965),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1997),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1964),
.B(n_1938),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1989),
.B(n_1939),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1996),
.A2(n_1881),
.B1(n_1901),
.B2(n_1848),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_1989),
.Y(n_2031)
);

OAI33xp33_ASAP7_75t_L g2032 ( 
.A1(n_1971),
.A2(n_1941),
.A3(n_1952),
.B1(n_1940),
.B2(n_1949),
.B3(n_1948),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1961),
.B(n_1938),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1986),
.Y(n_2034)
);

AND2x4_ASAP7_75t_SL g2035 ( 
.A(n_1986),
.B(n_1881),
.Y(n_2035)
);

NOR2x1_ASAP7_75t_L g2036 ( 
.A(n_1986),
.B(n_1881),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1982),
.B(n_1939),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1975),
.B(n_1939),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1992),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1977),
.Y(n_2040)
);

AND2x4_ASAP7_75t_L g2041 ( 
.A(n_1963),
.B(n_1953),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_1975),
.B(n_1915),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1965),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1960),
.B(n_1888),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1987),
.Y(n_2045)
);

AOI21xp33_ASAP7_75t_L g2046 ( 
.A1(n_2008),
.A2(n_1994),
.B(n_1986),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2008),
.B(n_2039),
.Y(n_2047)
);

AOI21xp33_ASAP7_75t_L g2048 ( 
.A1(n_2018),
.A2(n_1990),
.B(n_1988),
.Y(n_2048)
);

OAI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_2022),
.A2(n_1880),
.B(n_2000),
.Y(n_2049)
);

AOI22xp5_ASAP7_75t_L g2050 ( 
.A1(n_2016),
.A2(n_1980),
.B1(n_1963),
.B2(n_1881),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_2039),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_2020),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_2027),
.B(n_2001),
.Y(n_2053)
);

AND2x4_ASAP7_75t_L g2054 ( 
.A(n_2025),
.B(n_2031),
.Y(n_2054)
);

INVx1_ASAP7_75t_SL g2055 ( 
.A(n_2023),
.Y(n_2055)
);

OAI21xp5_ASAP7_75t_SL g2056 ( 
.A1(n_2030),
.A2(n_1980),
.B(n_1963),
.Y(n_2056)
);

OAI322xp33_ASAP7_75t_L g2057 ( 
.A1(n_2012),
.A2(n_1978),
.A3(n_2003),
.B1(n_1974),
.B2(n_2005),
.C1(n_1984),
.C2(n_1979),
.Y(n_2057)
);

OAI32xp33_ASAP7_75t_L g2058 ( 
.A1(n_2028),
.A2(n_2003),
.A3(n_1903),
.B1(n_1969),
.B2(n_1876),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_2013),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2013),
.Y(n_2060)
);

AOI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_2022),
.A2(n_1980),
.B1(n_1969),
.B2(n_1995),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2014),
.Y(n_2062)
);

AOI21xp33_ASAP7_75t_L g2063 ( 
.A1(n_2022),
.A2(n_1981),
.B(n_1973),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_2014),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2015),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2015),
.Y(n_2066)
);

AOI21xp33_ASAP7_75t_L g2067 ( 
.A1(n_2022),
.A2(n_1981),
.B(n_1973),
.Y(n_2067)
);

AOI22xp5_ASAP7_75t_L g2068 ( 
.A1(n_2025),
.A2(n_1995),
.B1(n_1901),
.B2(n_1953),
.Y(n_2068)
);

OAI221xp5_ASAP7_75t_L g2069 ( 
.A1(n_2036),
.A2(n_1750),
.B1(n_1787),
.B2(n_1901),
.C(n_1756),
.Y(n_2069)
);

AOI22xp33_ASAP7_75t_L g2070 ( 
.A1(n_2032),
.A2(n_2031),
.B1(n_2033),
.B2(n_2035),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2011),
.B(n_1995),
.Y(n_2071)
);

OAI22xp33_ASAP7_75t_L g2072 ( 
.A1(n_2023),
.A2(n_1752),
.B1(n_1822),
.B2(n_1828),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2019),
.Y(n_2073)
);

AOI211xp5_ASAP7_75t_L g2074 ( 
.A1(n_2009),
.A2(n_1765),
.B(n_1761),
.C(n_1985),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2019),
.Y(n_2075)
);

AND2x2_ASAP7_75t_L g2076 ( 
.A(n_2051),
.B(n_2011),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2059),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2071),
.B(n_2029),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2054),
.B(n_2029),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_SL g2080 ( 
.A(n_2072),
.B(n_2017),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_2054),
.B(n_2037),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2049),
.A2(n_2037),
.B1(n_2041),
.B2(n_2035),
.Y(n_2082)
);

NAND3xp33_ASAP7_75t_L g2083 ( 
.A(n_2047),
.B(n_2034),
.C(n_2021),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2052),
.B(n_2042),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2070),
.B(n_2042),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_2053),
.B(n_1799),
.Y(n_2086)
);

NAND3xp33_ASAP7_75t_L g2087 ( 
.A(n_2070),
.B(n_2034),
.C(n_2021),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2060),
.Y(n_2088)
);

XNOR2x1_ASAP7_75t_L g2089 ( 
.A(n_2050),
.B(n_2023),
.Y(n_2089)
);

OAI21xp5_ASAP7_75t_L g2090 ( 
.A1(n_2069),
.A2(n_2034),
.B(n_2010),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2062),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2064),
.Y(n_2092)
);

AOI222xp33_ASAP7_75t_SL g2093 ( 
.A1(n_2055),
.A2(n_2045),
.B1(n_2040),
.B2(n_2043),
.C1(n_2026),
.C2(n_1985),
.Y(n_2093)
);

OA21x2_ASAP7_75t_L g2094 ( 
.A1(n_2063),
.A2(n_2043),
.B(n_2026),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2065),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2066),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_2061),
.Y(n_2097)
);

AOI22xp5_ASAP7_75t_L g2098 ( 
.A1(n_2069),
.A2(n_2010),
.B1(n_2009),
.B2(n_2007),
.Y(n_2098)
);

OAI22xp5_ASAP7_75t_SL g2099 ( 
.A1(n_2087),
.A2(n_1799),
.B1(n_2074),
.B2(n_2073),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_2094),
.Y(n_2100)
);

OAI32xp33_ASAP7_75t_L g2101 ( 
.A1(n_2080),
.A2(n_2046),
.A3(n_2048),
.B1(n_2067),
.B2(n_2075),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2077),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2077),
.Y(n_2103)
);

AOI21xp33_ASAP7_75t_L g2104 ( 
.A1(n_2089),
.A2(n_2056),
.B(n_2058),
.Y(n_2104)
);

NAND4xp25_ASAP7_75t_L g2105 ( 
.A(n_2082),
.B(n_2068),
.C(n_2041),
.D(n_2040),
.Y(n_2105)
);

AOI21xp33_ASAP7_75t_L g2106 ( 
.A1(n_2089),
.A2(n_2072),
.B(n_2045),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2092),
.Y(n_2107)
);

INVx1_ASAP7_75t_SL g2108 ( 
.A(n_2081),
.Y(n_2108)
);

INVx1_ASAP7_75t_SL g2109 ( 
.A(n_2081),
.Y(n_2109)
);

AOI222xp33_ASAP7_75t_L g2110 ( 
.A1(n_2085),
.A2(n_2057),
.B1(n_2007),
.B2(n_2041),
.C1(n_2038),
.C2(n_1993),
.Y(n_2110)
);

INVxp67_ASAP7_75t_L g2111 ( 
.A(n_2076),
.Y(n_2111)
);

OAI31xp33_ASAP7_75t_SL g2112 ( 
.A1(n_2090),
.A2(n_2007),
.A3(n_2038),
.B(n_1765),
.Y(n_2112)
);

XNOR2xp5_ASAP7_75t_L g2113 ( 
.A(n_2076),
.B(n_1759),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_2079),
.B(n_2024),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2100),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2108),
.B(n_2097),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2109),
.Y(n_2117)
);

NOR3xp33_ASAP7_75t_L g2118 ( 
.A(n_2101),
.B(n_2083),
.C(n_2111),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2100),
.B(n_2088),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2114),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2102),
.Y(n_2121)
);

A2O1A1Ixp33_ASAP7_75t_L g2122 ( 
.A1(n_2104),
.A2(n_2098),
.B(n_2097),
.C(n_2086),
.Y(n_2122)
);

NOR3xp33_ASAP7_75t_L g2123 ( 
.A(n_2099),
.B(n_2084),
.C(n_2091),
.Y(n_2123)
);

NOR3xp33_ASAP7_75t_L g2124 ( 
.A(n_2105),
.B(n_2095),
.C(n_2092),
.Y(n_2124)
);

NOR3xp33_ASAP7_75t_L g2125 ( 
.A(n_2106),
.B(n_2096),
.C(n_2095),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2103),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2107),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2113),
.B(n_2079),
.Y(n_2128)
);

NOR2x1_ASAP7_75t_L g2129 ( 
.A(n_2113),
.B(n_2094),
.Y(n_2129)
);

NAND3x1_ASAP7_75t_L g2130 ( 
.A(n_2129),
.B(n_2112),
.C(n_2096),
.Y(n_2130)
);

O2A1O1Ixp5_ASAP7_75t_L g2131 ( 
.A1(n_2115),
.A2(n_2078),
.B(n_2093),
.C(n_2094),
.Y(n_2131)
);

AOI221xp5_ASAP7_75t_L g2132 ( 
.A1(n_2118),
.A2(n_2078),
.B1(n_2110),
.B2(n_2094),
.C(n_2044),
.Y(n_2132)
);

INVx1_ASAP7_75t_SL g2133 ( 
.A(n_2128),
.Y(n_2133)
);

AOI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_2124),
.A2(n_2125),
.B1(n_2122),
.B2(n_2123),
.C(n_2116),
.Y(n_2134)
);

AOI22xp5_ASAP7_75t_L g2135 ( 
.A1(n_2117),
.A2(n_2044),
.B1(n_1956),
.B2(n_1953),
.Y(n_2135)
);

OAI31xp33_ASAP7_75t_L g2136 ( 
.A1(n_2119),
.A2(n_2024),
.A3(n_1953),
.B(n_1956),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2120),
.A2(n_2006),
.B1(n_1993),
.B2(n_1753),
.Y(n_2137)
);

AOI221xp5_ASAP7_75t_L g2138 ( 
.A1(n_2134),
.A2(n_2132),
.B1(n_2131),
.B2(n_2133),
.C(n_2119),
.Y(n_2138)
);

AOI221x1_ASAP7_75t_SL g2139 ( 
.A1(n_2130),
.A2(n_2127),
.B1(n_2126),
.B2(n_2121),
.C(n_2006),
.Y(n_2139)
);

NOR3xp33_ASAP7_75t_L g2140 ( 
.A(n_2135),
.B(n_1749),
.C(n_1735),
.Y(n_2140)
);

XOR2x2_ASAP7_75t_L g2141 ( 
.A(n_2137),
.B(n_1735),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2136),
.B(n_1956),
.Y(n_2142)
);

O2A1O1Ixp33_ASAP7_75t_L g2143 ( 
.A1(n_2131),
.A2(n_1956),
.B(n_1896),
.C(n_1892),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2131),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_R g2145 ( 
.A(n_2133),
.B(n_1745),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2144),
.Y(n_2146)
);

OAI21xp5_ASAP7_75t_L g2147 ( 
.A1(n_2138),
.A2(n_1931),
.B(n_1933),
.Y(n_2147)
);

INVx3_ASAP7_75t_SL g2148 ( 
.A(n_2141),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2139),
.Y(n_2149)
);

OR2x2_ASAP7_75t_L g2150 ( 
.A(n_2142),
.B(n_1947),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2143),
.B(n_1931),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2145),
.Y(n_2152)
);

NAND4xp25_ASAP7_75t_L g2153 ( 
.A(n_2146),
.B(n_2140),
.C(n_1757),
.D(n_1780),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2148),
.B(n_1933),
.Y(n_2154)
);

AND2x2_ASAP7_75t_L g2155 ( 
.A(n_2147),
.B(n_1917),
.Y(n_2155)
);

AND2x2_ASAP7_75t_L g2156 ( 
.A(n_2155),
.B(n_2147),
.Y(n_2156)
);

CKINVDCx20_ASAP7_75t_R g2157 ( 
.A(n_2156),
.Y(n_2157)
);

OAI21x1_ASAP7_75t_L g2158 ( 
.A1(n_2157),
.A2(n_2149),
.B(n_2152),
.Y(n_2158)
);

OAI22x1_ASAP7_75t_SL g2159 ( 
.A1(n_2157),
.A2(n_2154),
.B1(n_2153),
.B2(n_2150),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2159),
.Y(n_2160)
);

OAI22x1_ASAP7_75t_L g2161 ( 
.A1(n_2158),
.A2(n_2151),
.B1(n_1946),
.B2(n_1952),
.Y(n_2161)
);

OAI221xp5_ASAP7_75t_SL g2162 ( 
.A1(n_2160),
.A2(n_1941),
.B1(n_1942),
.B2(n_1949),
.C(n_1948),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2161),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_2163),
.B(n_1947),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2164),
.Y(n_2165)
);

INVx1_ASAP7_75t_L g2166 ( 
.A(n_2165),
.Y(n_2166)
);

OAI221xp5_ASAP7_75t_R g2167 ( 
.A1(n_2166),
.A2(n_2162),
.B1(n_1913),
.B2(n_1946),
.C(n_1940),
.Y(n_2167)
);

AOI211xp5_ASAP7_75t_L g2168 ( 
.A1(n_2167),
.A2(n_1758),
.B(n_1737),
.C(n_1739),
.Y(n_2168)
);


endmodule