module fake_jpeg_30827_n_136 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_136);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx4f_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_0),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_60),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_65),
.A2(n_60),
.B1(n_49),
.B2(n_46),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_74),
.Y(n_93)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_53),
.B1(n_60),
.B2(n_45),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_55),
.B1(n_20),
.B2(n_26),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_52),
.B1(n_59),
.B2(n_54),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_52),
.B1(n_51),
.B2(n_58),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_77),
.C(n_2),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_57),
.B1(n_50),
.B2(n_48),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_3),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_76),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_85),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_106)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_84),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_1),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_1),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_91),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_5),
.Y(n_107)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_28),
.C(n_42),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_104),
.C(n_105),
.Y(n_117)
);

OAI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_18),
.B(n_41),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_87),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_93),
.B(n_17),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_16),
.C(n_40),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_98),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_43),
.B1(n_29),
.B2(n_30),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_110),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_96),
.A2(n_94),
.B1(n_33),
.B2(n_35),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_122),
.B(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_115),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_10),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_15),
.C(n_31),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_105),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_12),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_103),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_122)
);

BUFx24_ASAP7_75t_SL g129 ( 
.A(n_126),
.Y(n_129)
);

OAI321xp33_ASAP7_75t_L g130 ( 
.A1(n_127),
.A2(n_101),
.A3(n_116),
.B1(n_104),
.B2(n_99),
.C(n_112),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_125),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_124),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_132),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_129),
.A3(n_128),
.B1(n_121),
.B2(n_113),
.C1(n_120),
.C2(n_126),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_117),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_117),
.Y(n_136)
);


endmodule