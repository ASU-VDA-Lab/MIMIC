module real_jpeg_29915_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_313, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_313;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_0),
.A2(n_64),
.B1(n_65),
.B2(n_136),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_0),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_0),
.A2(n_48),
.B1(n_51),
.B2(n_136),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_136),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_0),
.A2(n_29),
.B1(n_30),
.B2(n_136),
.Y(n_250)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_1),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_2),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_2),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_2),
.A2(n_34),
.B1(n_35),
.B2(n_70),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_2),
.A2(n_48),
.B1(n_51),
.B2(n_70),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_3),
.B(n_35),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g152 ( 
.A1(n_3),
.A2(n_35),
.B(n_43),
.C(n_150),
.D(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_32),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_3),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_83),
.B(n_167),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_30),
.B(n_31),
.C(n_198),
.D(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_30),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_3),
.A2(n_29),
.B(n_62),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_182),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_34),
.B1(n_35),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_4),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_4),
.A2(n_48),
.B1(n_51),
.B2(n_162),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_162),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_4),
.A2(n_64),
.B1(n_65),
.B2(n_162),
.Y(n_267)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_5),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_7),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_7),
.A2(n_48),
.B1(n_51),
.B2(n_67),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_7),
.A2(n_34),
.B1(n_35),
.B2(n_67),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_8),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_34),
.B1(n_35),
.B2(n_98),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_8),
.A2(n_48),
.B1(n_51),
.B2(n_98),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_98),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_34),
.B1(n_35),
.B2(n_54),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_10),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_54),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_35),
.B(n_44),
.C(n_47),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_40),
.B1(n_48),
.B2(n_51),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_15),
.A2(n_28),
.B1(n_34),
.B2(n_35),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_15),
.A2(n_28),
.B1(n_64),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_15),
.A2(n_28),
.B1(n_48),
.B2(n_51),
.Y(n_237)
);

INVx11_ASAP7_75t_SL g50 ( 
.A(n_16),
.Y(n_50)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_114),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_113),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_99),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_21),
.B(n_99),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_80),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_73),
.Y(n_140)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_57),
.B2(n_71),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_41),
.B1(n_55),
.B2(n_56),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_26),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_26),
.B(n_56),
.C(n_57),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_39),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_27),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_77)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_29),
.A2(n_30),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_29),
.A2(n_35),
.A3(n_198),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_31),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_31),
.A2(n_32),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_34),
.Y(n_35)
);

AOI32xp33_ASAP7_75t_L g149 ( 
.A1(n_34),
.A2(n_46),
.A3(n_51),
.B1(n_150),
.B2(n_151),
.Y(n_149)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_34),
.B(n_36),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_36),
.Y(n_209)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_39),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_41),
.A2(n_56),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_52),
.B(n_53),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_42),
.A2(n_52),
.B1(n_93),
.B2(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_42),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_42),
.A2(n_52),
.B1(n_130),
.B2(n_253),
.Y(n_272)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_47),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_43),
.A2(n_47),
.B1(n_75),
.B2(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_43),
.B(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_43),
.A2(n_47),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_45),
.B(n_48),
.Y(n_151)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2x1_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_51),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_52),
.B(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_52),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_52),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_52),
.A2(n_163),
.B(n_253),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_53),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_57),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_71),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_68),
.B1(n_69),
.B2(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_58),
.A2(n_134),
.B(n_137),
.Y(n_133)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_59),
.B(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_59),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_59),
.A2(n_60),
.B1(n_135),
.B2(n_267),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_60),
.B(n_97),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_61),
.A2(n_64),
.B(n_182),
.C(n_240),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_64),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_68),
.B(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_68),
.B(n_182),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_68),
.A2(n_96),
.B(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g122 ( 
.A1(n_73),
.A2(n_74),
.B(n_77),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_79),
.A2(n_108),
.B1(n_110),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_80),
.A2(n_81),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_89),
.B(n_94),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_82),
.A2(n_94),
.B1(n_95),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_82),
.A2(n_90),
.B1(n_91),
.B2(n_120),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_85),
.B(n_88),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_88),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_83),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_83),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_83),
.B(n_169),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_83),
.A2(n_85),
.B1(n_207),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_83),
.A2(n_87),
.B1(n_127),
.B2(n_271),
.Y(n_270)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_85),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_85),
.A2(n_174),
.B(n_184),
.Y(n_183)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g128 ( 
.A(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_86),
.B(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_86),
.A2(n_185),
.B(n_206),
.Y(n_205)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_87),
.B(n_182),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_112),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_108),
.A2(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_110),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_110),
.A2(n_132),
.B(n_217),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_141),
.B(n_311),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_138),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_116),
.B(n_138),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_123),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_299)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_123),
.B(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.C(n_133),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_124),
.A2(n_125),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_126),
.B(n_129),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_131),
.B(n_133),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_137),
.Y(n_245)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI321xp33_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_291),
.A3(n_300),
.B1(n_305),
.B2(n_310),
.C(n_313),
.Y(n_141)
);

NOR3xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_255),
.C(n_287),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_229),
.B(n_254),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_212),
.B(n_228),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_193),
.B(n_211),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_170),
.B(n_192),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_148),
.B(n_155),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_152),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_154),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_160),
.C(n_165),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_166),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_179),
.B(n_191),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_178),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_172),
.B(n_178),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_175),
.A2(n_177),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_186),
.B(n_190),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_183),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_194),
.B(n_195),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_196),
.B(n_213),
.Y(n_228)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_201),
.CI(n_204),
.CON(n_196),
.SN(n_196)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_199),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_203),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_224),
.C(n_225),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_220),
.C(n_221),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_222),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_231),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_242),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_234),
.C(n_242),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_235),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_237),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_241),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_248),
.C(n_251),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_256),
.A2(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_274),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_257),
.B(n_274),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_269),
.C(n_273),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_261),
.C(n_268),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_265),
.B2(n_268),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_265),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_273),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_272),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_274)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_275),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_276),
.B(n_283),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_283),
.C(n_286),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_280),
.C(n_281),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_289),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_298),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_298),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.C(n_297),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_301),
.A2(n_306),
.B(n_309),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_303),
.Y(n_309)
);


endmodule