module fake_netlist_6_4829_n_171 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_25, n_171);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_25;

output n_171;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_102;
wire n_87;
wire n_32;
wire n_85;
wire n_99;
wire n_130;
wire n_66;
wire n_84;
wire n_78;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_81;
wire n_59;
wire n_76;
wire n_36;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_107;
wire n_71;
wire n_74;
wire n_123;
wire n_136;
wire n_72;
wire n_89;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_35;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_31;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVxp67_ASAP7_75t_SL g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVxp67_ASAP7_75t_SL g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_28),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_46),
.B1(n_37),
.B2(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_32),
.B(n_3),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

OA21x2_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_3),
.B(n_4),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_34),
.B(n_5),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_54),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_33),
.B1(n_44),
.B2(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_49),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_67),
.Y(n_83)
);

OAI221xp5_ASAP7_75t_L g84 ( 
.A1(n_59),
.A2(n_38),
.B1(n_42),
.B2(n_43),
.C(n_50),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_50),
.Y(n_86)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_62),
.Y(n_95)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_88),
.B(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_86),
.B(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_77),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_69),
.B1(n_61),
.B2(n_63),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_74),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_83),
.A2(n_44),
.B1(n_33),
.B2(n_73),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_83),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_91),
.B(n_90),
.Y(n_105)
);

AND2x4_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_85),
.Y(n_108)
);

NOR2xp67_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_81),
.Y(n_109)
);

AND2x4_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_71),
.Y(n_110)
);

OR2x6_ASAP7_75t_SL g111 ( 
.A(n_103),
.B(n_43),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_106),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_99),
.B1(n_98),
.B2(n_87),
.Y(n_113)
);

AO32x2_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_99),
.A3(n_87),
.B1(n_96),
.B2(n_69),
.Y(n_114)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_94),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_104),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_87),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_116),
.A2(n_112),
.B(n_110),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_108),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_84),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_107),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_118),
.B(n_113),
.Y(n_126)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_118),
.B(n_105),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_120),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_115),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_107),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_114),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_125),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_128),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_114),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_129),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_130),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_129),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_140),
.B(n_126),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_124),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_143),
.B(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_138),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_138),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_146),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_147),
.B(n_145),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_128),
.B1(n_127),
.B2(n_124),
.Y(n_155)
);

AOI221x1_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_68),
.B1(n_66),
.B2(n_137),
.C(n_70),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_131),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_137),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_153),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_135),
.B(n_134),
.Y(n_161)
);

OAI211xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_75),
.B(n_10),
.C(n_9),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_161),
.A2(n_135),
.B1(n_133),
.B2(n_132),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_133),
.C(n_78),
.Y(n_165)
);

AOI322xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_10),
.A3(n_133),
.B1(n_110),
.B2(n_78),
.C1(n_89),
.C2(n_14),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_89),
.B1(n_110),
.B2(n_93),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_SL g168 ( 
.A(n_166),
.B(n_16),
.C(n_17),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_110),
.C(n_93),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_168),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_169),
.B(n_164),
.C(n_167),
.Y(n_171)
);


endmodule