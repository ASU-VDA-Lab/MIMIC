module fake_netlist_5_391_n_1494 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_376, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_378, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_372, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_373, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_375, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_371, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_377, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1494);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_376;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_378;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_372;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_375;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_371;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1494;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_1483;
wire n_1314;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_696;
wire n_550;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_851;
wire n_615;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1233;
wire n_526;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_1163;
wire n_906;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_141),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_83),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_97),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_151),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_168),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_350),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_374),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_59),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_288),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_287),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_80),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_11),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_226),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_5),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_260),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_231),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_33),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_55),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_272),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_153),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_117),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_198),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_94),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_376),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_222),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_46),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_266),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_225),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_180),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_183),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_378),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_297),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_277),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_305),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_100),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_14),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_377),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_111),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_337),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_148),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_241),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_216),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_108),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_17),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_306),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_40),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_301),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_162),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_317),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_133),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_293),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_65),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_357),
.Y(n_432)
);

INVxp67_ASAP7_75t_SL g433 ( 
.A(n_320),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_167),
.Y(n_434)
);

BUFx8_ASAP7_75t_SL g435 ( 
.A(n_77),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_192),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_258),
.Y(n_437)
);

BUFx3_ASAP7_75t_L g438 ( 
.A(n_228),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_275),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_307),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_159),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_45),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_223),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_324),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_191),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_21),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_179),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_9),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_318),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_303),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_146),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_237),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_158),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_250),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_359),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_369),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_234),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_2),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_373),
.Y(n_459)
);

BUFx5_ASAP7_75t_L g460 ( 
.A(n_81),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_285),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_155),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_58),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_177),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_219),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_217),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_274),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_143),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_215),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_299),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_365),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_101),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_334),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_355),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_344),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_62),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_259),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_11),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_63),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_321),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_92),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_208),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_67),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_181),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_138),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_120),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_327),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_170),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_109),
.Y(n_489)
);

INVx4_ASAP7_75t_R g490 ( 
.A(n_224),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_171),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_343),
.Y(n_492)
);

BUFx10_ASAP7_75t_L g493 ( 
.A(n_302),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_22),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_98),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_322),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_84),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_351),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_25),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_356),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_340),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_21),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_332),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_353),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_60),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_67),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_113),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_76),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_45),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_326),
.Y(n_510)
);

INVx2_ASAP7_75t_SL g511 ( 
.A(n_367),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_184),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_48),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_319),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_121),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_118),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_206),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_210),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_41),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_131),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_262),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_103),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_161),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_126),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_227),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_16),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_235),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_130),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_174),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_116),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_0),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_129),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_119),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_323),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_54),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_366),
.Y(n_536)
);

CKINVDCx16_ASAP7_75t_R g537 ( 
.A(n_88),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_333),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_349),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_14),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_341),
.Y(n_541)
);

INVx1_ASAP7_75t_SL g542 ( 
.A(n_214),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_18),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_165),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_347),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_265),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g547 ( 
.A(n_361),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_104),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_46),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_295),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_99),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_127),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_246),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_0),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_76),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_182),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_281),
.Y(n_557)
);

BUFx2_ASAP7_75t_L g558 ( 
.A(n_105),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_279),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_19),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_29),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_147),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_201),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_230),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_382),
.B(n_1),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_409),
.Y(n_566)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_382),
.B(n_1),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_554),
.B(n_2),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_554),
.B(n_3),
.Y(n_569)
);

BUFx12f_ASAP7_75t_L g570 ( 
.A(n_386),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_513),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_448),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_397),
.B(n_3),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_448),
.Y(n_574)
);

CKINVDCx6p67_ASAP7_75t_R g575 ( 
.A(n_386),
.Y(n_575)
);

BUFx12f_ASAP7_75t_L g576 ( 
.A(n_386),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_435),
.Y(n_577)
);

BUFx8_ASAP7_75t_SL g578 ( 
.A(n_435),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_409),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g580 ( 
.A(n_409),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_397),
.B(n_4),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_448),
.B(n_4),
.Y(n_582)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_449),
.Y(n_583)
);

BUFx8_ASAP7_75t_SL g584 ( 
.A(n_390),
.Y(n_584)
);

XNOR2x1_ASAP7_75t_L g585 ( 
.A(n_392),
.B(n_5),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_448),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_396),
.Y(n_587)
);

INVx3_ASAP7_75t_L g588 ( 
.A(n_404),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_425),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_409),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_454),
.B(n_547),
.Y(n_591)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_465),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_442),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_460),
.Y(n_594)
);

INVx5_ASAP7_75t_L g595 ( 
.A(n_465),
.Y(n_595)
);

BUFx8_ASAP7_75t_SL g596 ( 
.A(n_558),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_465),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_417),
.B(n_6),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_476),
.Y(n_599)
);

BUFx12f_ASAP7_75t_L g600 ( 
.A(n_493),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_460),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_404),
.Y(n_602)
);

INVx5_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g604 ( 
.A(n_493),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_431),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_454),
.B(n_6),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_438),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_438),
.B(n_7),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_460),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_518),
.B(n_7),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_529),
.B(n_417),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_529),
.B(n_440),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_551),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_493),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_551),
.Y(n_615)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_551),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_551),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_536),
.B(n_8),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_440),
.B(n_8),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_498),
.B(n_532),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_469),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_498),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_532),
.B(n_9),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_541),
.B(n_511),
.Y(n_624)
);

INVx5_ASAP7_75t_L g625 ( 
.A(n_514),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_460),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_431),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_541),
.B(n_10),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_543),
.B(n_10),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_381),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_543),
.B(n_385),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_387),
.B(n_12),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_537),
.B(n_12),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_388),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_407),
.B(n_13),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_542),
.B(n_13),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_460),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_389),
.B(n_15),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_391),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_433),
.B(n_15),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_499),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_460),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_509),
.Y(n_643)
);

BUFx2_ASAP7_75t_L g644 ( 
.A(n_395),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_460),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_519),
.B(n_16),
.Y(n_646)
);

INVx5_ASAP7_75t_L g647 ( 
.A(n_490),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_379),
.Y(n_648)
);

BUFx12f_ASAP7_75t_L g649 ( 
.A(n_414),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_394),
.B(n_17),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_555),
.B(n_18),
.Y(n_651)
);

AND2x4_ASAP7_75t_L g652 ( 
.A(n_410),
.B(n_19),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_560),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_412),
.B(n_20),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_423),
.B(n_20),
.Y(n_655)
);

BUFx8_ASAP7_75t_SL g656 ( 
.A(n_398),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_413),
.B(n_22),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_380),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_383),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_415),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_420),
.B(n_23),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_384),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_428),
.B(n_23),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_429),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_393),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_574),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_572),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_591),
.B(n_662),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_622),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_647),
.B(n_399),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_614),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_586),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_611),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_622),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_SL g675 ( 
.A1(n_571),
.A2(n_458),
.B1(n_463),
.B2(n_446),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_611),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_665),
.B(n_441),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_610),
.A2(n_479),
.B1(n_483),
.B2(n_478),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_586),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_621),
.B(n_447),
.Y(n_680)
);

AO22x2_ASAP7_75t_L g681 ( 
.A1(n_610),
.A2(n_456),
.B1(n_457),
.B2(n_453),
.Y(n_681)
);

OAI22xp33_ASAP7_75t_R g682 ( 
.A1(n_571),
.A2(n_462),
.B1(n_466),
.B2(n_459),
.Y(n_682)
);

OAI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_631),
.A2(n_619),
.B1(n_628),
.B2(n_598),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_SL g684 ( 
.A1(n_631),
.A2(n_480),
.B1(n_487),
.B2(n_473),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_585),
.A2(n_416),
.B1(n_421),
.B2(n_400),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_647),
.B(n_401),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_647),
.B(n_402),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_566),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_647),
.B(n_403),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_566),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_SL g691 ( 
.A1(n_598),
.A2(n_491),
.B1(n_492),
.B2(n_489),
.Y(n_691)
);

AO22x1_ASAP7_75t_L g692 ( 
.A1(n_573),
.A2(n_581),
.B1(n_623),
.B2(n_569),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_583),
.B(n_494),
.Y(n_693)
);

NOR2x1p5_ASAP7_75t_L g694 ( 
.A(n_600),
.B(n_502),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_640),
.A2(n_506),
.B1(n_508),
.B2(n_505),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_644),
.B(n_405),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_L g697 ( 
.A1(n_640),
.A2(n_531),
.B1(n_535),
.B2(n_526),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_566),
.Y(n_698)
);

OAI22xp33_ASAP7_75t_SL g699 ( 
.A1(n_619),
.A2(n_628),
.B1(n_661),
.B2(n_654),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_579),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_622),
.Y(n_701)
);

AO22x2_ASAP7_75t_L g702 ( 
.A1(n_573),
.A2(n_496),
.B1(n_500),
.B2(n_495),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_579),
.Y(n_703)
);

OA22x2_ASAP7_75t_L g704 ( 
.A1(n_643),
.A2(n_549),
.B1(n_561),
.B2(n_540),
.Y(n_704)
);

BUFx6f_ASAP7_75t_SL g705 ( 
.A(n_581),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_607),
.B(n_406),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_629),
.A2(n_646),
.B1(n_651),
.B2(n_643),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_565),
.B(n_567),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_SL g709 ( 
.A1(n_654),
.A2(n_530),
.B1(n_533),
.B2(n_512),
.Y(n_709)
);

XNOR2xp5_ASAP7_75t_L g710 ( 
.A(n_577),
.B(n_426),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_605),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_579),
.Y(n_712)
);

OAI22xp33_ASAP7_75t_L g713 ( 
.A1(n_661),
.A2(n_437),
.B1(n_455),
.B2(n_434),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_629),
.A2(n_557),
.B1(n_538),
.B2(n_411),
.Y(n_714)
);

OAI22xp33_ASAP7_75t_L g715 ( 
.A1(n_575),
.A2(n_548),
.B1(n_525),
.B2(n_418),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_606),
.B(n_408),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_605),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_646),
.A2(n_651),
.B1(n_635),
.B2(n_636),
.Y(n_718)
);

AO22x2_ASAP7_75t_L g719 ( 
.A1(n_623),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_635),
.A2(n_422),
.B1(n_424),
.B2(n_419),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_587),
.Y(n_721)
);

AO22x2_ASAP7_75t_L g722 ( 
.A1(n_618),
.A2(n_27),
.B1(n_24),
.B2(n_26),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_580),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_636),
.A2(n_430),
.B1(n_432),
.B2(n_427),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_580),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_633),
.A2(n_439),
.B1(n_443),
.B2(n_436),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_608),
.B(n_444),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_604),
.A2(n_450),
.B1(n_451),
.B2(n_445),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_580),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_590),
.Y(n_730)
);

OAI22xp33_ASAP7_75t_L g731 ( 
.A1(n_570),
.A2(n_461),
.B1(n_464),
.B2(n_452),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_SL g732 ( 
.A1(n_568),
.A2(n_468),
.B1(n_470),
.B2(n_467),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_590),
.Y(n_733)
);

OAI22xp33_ASAP7_75t_L g734 ( 
.A1(n_576),
.A2(n_472),
.B1(n_474),
.B2(n_471),
.Y(n_734)
);

XNOR2xp5_ASAP7_75t_L g735 ( 
.A(n_655),
.B(n_27),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_590),
.Y(n_736)
);

AO22x2_ASAP7_75t_L g737 ( 
.A1(n_632),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_589),
.Y(n_738)
);

BUFx10_ASAP7_75t_L g739 ( 
.A(n_612),
.Y(n_739)
);

OAI22xp33_ASAP7_75t_L g740 ( 
.A1(n_638),
.A2(n_477),
.B1(n_481),
.B2(n_475),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_593),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_621),
.B(n_482),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_621),
.B(n_484),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_656),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_599),
.Y(n_745)
);

AO22x2_ASAP7_75t_L g746 ( 
.A1(n_632),
.A2(n_652),
.B1(n_612),
.B2(n_624),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_624),
.B(n_485),
.Y(n_747)
);

AOI22xp5_ASAP7_75t_L g748 ( 
.A1(n_638),
.A2(n_488),
.B1(n_497),
.B2(n_486),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_650),
.A2(n_663),
.B1(n_657),
.B2(n_569),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_592),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_721),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_749),
.B(n_648),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_718),
.B(n_648),
.Y(n_753)
);

AND2x4_ASAP7_75t_L g754 ( 
.A(n_706),
.B(n_652),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_738),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_741),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_711),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_744),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_745),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_669),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_674),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_701),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_725),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_725),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_673),
.B(n_649),
.Y(n_765)
);

XOR2xp5_ASAP7_75t_L g766 ( 
.A(n_710),
.B(n_501),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_733),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_733),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_708),
.B(n_594),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_673),
.B(n_620),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_699),
.B(n_621),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_688),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_699),
.B(n_625),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_690),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_698),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_700),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_676),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_703),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_712),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_723),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_668),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_729),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_730),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_736),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_750),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_667),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_717),
.B(n_653),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_671),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_672),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_716),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_683),
.B(n_625),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_679),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_666),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_676),
.B(n_620),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_739),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_739),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_746),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_746),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_747),
.Y(n_799)
);

XOR2xp5_ASAP7_75t_L g800 ( 
.A(n_685),
.B(n_503),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_727),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_683),
.B(n_601),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_692),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_677),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_705),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_722),
.B(n_578),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_702),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_705),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_702),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_696),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_681),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_720),
.B(n_648),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_681),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_680),
.Y(n_814)
);

XNOR2xp5_ASAP7_75t_L g815 ( 
.A(n_685),
.B(n_584),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_670),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_693),
.Y(n_817)
);

XNOR2x1_ASAP7_75t_L g818 ( 
.A(n_735),
.B(n_596),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_686),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_724),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_678),
.B(n_625),
.Y(n_821)
);

XOR2xp5_ASAP7_75t_L g822 ( 
.A(n_704),
.B(n_504),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_687),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_707),
.B(n_625),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_724),
.B(n_588),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_689),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_691),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_726),
.B(n_641),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_691),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_709),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_707),
.B(n_609),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_709),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_684),
.B(n_626),
.Y(n_833)
);

INVxp67_ASAP7_75t_SL g834 ( 
.A(n_684),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_732),
.B(n_648),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_743),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_719),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_719),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_737),
.Y(n_839)
);

INVxp33_ASAP7_75t_L g840 ( 
.A(n_675),
.Y(n_840)
);

XNOR2x1_ASAP7_75t_L g841 ( 
.A(n_722),
.B(n_28),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_817),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_769),
.Y(n_843)
);

AND2x4_ASAP7_75t_SL g844 ( 
.A(n_777),
.B(n_726),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_769),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_785),
.Y(n_846)
);

OR2x2_ASAP7_75t_SL g847 ( 
.A(n_807),
.B(n_682),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_826),
.B(n_732),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_793),
.Y(n_849)
);

AND2x4_ASAP7_75t_SL g850 ( 
.A(n_777),
.B(n_748),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_785),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_751),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_755),
.Y(n_853)
);

AND2x2_ASAP7_75t_SL g854 ( 
.A(n_752),
.B(n_568),
.Y(n_854)
);

INVx6_ASAP7_75t_L g855 ( 
.A(n_785),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_797),
.B(n_694),
.Y(n_856)
);

OAI21xp5_ASAP7_75t_L g857 ( 
.A1(n_802),
.A2(n_753),
.B(n_831),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_786),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_802),
.A2(n_748),
.B(n_714),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_781),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_788),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_770),
.B(n_737),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_756),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_789),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_759),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_787),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_787),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_794),
.B(n_588),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_798),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_804),
.B(n_602),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_758),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_831),
.A2(n_714),
.B(n_740),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_790),
.B(n_713),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_757),
.B(n_602),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_778),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_820),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_757),
.B(n_627),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_792),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_760),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_825),
.B(n_627),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_761),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_772),
.Y(n_882)
);

NAND2x1p5_ASAP7_75t_L g883 ( 
.A(n_803),
.B(n_592),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_790),
.B(n_742),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_796),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_765),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_774),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_754),
.B(n_582),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_810),
.B(n_695),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_795),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_762),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_836),
.B(n_658),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_824),
.B(n_658),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_824),
.B(n_658),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_775),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_776),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_754),
.B(n_582),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_779),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_811),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_780),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_816),
.B(n_658),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_834),
.A2(n_697),
.B1(n_715),
.B2(n_728),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_819),
.B(n_659),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_782),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_783),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_784),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_763),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_764),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_834),
.A2(n_731),
.B1(n_734),
.B2(n_675),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_767),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_801),
.B(n_650),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_823),
.B(n_659),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_813),
.Y(n_913)
);

AND2x6_ASAP7_75t_L g914 ( 
.A(n_827),
.B(n_657),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_814),
.B(n_663),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_768),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_799),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_771),
.B(n_659),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_833),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_771),
.B(n_507),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_829),
.Y(n_921)
);

AND2x2_ASAP7_75t_SL g922 ( 
.A(n_812),
.B(n_637),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_828),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_833),
.Y(n_924)
);

BUFx4_ASAP7_75t_SL g925 ( 
.A(n_806),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_830),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_773),
.A2(n_642),
.B(n_515),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_832),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_773),
.A2(n_791),
.B(n_835),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_791),
.B(n_659),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_809),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_828),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_805),
.B(n_510),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_835),
.Y(n_934)
);

AND2x2_ASAP7_75t_SL g935 ( 
.A(n_821),
.B(n_630),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_821),
.B(n_630),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_808),
.B(n_516),
.Y(n_937)
);

AND2x2_ASAP7_75t_SL g938 ( 
.A(n_838),
.B(n_630),
.Y(n_938)
);

BUFx5_ASAP7_75t_L g939 ( 
.A(n_839),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_837),
.B(n_634),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_837),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_928),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_851),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_858),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_851),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_928),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_907),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_851),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_923),
.B(n_885),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_860),
.Y(n_950)
);

INVxp67_ASAP7_75t_L g951 ( 
.A(n_911),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_851),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_871),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_843),
.B(n_840),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_870),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_843),
.B(n_822),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_861),
.B(n_806),
.Y(n_957)
);

OR2x6_ASAP7_75t_L g958 ( 
.A(n_861),
.B(n_806),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_885),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_921),
.B(n_800),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_845),
.B(n_517),
.Y(n_961)
);

INVx4_ASAP7_75t_L g962 ( 
.A(n_855),
.Y(n_962)
);

INVx1_ASAP7_75t_SL g963 ( 
.A(n_842),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_858),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_845),
.B(n_520),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_941),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_907),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_849),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_932),
.B(n_79),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_849),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_864),
.Y(n_971)
);

BUFx2_ASAP7_75t_L g972 ( 
.A(n_842),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_866),
.B(n_82),
.Y(n_973)
);

BUFx3_ASAP7_75t_L g974 ( 
.A(n_871),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_890),
.B(n_841),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_856),
.B(n_815),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_867),
.B(n_85),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_919),
.B(n_521),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_919),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_864),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_941),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_921),
.B(n_766),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_924),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_924),
.B(n_522),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_857),
.B(n_523),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_880),
.B(n_818),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_899),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_934),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_874),
.B(n_634),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_922),
.B(n_524),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_926),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_879),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_922),
.B(n_527),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_847),
.B(n_634),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_855),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_917),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_931),
.B(n_852),
.Y(n_997)
);

INVx6_ASAP7_75t_L g998 ( 
.A(n_856),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_934),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_SL g1000 ( 
.A(n_876),
.B(n_528),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_908),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_854),
.B(n_534),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_877),
.B(n_539),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_899),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_854),
.B(n_544),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_SL g1006 ( 
.A(n_876),
.B(n_545),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_890),
.B(n_592),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_868),
.B(n_639),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_908),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_913),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_934),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_915),
.B(n_639),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_853),
.B(n_863),
.Y(n_1013)
);

AND2x6_ASAP7_75t_L g1014 ( 
.A(n_934),
.B(n_613),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_933),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_889),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_981),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_950),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_953),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_SL g1020 ( 
.A1(n_1002),
.A2(n_873),
.B1(n_935),
.B2(n_850),
.Y(n_1020)
);

INVx1_ASAP7_75t_SL g1021 ( 
.A(n_963),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_981),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1016),
.B(n_884),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_981),
.Y(n_1024)
);

INVx2_ASAP7_75t_SL g1025 ( 
.A(n_998),
.Y(n_1025)
);

BUFx4f_ASAP7_75t_L g1026 ( 
.A(n_1015),
.Y(n_1026)
);

INVx5_ASAP7_75t_L g1027 ( 
.A(n_945),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_996),
.B(n_865),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_972),
.Y(n_1029)
);

AOI22xp33_ASAP7_75t_L g1030 ( 
.A1(n_979),
.A2(n_872),
.B1(n_859),
.B2(n_929),
.Y(n_1030)
);

CKINVDCx14_ASAP7_75t_R g1031 ( 
.A(n_974),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_959),
.Y(n_1032)
);

BUFx8_ASAP7_75t_SL g1033 ( 
.A(n_976),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_945),
.Y(n_1034)
);

INVx6_ASAP7_75t_L g1035 ( 
.A(n_959),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_994),
.Y(n_1036)
);

BUFx4f_ASAP7_75t_L g1037 ( 
.A(n_988),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_959),
.Y(n_1038)
);

NAND2x1p5_ASAP7_75t_L g1039 ( 
.A(n_988),
.B(n_846),
.Y(n_1039)
);

BUFx6f_ASAP7_75t_L g1040 ( 
.A(n_945),
.Y(n_1040)
);

OR2x6_ASAP7_75t_L g1041 ( 
.A(n_957),
.B(n_869),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_979),
.Y(n_1042)
);

INVxp33_ASAP7_75t_L g1043 ( 
.A(n_956),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_987),
.Y(n_1044)
);

INVx5_ASAP7_75t_L g1045 ( 
.A(n_948),
.Y(n_1045)
);

BUFx6f_ASAP7_75t_L g1046 ( 
.A(n_948),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_983),
.Y(n_1047)
);

INVx8_ASAP7_75t_L g1048 ( 
.A(n_948),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_988),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_999),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_983),
.Y(n_1051)
);

INVx6_ASAP7_75t_L g1052 ( 
.A(n_962),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_999),
.Y(n_1053)
);

INVx1_ASAP7_75t_SL g1054 ( 
.A(n_1004),
.Y(n_1054)
);

BUFx5_ASAP7_75t_L g1055 ( 
.A(n_942),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_999),
.Y(n_1056)
);

BUFx4f_ASAP7_75t_L g1057 ( 
.A(n_1011),
.Y(n_1057)
);

AND2x2_ASAP7_75t_L g1058 ( 
.A(n_1012),
.B(n_873),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_947),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_951),
.B(n_862),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_1011),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_1011),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_966),
.Y(n_1063)
);

INVx4_ASAP7_75t_L g1064 ( 
.A(n_962),
.Y(n_1064)
);

CKINVDCx16_ASAP7_75t_R g1065 ( 
.A(n_1000),
.Y(n_1065)
);

BUFx3_ASAP7_75t_L g1066 ( 
.A(n_998),
.Y(n_1066)
);

BUFx12f_ASAP7_75t_L g1067 ( 
.A(n_957),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_1010),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_949),
.Y(n_1069)
);

BUFx6f_ASAP7_75t_L g1070 ( 
.A(n_943),
.Y(n_1070)
);

BUFx3_ASAP7_75t_L g1071 ( 
.A(n_949),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_947),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_975),
.Y(n_1073)
);

INVx3_ASAP7_75t_L g1074 ( 
.A(n_943),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_958),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_967),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_995),
.B(n_846),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_952),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_986),
.Y(n_1079)
);

INVx3_ASAP7_75t_SL g1080 ( 
.A(n_976),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_1044),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1059),
.Y(n_1082)
);

AOI22xp33_ASAP7_75t_SL g1083 ( 
.A1(n_1065),
.A2(n_960),
.B1(n_1006),
.B2(n_850),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_1058),
.B(n_954),
.Y(n_1084)
);

CKINVDCx20_ASAP7_75t_R g1085 ( 
.A(n_1031),
.Y(n_1085)
);

CKINVDCx14_ASAP7_75t_R g1086 ( 
.A(n_1031),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_1054),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1020),
.A2(n_982),
.B1(n_909),
.B2(n_1005),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1059),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1020),
.A2(n_935),
.B1(n_914),
.B2(n_902),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1030),
.A2(n_991),
.B1(n_848),
.B2(n_889),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_1040),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1030),
.A2(n_914),
.B1(n_920),
.B2(n_1013),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1063),
.Y(n_1094)
);

AOI22xp33_ASAP7_75t_L g1095 ( 
.A1(n_1043),
.A2(n_914),
.B1(n_920),
.B2(n_1013),
.Y(n_1095)
);

CKINVDCx20_ASAP7_75t_R g1096 ( 
.A(n_1018),
.Y(n_1096)
);

INVx6_ASAP7_75t_L g1097 ( 
.A(n_1035),
.Y(n_1097)
);

BUFx4_ASAP7_75t_R g1098 ( 
.A(n_1033),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1042),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_SL g1100 ( 
.A1(n_1079),
.A2(n_844),
.B1(n_886),
.B2(n_990),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1072),
.Y(n_1101)
);

CKINVDCx11_ASAP7_75t_R g1102 ( 
.A(n_1029),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1043),
.A2(n_914),
.B1(n_888),
.B2(n_897),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1042),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_1018),
.Y(n_1105)
);

OAI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1036),
.A2(n_955),
.B1(n_993),
.B2(n_958),
.Y(n_1106)
);

INVx6_ASAP7_75t_L g1107 ( 
.A(n_1035),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_1060),
.A2(n_914),
.B1(n_888),
.B2(n_897),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1047),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1029),
.Y(n_1110)
);

CKINVDCx11_ASAP7_75t_R g1111 ( 
.A(n_1080),
.Y(n_1111)
);

BUFx10_ASAP7_75t_L g1112 ( 
.A(n_1028),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_1028),
.A2(n_844),
.B1(n_969),
.B2(n_973),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1047),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1040),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_1072),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1076),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1051),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1023),
.A2(n_942),
.B1(n_946),
.B2(n_969),
.Y(n_1119)
);

BUFx3_ASAP7_75t_L g1120 ( 
.A(n_1019),
.Y(n_1120)
);

AOI22xp33_ASAP7_75t_L g1121 ( 
.A1(n_1041),
.A2(n_977),
.B1(n_973),
.B2(n_985),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1041),
.A2(n_977),
.B1(n_927),
.B2(n_997),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_1021),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1051),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1076),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1079),
.A2(n_1008),
.B1(n_1003),
.B2(n_997),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_1041),
.A2(n_989),
.B1(n_992),
.B2(n_944),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1037),
.A2(n_946),
.B1(n_938),
.B2(n_913),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1069),
.B(n_961),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1073),
.B(n_1068),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1062),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_1040),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_1071),
.B(n_938),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_1037),
.A2(n_964),
.B1(n_940),
.B2(n_967),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1062),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1071),
.A2(n_970),
.B1(n_971),
.B2(n_968),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1032),
.B(n_965),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1057),
.A2(n_1001),
.B1(n_1009),
.B2(n_936),
.Y(n_1138)
);

CKINVDCx11_ASAP7_75t_R g1139 ( 
.A(n_1080),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1055),
.Y(n_1140)
);

INVx6_ASAP7_75t_L g1141 ( 
.A(n_1035),
.Y(n_1141)
);

INVx1_ASAP7_75t_SL g1142 ( 
.A(n_1019),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1088),
.A2(n_1075),
.B1(n_1067),
.B2(n_937),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1090),
.A2(n_937),
.B(n_933),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1083),
.A2(n_984),
.B(n_978),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1100),
.A2(n_1075),
.B1(n_879),
.B2(n_891),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_SL g1147 ( 
.A1(n_1096),
.A2(n_1025),
.B1(n_1066),
.B2(n_1038),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1091),
.A2(n_881),
.B1(n_891),
.B2(n_878),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1091),
.A2(n_881),
.B1(n_980),
.B2(n_898),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1094),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1092),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_SL g1152 ( 
.A1(n_1126),
.A2(n_894),
.B(n_893),
.Y(n_1152)
);

AOI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1108),
.A2(n_887),
.B1(n_904),
.B2(n_900),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1099),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1103),
.A2(n_905),
.B1(n_895),
.B2(n_896),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_SL g1156 ( 
.A1(n_1142),
.A2(n_1026),
.B1(n_1057),
.B2(n_1066),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1106),
.A2(n_1093),
.B1(n_1095),
.B2(n_1084),
.Y(n_1157)
);

NOR2x1_ASAP7_75t_L g1158 ( 
.A(n_1105),
.B(n_1064),
.Y(n_1158)
);

AOI222xp33_ASAP7_75t_L g1159 ( 
.A1(n_1142),
.A2(n_1026),
.B1(n_869),
.B2(n_1001),
.C1(n_1009),
.C2(n_916),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1082),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1092),
.Y(n_1161)
);

BUFx12f_ASAP7_75t_L g1162 ( 
.A(n_1102),
.Y(n_1162)
);

NAND2xp33_ASAP7_75t_SL g1163 ( 
.A(n_1085),
.B(n_1064),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1121),
.A2(n_895),
.B1(n_906),
.B2(n_896),
.Y(n_1164)
);

AOI222xp33_ASAP7_75t_L g1165 ( 
.A1(n_1087),
.A2(n_910),
.B1(n_550),
.B2(n_552),
.C1(n_553),
.C2(n_556),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_1123),
.A2(n_906),
.B1(n_930),
.B2(n_918),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1122),
.A2(n_882),
.B1(n_1033),
.B2(n_903),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1113),
.A2(n_1052),
.B1(n_1038),
.B2(n_1032),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_SL g1169 ( 
.A1(n_1086),
.A2(n_1120),
.B1(n_1128),
.B2(n_1133),
.Y(n_1169)
);

AOI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_1129),
.A2(n_901),
.B1(n_912),
.B2(n_892),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1127),
.A2(n_1052),
.B1(n_1022),
.B2(n_1024),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1092),
.Y(n_1172)
);

INVx5_ASAP7_75t_SL g1173 ( 
.A(n_1115),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_1115),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1137),
.A2(n_882),
.B1(n_1017),
.B2(n_875),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_1119),
.A2(n_875),
.B1(n_1014),
.B2(n_1055),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_1119),
.A2(n_1052),
.B1(n_1007),
.B2(n_883),
.Y(n_1177)
);

OAI22xp5_ASAP7_75t_L g1178 ( 
.A1(n_1081),
.A2(n_883),
.B1(n_1034),
.B2(n_1027),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1130),
.B(n_939),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1081),
.B(n_939),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1104),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1128),
.A2(n_1027),
.B1(n_1045),
.B2(n_1034),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1136),
.A2(n_1027),
.B1(n_1045),
.B2(n_1034),
.Y(n_1183)
);

OAI222xp33_ASAP7_75t_L g1184 ( 
.A1(n_1134),
.A2(n_1131),
.B1(n_1135),
.B2(n_1138),
.C1(n_1114),
.C2(n_1118),
.Y(n_1184)
);

AOI22xp33_ASAP7_75t_L g1185 ( 
.A1(n_1111),
.A2(n_1014),
.B1(n_1055),
.B2(n_1050),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1089),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1109),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1112),
.B(n_1101),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_L g1189 ( 
.A(n_1097),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1112),
.B(n_1050),
.Y(n_1190)
);

AOI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_1139),
.A2(n_1014),
.B1(n_1055),
.B2(n_1056),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1110),
.A2(n_1014),
.B1(n_1055),
.B2(n_1056),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1115),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1116),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1134),
.A2(n_1055),
.B1(n_939),
.B2(n_1074),
.Y(n_1195)
);

BUFx12f_ASAP7_75t_L g1196 ( 
.A(n_1097),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1138),
.A2(n_939),
.B1(n_1078),
.B2(n_1074),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1117),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1124),
.A2(n_939),
.B1(n_1078),
.B2(n_1070),
.Y(n_1199)
);

BUFx8_ASAP7_75t_L g1200 ( 
.A(n_1098),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1125),
.Y(n_1201)
);

BUFx12f_ASAP7_75t_L g1202 ( 
.A(n_1097),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1107),
.A2(n_939),
.B1(n_1070),
.B2(n_1053),
.Y(n_1203)
);

CKINVDCx11_ASAP7_75t_R g1204 ( 
.A(n_1132),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1132),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1107),
.A2(n_925),
.B1(n_1034),
.B2(n_1027),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1132),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1140),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_L g1209 ( 
.A(n_1107),
.B(n_660),
.C(n_639),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1141),
.A2(n_1070),
.B1(n_1053),
.B2(n_1061),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1141),
.A2(n_925),
.B1(n_1045),
.B2(n_1049),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1141),
.A2(n_1045),
.B(n_1077),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1082),
.Y(n_1213)
);

OAI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1088),
.A2(n_1077),
.B1(n_1039),
.B2(n_995),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1088),
.A2(n_1039),
.B1(n_1061),
.B2(n_1049),
.Y(n_1215)
);

NAND3xp33_ASAP7_75t_L g1216 ( 
.A(n_1088),
.B(n_664),
.C(n_660),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1088),
.A2(n_1070),
.B1(n_1049),
.B2(n_1061),
.Y(n_1217)
);

INVx5_ASAP7_75t_SL g1218 ( 
.A(n_1092),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1094),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1157),
.B(n_1049),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1169),
.A2(n_559),
.B1(n_562),
.B2(n_546),
.Y(n_1221)
);

HB1xp67_ASAP7_75t_L g1222 ( 
.A(n_1150),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1143),
.A2(n_564),
.B1(n_563),
.B2(n_1061),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1154),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_SL g1225 ( 
.A1(n_1216),
.A2(n_1048),
.B1(n_1046),
.B2(n_1040),
.Y(n_1225)
);

AOI222xp33_ASAP7_75t_L g1226 ( 
.A1(n_1144),
.A2(n_660),
.B1(n_664),
.B2(n_645),
.C1(n_33),
.C2(n_34),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1144),
.A2(n_855),
.B1(n_1048),
.B2(n_664),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1146),
.A2(n_952),
.B1(n_1046),
.B2(n_1048),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1167),
.A2(n_1046),
.B1(n_645),
.B2(n_615),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1165),
.A2(n_1046),
.B1(n_645),
.B2(n_615),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1156),
.A2(n_1211),
.B1(n_1217),
.B2(n_1206),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1216),
.A2(n_645),
.B1(n_615),
.B2(n_616),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_SL g1233 ( 
.A1(n_1182),
.A2(n_616),
.B1(n_617),
.B2(n_613),
.Y(n_1233)
);

OAI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1185),
.A2(n_616),
.B1(n_617),
.B2(n_613),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1181),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1166),
.A2(n_617),
.B1(n_597),
.B2(n_603),
.Y(n_1236)
);

OAI222xp33_ASAP7_75t_L g1237 ( 
.A1(n_1191),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.C1(n_34),
.C2(n_35),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1145),
.B(n_31),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1145),
.B(n_32),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1159),
.A2(n_597),
.B1(n_603),
.B2(n_595),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1159),
.B(n_35),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1163),
.A2(n_597),
.B1(n_603),
.B2(n_595),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1158),
.A2(n_597),
.B1(n_603),
.B2(n_595),
.Y(n_1243)
);

OAI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1170),
.A2(n_595),
.B1(n_38),
.B2(n_36),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1160),
.B(n_36),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1153),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1164),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1186),
.B(n_41),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1147),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1187),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1152),
.B(n_42),
.C(n_43),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1194),
.B(n_44),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1201),
.B(n_47),
.Y(n_1253)
);

OAI222xp33_ASAP7_75t_L g1254 ( 
.A1(n_1215),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.C1(n_50),
.C2(n_51),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1192),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1214),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1148),
.A2(n_52),
.B1(n_53),
.B2(n_55),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1175),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1155),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1177),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1219),
.B(n_61),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1198),
.Y(n_1262)
);

AO21x1_ASAP7_75t_SL g1263 ( 
.A1(n_1184),
.A2(n_63),
.B(n_64),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1189),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1168),
.A2(n_1188),
.B1(n_1149),
.B2(n_1171),
.Y(n_1265)
);

OAI221xp5_ASAP7_75t_L g1266 ( 
.A1(n_1152),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1213),
.B(n_66),
.Y(n_1267)
);

OAI211xp5_ASAP7_75t_L g1268 ( 
.A1(n_1180),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1179),
.B(n_69),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1208),
.B(n_70),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1200),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1162),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1190),
.B(n_74),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1197),
.A2(n_74),
.B1(n_75),
.B2(n_77),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1200),
.A2(n_75),
.B1(n_78),
.B2(n_86),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1195),
.A2(n_78),
.B1(n_87),
.B2(n_89),
.Y(n_1276)
);

OAI222xp33_ASAP7_75t_L g1277 ( 
.A1(n_1178),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.C1(n_95),
.C2(n_96),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1212),
.B(n_102),
.C(n_106),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1176),
.A2(n_107),
.B1(n_110),
.B2(n_112),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1209),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1183),
.A2(n_114),
.B1(n_115),
.B2(n_122),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1207),
.B(n_1205),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1196),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1202),
.A2(n_128),
.B1(n_132),
.B2(n_134),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1204),
.A2(n_135),
.B1(n_136),
.B2(n_137),
.Y(n_1285)
);

OAI222xp33_ASAP7_75t_L g1286 ( 
.A1(n_1199),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.C1(n_144),
.C2(n_145),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1222),
.B(n_1151),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_SL g1288 ( 
.A(n_1226),
.B(n_1209),
.Y(n_1288)
);

NOR3xp33_ASAP7_75t_L g1289 ( 
.A(n_1266),
.B(n_1172),
.C(n_1151),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1251),
.A2(n_1189),
.B1(n_1210),
.B2(n_1203),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1224),
.Y(n_1291)
);

NAND2xp33_ASAP7_75t_L g1292 ( 
.A(n_1238),
.B(n_1161),
.Y(n_1292)
);

NAND3xp33_ASAP7_75t_L g1293 ( 
.A(n_1239),
.B(n_1174),
.C(n_1161),
.Y(n_1293)
);

OA21x2_ASAP7_75t_L g1294 ( 
.A1(n_1280),
.A2(n_1227),
.B(n_1224),
.Y(n_1294)
);

OAI22xp5_ASAP7_75t_L g1295 ( 
.A1(n_1249),
.A2(n_1218),
.B1(n_1173),
.B2(n_1193),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1262),
.B(n_1172),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1262),
.B(n_1193),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1271),
.A2(n_1174),
.B(n_1161),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1250),
.B(n_1174),
.Y(n_1299)
);

OAI221xp5_ASAP7_75t_SL g1300 ( 
.A1(n_1272),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.C(n_154),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1250),
.B(n_1173),
.Y(n_1301)
);

NOR2xp33_ASAP7_75t_L g1302 ( 
.A(n_1269),
.B(n_1173),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1235),
.B(n_1218),
.Y(n_1303)
);

OAI221xp5_ASAP7_75t_L g1304 ( 
.A1(n_1275),
.A2(n_156),
.B1(n_157),
.B2(n_160),
.C(n_163),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1235),
.B(n_1218),
.Y(n_1305)
);

AOI211xp5_ASAP7_75t_L g1306 ( 
.A1(n_1244),
.A2(n_164),
.B(n_166),
.C(n_169),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1253),
.B(n_172),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1261),
.B(n_1270),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1253),
.B(n_1261),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1241),
.B(n_173),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1265),
.B(n_175),
.Y(n_1311)
);

NAND3xp33_ASAP7_75t_L g1312 ( 
.A(n_1268),
.B(n_176),
.C(n_178),
.Y(n_1312)
);

NAND3xp33_ASAP7_75t_L g1313 ( 
.A(n_1256),
.B(n_185),
.C(n_186),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1260),
.A2(n_1246),
.B1(n_1257),
.B2(n_1247),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1270),
.B(n_187),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1220),
.B(n_188),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1282),
.B(n_1245),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1254),
.A2(n_189),
.B(n_190),
.Y(n_1318)
);

OAI21xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1237),
.A2(n_193),
.B(n_194),
.Y(n_1319)
);

OAI221xp5_ASAP7_75t_SL g1320 ( 
.A1(n_1221),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1273),
.B(n_200),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1264),
.B(n_375),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1248),
.B(n_202),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1231),
.A2(n_372),
.B1(n_204),
.B2(n_205),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1252),
.B(n_203),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1280),
.Y(n_1326)
);

AND2x2_ASAP7_75t_SL g1327 ( 
.A(n_1240),
.B(n_207),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1229),
.A2(n_209),
.B(n_211),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1267),
.B(n_1264),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1230),
.B(n_212),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1263),
.B(n_371),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1274),
.B(n_213),
.Y(n_1332)
);

NAND4xp25_ASAP7_75t_L g1333 ( 
.A(n_1259),
.B(n_218),
.C(n_220),
.D(n_221),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1255),
.B(n_229),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1225),
.B(n_232),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1258),
.B(n_233),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1263),
.B(n_370),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1223),
.B(n_236),
.Y(n_1338)
);

OA211x2_ASAP7_75t_L g1339 ( 
.A1(n_1278),
.A2(n_238),
.B(n_239),
.C(n_240),
.Y(n_1339)
);

OAI211xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1276),
.A2(n_1281),
.B(n_1285),
.C(n_1284),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1279),
.B(n_242),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1308),
.B(n_1309),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1288),
.A2(n_1311),
.B1(n_1314),
.B2(n_1327),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1326),
.B(n_1234),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1326),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1288),
.A2(n_1277),
.B(n_1242),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1317),
.B(n_1236),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1291),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1287),
.B(n_1232),
.Y(n_1349)
);

NAND4xp25_ASAP7_75t_L g1350 ( 
.A(n_1293),
.B(n_1283),
.C(n_1233),
.D(n_1228),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1296),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1329),
.B(n_1243),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1301),
.B(n_243),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1297),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1311),
.A2(n_1286),
.B1(n_245),
.B2(n_247),
.Y(n_1355)
);

NAND3xp33_ASAP7_75t_L g1356 ( 
.A(n_1306),
.B(n_244),
.C(n_248),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1292),
.B(n_249),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1294),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1305),
.B(n_251),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_L g1360 ( 
.A(n_1292),
.B(n_252),
.Y(n_1360)
);

NOR2x1_ASAP7_75t_L g1361 ( 
.A(n_1299),
.B(n_253),
.Y(n_1361)
);

NAND3xp33_ASAP7_75t_L g1362 ( 
.A(n_1312),
.B(n_254),
.C(n_255),
.Y(n_1362)
);

NOR2x1_ASAP7_75t_L g1363 ( 
.A(n_1303),
.B(n_256),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1302),
.B(n_257),
.Y(n_1364)
);

NOR2x1_ASAP7_75t_L g1365 ( 
.A(n_1302),
.B(n_261),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1294),
.B(n_263),
.Y(n_1366)
);

NOR3xp33_ASAP7_75t_L g1367 ( 
.A(n_1318),
.B(n_264),
.C(n_267),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1294),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1321),
.B(n_268),
.Y(n_1369)
);

NAND2x1_ASAP7_75t_L g1370 ( 
.A(n_1289),
.B(n_269),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1289),
.Y(n_1371)
);

AND2x4_ASAP7_75t_L g1372 ( 
.A(n_1322),
.B(n_270),
.Y(n_1372)
);

NAND4xp25_ASAP7_75t_L g1373 ( 
.A(n_1310),
.B(n_271),
.C(n_273),
.D(n_276),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1331),
.B(n_278),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1316),
.B(n_280),
.Y(n_1375)
);

AOI221xp5_ASAP7_75t_L g1376 ( 
.A1(n_1319),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.C(n_286),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1314),
.A2(n_289),
.B1(n_290),
.B2(n_291),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1315),
.Y(n_1378)
);

NOR4xp25_ASAP7_75t_L g1379 ( 
.A(n_1343),
.B(n_1298),
.C(n_1300),
.D(n_1320),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1348),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1342),
.B(n_1351),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1345),
.B(n_1307),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1345),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1354),
.Y(n_1384)
);

XNOR2x2_ASAP7_75t_L g1385 ( 
.A(n_1371),
.B(n_1333),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1358),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1358),
.B(n_1337),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1368),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1366),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1378),
.B(n_1323),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1344),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1364),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1349),
.Y(n_1393)
);

NOR4xp25_ASAP7_75t_L g1394 ( 
.A(n_1343),
.B(n_1340),
.C(n_1304),
.D(n_1295),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1352),
.B(n_1325),
.Y(n_1395)
);

XNOR2xp5_ASAP7_75t_L g1396 ( 
.A(n_1365),
.B(n_1324),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1347),
.Y(n_1397)
);

NAND4xp75_ASAP7_75t_L g1398 ( 
.A(n_1376),
.B(n_1339),
.C(n_1327),
.D(n_1335),
.Y(n_1398)
);

NAND4xp75_ASAP7_75t_L g1399 ( 
.A(n_1363),
.B(n_1334),
.C(n_1341),
.D(n_1338),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1393),
.B(n_1353),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1393),
.B(n_1346),
.Y(n_1401)
);

AOI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1398),
.A2(n_1367),
.B1(n_1346),
.B2(n_1356),
.Y(n_1402)
);

CKINVDCx16_ASAP7_75t_R g1403 ( 
.A(n_1392),
.Y(n_1403)
);

INVxp67_ASAP7_75t_L g1404 ( 
.A(n_1397),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_SL g1405 ( 
.A(n_1399),
.B(n_1367),
.Y(n_1405)
);

INVxp67_ASAP7_75t_L g1406 ( 
.A(n_1391),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1380),
.Y(n_1407)
);

XNOR2xp5_ASAP7_75t_L g1408 ( 
.A(n_1396),
.B(n_1359),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_L g1409 ( 
.A(n_1395),
.B(n_1370),
.Y(n_1409)
);

XOR2x2_ASAP7_75t_L g1410 ( 
.A(n_1385),
.B(n_1377),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1384),
.B(n_1357),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1388),
.Y(n_1412)
);

XOR2x2_ASAP7_75t_L g1413 ( 
.A(n_1385),
.B(n_1396),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1388),
.Y(n_1414)
);

OA22x2_ASAP7_75t_L g1415 ( 
.A1(n_1402),
.A2(n_1387),
.B1(n_1391),
.B2(n_1389),
.Y(n_1415)
);

OA22x2_ASAP7_75t_L g1416 ( 
.A1(n_1413),
.A2(n_1387),
.B1(n_1381),
.B2(n_1374),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1412),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1406),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1414),
.Y(n_1419)
);

OAI22x1_ASAP7_75t_L g1420 ( 
.A1(n_1408),
.A2(n_1383),
.B1(n_1390),
.B2(n_1382),
.Y(n_1420)
);

XOR2x2_ASAP7_75t_L g1421 ( 
.A(n_1410),
.B(n_1390),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1407),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_SL g1423 ( 
.A1(n_1405),
.A2(n_1357),
.B1(n_1360),
.B2(n_1379),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1403),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1400),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1401),
.Y(n_1426)
);

OA22x2_ASAP7_75t_L g1427 ( 
.A1(n_1404),
.A2(n_1394),
.B1(n_1386),
.B2(n_1383),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1411),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1405),
.A2(n_1377),
.B1(n_1355),
.B2(n_1373),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1411),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1422),
.Y(n_1431)
);

BUFx2_ASAP7_75t_L g1432 ( 
.A(n_1424),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1418),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1425),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1423),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1427),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1428),
.Y(n_1437)
);

HB1xp67_ASAP7_75t_L g1438 ( 
.A(n_1420),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1417),
.Y(n_1439)
);

AO22x1_ASAP7_75t_L g1440 ( 
.A1(n_1435),
.A2(n_1423),
.B1(n_1427),
.B2(n_1421),
.Y(n_1440)
);

AO22x2_ASAP7_75t_L g1441 ( 
.A1(n_1436),
.A2(n_1433),
.B1(n_1434),
.B2(n_1431),
.Y(n_1441)
);

OA22x2_ASAP7_75t_L g1442 ( 
.A1(n_1438),
.A2(n_1429),
.B1(n_1430),
.B2(n_1426),
.Y(n_1442)
);

OAI22x1_ASAP7_75t_L g1443 ( 
.A1(n_1432),
.A2(n_1429),
.B1(n_1409),
.B2(n_1430),
.Y(n_1443)
);

NAND4xp25_ASAP7_75t_SL g1444 ( 
.A(n_1433),
.B(n_1415),
.C(n_1355),
.D(n_1416),
.Y(n_1444)
);

AOI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1436),
.A2(n_1415),
.B1(n_1419),
.B2(n_1360),
.Y(n_1445)
);

OA22x2_ASAP7_75t_L g1446 ( 
.A1(n_1445),
.A2(n_1432),
.B1(n_1434),
.B2(n_1437),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1441),
.Y(n_1447)
);

A2O1A1Ixp33_ASAP7_75t_SL g1448 ( 
.A1(n_1444),
.A2(n_1439),
.B(n_1375),
.C(n_1369),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1442),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_SL g1450 ( 
.A1(n_1440),
.A2(n_1382),
.B(n_1290),
.C(n_1362),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1443),
.Y(n_1451)
);

AOI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1449),
.A2(n_1372),
.B1(n_1350),
.B2(n_1361),
.Y(n_1452)
);

INVxp67_ASAP7_75t_SL g1453 ( 
.A(n_1447),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1446),
.A2(n_1372),
.B1(n_1313),
.B2(n_1381),
.Y(n_1454)
);

NOR2x1_ASAP7_75t_L g1455 ( 
.A(n_1451),
.B(n_1336),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1450),
.A2(n_1332),
.B1(n_1330),
.B2(n_1328),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1448),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1447),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1453),
.B(n_292),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1458),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1455),
.Y(n_1461)
);

NOR2x1_ASAP7_75t_L g1462 ( 
.A(n_1457),
.B(n_294),
.Y(n_1462)
);

INVxp67_ASAP7_75t_SL g1463 ( 
.A(n_1454),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1452),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_SL g1465 ( 
.A1(n_1460),
.A2(n_1456),
.B(n_298),
.C(n_300),
.Y(n_1465)
);

AND4x1_ASAP7_75t_L g1466 ( 
.A(n_1462),
.B(n_296),
.C(n_304),
.D(n_308),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1459),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1463),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_1468)
);

OAI22xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1463),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1467),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1466),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1469),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1468),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1465),
.A2(n_1464),
.B1(n_1461),
.B2(n_325),
.Y(n_1474)
);

HB1xp67_ASAP7_75t_L g1475 ( 
.A(n_1471),
.Y(n_1475)
);

HB1xp67_ASAP7_75t_L g1476 ( 
.A(n_1472),
.Y(n_1476)
);

CKINVDCx16_ASAP7_75t_R g1477 ( 
.A(n_1473),
.Y(n_1477)
);

AOI31xp33_ASAP7_75t_L g1478 ( 
.A1(n_1470),
.A2(n_315),
.A3(n_316),
.B(n_328),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1474),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1477),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1475),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1476),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1479),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1478),
.Y(n_1484)
);

AOI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1480),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1481),
.A2(n_335),
.B1(n_336),
.B2(n_338),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1482),
.A2(n_339),
.B1(n_342),
.B2(n_345),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1486),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1485),
.Y(n_1489)
);

AOI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1489),
.A2(n_1483),
.B1(n_1484),
.B2(n_1487),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1488),
.A2(n_346),
.B1(n_348),
.B2(n_352),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1490),
.Y(n_1492)
);

AOI221xp5_ASAP7_75t_L g1493 ( 
.A1(n_1492),
.A2(n_1491),
.B1(n_358),
.B2(n_360),
.C(n_362),
.Y(n_1493)
);

AOI211xp5_ASAP7_75t_L g1494 ( 
.A1(n_1493),
.A2(n_354),
.B(n_363),
.C(n_364),
.Y(n_1494)
);


endmodule