module fake_jpeg_21891_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_1),
.Y(n_41)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_36),
.B1(n_22),
.B2(n_14),
.Y(n_40)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_37),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g38 ( 
.A1(n_32),
.A2(n_26),
.B1(n_25),
.B2(n_17),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_25),
.B1(n_17),
.B2(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_44),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_13),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_19),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_53),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_23),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_52),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_31),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_54),
.A2(n_35),
.B1(n_34),
.B2(n_45),
.Y(n_77)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_60),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_58),
.B(n_15),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_33),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_38),
.Y(n_69)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_48),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_78),
.B(n_47),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_37),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_43),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_63),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_58),
.C(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_77),
.A2(n_36),
.B1(n_28),
.B2(n_43),
.Y(n_90)
);

HAxp5_ASAP7_75t_SL g78 ( 
.A(n_59),
.B(n_48),
.CON(n_78),
.SN(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_64),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_80),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_59),
.C(n_60),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_65),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_53),
.C(n_51),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_85),
.B(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_90),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_47),
.B1(n_28),
.B2(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_105),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_96),
.A2(n_103),
.B(n_84),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_75),
.B(n_66),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_78),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_73),
.Y(n_102)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_85),
.B(n_66),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

AOI321xp33_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_114),
.A3(n_101),
.B1(n_24),
.B2(n_23),
.C(n_13),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_103),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_83),
.C(n_67),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_112),
.C(n_55),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_67),
.C(n_68),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_115),
.A2(n_101),
.B1(n_104),
.B2(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_117),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_122),
.C(n_111),
.Y(n_123)
);

NOR3xp33_ASAP7_75t_SL g120 ( 
.A(n_114),
.B(n_15),
.C(n_24),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_21),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_123),
.B(n_125),
.C(n_126),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_112),
.C(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_55),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_62),
.C(n_49),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_121),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_128),
.A2(n_9),
.B1(n_6),
.B2(n_8),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_129),
.B(n_131),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_124),
.A2(n_120),
.B1(n_30),
.B2(n_3),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_1),
.A3(n_2),
.B1(n_11),
.B2(n_30),
.C1(n_129),
.C2(n_124),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.C(n_2),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.C(n_30),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_133),
.Y(n_137)
);


endmodule