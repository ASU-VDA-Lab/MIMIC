module fake_aes_11800_n_342 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_342);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_342;
wire n_117;
wire n_185;
wire n_284;
wire n_278;
wire n_114;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_252;
wire n_152;
wire n_113;
wire n_206;
wire n_288;
wire n_296;
wire n_157;
wire n_202;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_163;
wire n_105;
wire n_227;
wire n_231;
wire n_298;
wire n_144;
wire n_183;
wire n_199;
wire n_100;
wire n_305;
wire n_228;
wire n_236;
wire n_340;
wire n_150;
wire n_301;
wire n_222;
wire n_234;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_119;
wire n_167;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_247;
wire n_304;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_243;
wire n_235;
wire n_331;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_153;
wire n_259;
wire n_308;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_107;
wire n_254;
wire n_262;
wire n_239;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_217;
wire n_139;
wire n_193;
wire n_273;
wire n_120;
wire n_245;
wire n_260;
wire n_201;
wire n_197;
wire n_317;
wire n_111;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_179;
wire n_315;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_136;
wire n_283;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_168;
wire n_134;
wire n_233;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_225;
wire n_220;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_103;
wire n_180;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_188;
wire n_127;
wire n_291;
wire n_170;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_138;
wire n_323;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_226;
wire n_159;
wire n_337;
wire n_176;
wire n_123;
wire n_223;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_164;
wire n_175;
wire n_145;
wire n_290;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_151;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g98 ( .A(n_43), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_82), .Y(n_99) );
INVx2_ASAP7_75t_SL g100 ( .A(n_84), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_96), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_77), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_42), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_58), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_85), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_47), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_31), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_87), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_45), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_94), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_95), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_75), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_56), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_6), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_34), .B(n_2), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_79), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_59), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_6), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_27), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_46), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_37), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_93), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_65), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_91), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_54), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_32), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_19), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_51), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_73), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_22), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_33), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_25), .Y(n_132) );
CKINVDCx14_ASAP7_75t_R g133 ( .A(n_78), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_29), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_26), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_57), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_90), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_36), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_88), .Y(n_139) );
INVxp33_ASAP7_75t_L g140 ( .A(n_81), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_66), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_61), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_62), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_70), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_80), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_60), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_23), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_11), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_44), .Y(n_149) );
BUFx5_ASAP7_75t_L g150 ( .A(n_64), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_48), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_40), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_49), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_53), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_89), .Y(n_155) );
INVxp67_ASAP7_75t_SL g156 ( .A(n_52), .Y(n_156) );
AND2x6_ASAP7_75t_L g157 ( .A(n_99), .B(n_17), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_107), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_109), .Y(n_159) );
AND2x6_ASAP7_75t_L g160 ( .A(n_101), .B(n_18), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_150), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_150), .Y(n_162) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_111), .B(n_97), .Y(n_163) );
BUFx8_ASAP7_75t_L g164 ( .A(n_100), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_98), .B(n_0), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_114), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_150), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_150), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_118), .B(n_1), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_110), .Y(n_171) );
AND2x6_ASAP7_75t_L g172 ( .A(n_169), .B(n_102), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_161), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_162), .Y(n_174) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_167), .B(n_150), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_168), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_158), .B(n_140), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_169), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_170), .B(n_126), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_166), .Y(n_180) );
INVx6_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_159), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_171), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_173), .B(n_163), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_174), .B(n_163), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_180), .B(n_165), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_176), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_184), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_178), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_182), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_175), .A2(n_160), .B(n_157), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_182), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_181), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_172), .B(n_157), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_172), .B(n_148), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_175), .B(n_103), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_179), .Y(n_198) );
NAND2xp33_ASAP7_75t_L g199 ( .A(n_183), .B(n_115), .Y(n_199) );
INVxp67_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_177), .B(n_133), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_192), .A2(n_156), .B(n_105), .Y(n_203) );
NOR2xp33_ASAP7_75t_R g204 ( .A(n_194), .B(n_153), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_200), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_195), .Y(n_206) );
CKINVDCx10_ASAP7_75t_R g207 ( .A(n_199), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_185), .A2(n_117), .B(n_116), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_190), .B(n_120), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_196), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_186), .A2(n_124), .B(n_121), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_187), .A2(n_127), .B(n_125), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_198), .A2(n_129), .B(n_128), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_202), .B(n_104), .Y(n_214) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_188), .A2(n_201), .B(n_197), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_201), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_SL g217 ( .A1(n_189), .A2(n_131), .B(n_132), .C(n_130), .Y(n_217) );
AO31x2_ASAP7_75t_L g218 ( .A1(n_211), .A2(n_134), .A3(n_136), .B(n_135), .Y(n_218) );
NOR2xp33_ASAP7_75t_R g219 ( .A(n_207), .B(n_106), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_204), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_215), .Y(n_221) );
AO31x2_ASAP7_75t_L g222 ( .A1(n_203), .A2(n_139), .A3(n_142), .B(n_141), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_216), .Y(n_223) );
NOR2xp67_ASAP7_75t_L g224 ( .A(n_205), .B(n_3), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_209), .Y(n_225) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_208), .A2(n_193), .B(n_191), .Y(n_226) );
O2A1O1Ixp5_ASAP7_75t_L g227 ( .A1(n_208), .A2(n_193), .B(n_146), .C(n_149), .Y(n_227) );
AO31x2_ASAP7_75t_L g228 ( .A1(n_213), .A2(n_147), .A3(n_152), .B(n_151), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_212), .A2(n_155), .B(n_154), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g230 ( .A1(n_210), .A2(n_112), .B1(n_113), .B2(n_108), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_214), .A2(n_122), .B(n_119), .Y(n_231) );
NOR2x1_ASAP7_75t_SL g232 ( .A(n_206), .B(n_123), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g233 ( .A1(n_217), .A2(n_5), .B(n_3), .C(n_4), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_225), .B(n_4), .Y(n_234) );
OAI21x1_ASAP7_75t_L g235 ( .A1(n_221), .A2(n_144), .B(n_159), .Y(n_235) );
OA21x2_ASAP7_75t_L g236 ( .A1(n_226), .A2(n_138), .B(n_137), .Y(n_236) );
NAND3xp33_ASAP7_75t_L g237 ( .A(n_233), .B(n_145), .C(n_143), .Y(n_237) );
BUFx8_ASAP7_75t_SL g238 ( .A(n_220), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_219), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_228), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_224), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_228), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_230), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_229), .A2(n_21), .B(n_20), .Y(n_244) );
AND2x2_ASAP7_75t_L g245 ( .A(n_222), .B(n_7), .Y(n_245) );
BUFx12f_ASAP7_75t_L g246 ( .A(n_232), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_231), .B(n_7), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_218), .Y(n_248) );
OR2x6_ASAP7_75t_L g249 ( .A(n_218), .B(n_8), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_227), .A2(n_9), .B(n_10), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_219), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_223), .Y(n_252) );
INVx3_ASAP7_75t_L g253 ( .A(n_246), .Y(n_253) );
BUFx2_ASAP7_75t_SL g254 ( .A(n_239), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_248), .Y(n_255) );
INVx5_ASAP7_75t_L g256 ( .A(n_249), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_238), .Y(n_257) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_240), .Y(n_258) );
AO21x1_ASAP7_75t_SL g259 ( .A1(n_250), .A2(n_12), .B(n_13), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_234), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_251), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_247), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_245), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_243), .B(n_14), .Y(n_265) );
CKINVDCx6p67_ASAP7_75t_R g266 ( .A(n_241), .Y(n_266) );
OR2x6_ASAP7_75t_L g267 ( .A(n_244), .B(n_15), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_236), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g269 ( .A1(n_237), .A2(n_16), .B(n_24), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_252), .Y(n_270) );
OA21x2_ASAP7_75t_L g271 ( .A1(n_235), .A2(n_28), .B(n_30), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_246), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_270), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_264), .B(n_35), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_258), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_262), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_253), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_265), .B(n_38), .Y(n_278) );
INVx3_ASAP7_75t_L g279 ( .A(n_256), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_260), .B(n_39), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_265), .B(n_41), .Y(n_282) );
INVx3_ASAP7_75t_L g283 ( .A(n_256), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_258), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_272), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_263), .Y(n_287) );
NOR2x1p5_ASAP7_75t_L g288 ( .A(n_266), .B(n_50), .Y(n_288) );
BUFx3_ASAP7_75t_L g289 ( .A(n_257), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_254), .B(n_92), .Y(n_290) );
NAND2x1_ASAP7_75t_L g291 ( .A(n_267), .B(n_55), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_259), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_267), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_268), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_267), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_269), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_261), .B(n_63), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_273), .Y(n_298) );
OR2x2_ASAP7_75t_L g299 ( .A(n_275), .B(n_271), .Y(n_299) );
INVx4_ASAP7_75t_L g300 ( .A(n_277), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_293), .B(n_295), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_276), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_284), .B(n_67), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_285), .B(n_68), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_294), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_287), .B(n_69), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_292), .B(n_71), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_296), .B(n_72), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_292), .B(n_74), .Y(n_310) );
AND2x6_ASAP7_75t_SL g311 ( .A(n_297), .B(n_76), .Y(n_311) );
NOR2x1_ASAP7_75t_L g312 ( .A(n_288), .B(n_83), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_279), .B(n_86), .Y(n_313) );
NAND2x1_ASAP7_75t_L g314 ( .A(n_300), .B(n_281), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_301), .B(n_281), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_307), .B(n_283), .Y(n_316) );
OR2x2_ASAP7_75t_L g317 ( .A(n_298), .B(n_289), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_300), .B(n_291), .Y(n_318) );
INVxp67_ASAP7_75t_SL g319 ( .A(n_299), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_302), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_305), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_312), .B(n_290), .Y(n_322) );
BUFx2_ASAP7_75t_L g323 ( .A(n_321), .Y(n_323) );
INVx2_ASAP7_75t_SL g324 ( .A(n_317), .Y(n_324) );
INVxp67_ASAP7_75t_L g325 ( .A(n_316), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_314), .B(n_308), .Y(n_326) );
OR2x2_ASAP7_75t_L g327 ( .A(n_323), .B(n_319), .Y(n_327) );
INVx3_ASAP7_75t_L g328 ( .A(n_326), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_326), .A2(n_322), .B1(n_318), .B2(n_315), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_SL g330 ( .A1(n_327), .A2(n_325), .B(n_324), .C(n_310), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_330), .A2(n_329), .B(n_328), .Y(n_331) );
INVx1_ASAP7_75t_SL g332 ( .A(n_331), .Y(n_332) );
NAND4xp25_ASAP7_75t_L g333 ( .A(n_332), .B(n_282), .C(n_278), .D(n_311), .Y(n_333) );
NOR2x1_ASAP7_75t_L g334 ( .A(n_333), .B(n_313), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_334), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_335), .B(n_320), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_336), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_337), .Y(n_338) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_338), .A2(n_303), .B1(n_304), .B2(n_280), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_339), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_340), .B(n_306), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_341), .A2(n_274), .B(n_309), .Y(n_342) );
endmodule