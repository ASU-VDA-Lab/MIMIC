module fake_jpeg_22267_n_321 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_41),
.A2(n_45),
.B1(n_18),
.B2(n_26),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_30),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g64 ( 
.A(n_49),
.B(n_35),
.CON(n_64),
.SN(n_64)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_53),
.Y(n_95)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_28),
.B1(n_26),
.B2(n_18),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_41),
.A2(n_28),
.B1(n_27),
.B2(n_21),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_21),
.B1(n_27),
.B2(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_63),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_62),
.A2(n_73),
.B1(n_82),
.B2(n_20),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_64),
.A2(n_74),
.B(n_90),
.C(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_49),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_65),
.B(n_69),
.Y(n_91)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_34),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_37),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_80),
.Y(n_102)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_79),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_20),
.B1(n_37),
.B2(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_33),
.B1(n_29),
.B2(n_22),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_44),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_29),
.Y(n_96)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_37),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_83),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_36),
.B1(n_25),
.B2(n_32),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_40),
.B(n_33),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_84),
.B(n_22),
.C(n_31),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_49),
.B(n_36),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_41),
.A2(n_32),
.B1(n_31),
.B2(n_19),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_24),
.A3(n_30),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_88),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_39),
.B(n_0),
.Y(n_90)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_66),
.Y(n_92)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_93),
.A2(n_115),
.B1(n_68),
.B2(n_61),
.Y(n_152)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_96),
.B(n_114),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_104),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_105),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_55),
.C(n_58),
.Y(n_139)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_89),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_116),
.B(n_122),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_117),
.Y(n_127)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_118),
.Y(n_135)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_121),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_90),
.B(n_30),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_60),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_126),
.B(n_52),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_80),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_131),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_80),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_57),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_136),
.C(n_97),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_71),
.B(n_63),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_95),
.B(n_110),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_71),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_139),
.B(n_153),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g140 ( 
.A(n_109),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_145),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_92),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_141),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_59),
.B1(n_64),
.B2(n_24),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_144),
.A2(n_154),
.B1(n_148),
.B2(n_139),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_51),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_156),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_103),
.B(n_51),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_155),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_30),
.B(n_72),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_155),
.B(n_125),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_99),
.B(n_107),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_30),
.B1(n_2),
.B2(n_3),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_106),
.A2(n_1),
.B(n_2),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_1),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_157),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_160),
.Y(n_200)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_161),
.B(n_164),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_162),
.A2(n_174),
.B(n_151),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_126),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_163),
.A2(n_166),
.B(n_172),
.Y(n_221)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_177),
.C(n_133),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_175),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_171),
.A2(n_191),
.B1(n_165),
.B2(n_183),
.Y(n_209)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_134),
.A2(n_92),
.B(n_120),
.C(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_173),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_131),
.A2(n_97),
.B(n_91),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_121),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_111),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_181),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_111),
.C(n_109),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_105),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_186),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_137),
.A2(n_100),
.B1(n_118),
.B2(n_113),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_158),
.B1(n_146),
.B2(n_133),
.Y(n_210)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_101),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_185),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_135),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_150),
.B(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_132),
.B(n_94),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_188),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_138),
.B(n_3),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_189),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_4),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_193),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_4),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_146),
.B1(n_137),
.B2(n_158),
.Y(n_194)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_173),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_198),
.B(n_204),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_180),
.Y(n_232)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_220),
.C(n_192),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_166),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_210),
.A2(n_215),
.B1(n_170),
.B2(n_190),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_135),
.B1(n_159),
.B2(n_149),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_129),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_178),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_149),
.B1(n_142),
.B2(n_7),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_216),
.B(n_217),
.Y(n_225)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_222),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_219),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_5),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_168),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_239),
.B1(n_211),
.B2(n_172),
.Y(n_253)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_228),
.A2(n_242),
.B1(n_245),
.B2(n_170),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_206),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_229),
.B(n_237),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_234),
.C(n_244),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_201),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_233),
.A2(n_225),
.B(n_236),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_221),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_204),
.A2(n_172),
.A3(n_162),
.B1(n_164),
.B2(n_169),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_241),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_207),
.Y(n_236)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_236),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_208),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_181),
.Y(n_241)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_167),
.C(n_177),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_232),
.B(n_209),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_256),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_221),
.B1(n_203),
.B2(n_217),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_255),
.B1(n_230),
.B2(n_239),
.Y(n_269)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_195),
.B(n_196),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_264),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_253),
.B(n_258),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_220),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_202),
.C(n_207),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_262),
.C(n_245),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_200),
.B1(n_219),
.B2(n_198),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_213),
.B1(n_178),
.B2(n_237),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_261),
.A2(n_235),
.B(n_212),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_233),
.C(n_202),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_228),
.A2(n_200),
.B1(n_214),
.B2(n_161),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_227),
.A2(n_196),
.B(n_212),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_238),
.Y(n_266)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_266),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_247),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_260),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_270),
.B(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_273),
.C(n_278),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_230),
.C(n_174),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_172),
.B1(n_242),
.B2(n_188),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_SL g275 ( 
.A(n_261),
.B(n_172),
.C(n_186),
.Y(n_275)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_259),
.CI(n_256),
.CON(n_289),
.SN(n_289)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_224),
.C(n_222),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_5),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_279),
.B(n_248),
.C(n_262),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_287),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_SL g282 ( 
.A1(n_267),
.A2(n_257),
.B(n_251),
.C(n_246),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_277),
.B1(n_268),
.B2(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_258),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_289),
.B(n_276),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_6),
.C(n_7),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_292),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_6),
.C(n_8),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_294),
.A2(n_284),
.B1(n_287),
.B2(n_289),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_295),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_271),
.B(n_280),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_9),
.B(n_10),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_288),
.A2(n_273),
.B1(n_271),
.B2(n_280),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_299),
.A2(n_282),
.B1(n_291),
.B2(n_11),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_283),
.B(n_6),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_301),
.Y(n_305)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_281),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_304),
.C(n_307),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_298),
.B(n_285),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_306),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_282),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_308),
.B(n_295),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_310),
.B(n_307),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_299),
.B(n_297),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_313),
.B(n_297),
.C(n_296),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_316),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_315),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_317),
.A2(n_312),
.B(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_318),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_11),
.Y(n_321)
);


endmodule