module fake_jpeg_15343_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_19),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_23),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_33),
.B(n_16),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_27),
.A2(n_16),
.B1(n_25),
.B2(n_14),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_20),
.B1(n_18),
.B2(n_17),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_43),
.Y(n_57)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_19),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_28),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_33),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_44),
.B(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_52),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_23),
.B(n_15),
.C(n_28),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_26),
.B(n_0),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_49),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_28),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_24),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_24),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_27),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_31),
.C(n_22),
.Y(n_71)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_63),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_0),
.B(n_30),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_30),
.B1(n_32),
.B2(n_22),
.Y(n_68)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_50),
.B(n_49),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_59),
.C(n_55),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_72),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_81),
.Y(n_85)
);

OAI21x1_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_66),
.B(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_46),
.B(n_48),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_80),
.A2(n_82),
.B(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_56),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_83),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_71),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_86),
.B(n_87),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_74),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_74),
.Y(n_88)
);

NAND4xp25_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_79),
.C(n_76),
.D(n_62),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_89),
.A2(n_92),
.B(n_80),
.C(n_78),
.D(n_66),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_91),
.A2(n_92),
.B(n_58),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g102 ( 
.A1(n_93),
.A2(n_95),
.A3(n_86),
.B1(n_57),
.B2(n_69),
.C(n_90),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_77),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_98),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_70),
.C(n_78),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_99),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_69),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_101),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_104),
.B(n_107),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_93),
.C(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

AOI322xp5_ASAP7_75t_L g112 ( 
.A1(n_109),
.A2(n_110),
.A3(n_63),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_6),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_106),
.B(n_100),
.Y(n_110)
);

NAND3xp33_ASAP7_75t_SL g111 ( 
.A(n_108),
.B(n_107),
.C(n_32),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_112),
.Y(n_113)
);

AOI322xp5_ASAP7_75t_L g114 ( 
.A1(n_113),
.A2(n_1),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.C1(n_47),
.C2(n_31),
.Y(n_114)
);


endmodule