module real_jpeg_28240_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_3),
.A2(n_7),
.B1(n_24),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_26),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_3),
.A2(n_20),
.B1(n_22),
.B2(n_26),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_26),
.B1(n_77),
.B2(n_84),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_57),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_6),
.A2(n_7),
.B1(n_24),
.B2(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_6),
.A2(n_29),
.B1(n_40),
.B2(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_6),
.A2(n_20),
.B1(n_22),
.B2(n_29),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_6),
.A2(n_8),
.B(n_20),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_SL g76 ( 
.A1(n_6),
.A2(n_7),
.B(n_36),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_6),
.A2(n_29),
.B1(n_77),
.B2(n_84),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g118 ( 
.A1(n_6),
.A2(n_41),
.B(n_56),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_6),
.B(n_19),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g23 ( 
.A1(n_7),
.A2(n_8),
.B1(n_21),
.B2(n_24),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_24),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_7),
.A2(n_29),
.B(n_65),
.C(n_66),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_8),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_9),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_101),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_12),
.B(n_99),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_70),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_13),
.B(n_70),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_53),
.C(n_61),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_14),
.A2(n_15),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_16),
.B(n_32),
.C(n_38),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_25),
.B1(n_27),
.B2(n_30),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_18),
.B(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_20),
.A2(n_22),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_20),
.A2(n_29),
.B(n_57),
.C(n_118),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_25),
.A2(n_30),
.B(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_29),
.A2(n_35),
.B(n_76),
.C(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_29),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_29),
.B(n_58),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_34),
.B(n_88),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_35),
.A2(n_36),
.B1(n_77),
.B2(n_84),
.Y(n_88)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_37),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_37),
.B(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_38),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_43),
.B(n_44),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_43),
.B1(n_46),
.B2(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_40),
.B(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_43),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_47),
.Y(n_69)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_53),
.A2(n_61),
.B1(n_62),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_53),
.A2(n_112),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_53),
.B(n_79),
.C(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_54),
.B(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_54),
.B(n_60),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_64),
.B1(n_67),
.B2(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_80),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_77),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_79),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_136),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_89),
.B1(n_97),
.B2(n_98),
.Y(n_80)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_104),
.C(n_108),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_94),
.A2(n_95),
.B1(n_104),
.B2(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_113),
.B(n_145),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_109),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_103),
.B(n_109),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_117),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_104),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_140),
.B(n_144),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_124),
.B(n_139),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_119),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_117),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_121),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_129),
.B(n_138),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_135),
.B(n_137),
.Y(n_129)
);

INVx5_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_142),
.Y(n_144)
);


endmodule