module fake_jpeg_24130_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_28),
.A2(n_26),
.B1(n_21),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_13),
.B1(n_26),
.B2(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_40),
.B(n_44),
.Y(n_70)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_27),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_20),
.Y(n_90)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_71),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_64),
.A2(n_54),
.B1(n_55),
.B2(n_46),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_26),
.B1(n_21),
.B2(n_13),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_24),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_27),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_75),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_21),
.B1(n_26),
.B2(n_13),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_77),
.B(n_94),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_25),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_80),
.B(n_98),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_49),
.B1(n_48),
.B2(n_41),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_85),
.A2(n_92),
.B1(n_72),
.B2(n_67),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_58),
.A2(n_22),
.B(n_45),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_86),
.A2(n_14),
.B(n_15),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_49),
.B1(n_48),
.B2(n_37),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_70),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_89),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_14),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_41),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_61),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_59),
.A2(n_46),
.B1(n_44),
.B2(n_54),
.Y(n_93)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_100),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_101),
.B(n_103),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_88),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_104),
.A2(n_112),
.B1(n_121),
.B2(n_108),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_61),
.C(n_14),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_114),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_107),
.A2(n_120),
.B(n_98),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_15),
.C(n_14),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_81),
.A2(n_15),
.B1(n_55),
.B2(n_57),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_111),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_90),
.B(n_74),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_74),
.C(n_66),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_102),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_60),
.B(n_35),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_84),
.A2(n_62),
.B(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_123),
.A2(n_128),
.B1(n_132),
.B2(n_145),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_133),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_125),
.A2(n_109),
.B1(n_106),
.B2(n_116),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_113),
.B(n_80),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_136),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_134),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_112),
.A2(n_85),
.B1(n_92),
.B2(n_87),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_92),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_79),
.B(n_89),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_138),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_79),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_143),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_16),
.B(n_24),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_118),
.C(n_119),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_115),
.B(n_27),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_140),
.B(n_115),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_16),
.B(n_25),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_110),
.Y(n_162)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_108),
.A2(n_82),
.B1(n_78),
.B2(n_96),
.Y(n_145)
);

XNOR2x2_ASAP7_75t_SL g146 ( 
.A(n_125),
.B(n_109),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_127),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_121),
.B1(n_117),
.B2(n_116),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_147),
.A2(n_149),
.B1(n_158),
.B2(n_168),
.Y(n_174)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_144),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_166),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_128),
.A2(n_104),
.B1(n_117),
.B2(n_114),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_145),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_150),
.B(n_155),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_154),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_156),
.A2(n_169),
.B(n_129),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_82),
.B1(n_78),
.B2(n_96),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_104),
.B1(n_117),
.B2(n_110),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_19),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_139),
.C(n_127),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_111),
.Y(n_165)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_137),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_19),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_122),
.A2(n_117),
.B1(n_118),
.B2(n_95),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_184),
.Y(n_204)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_187),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_135),
.C(n_124),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_146),
.A2(n_131),
.B1(n_142),
.B2(n_138),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_179),
.A2(n_147),
.B1(n_167),
.B2(n_151),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_133),
.C(n_134),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_157),
.A2(n_101),
.B1(n_96),
.B2(n_95),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_164),
.B1(n_166),
.B2(n_152),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_20),
.A3(n_19),
.B1(n_51),
.B2(n_69),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_193),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_159),
.B(n_156),
.C(n_160),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_162),
.C(n_155),
.Y(n_203)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_51),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_190),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_150),
.A2(n_25),
.B1(n_23),
.B2(n_17),
.Y(n_191)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_179),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_168),
.B(n_149),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_198),
.A2(n_190),
.B(n_7),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_199),
.A2(n_201),
.B(n_194),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_164),
.B1(n_152),
.B2(n_169),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_192),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_193),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_208),
.C(n_213),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_19),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_6),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_23),
.C(n_17),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_177),
.A2(n_23),
.B1(n_17),
.B2(n_20),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_209),
.A2(n_183),
.B1(n_174),
.B2(n_173),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_181),
.B(n_175),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_211),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_20),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_212),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_0),
.C(n_1),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_230),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_213),
.B(n_203),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_217),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_186),
.B1(n_185),
.B2(n_171),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_218),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_210),
.B(n_172),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_222),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_189),
.C(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_226),
.C(n_227),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_223),
.B(n_224),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_207),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_197),
.B(n_208),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_0),
.C(n_1),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_6),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_228),
.B(n_0),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_216),
.A2(n_198),
.B(n_194),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_232),
.A2(n_238),
.B(n_240),
.Y(n_255)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_235),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_210),
.C(n_204),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_5),
.C(n_11),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_204),
.B(n_206),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_225),
.B(n_226),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_241),
.A2(n_227),
.B(n_8),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_7),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_244),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_215),
.B(n_7),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g247 ( 
.A(n_236),
.B(n_229),
.Y(n_247)
);

OAI21x1_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_259),
.B(n_4),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_215),
.B1(n_217),
.B2(n_219),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_252),
.C(n_254),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_234),
.B(n_10),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_0),
.C(n_1),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_256),
.B(n_239),
.C(n_10),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_232),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_257),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_245),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_258),
.B(n_256),
.Y(n_261)
);

NOR2x1_ASAP7_75t_SL g259 ( 
.A(n_233),
.B(n_12),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_262),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_261),
.B(n_9),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_237),
.Y(n_262)
);

AOI21x1_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_255),
.B(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_247),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_268),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_253),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_269),
.A2(n_254),
.B(n_248),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_263),
.Y(n_279)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_255),
.B(n_252),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_273),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_9),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_276),
.A2(n_263),
.B(n_266),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.C(n_281),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_280),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_283),
.Y(n_284)
);

OAI321xp33_ASAP7_75t_L g285 ( 
.A1(n_284),
.A2(n_277),
.A3(n_282),
.B1(n_274),
.B2(n_12),
.C(n_9),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_12),
.C(n_9),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_11),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_11),
.Y(n_288)
);


endmodule