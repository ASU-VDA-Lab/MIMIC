module fake_netlist_1_2400_n_26 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_3), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_8), .Y(n_12) );
BUFx16f_ASAP7_75t_R g13 ( .A(n_7), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_9), .Y(n_14) );
OA22x2_ASAP7_75t_L g15 ( .A1(n_11), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_11), .B(n_0), .Y(n_16) );
HB1xp67_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_15), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_17), .B(n_13), .Y(n_19) );
AOI21xp33_ASAP7_75t_SL g20 ( .A1(n_19), .A2(n_1), .B(n_10), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
BUFx6f_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
OAI22xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_19), .B1(n_18), .B2(n_12), .Y(n_24) );
OA22x2_ASAP7_75t_L g25 ( .A1(n_22), .A2(n_14), .B1(n_5), .B2(n_6), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_4), .B1(n_22), .B2(n_24), .Y(n_26) );
endmodule