module real_jpeg_23650_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_1),
.A2(n_37),
.B1(n_40),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_1),
.A2(n_46),
.B1(n_64),
.B2(n_65),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_63),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_3),
.Y(n_77)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_37),
.B1(n_40),
.B2(n_55),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_6),
.A2(n_55),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_6),
.A2(n_55),
.B1(n_64),
.B2(n_65),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_7),
.A2(n_27),
.B1(n_37),
.B2(n_40),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_7),
.A2(n_27),
.B1(n_48),
.B2(n_49),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_7),
.A2(n_27),
.B1(n_64),
.B2(n_65),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_8),
.A2(n_64),
.B1(n_65),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_8),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_69),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_11),
.B(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_11),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_11),
.B(n_36),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_11),
.B(n_49),
.C(n_51),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_37),
.B1(n_40),
.B2(n_157),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_11),
.B(n_105),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_11),
.A2(n_48),
.B1(n_49),
.B2(n_157),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_11),
.B(n_64),
.C(n_77),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_11),
.A2(n_66),
.B(n_218),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_13),
.A2(n_29),
.B1(n_34),
.B2(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_13),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_13),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_13),
.A2(n_42),
.B1(n_64),
.B2(n_65),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_14),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_14),
.A2(n_64),
.B1(n_65),
.B2(n_82),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_14),
.A2(n_37),
.B1(n_40),
.B2(n_82),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_15),
.A2(n_64),
.B1(n_65),
.B2(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_15),
.Y(n_86)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_16),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_16),
.A2(n_108),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_142),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_140),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_119),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_20),
.B(n_119),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.C(n_93),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_21),
.A2(n_22),
.B1(n_83),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_25),
.B(n_43),
.C(n_59),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_36),
.B2(n_41),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_26),
.Y(n_95)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_29),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_30),
.B(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_30),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_30),
.A2(n_137),
.B(n_156),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_35),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_32),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g118 ( 
.A(n_32),
.B(n_37),
.Y(n_118)
);

AOI32xp33_ASAP7_75t_L g114 ( 
.A1(n_33),
.A2(n_34),
.A3(n_40),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_34),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_35),
.A2(n_95),
.B(n_96),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_35),
.B(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_40),
.B1(n_51),
.B2(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_37),
.B(n_181),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_41),
.Y(n_134)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_53),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_45),
.A2(n_47),
.B1(n_57),
.B2(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_47),
.A2(n_53),
.B(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_49),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_49),
.B(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_54),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_56),
.A2(n_103),
.B1(n_105),
.B2(n_150),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_102),
.B(n_104),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_57),
.A2(n_104),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_73),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_60),
.B(n_73),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_66),
.B1(n_68),
.B2(n_70),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_62),
.A2(n_108),
.B1(n_109),
.B2(n_111),
.Y(n_107)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_67),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_65),
.B(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_66),
.A2(n_70),
.B(n_85),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_66),
.A2(n_110),
.B1(n_112),
.B2(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_66),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_66),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_72),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_72),
.B(n_157),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_74),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_74),
.A2(n_206),
.B(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_75),
.A2(n_89),
.B1(n_90),
.B2(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_75),
.B(n_154),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_75),
.A2(n_90),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_79),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_79),
.A2(n_80),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_79),
.A2(n_153),
.B(n_191),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_79),
.B(n_157),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_83),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_87),
.B1(n_91),
.B2(n_92),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_84),
.B(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_90),
.B(n_154),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_93),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.C(n_106),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_94),
.B(n_101),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g156 ( 
.A1(n_100),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_106),
.B(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_114),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_112),
.A2(n_231),
.B(n_239),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_115),
.Y(n_158)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_139),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_125),
.B2(n_126),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_130),
.B2(n_138),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_133),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B(n_136),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_173),
.B(n_260),
.C(n_265),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_167),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_167),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_159),
.C(n_160),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_145),
.A2(n_146),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_155),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_151),
.C(n_155),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_159),
.B(n_160),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_165),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_200),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_166),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_168),
.B(n_171),
.C(n_172),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_254),
.B(n_259),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_207),
.B(n_253),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_196),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_178),
.B(n_196),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_189),
.C(n_193),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_179),
.B(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_182),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_184),
.B(n_187),
.Y(n_182)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_187),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_189),
.A2(n_193),
.B1(n_194),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_189),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_192),
.Y(n_205)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_203),
.C(n_204),
.Y(n_258)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_247),
.B(n_252),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_227),
.B(n_246),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_221),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_221),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_251)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_217),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_225),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_235),
.B(n_245),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_244),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_251),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_258),
.Y(n_259)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);


endmodule