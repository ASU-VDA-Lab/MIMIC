module fake_jpeg_14408_n_272 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_272);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_272;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_39),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_6),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_40),
.B(n_42),
.Y(n_74)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_6),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_27),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_6),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_52),
.Y(n_63)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_29),
.A2(n_0),
.B(n_1),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_30),
.B(n_7),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_22),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_1),
.Y(n_62)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_59),
.A2(n_61),
.B1(n_69),
.B2(n_72),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_62),
.B(n_63),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_28),
.B1(n_15),
.B2(n_25),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_68),
.A2(n_75),
.B1(n_91),
.B2(n_51),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_39),
.A2(n_17),
.B1(n_32),
.B2(n_27),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_17),
.B1(n_32),
.B2(n_15),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_23),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_100),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_15),
.B1(n_17),
.B2(n_19),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_41),
.A2(n_32),
.B1(n_23),
.B2(n_21),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_79),
.B1(n_5),
.B2(n_12),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_21),
.B1(n_20),
.B2(n_16),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_30),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_80),
.B(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_35),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_19),
.B1(n_16),
.B2(n_26),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_34),
.B1(n_10),
.B2(n_4),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_37),
.Y(n_93)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_93),
.Y(n_128)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_43),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_97),
.A2(n_98),
.B1(n_44),
.B2(n_51),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_43),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_14),
.Y(n_99)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_99),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_2),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_95),
.B(n_54),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_102),
.Y(n_163)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_104),
.A2(n_105),
.B1(n_114),
.B2(n_115),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_55),
.B1(n_48),
.B2(n_45),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_121),
.B1(n_125),
.B2(n_96),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_55),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_112),
.C(n_123),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_48),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_58),
.B1(n_34),
.B2(n_3),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_SL g115 ( 
.A1(n_85),
.A2(n_58),
.B(n_9),
.C(n_10),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_83),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_73),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_122),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_12),
.B1(n_13),
.B2(n_100),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_76),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_13),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_124),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_13),
.B1(n_89),
.B2(n_86),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_92),
.A2(n_76),
.B1(n_70),
.B2(n_84),
.Y(n_129)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_106),
.A3(n_113),
.B1(n_115),
.B2(n_90),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_66),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g131 ( 
.A(n_62),
.B(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_131),
.B(n_112),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_84),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_144),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_136),
.B(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_137),
.A2(n_149),
.B1(n_164),
.B2(n_163),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_70),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_60),
.B(n_74),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_145),
.A2(n_123),
.B(n_102),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_74),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_149),
.A2(n_103),
.B1(n_129),
.B2(n_132),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_94),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_83),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_162),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_60),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_121),
.C(n_102),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_109),
.B(n_90),
.C(n_66),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_158),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_109),
.B(n_96),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_159),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_65),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_103),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_161),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_65),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_78),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_78),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_111),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_167),
.A2(n_135),
.B(n_147),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_104),
.B1(n_107),
.B2(n_105),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_168),
.A2(n_179),
.B1(n_189),
.B2(n_190),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_107),
.B1(n_115),
.B2(n_129),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_184),
.B1(n_187),
.B2(n_192),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_174),
.C(n_187),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_179),
.B(n_167),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_144),
.A2(n_129),
.B1(n_86),
.B2(n_117),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_183),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_153),
.B(n_111),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_185),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_118),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_156),
.A2(n_71),
.B1(n_117),
.B2(n_162),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_133),
.B(n_71),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_156),
.A2(n_152),
.B1(n_139),
.B2(n_163),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_156),
.A2(n_137),
.B1(n_149),
.B2(n_139),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_140),
.A2(n_150),
.B1(n_143),
.B2(n_145),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_191),
.A2(n_189),
.B1(n_168),
.B2(n_173),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_141),
.A2(n_142),
.B1(n_158),
.B2(n_146),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_140),
.B1(n_135),
.B2(n_160),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_198),
.B(n_203),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_134),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_134),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_200),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_172),
.B(n_135),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_166),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_186),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_206),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_181),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_183),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_165),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_147),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_176),
.C(n_182),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_173),
.B1(n_171),
.B2(n_170),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_177),
.B1(n_188),
.B2(n_210),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_214),
.A2(n_170),
.B1(n_169),
.B2(n_185),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_225),
.C(n_226),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_229),
.B1(n_206),
.B2(n_203),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_212),
.B(n_169),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_180),
.C(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_231),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_195),
.A2(n_214),
.B1(n_204),
.B2(n_197),
.Y(n_231)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_236),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_221),
.B(n_196),
.Y(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_210),
.B1(n_213),
.B2(n_227),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_223),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_238),
.A2(n_228),
.B1(n_224),
.B2(n_216),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_218),
.B(n_196),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_240),
.B(n_242),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_201),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_198),
.B(n_193),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_220),
.B(n_205),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_227),
.B(n_198),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_233),
.B(n_217),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_236),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_246),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_225),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_237),
.A2(n_230),
.B(n_226),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_248),
.B(n_235),
.Y(n_255)
);

O2A1O1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_195),
.B(n_229),
.C(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_249),
.A2(n_232),
.B1(n_240),
.B2(n_199),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_250),
.B(n_224),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_254),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_255),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_235),
.B(n_249),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_258),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_244),
.A2(n_232),
.B1(n_228),
.B2(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_251),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_259),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_253),
.B(n_243),
.C(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_247),
.C(n_219),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_260),
.A2(n_258),
.B(n_257),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_263),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_262),
.C(n_247),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_268),
.C(n_261),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_269),
.A2(n_266),
.B(n_208),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_209),
.B(n_200),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_207),
.Y(n_272)
);


endmodule