module fake_jpeg_11171_n_302 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_302);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_302;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_23),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_48),
.B(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_23),
.Y(n_50)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g93 ( 
.A(n_53),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_56),
.B(n_57),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_61),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_43),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_71),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_41),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_31),
.C(n_34),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_42),
.C(n_19),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_30),
.B1(n_34),
.B2(n_27),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_25),
.B1(n_26),
.B2(n_17),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_43),
.Y(n_76)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_78),
.B(n_83),
.Y(n_110)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_47),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_34),
.B1(n_27),
.B2(n_33),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_100),
.B1(n_105),
.B2(n_55),
.Y(n_107)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_29),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_34),
.B1(n_19),
.B2(n_26),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_85),
.A2(n_86),
.B1(n_95),
.B2(n_98),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_22),
.B1(n_28),
.B2(n_20),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_88),
.B(n_10),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_61),
.A2(n_32),
.B(n_21),
.C(n_20),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_90),
.A2(n_104),
.B(n_69),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_51),
.A2(n_24),
.B1(n_18),
.B2(n_32),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_97),
.B(n_102),
.Y(n_132)
);

AO22x2_ASAP7_75t_SL g98 ( 
.A1(n_53),
.A2(n_38),
.B1(n_24),
.B2(n_18),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_55),
.B1(n_65),
.B2(n_67),
.Y(n_117)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_69),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_51),
.A2(n_24),
.B1(n_18),
.B2(n_21),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_28),
.B1(n_38),
.B2(n_2),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_0),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_38),
.B(n_1),
.C(n_3),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_60),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_107),
.B(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_85),
.C(n_96),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_87),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_117),
.B1(n_122),
.B2(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_97),
.B(n_62),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_125),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_55),
.B(n_47),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_96),
.B(n_106),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_60),
.B1(n_59),
.B2(n_47),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_92),
.B(n_59),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_78),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_103),
.A2(n_70),
.B1(n_49),
.B2(n_9),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_102),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_76),
.B(n_70),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_83),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_87),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_134),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_87),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_135),
.B(n_159),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_90),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_136),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_74),
.B1(n_76),
.B2(n_98),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_139),
.A2(n_142),
.B1(n_160),
.B2(n_162),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

AO21x2_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_104),
.B(n_93),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_84),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_149),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_83),
.B(n_93),
.C(n_100),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_79),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_154),
.C(n_165),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_91),
.C(n_94),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_111),
.B(n_82),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_151),
.Y(n_190)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_107),
.A2(n_95),
.B1(n_77),
.B2(n_89),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_163),
.B1(n_127),
.B2(n_134),
.Y(n_168)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_158),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_99),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_81),
.B1(n_77),
.B2(n_106),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_110),
.A2(n_49),
.B1(n_8),
.B2(n_11),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_132),
.A2(n_49),
.B1(n_8),
.B2(n_11),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_0),
.B(n_1),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_111),
.B(n_6),
.C(n_14),
.Y(n_165)
);

BUFx10_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_166),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_133),
.B1(n_130),
.B2(n_122),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_167),
.A2(n_173),
.B1(n_181),
.B2(n_146),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_168),
.B(n_190),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_172),
.B(n_185),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_133),
.B1(n_108),
.B2(n_112),
.Y(n_173)
);

AOI22x1_ASAP7_75t_L g177 ( 
.A1(n_161),
.A2(n_121),
.B1(n_114),
.B2(n_115),
.Y(n_177)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_108),
.B1(n_124),
.B2(n_115),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_180),
.A2(n_139),
.B1(n_142),
.B2(n_145),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_124),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_154),
.C(n_156),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_137),
.C(n_161),
.Y(n_200)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_7),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_193),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_114),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_189),
.Y(n_203)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_137),
.B(n_108),
.C(n_6),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_142),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_15),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_13),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_195),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_163),
.B(n_7),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_204),
.C(n_206),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_202),
.A2(n_162),
.B1(n_171),
.B2(n_189),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_184),
.Y(n_204)
);

XOR2x1_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_136),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_177),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_169),
.Y(n_208)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_164),
.B(n_136),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_213),
.B(n_191),
.Y(n_227)
);

BUFx24_ASAP7_75t_SL g211 ( 
.A(n_170),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_178),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_182),
.A2(n_142),
.B(n_147),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_217),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_167),
.B1(n_182),
.B2(n_173),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_216),
.B(n_218),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_179),
.B(n_140),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_175),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_174),
.B(n_140),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_219),
.B(n_182),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_190),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_221),
.A2(n_196),
.B1(n_216),
.B2(n_215),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_223),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_235),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_178),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_228),
.C(n_234),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_232),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_177),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_191),
.B(n_176),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_202),
.A2(n_168),
.B1(n_142),
.B2(n_187),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_233),
.A2(n_239),
.B1(n_209),
.B2(n_205),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_143),
.C(n_166),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_212),
.B(n_176),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_158),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_238),
.B(n_241),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_222),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_243),
.Y(n_259)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_207),
.B1(n_196),
.B2(n_220),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_248),
.B1(n_230),
.B2(n_234),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_231),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_249),
.A2(n_256),
.B1(n_229),
.B2(n_222),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_253),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_218),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_231),
.B(n_201),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_230),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_240),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_233),
.A2(n_214),
.B1(n_198),
.B2(n_210),
.Y(n_256)
);

NAND4xp25_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_166),
.C(n_232),
.D(n_227),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_265),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_228),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_261),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_262),
.A2(n_270),
.B1(n_257),
.B2(n_254),
.Y(n_272)
);

FAx1_ASAP7_75t_SL g264 ( 
.A(n_247),
.B(n_224),
.CI(n_226),
.CON(n_264),
.SN(n_264)
);

A2O1A1O1Ixp25_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_245),
.B(n_262),
.C(n_268),
.D(n_250),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_230),
.C(n_166),
.Y(n_265)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_266),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_240),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_243),
.C(n_252),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_256),
.C(n_245),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_251),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_267),
.A2(n_244),
.B(n_257),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_259),
.B1(n_264),
.B2(n_229),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_260),
.C(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_274),
.B(n_278),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_277),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_203),
.C(n_242),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g281 ( 
.A(n_263),
.Y(n_281)
);

AOI21xp33_ASAP7_75t_L g284 ( 
.A1(n_281),
.A2(n_143),
.B(n_264),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_274),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_284),
.B(n_275),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_279),
.A2(n_266),
.B1(n_171),
.B2(n_12),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_286),
.A2(n_12),
.B(n_3),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_273),
.B1(n_280),
.B2(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_290),
.Y(n_294)
);

NAND4xp25_ASAP7_75t_SL g291 ( 
.A(n_287),
.B(n_12),
.C(n_1),
.D(n_3),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_0),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_292),
.A2(n_293),
.B(n_282),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_295),
.B(n_296),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_294),
.A2(n_285),
.B(n_291),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_298),
.Y(n_299)
);

AO22x1_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_285),
.B1(n_297),
.B2(n_4),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_300),
.A2(n_4),
.B1(n_5),
.B2(n_195),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_301),
.A2(n_4),
.B(n_5),
.Y(n_302)
);


endmodule