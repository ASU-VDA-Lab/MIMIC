module fake_jpeg_30261_n_126 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_37),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx4f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_1),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_61),
.Y(n_72)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_2),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_50),
.B1(n_51),
.B2(n_42),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_42),
.B1(n_51),
.B2(n_49),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_69),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_58),
.A2(n_47),
.B1(n_43),
.B2(n_53),
.Y(n_67)
);

OAI32xp33_ASAP7_75t_L g87 ( 
.A1(n_67),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_3),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_68),
.B(n_7),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_49),
.B1(n_48),
.B2(n_52),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_48),
.B1(n_45),
.B2(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_74),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_41),
.B1(n_22),
.B2(n_23),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_72),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_76),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_5),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_6),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_77),
.B(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_70),
.B(n_6),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_86),
.B(n_88),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_21),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_8),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_95),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_82),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_105),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_82),
.B(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_12),
.C(n_13),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_99),
.C(n_31),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_16),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_100),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_101),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_107),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_110),
.C(n_105),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_33),
.Y(n_110)
);

AND2x4_ASAP7_75t_SL g113 ( 
.A(n_98),
.B(n_34),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_114),
.B(n_90),
.Y(n_118)
);

NAND2x1p5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_35),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_116),
.B(n_118),
.Y(n_120)
);

NOR4xp25_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_113),
.C(n_111),
.D(n_92),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_115),
.C(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_120),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_94),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_100),
.B(n_112),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_104),
.B1(n_97),
.B2(n_91),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_36),
.Y(n_126)
);


endmodule