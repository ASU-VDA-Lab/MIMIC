module fake_jpeg_1278_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_4),
.B(n_1),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_0),
.Y(n_10)
);

INVx6_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx13_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx5_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g18 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_10),
.B1(n_8),
.B2(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_0),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_3),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_23),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_SL g23 ( 
.A(n_12),
.B(n_3),
.C(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_28),
.B1(n_14),
.B2(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_19),
.A2(n_16),
.B(n_10),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_33),
.B(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_17),
.B(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_25),
.A2(n_20),
.B1(n_24),
.B2(n_21),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_40),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_9),
.B1(n_15),
.B2(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_34),
.A2(n_30),
.B(n_29),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_46),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_29),
.C(n_9),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_32),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_37),
.C(n_35),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.C(n_51),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_35),
.C(n_40),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_43),
.B(n_39),
.C(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_54),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_36),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_12),
.B(n_14),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_56),
.A2(n_55),
.B(n_57),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_53),
.B(n_6),
.Y(n_59)
);


endmodule