module fake_netlist_6_2657_n_19665 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_19665);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_19665;

wire n_5643;
wire n_18652;
wire n_2817;
wire n_18318;
wire n_2576;
wire n_1674;
wire n_16664;
wire n_19057;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_1212;
wire n_208;
wire n_4251;
wire n_11111;
wire n_7933;
wire n_578;
wire n_4395;
wire n_19613;
wire n_1061;
wire n_16335;
wire n_5653;
wire n_4978;
wire n_13125;
wire n_3088;
wire n_8186;
wire n_6725;
wire n_6126;
wire n_4699;
wire n_17647;
wire n_8899;
wire n_5345;
wire n_17634;
wire n_10053;
wire n_1930;
wire n_8534;
wire n_3376;
wire n_4868;
wire n_10020;
wire n_17991;
wire n_15665;
wire n_19382;
wire n_1555;
wire n_17735;
wire n_19161;
wire n_7161;
wire n_19232;
wire n_830;
wire n_7868;
wire n_15764;
wire n_5725;
wire n_447;
wire n_5229;
wire n_3427;
wire n_18903;
wire n_18105;
wire n_5101;
wire n_3071;
wire n_8561;
wire n_14998;
wire n_14944;
wire n_11954;
wire n_19220;
wire n_14341;
wire n_10392;
wire n_15074;
wire n_5545;
wire n_2321;
wire n_15253;
wire n_4501;
wire n_9626;
wire n_5598;
wire n_19097;
wire n_15898;
wire n_18013;
wire n_7389;
wire n_10719;
wire n_5259;
wire n_6913;
wire n_10015;
wire n_6948;
wire n_3929;
wire n_3048;
wire n_9362;
wire n_7516;
wire n_7401;
wire n_12767;
wire n_16095;
wire n_18502;
wire n_5930;
wire n_9658;
wire n_1971;
wire n_5354;
wire n_8426;
wire n_5908;
wire n_953;
wire n_3664;
wire n_13681;
wire n_5420;
wire n_17209;
wire n_6243;
wire n_4414;
wire n_6585;
wire n_16553;
wire n_18122;
wire n_2625;
wire n_11543;
wire n_4646;
wire n_7651;
wire n_2843;
wire n_3760;
wire n_14662;
wire n_13247;
wire n_16286;
wire n_7956;
wire n_7369;
wire n_16549;
wire n_15421;
wire n_5136;
wire n_15964;
wire n_5638;
wire n_9100;
wire n_6784;
wire n_18310;
wire n_10868;
wire n_9067;
wire n_6323;
wire n_17847;
wire n_14431;
wire n_17478;
wire n_13515;
wire n_6110;
wire n_1967;
wire n_11684;
wire n_16324;
wire n_14410;
wire n_15800;
wire n_9400;
wire n_1911;
wire n_13139;
wire n_7774;
wire n_15600;
wire n_16267;
wire n_6951;
wire n_15899;
wire n_279;
wire n_18317;
wire n_2735;
wire n_13729;
wire n_4671;
wire n_18709;
wire n_14813;
wire n_4314;
wire n_18002;
wire n_323;
wire n_14628;
wire n_8421;
wire n_1381;
wire n_331;
wire n_2093;
wire n_18863;
wire n_17854;
wire n_10114;
wire n_10357;
wire n_15762;
wire n_2770;
wire n_16351;
wire n_15883;
wire n_17706;
wire n_8389;
wire n_2917;
wire n_13711;
wire n_16721;
wire n_12742;
wire n_3923;
wire n_11768;
wire n_9267;
wire n_939;
wire n_19401;
wire n_9652;
wire n_5493;
wire n_8849;
wire n_9059;
wire n_15332;
wire n_5346;
wire n_5252;
wire n_3446;
wire n_18445;
wire n_5309;
wire n_1895;
wire n_4698;
wire n_16254;
wire n_7564;
wire n_3859;
wire n_14989;
wire n_17564;
wire n_10204;
wire n_6383;
wire n_3397;
wire n_18669;
wire n_11637;
wire n_3575;
wire n_8151;
wire n_2469;
wire n_9038;
wire n_16004;
wire n_8748;
wire n_13984;
wire n_5452;
wire n_6794;
wire n_18608;
wire n_8718;
wire n_2764;
wire n_9935;
wire n_6990;
wire n_14288;
wire n_14824;
wire n_18699;
wire n_8223;
wire n_4856;
wire n_3492;
wire n_9135;
wire n_16800;
wire n_13771;
wire n_18644;
wire n_11295;
wire n_4291;
wire n_13960;
wire n_5532;
wire n_5897;
wire n_2434;
wire n_9070;
wire n_11708;
wire n_15629;
wire n_14401;
wire n_10827;
wire n_3247;
wire n_5922;
wire n_14922;
wire n_12158;
wire n_7823;
wire n_7569;
wire n_7062;
wire n_9477;
wire n_14769;
wire n_355;
wire n_8577;
wire n_14961;
wire n_8594;
wire n_8428;
wire n_9829;
wire n_13341;
wire n_2254;
wire n_5058;
wire n_10685;
wire n_1926;
wire n_17139;
wire n_15185;
wire n_12083;
wire n_12014;
wire n_14803;
wire n_19270;
wire n_1747;
wire n_16035;
wire n_10607;
wire n_15490;
wire n_18033;
wire n_5042;
wire n_19569;
wire n_8164;
wire n_4072;
wire n_835;
wire n_928;
wire n_15100;
wire n_10368;
wire n_19137;
wire n_9088;
wire n_10183;
wire n_17161;
wire n_6952;
wire n_11464;
wire n_19421;
wire n_3997;
wire n_14878;
wire n_15046;
wire n_2468;
wire n_5144;
wire n_10383;
wire n_2096;
wire n_3968;
wire n_4466;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_13550;
wire n_17601;
wire n_13348;
wire n_2812;
wire n_10724;
wire n_16398;
wire n_19396;
wire n_9988;
wire n_7009;
wire n_2136;
wire n_2409;
wire n_3834;
wire n_11553;
wire n_12795;
wire n_2075;
wire n_10876;
wire n_18780;
wire n_9137;
wire n_11180;
wire n_14043;
wire n_18820;
wire n_3192;
wire n_8995;
wire n_1546;
wire n_4394;
wire n_6010;
wire n_3352;
wire n_8711;
wire n_12505;
wire n_18602;
wire n_2150;
wire n_4082;
wire n_1420;
wire n_13721;
wire n_18430;
wire n_10820;
wire n_13514;
wire n_8306;
wire n_7488;
wire n_2558;
wire n_13194;
wire n_8887;
wire n_18677;
wire n_16183;
wire n_4289;
wire n_11866;
wire n_11450;
wire n_13575;
wire n_12522;
wire n_15659;
wire n_1487;
wire n_9578;
wire n_13109;
wire n_7438;
wire n_16631;
wire n_14355;
wire n_7337;
wire n_9489;
wire n_14123;
wire n_5957;
wire n_10728;
wire n_6357;
wire n_925;
wire n_6800;
wire n_18962;
wire n_4322;
wire n_10655;
wire n_9797;
wire n_1249;
wire n_2693;
wire n_8332;
wire n_9478;
wire n_2767;
wire n_11379;
wire n_16627;
wire n_19571;
wire n_19659;
wire n_10670;
wire n_5929;
wire n_5787;
wire n_11981;
wire n_19181;
wire n_9351;
wire n_5445;
wire n_14556;
wire n_6839;
wire n_532;
wire n_173;
wire n_9189;
wire n_413;
wire n_18888;
wire n_16528;
wire n_2170;
wire n_4156;
wire n_14701;
wire n_7098;
wire n_16587;
wire n_18936;
wire n_3158;
wire n_1788;
wire n_8921;
wire n_9356;
wire n_15880;
wire n_16499;
wire n_1835;
wire n_5076;
wire n_18328;
wire n_5870;
wire n_9175;
wire n_6508;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_10959;
wire n_6809;
wire n_11233;
wire n_4310;
wire n_7782;
wire n_5212;
wire n_13385;
wire n_2689;
wire n_1473;
wire n_6636;
wire n_5286;
wire n_16339;
wire n_1246;
wire n_4528;
wire n_899;
wire n_13992;
wire n_17429;
wire n_19103;
wire n_13790;
wire n_4914;
wire n_499;
wire n_3418;
wire n_705;
wire n_1004;
wire n_10624;
wire n_13304;
wire n_14633;
wire n_15699;
wire n_11900;
wire n_2297;
wire n_5901;
wire n_6538;
wire n_5599;
wire n_12883;
wire n_5324;
wire n_2103;
wire n_8983;
wire n_10422;
wire n_3770;
wire n_9818;
wire n_4402;
wire n_927;
wire n_16503;
wire n_18974;
wire n_12367;
wire n_17360;
wire n_5009;
wire n_13526;
wire n_12563;
wire n_7243;
wire n_13321;
wire n_15042;
wire n_15519;
wire n_14722;
wire n_13427;
wire n_4627;
wire n_4079;
wire n_9909;
wire n_19607;
wire n_8620;
wire n_19204;
wire n_15264;
wire n_13270;
wire n_10052;
wire n_10109;
wire n_18151;
wire n_3390;
wire n_19582;
wire n_10448;
wire n_11196;
wire n_16239;
wire n_11963;
wire n_16334;
wire n_8424;
wire n_9571;
wire n_2137;
wire n_16003;
wire n_4798;
wire n_2532;
wire n_12655;
wire n_7941;
wire n_16096;
wire n_18628;
wire n_11483;
wire n_15067;
wire n_19591;
wire n_19345;
wire n_5089;
wire n_13356;
wire n_2849;
wire n_14912;
wire n_1398;
wire n_884;
wire n_19177;
wire n_731;
wire n_8907;
wire n_11080;
wire n_958;
wire n_5137;
wire n_17557;
wire n_14079;
wire n_15168;
wire n_9894;
wire n_8324;
wire n_15411;
wire n_10906;
wire n_6380;
wire n_9441;
wire n_7913;
wire n_15144;
wire n_5288;
wire n_3606;
wire n_819;
wire n_14224;
wire n_2788;
wire n_10380;
wire n_6449;
wire n_18687;
wire n_6461;
wire n_3892;
wire n_18273;
wire n_4069;
wire n_14682;
wire n_2748;
wire n_5194;
wire n_1834;
wire n_9033;
wire n_2331;
wire n_15031;
wire n_12933;
wire n_15718;
wire n_9537;
wire n_11297;
wire n_14635;
wire n_17076;
wire n_13893;
wire n_5947;
wire n_1877;
wire n_2030;
wire n_11946;
wire n_9443;
wire n_9996;
wire n_14950;
wire n_7800;
wire n_13795;
wire n_3026;
wire n_17501;
wire n_14547;
wire n_15416;
wire n_221;
wire n_3847;
wire n_2552;
wire n_17942;
wire n_18735;
wire n_9938;
wire n_7261;
wire n_9023;
wire n_14415;
wire n_11818;
wire n_16298;
wire n_18739;
wire n_6773;
wire n_13569;
wire n_18042;
wire n_7455;
wire n_19105;
wire n_2160;
wire n_9201;
wire n_6531;
wire n_10952;
wire n_2131;
wire n_13628;
wire n_18958;
wire n_9559;
wire n_11803;
wire n_15738;
wire n_16301;
wire n_8015;
wire n_18507;
wire n_1933;
wire n_19102;
wire n_15613;
wire n_14786;
wire n_4411;
wire n_9184;
wire n_13585;
wire n_18418;
wire n_18472;
wire n_8024;
wire n_12562;
wire n_18396;
wire n_4180;
wire n_16531;
wire n_3354;
wire n_11090;
wire n_19035;
wire n_5740;
wire n_5820;
wire n_13266;
wire n_13957;
wire n_9403;
wire n_9875;
wire n_5180;
wire n_2049;
wire n_5182;
wire n_11561;
wire n_5534;
wire n_8003;
wire n_8785;
wire n_3566;
wire n_17826;
wire n_2829;
wire n_8692;
wire n_6889;
wire n_16142;
wire n_9183;
wire n_3804;
wire n_4207;
wire n_14326;
wire n_5196;
wire n_16381;
wire n_10852;
wire n_4470;
wire n_9529;
wire n_3901;
wire n_465;
wire n_11425;
wire n_4704;
wire n_2142;
wire n_4596;
wire n_6478;
wire n_820;
wire n_6100;
wire n_6516;
wire n_17845;
wire n_6977;
wire n_16854;
wire n_17542;
wire n_7660;
wire n_2263;
wire n_6911;
wire n_6599;
wire n_6522;
wire n_17189;
wire n_5660;
wire n_2756;
wire n_5334;
wire n_9347;
wire n_807;
wire n_4761;
wire n_18879;
wire n_16395;
wire n_13603;
wire n_6207;
wire n_6931;
wire n_7948;
wire n_238;
wire n_9082;
wire n_1595;
wire n_8685;
wire n_6963;
wire n_16252;
wire n_4932;
wire n_19358;
wire n_5456;
wire n_10618;
wire n_9594;
wire n_7837;
wire n_19531;
wire n_9445;
wire n_7627;
wire n_9803;
wire n_16698;
wire n_17041;
wire n_7601;
wire n_3195;
wire n_6346;
wire n_4274;
wire n_15729;
wire n_17519;
wire n_5386;
wire n_14737;
wire n_11676;
wire n_12266;
wire n_2595;
wire n_16949;
wire n_12287;
wire n_13485;
wire n_12991;
wire n_11134;
wire n_13735;
wire n_8886;
wire n_7211;
wire n_10933;
wire n_5618;
wire n_8506;
wire n_2264;
wire n_6494;
wire n_16365;
wire n_11548;
wire n_13041;
wire n_17037;
wire n_13154;
wire n_7822;
wire n_6453;
wire n_9307;
wire n_10762;
wire n_11342;
wire n_7785;
wire n_1891;
wire n_1213;
wire n_2235;
wire n_11266;
wire n_5082;
wire n_5338;
wire n_12479;
wire n_8352;
wire n_18941;
wire n_10360;
wire n_9450;
wire n_2298;
wire n_490;
wire n_3594;
wire n_5689;
wire n_16777;
wire n_4165;
wire n_12454;
wire n_8143;
wire n_10480;
wire n_4626;
wire n_4144;
wire n_12537;
wire n_17183;
wire n_9693;
wire n_17582;
wire n_12921;
wire n_2169;
wire n_13567;
wire n_11957;
wire n_10633;
wire n_13686;
wire n_13645;
wire n_16753;
wire n_12215;
wire n_18473;
wire n_9880;
wire n_12467;
wire n_6329;
wire n_11607;
wire n_11546;
wire n_15259;
wire n_16946;
wire n_15460;
wire n_330;
wire n_7158;
wire n_1406;
wire n_13400;
wire n_9905;
wire n_18717;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_13331;
wire n_9456;
wire n_7044;
wire n_9710;
wire n_8623;
wire n_11113;
wire n_18593;
wire n_2518;
wire n_17769;
wire n_19193;
wire n_13812;
wire n_14970;
wire n_7838;
wire n_4842;
wire n_204;
wire n_482;
wire n_4135;
wire n_16969;
wire n_1845;
wire n_12731;
wire n_7518;
wire n_2798;
wire n_6147;
wire n_9199;
wire n_13544;
wire n_7791;
wire n_2753;
wire n_2007;
wire n_2039;
wire n_18172;
wire n_12616;
wire n_1544;
wire n_18333;
wire n_3437;
wire n_4111;
wire n_14375;
wire n_12653;
wire n_533;
wire n_7146;
wire n_18081;
wire n_16580;
wire n_18498;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_12587;
wire n_10747;
wire n_13110;
wire n_16628;
wire n_2973;
wire n_9422;
wire n_18344;
wire n_5218;
wire n_12348;
wire n_3665;
wire n_16929;
wire n_273;
wire n_16099;
wire n_15590;
wire n_10843;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_16869;
wire n_3174;
wire n_10997;
wire n_1948;
wire n_9010;
wire n_13707;
wire n_15241;
wire n_19640;
wire n_6073;
wire n_19157;
wire n_6331;
wire n_13498;
wire n_2283;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_18289;
wire n_11408;
wire n_4196;
wire n_2056;
wire n_13183;
wire n_12519;
wire n_17184;
wire n_4902;
wire n_6405;
wire n_7580;
wire n_14077;
wire n_13007;
wire n_2680;
wire n_10112;
wire n_7304;
wire n_3713;
wire n_1931;
wire n_502;
wire n_1257;
wire n_3197;
wire n_7223;
wire n_14868;
wire n_7833;
wire n_5512;
wire n_9297;
wire n_2398;
wire n_6206;
wire n_9068;
wire n_8136;
wire n_5033;
wire n_9808;
wire n_18534;
wire n_2695;
wire n_4035;
wire n_7445;
wire n_11086;
wire n_6529;
wire n_1949;
wire n_3759;
wire n_4516;
wire n_1804;
wire n_11710;
wire n_251;
wire n_10253;
wire n_6290;
wire n_6025;
wire n_1337;
wire n_6455;
wire n_15277;
wire n_18435;
wire n_13804;
wire n_12455;
wire n_13099;
wire n_4492;
wire n_19524;
wire n_18516;
wire n_5607;
wire n_7695;
wire n_7179;
wire n_7122;
wire n_12157;
wire n_5999;
wire n_6203;
wire n_15806;
wire n_13064;
wire n_7630;
wire n_16246;
wire n_8643;
wire n_15660;
wire n_15357;
wire n_10821;
wire n_8565;
wire n_13648;
wire n_4542;
wire n_6892;
wire n_4462;
wire n_15722;
wire n_14181;
wire n_15278;
wire n_18054;
wire n_13338;
wire n_6685;
wire n_11639;
wire n_4931;
wire n_14213;
wire n_17320;
wire n_17885;
wire n_7051;
wire n_8477;
wire n_9793;
wire n_11692;
wire n_15054;
wire n_14842;
wire n_13115;
wire n_1291;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_5911;
wire n_11601;
wire n_11971;
wire n_2122;
wire n_12314;
wire n_3503;
wire n_1065;
wire n_11116;
wire n_12604;
wire n_13305;
wire n_1255;
wire n_8876;
wire n_5124;
wire n_19017;
wire n_3951;
wire n_9359;
wire n_14189;
wire n_3874;
wire n_15761;
wire n_5123;
wire n_8060;
wire n_3027;
wire n_4083;
wire n_11124;
wire n_6392;
wire n_182;
wire n_17470;
wire n_15301;
wire n_7351;
wire n_9352;
wire n_2746;
wire n_389;
wire n_7608;
wire n_17053;
wire n_15567;
wire n_6832;
wire n_7394;
wire n_13202;
wire n_15350;
wire n_13638;
wire n_4171;
wire n_17948;
wire n_14392;
wire n_19347;
wire n_7027;
wire n_1105;
wire n_7992;
wire n_6912;
wire n_10330;
wire n_1461;
wire n_8276;
wire n_2076;
wire n_3567;
wire n_11465;
wire n_8027;
wire n_4705;
wire n_3807;
wire n_17808;
wire n_11265;
wire n_11125;
wire n_1114;
wire n_17244;
wire n_7783;
wire n_13220;
wire n_10276;
wire n_191;
wire n_8978;
wire n_10594;
wire n_8245;
wire n_15072;
wire n_12910;
wire n_18725;
wire n_18215;
wire n_8454;
wire n_2881;
wire n_1116;
wire n_8891;
wire n_1219;
wire n_11690;
wire n_18719;
wire n_19142;
wire n_16194;
wire n_3897;
wire n_5591;
wire n_11373;
wire n_3372;
wire n_6403;
wire n_7947;
wire n_1221;
wire n_16826;
wire n_6491;
wire n_19519;
wire n_16321;
wire n_14072;
wire n_17120;
wire n_11412;
wire n_13039;
wire n_13130;
wire n_10441;
wire n_19500;
wire n_17237;
wire n_5518;
wire n_15671;
wire n_9124;
wire n_6661;
wire n_13719;
wire n_8847;
wire n_14548;
wire n_19099;
wire n_4068;
wire n_10841;
wire n_16076;
wire n_12313;
wire n_18071;
wire n_2743;
wire n_4766;
wire n_14661;
wire n_8356;
wire n_6136;
wire n_16384;
wire n_16416;
wire n_3378;
wire n_15305;
wire n_15588;
wire n_3745;
wire n_8888;
wire n_11810;
wire n_14267;
wire n_5357;
wire n_3523;
wire n_2222;
wire n_13062;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_14130;
wire n_14930;
wire n_5541;
wire n_10576;
wire n_16596;
wire n_334;
wire n_6668;
wire n_2999;
wire n_15548;
wire n_1239;
wire n_3697;
wire n_16714;
wire n_19168;
wire n_2408;
wire n_6859;
wire n_18752;
wire n_13752;
wire n_10237;
wire n_19484;
wire n_13596;
wire n_12889;
wire n_18092;
wire n_12050;
wire n_12922;
wire n_12250;
wire n_9515;
wire n_6971;
wire n_17957;
wire n_9642;
wire n_393;
wire n_14231;
wire n_12385;
wire n_13219;
wire n_5673;
wire n_5443;
wire n_17449;
wire n_6351;
wire n_9382;
wire n_16392;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_19207;
wire n_13295;
wire n_3936;
wire n_1349;
wire n_16906;
wire n_18194;
wire n_17693;
wire n_6829;
wire n_2723;
wire n_17981;
wire n_3496;
wire n_13160;
wire n_15249;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_17337;
wire n_10708;
wire n_13818;
wire n_15024;
wire n_8803;
wire n_3239;
wire n_4062;
wire n_3902;
wire n_18478;
wire n_4396;
wire n_9706;
wire n_3101;
wire n_15174;
wire n_17904;
wire n_3374;
wire n_10387;
wire n_13764;
wire n_19408;
wire n_1552;
wire n_11224;
wire n_8790;
wire n_15569;
wire n_4293;
wire n_10219;
wire n_1031;
wire n_11924;
wire n_15193;
wire n_9591;
wire n_6137;
wire n_14833;
wire n_10364;
wire n_11422;
wire n_8338;
wire n_4412;
wire n_14480;
wire n_12489;
wire n_8491;
wire n_2217;
wire n_4781;
wire n_16610;
wire n_9283;
wire n_19299;
wire n_12030;
wire n_206;
wire n_633;
wire n_12565;
wire n_15236;
wire n_1040;
wire n_3059;
wire n_14098;
wire n_14482;
wire n_9468;
wire n_17174;
wire n_14223;
wire n_15962;
wire n_5424;
wire n_12415;
wire n_3017;
wire n_1805;
wire n_17332;
wire n_10559;
wire n_13173;
wire n_15355;
wire n_15945;
wire n_14848;
wire n_18548;
wire n_7154;
wire n_16232;
wire n_8304;
wire n_19644;
wire n_19012;
wire n_11418;
wire n_6655;
wire n_19187;
wire n_3274;
wire n_9958;
wire n_14544;
wire n_4457;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_16122;
wire n_722;
wire n_5613;
wire n_18852;
wire n_14604;
wire n_14735;
wire n_2223;
wire n_1621;
wire n_19572;
wire n_13101;
wire n_6786;
wire n_8315;
wire n_16446;
wire n_15885;
wire n_17528;
wire n_18964;
wire n_11040;
wire n_11754;
wire n_14916;
wire n_9756;
wire n_4762;
wire n_192;
wire n_13748;
wire n_11672;
wire n_3113;
wire n_10353;
wire n_10847;
wire n_10451;
wire n_1458;
wire n_15801;
wire n_17778;
wire n_5303;
wire n_12240;
wire n_12003;
wire n_7496;
wire n_223;
wire n_4154;
wire n_12165;
wire n_10866;
wire n_18127;
wire n_9940;
wire n_6200;
wire n_4504;
wire n_14600;
wire n_3844;
wire n_1237;
wire n_11763;
wire n_15010;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_18730;
wire n_10653;
wire n_8535;
wire n_11587;
wire n_6373;
wire n_12280;
wire n_13461;
wire n_12492;
wire n_19535;
wire n_16282;
wire n_17011;
wire n_2243;
wire n_4898;
wire n_5601;
wire n_13188;
wire n_4819;
wire n_17639;
wire n_7131;
wire n_9586;
wire n_8909;
wire n_3332;
wire n_18977;
wire n_16356;
wire n_11843;
wire n_2570;
wire n_14614;
wire n_4645;
wire n_11629;
wire n_15147;
wire n_9554;
wire n_18246;
wire n_5635;
wire n_17180;
wire n_5091;
wire n_6546;
wire n_4302;
wire n_15927;
wire n_3395;
wire n_7060;
wire n_19439;
wire n_13217;
wire n_5363;
wire n_4178;
wire n_5165;
wire n_16332;
wire n_1711;
wire n_14397;
wire n_17971;
wire n_10853;
wire n_13802;
wire n_18559;
wire n_7761;
wire n_10338;
wire n_12978;
wire n_1422;
wire n_15668;
wire n_15137;
wire n_8496;
wire n_1842;
wire n_12476;
wire n_8568;
wire n_516;
wire n_8852;
wire n_18423;
wire n_12023;
wire n_17655;
wire n_8637;
wire n_2703;
wire n_6168;
wire n_16225;
wire n_16677;
wire n_4606;
wire n_13413;
wire n_6450;
wire n_15153;
wire n_13203;
wire n_2058;
wire n_2660;
wire n_19128;
wire n_14462;
wire n_8456;
wire n_4962;
wire n_4563;
wire n_7137;
wire n_14933;
wire n_5056;
wire n_9920;
wire n_12598;
wire n_9039;
wire n_11854;
wire n_8573;
wire n_2124;
wire n_19070;
wire n_5336;
wire n_5447;
wire n_18623;
wire n_17389;
wire n_7743;
wire n_13230;
wire n_6179;
wire n_19230;
wire n_9125;
wire n_9139;
wire n_17941;
wire n_5747;
wire n_12733;
wire n_13750;
wire n_8775;
wire n_14104;
wire n_808;
wire n_18695;
wire n_14684;
wire n_5753;
wire n_12245;
wire n_15713;
wire n_1193;
wire n_18124;
wire n_14572;
wire n_9972;
wire n_6083;
wire n_12909;
wire n_6434;
wire n_551;
wire n_9157;
wire n_16417;
wire n_3884;
wire n_17880;
wire n_9324;
wire n_5808;
wire n_8807;
wire n_6933;
wire n_8521;
wire n_6547;
wire n_5193;
wire n_9442;
wire n_1481;
wire n_19374;
wire n_6984;
wire n_18394;
wire n_17392;
wire n_10763;
wire n_9957;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_17586;
wire n_5961;
wire n_18757;
wire n_6507;
wire n_9313;
wire n_6687;
wire n_9173;
wire n_6690;
wire n_7412;
wire n_12144;
wire n_9160;
wire n_219;
wire n_9974;
wire n_19365;
wire n_12129;
wire n_14753;
wire n_13658;
wire n_5533;
wire n_14671;
wire n_4257;
wire n_16454;
wire n_17977;
wire n_18441;
wire n_13572;
wire n_15547;
wire n_12032;
wire n_4720;
wire n_14674;
wire n_3857;
wire n_243;
wire n_1873;
wire n_19496;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_12835;
wire n_10129;
wire n_16089;
wire n_1330;
wire n_7523;
wire n_8654;
wire n_2876;
wire n_14229;
wire n_15060;
wire n_11241;
wire n_15520;
wire n_5953;
wire n_14188;
wire n_11508;
wire n_7141;
wire n_5198;
wire n_16139;
wire n_5718;
wire n_6505;
wire n_1663;
wire n_12636;
wire n_4172;
wire n_3403;
wire n_11227;
wire n_1107;
wire n_3294;
wire n_6001;
wire n_11218;
wire n_4502;
wire n_318;
wire n_10195;
wire n_13722;
wire n_3490;
wire n_4849;
wire n_277;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_12938;
wire n_13057;
wire n_8367;
wire n_7367;
wire n_3581;
wire n_16439;
wire n_6023;
wire n_14897;
wire n_19251;
wire n_12173;
wire n_6905;
wire n_17520;
wire n_15925;
wire n_18255;
wire n_19275;
wire n_7368;
wire n_429;
wire n_5553;
wire n_8011;
wire n_4066;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_15141;
wire n_12411;
wire n_10280;
wire n_4004;
wire n_5404;
wire n_18634;
wire n_4292;
wire n_8570;
wire n_6163;
wire n_7628;
wire n_9074;
wire n_5549;
wire n_9408;
wire n_267;
wire n_6553;
wire n_1124;
wire n_1624;
wire n_19190;
wire n_12568;
wire n_3280;
wire n_16163;
wire n_13478;
wire n_18256;
wire n_12970;
wire n_1515;
wire n_8902;
wire n_14295;
wire n_7557;
wire n_593;
wire n_7128;
wire n_14367;
wire n_637;
wire n_13915;
wire n_7594;
wire n_15057;
wire n_19479;
wire n_16300;
wire n_19236;
wire n_18288;
wire n_10504;
wire n_2525;
wire n_7788;
wire n_13783;
wire n_5154;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_3889;
wire n_2687;
wire n_2887;
wire n_2194;
wire n_5637;
wire n_1987;
wire n_7586;
wire n_968;
wire n_7767;
wire n_8294;
wire n_12279;
wire n_9419;
wire n_16402;
wire n_13705;
wire n_17986;
wire n_17771;
wire n_9277;
wire n_9257;
wire n_17773;
wire n_2391;
wire n_2431;
wire n_17070;
wire n_5843;
wire n_9159;
wire n_8170;
wire n_11558;
wire n_18515;
wire n_7744;
wire n_10595;
wire n_7748;
wire n_6827;
wire n_18914;
wire n_11073;
wire n_1208;
wire n_1072;
wire n_815;
wire n_7485;
wire n_18867;
wire n_11974;
wire n_12881;
wire n_15736;
wire n_14986;
wire n_14920;
wire n_8671;
wire n_19196;
wire n_15313;
wire n_284;
wire n_3436;
wire n_9671;
wire n_1026;
wire n_289;
wire n_14994;
wire n_10080;
wire n_16505;
wire n_12228;
wire n_10570;
wire n_16120;
wire n_12929;
wire n_16065;
wire n_685;
wire n_3240;
wire n_15075;
wire n_12261;
wire n_18007;
wire n_12106;
wire n_5333;
wire n_5594;
wire n_12291;
wire n_14510;
wire n_12124;
wire n_11755;
wire n_9510;
wire n_18055;
wire n_13497;
wire n_15406;
wire n_19529;
wire n_14396;
wire n_2517;
wire n_2713;
wire n_11918;
wire n_11748;
wire n_12433;
wire n_5000;
wire n_5551;
wire n_8701;
wire n_16810;
wire n_6499;
wire n_18158;
wire n_12217;
wire n_15922;
wire n_12097;
wire n_5257;
wire n_8097;
wire n_13851;
wire n_9679;
wire n_8645;
wire n_13272;
wire n_18954;
wire n_4688;
wire n_4058;
wire n_3082;
wire n_4848;
wire n_16411;
wire n_19507;
wire n_156;
wire n_16717;
wire n_8824;
wire n_11673;
wire n_2407;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_6276;
wire n_10499;
wire n_8340;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_2667;
wire n_18425;
wire n_1571;
wire n_2948;
wire n_8455;
wire n_7208;
wire n_13613;
wire n_947;
wire n_12185;
wire n_9770;
wire n_1992;
wire n_11417;
wire n_7406;
wire n_8681;
wire n_16044;
wire n_18656;
wire n_3140;
wire n_4749;
wire n_9592;
wire n_5155;
wire n_17507;
wire n_9180;
wire n_10922;
wire n_926;
wire n_19013;
wire n_10718;
wire n_1698;
wire n_4100;
wire n_13821;
wire n_19198;
wire n_13712;
wire n_9625;
wire n_777;
wire n_15041;
wire n_4085;
wire n_15393;
wire n_4464;
wire n_14144;
wire n_6851;
wire n_6460;
wire n_19429;
wire n_4659;
wire n_5217;
wire n_6650;
wire n_8221;
wire n_11682;
wire n_15595;
wire n_8255;
wire n_15081;
wire n_8461;
wire n_6368;
wire n_1857;
wire n_16474;
wire n_6583;
wire n_4889;
wire n_4866;
wire n_3638;
wire n_16940;
wire n_4816;
wire n_17419;
wire n_12520;
wire n_2110;
wire n_1659;
wire n_3393;
wire n_17134;
wire n_3451;
wire n_11459;
wire n_4937;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_12436;
wire n_8792;
wire n_16344;
wire n_2053;
wire n_12808;
wire n_4222;
wire n_18275;
wire n_2710;
wire n_6064;
wire n_1966;
wire n_13801;
wire n_5793;
wire n_19286;
wire n_8523;
wire n_12143;
wire n_4976;
wire n_13879;
wire n_5578;
wire n_18064;
wire n_231;
wire n_1457;
wire n_1993;
wire n_11806;
wire n_2617;
wire n_1466;
wire n_11050;
wire n_5207;
wire n_17714;
wire n_5676;
wire n_1893;
wire n_4665;
wire n_11484;
wire n_2387;
wire n_19483;
wire n_2846;
wire n_19183;
wire n_10295;
wire n_1980;
wire n_5464;
wire n_2237;
wire n_10336;
wire n_4362;
wire n_7716;
wire n_17903;
wire n_8954;
wire n_12212;
wire n_7540;
wire n_775;
wire n_13231;
wire n_12624;
wire n_1531;
wire n_453;
wire n_8552;
wire n_17412;
wire n_7558;
wire n_4261;
wire n_8373;
wire n_13165;
wire n_426;
wire n_3986;
wire n_12151;
wire n_17407;
wire n_15204;
wire n_2556;
wire n_4747;
wire n_5251;
wire n_18284;
wire n_9970;
wire n_11365;
wire n_18138;
wire n_3175;
wire n_17016;
wire n_16081;
wire n_5475;
wire n_15341;
wire n_4448;
wire n_1096;
wire n_15477;
wire n_6233;
wire n_6377;
wire n_12402;
wire n_17959;
wire n_18782;
wire n_688;
wire n_1077;
wire n_4132;
wire n_10361;
wire n_1437;
wire n_7143;
wire n_10424;
wire n_8965;
wire n_4355;
wire n_18454;
wire n_2276;
wire n_13476;
wire n_2803;
wire n_379;
wire n_18399;
wire n_12162;
wire n_3202;
wire n_602;
wire n_17087;
wire n_7497;
wire n_4655;
wire n_11829;
wire n_11517;
wire n_7793;
wire n_16102;
wire n_587;
wire n_16274;
wire n_3554;
wire n_6991;
wire n_10556;
wire n_13776;
wire n_7248;
wire n_7204;
wire n_15835;
wire n_12852;
wire n_10567;
wire n_7578;
wire n_3462;
wire n_13343;
wire n_7654;
wire n_5132;
wire n_17339;
wire n_10230;
wire n_12675;
wire n_5627;
wire n_5774;
wire n_13907;
wire n_4846;
wire n_2984;
wire n_5187;
wire n_12821;
wire n_14782;
wire n_4024;
wire n_18756;
wire n_7120;
wire n_6335;
wire n_8728;
wire n_12837;
wire n_8386;
wire n_14070;
wire n_14330;
wire n_13491;
wire n_4860;
wire n_18654;
wire n_15748;
wire n_3414;
wire n_17995;
wire n_14235;
wire n_6173;
wire n_14851;
wire n_18012;
wire n_10058;
wire n_16471;
wire n_2563;
wire n_19434;
wire n_4989;
wire n_7757;
wire n_1683;
wire n_17539;
wire n_280;
wire n_6630;
wire n_1187;
wire n_4558;
wire n_16560;
wire n_8396;
wire n_6612;
wire n_6606;
wire n_13450;
wire n_3550;
wire n_19533;
wire n_14178;
wire n_5508;
wire n_12907;
wire n_15500;
wire n_14891;
wire n_17051;
wire n_11917;
wire n_6158;
wire n_9318;
wire n_9028;
wire n_17217;
wire n_4328;
wire n_8020;
wire n_1057;
wire n_9374;
wire n_2785;
wire n_2636;
wire n_13634;
wire n_18027;
wire n_10413;
wire n_3399;
wire n_19268;
wire n_1611;
wire n_2740;
wire n_17786;
wire n_4808;
wire n_5767;
wire n_1589;
wire n_12708;
wire n_4712;
wire n_10369;
wire n_2309;
wire n_6821;
wire n_5462;
wire n_9983;
wire n_6688;
wire n_8580;
wire n_9993;
wire n_3533;
wire n_13622;
wire n_4725;
wire n_11207;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3132;
wire n_16951;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_14794;
wire n_17684;
wire n_9237;
wire n_13931;
wire n_14404;
wire n_6557;
wire n_18302;
wire n_6753;
wire n_18164;
wire n_17151;
wire n_7341;
wire n_4908;
wire n_12088;
wire n_15423;
wire n_14377;
wire n_6639;
wire n_12508;
wire n_12096;
wire n_5150;
wire n_8832;
wire n_3819;
wire n_2050;
wire n_19412;
wire n_19399;
wire n_2164;
wire n_11098;
wire n_15815;
wire n_5179;
wire n_7957;
wire n_10938;
wire n_6627;
wire n_17147;
wire n_3544;
wire n_2904;
wire n_18019;
wire n_10927;
wire n_4616;
wire n_4982;
wire n_370;
wire n_8592;
wire n_11204;
wire n_6190;
wire n_1979;
wire n_2738;
wire n_16920;
wire n_12701;
wire n_10578;
wire n_4323;
wire n_16199;
wire n_19113;
wire n_6615;
wire n_17331;
wire n_2342;
wire n_2167;
wire n_7294;
wire n_4017;
wire n_11811;
wire n_13745;
wire n_10569;
wire n_2541;
wire n_8622;
wire n_2940;
wire n_4739;
wire n_15367;
wire n_19095;
wire n_8104;
wire n_2768;
wire n_18511;
wire n_17428;
wire n_4298;
wire n_2314;
wire n_10746;
wire n_9188;
wire n_16407;
wire n_18009;
wire n_4644;
wire n_19002;
wire n_8779;
wire n_5503;
wire n_5945;
wire n_11714;
wire n_10697;
wire n_16179;
wire n_2390;
wire n_15070;
wire n_1343;
wire n_2734;
wire n_7250;
wire n_8762;
wire n_17503;
wire n_18365;
wire n_17358;
wire n_1900;
wire n_3381;
wire n_13419;
wire n_9207;
wire n_11860;
wire n_17057;
wire n_10926;
wire n_8897;
wire n_11503;
wire n_17104;
wire n_4672;
wire n_8376;
wire n_18271;
wire n_2939;
wire n_18998;
wire n_5749;
wire n_1672;
wire n_15640;
wire n_6271;
wire n_15683;
wire n_16202;
wire n_4598;
wire n_8599;
wire n_13460;
wire n_15451;
wire n_5993;
wire n_15233;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_9418;
wire n_8616;
wire n_13105;
wire n_14467;
wire n_14789;
wire n_13076;
wire n_15526;
wire n_12950;
wire n_8628;
wire n_15150;
wire n_13028;
wire n_8547;
wire n_4424;
wire n_7113;
wire n_1751;
wire n_10433;
wire n_285;
wire n_9116;
wire n_14096;
wire n_11983;
wire n_10839;
wire n_11813;
wire n_3506;
wire n_1928;
wire n_14583;
wire n_4317;
wire n_14893;
wire n_8275;
wire n_6198;
wire n_5418;
wire n_18270;
wire n_6762;
wire n_4088;
wire n_3711;
wire n_9035;
wire n_729;
wire n_16960;
wire n_3642;
wire n_14915;
wire n_4650;
wire n_17780;
wire n_438;
wire n_17075;
wire n_2874;
wire n_1200;
wire n_4967;
wire n_9678;
wire n_8247;
wire n_6577;
wire n_12956;
wire n_17373;
wire n_14856;
wire n_15235;
wire n_4912;
wire n_9284;
wire n_5086;
wire n_4735;
wire n_187;
wire n_3300;
wire n_2978;
wire n_15711;
wire n_1050;
wire n_5170;
wire n_7604;
wire n_3515;
wire n_1150;
wire n_9606;
wire n_17018;
wire n_13459;
wire n_1023;
wire n_1118;
wire n_14268;
wire n_194;
wire n_2949;
wire n_10297;
wire n_12553;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_14127;
wire n_440;
wire n_3806;
wire n_8827;
wire n_2931;
wire n_3866;
wire n_17937;
wire n_9549;
wire n_14894;
wire n_12866;
wire n_17801;
wire n_4157;
wire n_6845;
wire n_9482;
wire n_3629;
wire n_969;
wire n_8877;
wire n_9412;
wire n_15561;
wire n_6321;
wire n_6819;
wire n_10136;
wire n_15148;
wire n_16457;
wire n_19560;
wire n_11356;
wire n_1379;
wire n_15955;
wire n_214;
wire n_8688;
wire n_4910;
wire n_3083;
wire n_10692;
wire n_14826;
wire n_16421;
wire n_15776;
wire n_11280;
wire n_14987;
wire n_8686;
wire n_12239;
wire n_17641;
wire n_3830;
wire n_8403;
wire n_11493;
wire n_17742;
wire n_3117;
wire n_8588;
wire n_15229;
wire n_11339;
wire n_15804;
wire n_5623;
wire n_15269;
wire n_10471;
wire n_2385;
wire n_4112;
wire n_3739;
wire n_14946;
wire n_18727;
wire n_15674;
wire n_4352;
wire n_17933;
wire n_8780;
wire n_17384;
wire n_7958;
wire n_18037;
wire n_4980;
wire n_11885;
wire n_1924;
wire n_15855;
wire n_3363;
wire n_10777;
wire n_3721;
wire n_16490;
wire n_7760;
wire n_13306;
wire n_9753;
wire n_8722;
wire n_16489;
wire n_19580;
wire n_8589;
wire n_3969;
wire n_7573;
wire n_6281;
wire n_7364;
wire n_5647;
wire n_13133;
wire n_4256;
wire n_4938;
wire n_8608;
wire n_12874;
wire n_11194;
wire n_10469;
wire n_11480;
wire n_445;
wire n_18650;
wire n_930;
wire n_9342;
wire n_18062;
wire n_2620;
wire n_9329;
wire n_1945;
wire n_5426;
wire n_19257;
wire n_17119;
wire n_9868;
wire n_1414;
wire n_7048;
wire n_944;
wire n_16491;
wire n_2744;
wire n_1011;
wire n_1566;
wire n_8145;
wire n_8928;
wire n_17638;
wire n_7682;
wire n_990;
wire n_18584;
wire n_12509;
wire n_6231;
wire n_14902;
wire n_6932;
wire n_13527;
wire n_7901;
wire n_870;
wire n_366;
wire n_5709;
wire n_7658;
wire n_10055;
wire n_10979;
wire n_3802;
wire n_6996;
wire n_15935;
wire n_17674;
wire n_376;
wire n_2111;
wire n_10408;
wire n_16180;
wire n_8572;
wire n_17182;
wire n_6337;
wire n_18212;
wire n_3643;
wire n_2425;
wire n_12936;
wire n_8227;
wire n_18424;
wire n_3060;
wire n_10482;
wire n_4105;
wire n_7405;
wire n_14151;
wire n_4926;
wire n_1518;
wire n_8314;
wire n_9386;
wire n_15120;
wire n_11121;
wire n_3038;
wire n_11270;
wire n_6310;
wire n_11689;
wire n_10003;
wire n_15601;
wire n_15936;
wire n_10321;
wire n_5310;
wire n_9661;
wire n_14284;
wire n_3863;
wire n_5722;
wire n_4640;
wire n_13232;
wire n_13001;
wire n_17377;
wire n_9901;
wire n_17334;
wire n_2805;
wire n_5593;
wire n_4769;
wire n_8934;
wire n_13059;
wire n_6365;
wire n_4628;
wire n_8407;
wire n_8567;
wire n_15455;
wire n_11288;
wire n_12772;
wire n_5237;
wire n_409;
wire n_11042;
wire n_10726;
wire n_16534;
wire n_19304;
wire n_4460;
wire n_4108;
wire n_14681;
wire n_11272;
wire n_14230;
wire n_5853;
wire n_8283;
wire n_5011;
wire n_14546;
wire n_9882;
wire n_16484;
wire n_10637;
wire n_9205;
wire n_17464;
wire n_7972;
wire n_1675;
wire n_13512;
wire n_7916;
wire n_9368;
wire n_13069;
wire n_12362;
wire n_19038;
wire n_6167;
wire n_13233;
wire n_18495;
wire n_8008;
wire n_18833;
wire n_13297;
wire n_2553;
wire n_6307;
wire n_149;
wire n_632;
wire n_2038;
wire n_7483;
wire n_14873;
wire n_9504;
wire n_14840;
wire n_16556;
wire n_6267;
wire n_5998;
wire n_17861;
wire n_6568;
wire n_19083;
wire n_7507;
wire n_7159;
wire n_18038;
wire n_6028;
wire n_1417;
wire n_16072;
wire n_14083;
wire n_681;
wire n_10189;
wire n_8697;
wire n_6813;
wire n_6669;
wire n_422;
wire n_8420;
wire n_8297;
wire n_3079;
wire n_10881;
wire n_13519;
wire n_16583;
wire n_15641;
wire n_16007;
wire n_17129;
wire n_4853;
wire n_8639;
wire n_16796;
wire n_16510;
wire n_531;
wire n_15892;
wire n_4272;
wire n_14049;
wire n_1025;
wire n_7562;
wire n_3111;
wire n_336;
wire n_12019;
wire n_8176;
wire n_14529;
wire n_17624;
wire n_16106;
wire n_10891;
wire n_9026;
wire n_10803;
wire n_13190;
wire n_6188;
wire n_5262;
wire n_4670;
wire n_4882;
wire n_11695;
wire n_17595;
wire n_4738;
wire n_8113;
wire n_18922;
wire n_15877;
wire n_1307;
wire n_11453;
wire n_19233;
wire n_17896;
wire n_19088;
wire n_5713;
wire n_16445;
wire n_168;
wire n_6318;
wire n_2353;
wire n_16997;
wire n_4099;
wire n_14690;
wire n_19252;
wire n_17356;
wire n_1738;
wire n_10290;
wire n_11862;
wire n_14839;
wire n_15409;
wire n_16207;
wire n_9433;
wire n_18568;
wire n_11660;
wire n_14249;
wire n_14241;
wire n_6604;
wire n_2386;
wire n_5373;
wire n_1724;
wire n_16101;
wire n_3708;
wire n_6391;
wire n_10284;
wire n_14446;
wire n_14719;
wire n_15575;
wire n_8522;
wire n_12971;
wire n_7942;
wire n_16599;
wire n_6473;
wire n_18620;
wire n_15696;
wire n_14558;
wire n_11318;
wire n_17198;
wire n_7725;
wire n_16950;
wire n_8626;
wire n_1393;
wire n_1867;
wire n_1603;
wire n_19277;
wire n_5466;
wire n_19475;
wire n_15095;
wire n_5955;
wire n_658;
wire n_1874;
wire n_11487;
wire n_2825;
wire n_8441;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_7778;
wire n_758;
wire n_2256;
wire n_4060;
wire n_8397;
wire n_5796;
wire n_17916;
wire n_8726;
wire n_17250;
wire n_770;
wire n_6958;
wire n_15417;
wire n_16615;
wire n_14667;
wire n_6523;
wire n_14713;
wire n_4687;
wire n_7531;
wire n_18686;
wire n_1404;
wire n_13214;
wire n_8615;
wire n_15975;
wire n_11062;
wire n_14202;
wire n_15859;
wire n_11933;
wire n_14554;
wire n_9887;
wire n_4600;
wire n_13211;
wire n_8316;
wire n_5829;
wire n_19654;
wire n_8057;
wire n_5191;
wire n_1231;
wire n_14874;
wire n_18198;
wire n_2370;
wire n_18550;
wire n_4253;
wire n_407;
wire n_913;
wire n_16824;
wire n_15098;
wire n_867;
wire n_16832;
wire n_13336;
wire n_1333;
wire n_2496;
wire n_16074;
wire n_3189;
wire n_19487;
wire n_18664;
wire n_13102;
wire n_4691;
wire n_12894;
wire n_10492;
wire n_15769;
wire n_4297;
wire n_9247;
wire n_17340;
wire n_8378;
wire n_2907;
wire n_577;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_9570;
wire n_5675;
wire n_12356;
wire n_2778;
wire n_19454;
wire n_11077;
wire n_1909;
wire n_5020;
wire n_9846;
wire n_13262;
wire n_1123;
wire n_10764;
wire n_18005;
wire n_18429;
wire n_9677;
wire n_3934;
wire n_4033;
wire n_6804;
wire n_6603;
wire n_17812;
wire n_3193;
wire n_7534;
wire n_8201;
wire n_4354;
wire n_16485;
wire n_14262;
wire n_9348;
wire n_1530;
wire n_8696;
wire n_938;
wire n_6396;
wire n_12630;
wire n_6890;
wire n_549;
wire n_4377;
wire n_12022;
wire n_905;
wire n_10741;
wire n_6109;
wire n_14727;
wire n_12425;
wire n_14762;
wire n_322;
wire n_689;
wire n_13507;
wire n_10915;
wire n_18290;
wire n_558;
wire n_3036;
wire n_7943;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_17133;
wire n_17729;
wire n_15410;
wire n_4511;
wire n_2908;
wire n_9707;
wire n_16002;
wire n_16258;
wire n_13594;
wire n_10680;
wire n_3599;
wire n_5543;
wire n_5885;
wire n_14228;
wire n_5356;
wire n_3772;
wire n_5458;
wire n_16131;
wire n_11473;
wire n_5038;
wire n_1760;
wire n_4585;
wire n_2664;
wire n_1722;
wire n_11726;
wire n_15944;
wire n_12574;
wire n_8833;
wire n_10142;
wire n_7828;
wire n_9918;
wire n_18643;
wire n_15932;
wire n_16345;
wire n_4427;
wire n_9390;
wire n_10069;
wire n_17325;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_2804;
wire n_2453;
wire n_18233;
wire n_5510;
wire n_5555;
wire n_13678;
wire n_12458;
wire n_19291;
wire n_6066;
wire n_14582;
wire n_6897;
wire n_13523;
wire n_9619;
wire n_11171;
wire n_15117;
wire n_4886;
wire n_9187;
wire n_2733;
wire n_16621;
wire n_13819;
wire n_15777;
wire n_14424;
wire n_18398;
wire n_14523;
wire n_11063;
wire n_18846;
wire n_9989;
wire n_8319;
wire n_4200;
wire n_3460;
wire n_12853;
wire n_12942;
wire n_9259;
wire n_3519;
wire n_12397;
wire n_16555;
wire n_15336;
wire n_14161;
wire n_6573;
wire n_16760;
wire n_7634;
wire n_5078;
wire n_13290;
wire n_13500;
wire n_11440;
wire n_16844;
wire n_10483;
wire n_17758;
wire n_4737;
wire n_4116;
wire n_7285;
wire n_11337;
wire n_12005;
wire n_11243;
wire n_8929;
wire n_9360;
wire n_18610;
wire n_9824;
wire n_342;
wire n_15089;
wire n_2658;
wire n_2665;
wire n_8233;
wire n_6130;
wire n_7273;
wire n_14750;
wire n_17939;
wire n_5976;
wire n_14074;
wire n_840;
wire n_2913;
wire n_12800;
wire n_2230;
wire n_1969;
wire n_1565;
wire n_16574;
wire n_15145;
wire n_17516;
wire n_8187;
wire n_9399;
wire n_15838;
wire n_15297;
wire n_13979;
wire n_9740;
wire n_615;
wire n_12947;
wire n_5371;
wire n_4651;
wire n_17178;
wire n_9764;
wire n_4854;
wire n_15160;
wire n_3789;
wire n_605;
wire n_12354;
wire n_7597;
wire n_12666;
wire n_14297;
wire n_17388;
wire n_16368;
wire n_12631;
wire n_1646;
wire n_19154;
wire n_14969;
wire n_14820;
wire n_10133;
wire n_18426;
wire n_18073;
wire n_6921;
wire n_14675;
wire n_18905;
wire n_9826;
wire n_3171;
wire n_3608;
wire n_11942;
wire n_15998;
wire n_3459;
wire n_19138;
wire n_6624;
wire n_6956;
wire n_12966;
wire n_15851;
wire n_15884;
wire n_5656;
wire n_5125;
wire n_7329;
wire n_14502;
wire n_14533;
wire n_5652;
wire n_17935;
wire n_10752;
wire n_18630;
wire n_10067;
wire n_18021;
wire n_10399;
wire n_12498;
wire n_656;
wire n_11010;
wire n_9590;
wire n_16017;
wire n_2717;
wire n_11588;
wire n_16346;
wire n_738;
wire n_13956;
wire n_3497;
wire n_7418;
wire n_6880;
wire n_19305;
wire n_3580;
wire n_12387;
wire n_9497;
wire n_13255;
wire n_15911;
wire n_2307;
wire n_3704;
wire n_684;
wire n_9219;
wire n_17376;
wire n_8028;
wire n_4280;
wire n_8914;
wire n_1181;
wire n_15276;
wire n_8391;
wire n_16343;
wire n_13749;
wire n_15552;
wire n_17722;
wire n_19370;
wire n_16228;
wire n_803;
wire n_1817;
wire n_12862;
wire n_13621;
wire n_8216;
wire n_2868;
wire n_16953;
wire n_2231;
wire n_3609;
wire n_9982;
wire n_7804;
wire n_18948;
wire n_12656;
wire n_8313;
wire n_14828;
wire n_7656;
wire n_19150;
wire n_8263;
wire n_6438;
wire n_11936;
wire n_19132;
wire n_10374;
wire n_7332;
wire n_10382;
wire n_18247;
wire n_4455;
wire n_8374;
wire n_13223;
wire n_13451;
wire n_4514;
wire n_13939;
wire n_18909;
wire n_13728;
wire n_4806;
wire n_7386;
wire n_17824;
wire n_11018;
wire n_10981;
wire n_16014;
wire n_2682;
wire n_13379;
wire n_13781;
wire n_19311;
wire n_5098;
wire n_17513;
wire n_10344;
wire n_5707;
wire n_14613;
wire n_19451;
wire n_11515;
wire n_17466;
wire n_3505;
wire n_15881;
wire n_7637;
wire n_16577;
wire n_10318;
wire n_4796;
wire n_4442;
wire n_18422;
wire n_2581;
wire n_18091;
wire n_12890;
wire n_3590;
wire n_5344;
wire n_954;
wire n_13994;
wire n_4419;
wire n_17060;
wire n_11972;
wire n_13484;
wire n_17298;
wire n_8460;
wire n_3327;
wire n_17468;
wire n_14593;
wire n_2701;
wire n_16013;
wire n_1080;
wire n_7409;
wire n_19266;
wire n_10735;
wire n_17153;
wire n_13807;
wire n_9825;
wire n_2784;
wire n_5494;
wire n_7444;
wire n_16942;
wire n_2421;
wire n_17569;
wire n_4387;
wire n_2618;
wire n_2464;
wire n_5128;
wire n_18661;
wire n_14033;
wire n_2224;
wire n_10393;
wire n_1092;
wire n_15221;
wire n_5467;
wire n_16090;
wire n_18467;
wire n_4890;
wire n_1784;
wire n_9045;
wire n_12281;
wire n_9373;
wire n_14337;
wire n_2929;
wire n_11809;
wire n_17994;
wire n_9967;
wire n_13553;
wire n_4236;
wire n_7187;
wire n_19039;
wire n_17063;
wire n_1831;
wire n_9182;
wire n_5079;
wire n_9365;
wire n_18960;
wire n_10909;
wire n_6336;
wire n_10083;
wire n_18891;
wire n_9224;
wire n_10347;
wire n_6541;
wire n_12410;
wire n_4706;
wire n_16327;
wire n_19238;
wire n_14707;
wire n_16043;
wire n_4622;
wire n_14612;
wire n_12294;
wire n_7603;
wire n_10667;
wire n_2732;
wire n_17688;
wire n_4206;
wire n_2249;
wire n_18794;
wire n_5835;
wire n_7979;
wire n_13382;
wire n_11675;
wire n_15543;
wire n_15906;
wire n_8657;
wire n_8296;
wire n_8006;
wire n_2955;
wire n_11083;
wire n_17418;
wire n_2158;
wire n_7866;
wire n_3367;
wire n_7205;
wire n_18283;
wire n_2202;
wire n_736;
wire n_11728;
wire n_2993;
wire n_4754;
wire n_11698;
wire n_4647;
wire n_9556;
wire n_8590;
wire n_16682;
wire n_4030;
wire n_1995;
wire n_17038;
wire n_15798;
wire n_4760;
wire n_11326;
wire n_6421;
wire n_11870;
wire n_7407;
wire n_6328;
wire n_11283;
wire n_11834;
wire n_6236;
wire n_13361;
wire n_17286;
wire n_4509;
wire n_15061;
wire n_2875;
wire n_1103;
wire n_6144;
wire n_11506;
wire n_13161;
wire n_10135;
wire n_144;
wire n_2219;
wire n_14010;
wire n_16413;
wire n_999;
wire n_4897;
wire n_15030;
wire n_18205;
wire n_9152;
wire n_3539;
wire n_16451;
wire n_19590;
wire n_8364;
wire n_3276;
wire n_15228;
wire n_15832;
wire n_10720;
wire n_10535;
wire n_19349;
wire n_17629;
wire n_17536;
wire n_3886;
wire n_6708;
wire n_11236;
wire n_18793;
wire n_4420;
wire n_892;
wire n_18529;
wire n_6242;
wire n_12379;
wire n_1468;
wire n_2855;
wire n_2156;
wire n_18222;
wire n_12932;
wire n_14078;
wire n_3548;
wire n_18985;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_14222;
wire n_16990;
wire n_3141;
wire n_5096;
wire n_1841;
wire n_12114;
wire n_10308;
wire n_11608;
wire n_14430;
wire n_1015;
wire n_10623;
wire n_4797;
wire n_6285;
wire n_4270;
wire n_16545;
wire n_19339;
wire n_13709;
wire n_4945;
wire n_17713;
wire n_5677;
wire n_9454;
wire n_10586;
wire n_8742;
wire n_12626;
wire n_11967;
wire n_15084;
wire n_9253;
wire n_13559;
wire n_8874;
wire n_5927;
wire n_15071;
wire n_11996;
wire n_9566;
wire n_11338;
wire n_13426;
wire n_1356;
wire n_4333;
wire n_18826;
wire n_7666;
wire n_11250;
wire n_15328;
wire n_1452;
wire n_2854;
wire n_7963;
wire n_6398;
wire n_8329;
wire n_302;
wire n_9503;
wire n_8270;
wire n_16051;
wire n_11738;
wire n_18196;
wire n_3217;
wire n_1983;
wire n_11522;
wire n_7737;
wire n_16569;
wire n_8614;
wire n_18459;
wire n_9568;
wire n_15621;
wire n_18411;
wire n_8816;
wire n_9119;
wire n_19337;
wire n_13529;
wire n_6224;
wire n_3279;
wire n_18293;
wire n_2402;
wire n_1081;
wire n_19616;
wire n_1084;
wire n_6614;
wire n_5912;
wire n_18395;
wire n_3501;
wire n_374;
wire n_12554;
wire n_8035;
wire n_12722;
wire n_6735;
wire n_17445;
wire n_10491;
wire n_921;
wire n_12037;
wire n_15371;
wire n_17572;
wire n_13453;
wire n_15080;
wire n_5265;
wire n_2257;
wire n_9943;
wire n_12391;
wire n_14242;
wire n_15622;
wire n_7152;
wire n_2200;
wire n_9575;
wire n_10409;
wire n_4548;
wire n_11822;
wire n_10521;
wire n_9610;
wire n_16483;
wire n_14016;
wire n_12323;
wire n_15566;
wire n_10527;
wire n_3115;
wire n_7570;
wire n_2084;
wire n_4875;
wire n_7817;
wire n_5682;
wire n_5387;
wire n_654;
wire n_11394;
wire n_2458;
wire n_3050;
wire n_9928;
wire n_11820;
wire n_13897;
wire n_2527;
wire n_14792;
wire n_16290;
wire n_14248;
wire n_8370;
wire n_164;
wire n_13300;
wire n_16296;
wire n_5681;
wire n_7566;
wire n_11940;
wire n_1271;
wire n_4901;
wire n_9217;
wire n_12901;
wire n_4040;
wire n_10518;
wire n_2406;
wire n_7617;
wire n_15170;
wire n_16936;
wire n_19262;
wire n_9771;
wire n_15774;
wire n_5316;
wire n_7718;
wire n_244;
wire n_13844;
wire n_19246;
wire n_7396;
wire n_282;
wire n_18543;
wire n_5703;
wire n_18930;
wire n_833;
wire n_523;
wire n_7998;
wire n_12432;
wire n_7561;
wire n_18349;
wire n_6810;
wire n_2196;
wire n_17010;
wire n_17040;
wire n_16130;
wire n_12879;
wire n_5564;
wire n_13746;
wire n_12559;
wire n_13508;
wire n_14660;
wire n_4530;
wire n_9899;
wire n_13004;
wire n_5406;
wire n_13479;
wire n_8277;
wire n_652;
wire n_18014;
wire n_1906;
wire n_14437;
wire n_4841;
wire n_1758;
wire n_13759;
wire n_5806;
wire n_4338;
wire n_10486;
wire n_306;
wire n_16613;
wire n_8724;
wire n_5738;
wire n_15938;
wire n_17216;
wire n_3151;
wire n_15146;
wire n_3779;
wire n_2388;
wire n_3984;
wire n_9995;
wire n_5710;
wire n_9076;
wire n_12351;
wire n_16360;
wire n_19146;
wire n_13359;
wire n_10372;
wire n_3558;
wire n_14867;
wire n_1984;
wire n_2236;
wire n_6044;
wire n_8867;
wire n_9491;
wire n_4326;
wire n_12702;
wire n_17811;
wire n_15188;
wire n_2834;
wire n_12439;
wire n_19478;
wire n_11008;
wire n_6125;
wire n_7314;
wire n_786;
wire n_14186;
wire n_7526;
wire n_17816;
wire n_5040;
wire n_14023;
wire n_17890;
wire n_10736;
wire n_19550;
wire n_11575;
wire n_7004;
wire n_14418;
wire n_8308;
wire n_18897;
wire n_151;
wire n_8165;
wire n_14283;
wire n_4788;
wire n_8400;
wire n_18177;
wire n_5977;
wire n_10446;
wire n_7879;
wire n_16372;
wire n_1908;
wire n_15958;
wire n_18853;
wire n_7696;
wire n_11570;
wire n_16567;
wire n_12952;
wire n_19096;
wire n_2045;
wire n_14795;
wire n_3687;
wire n_2216;
wire n_19318;
wire n_3621;
wire n_16425;
wire n_16769;
wire n_10603;
wire n_12004;
wire n_8217;
wire n_6962;
wire n_12830;
wire n_8858;
wire n_7246;
wire n_10255;
wire n_2719;
wire n_11490;
wire n_8689;
wire n_10113;
wire n_15086;
wire n_680;
wire n_3339;
wire n_10188;
wire n_6853;
wire n_10686;
wire n_9841;
wire n_8743;
wire n_7087;
wire n_8753;
wire n_6191;
wire n_4741;
wire n_16838;
wire n_10974;
wire n_11067;
wire n_8627;
wire n_13659;
wire n_12034;
wire n_16586;
wire n_1399;
wire n_16056;
wire n_13303;
wire n_6894;
wire n_13346;
wire n_13702;
wire n_9179;
wire n_2358;
wire n_15894;
wire n_8752;
wire n_2186;
wire n_18237;
wire n_3034;
wire n_4408;
wire n_18367;
wire n_10937;
wire n_643;
wire n_12134;
wire n_400;
wire n_12449;
wire n_2814;
wire n_16399;
wire n_789;
wire n_327;
wire n_6284;
wire n_10167;
wire n_12524;
wire n_18113;
wire n_6883;
wire n_12963;
wire n_10428;
wire n_16860;
wire n_17869;
wire n_19199;
wire n_18682;
wire n_12366;
wire n_747;
wire n_14951;
wire n_11068;
wire n_11035;
wire n_5495;
wire n_535;
wire n_19148;
wire n_12729;
wire n_13292;
wire n_12198;
wire n_9420;
wire n_3851;
wire n_16995;
wire n_14336;
wire n_10079;
wire n_7825;
wire n_7212;
wire n_19436;
wire n_6966;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_6035;
wire n_1652;
wire n_15435;
wire n_8634;
wire n_9531;
wire n_12605;
wire n_1258;
wire n_2438;
wire n_6253;
wire n_2914;
wire n_12828;
wire n_10258;
wire n_5786;
wire n_14960;
wire n_8532;
wire n_19109;
wire n_12661;
wire n_10588;
wire n_8991;
wire n_8065;
wire n_3100;
wire n_11140;
wire n_3573;
wire n_17882;
wire n_17677;
wire n_8518;
wire n_197;
wire n_18226;
wire n_13017;
wire n_1083;
wire n_16884;
wire n_15199;
wire n_18153;
wire n_1721;
wire n_9812;
wire n_1737;
wire n_15419;
wire n_752;
wire n_7361;
wire n_9949;
wire n_1028;
wire n_14889;
wire n_7228;
wire n_9576;
wire n_5872;
wire n_1973;
wire n_3181;
wire n_6338;
wire n_15267;
wire n_19366;
wire n_1500;
wire n_3699;
wire n_854;
wire n_4913;
wire n_6266;
wire n_14796;
wire n_2242;
wire n_19125;
wire n_11364;
wire n_12790;
wire n_4266;
wire n_8632;
wire n_2466;
wire n_19069;
wire n_17397;
wire n_7018;
wire n_5873;
wire n_7975;
wire n_10009;
wire n_9279;
wire n_11902;
wire n_924;
wire n_16782;
wire n_11993;
wire n_2318;
wire n_10443;
wire n_3170;
wire n_17317;
wire n_12813;
wire n_13534;
wire n_3304;
wire n_4968;
wire n_10384;
wire n_5085;
wire n_5736;
wire n_2433;
wire n_829;
wire n_7978;
wire n_10293;
wire n_17422;
wire n_12312;
wire n_10074;
wire n_13097;
wire n_17850;
wire n_15786;
wire n_4208;
wire n_9632;
wire n_12256;
wire n_11812;
wire n_9711;
wire n_9431;
wire n_4779;
wire n_14650;
wire n_18068;
wire n_481;
wire n_14610;
wire n_997;
wire n_11505;
wire n_4437;
wire n_7316;
wire n_17938;
wire n_1306;
wire n_3264;
wire n_18955;
wire n_7103;
wire n_14601;
wire n_436;
wire n_11363;
wire n_15794;
wire n_17066;
wire n_2426;
wire n_2478;
wire n_14645;
wire n_1133;
wire n_4642;
wire n_11151;
wire n_15825;
wire n_10716;
wire n_10664;
wire n_2578;
wire n_3709;
wire n_11434;
wire n_3738;
wire n_6873;
wire n_4186;
wire n_8494;
wire n_5812;
wire n_12468;
wire n_9429;
wire n_8544;
wire n_19536;
wire n_4998;
wire n_10749;
wire n_3330;
wire n_8788;
wire n_10992;
wire n_19380;
wire n_1629;
wire n_10160;
wire n_10560;
wire n_7404;
wire n_13171;
wire n_12857;
wire n_18615;
wire n_1260;
wire n_309;
wire n_9854;
wire n_14854;
wire n_812;
wire n_15266;
wire n_1006;
wire n_7271;
wire n_9713;
wire n_16501;
wire n_257;
wire n_19264;
wire n_1311;
wire n_10300;
wire n_9588;
wire n_14218;
wire n_15107;
wire n_6842;
wire n_13876;
wire n_4803;
wire n_18935;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_14487;
wire n_9127;
wire n_5996;
wire n_16767;
wire n_9869;
wire n_315;
wire n_14449;
wire n_17094;
wire n_12885;
wire n_2579;
wire n_15539;
wire n_2105;
wire n_9715;
wire n_17112;
wire n_8618;
wire n_18916;
wire n_3387;
wire n_12108;
wire n_7535;
wire n_11531;
wire n_19450;
wire n_9407;
wire n_2912;
wire n_14476;
wire n_3409;
wire n_15244;
wire n_2320;
wire n_19574;
wire n_11824;
wire n_1259;
wire n_6957;
wire n_9361;
wire n_13976;
wire n_16578;
wire n_18949;
wire n_13579;
wire n_11566;
wire n_17452;
wire n_16650;
wire n_14639;
wire n_8990;
wire n_17067;
wire n_6444;
wire n_19170;
wire n_226;
wire n_7944;
wire n_19235;
wire n_11374;
wire n_8647;
wire n_15857;
wire n_2003;
wire n_7016;
wire n_10782;
wire n_13557;
wire n_3301;
wire n_16709;
wire n_6379;
wire n_15589;
wire n_17491;
wire n_2324;
wire n_17757;
wire n_12754;
wire n_245;
wire n_13583;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_17333;
wire n_19043;
wire n_2847;
wire n_17749;
wire n_16658;
wire n_4050;
wire n_13455;
wire n_883;
wire n_19136;
wire n_6232;
wire n_9132;
wire n_1032;
wire n_10861;
wire n_17035;
wire n_8879;
wire n_1099;
wire n_19639;
wire n_11203;
wire n_16157;
wire n_11159;
wire n_8052;
wire n_2211;
wire n_6362;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_9332;
wire n_17097;
wire n_369;
wire n_16765;
wire n_11030;
wire n_4179;
wire n_1285;
wire n_6326;
wire n_10073;
wire n_14619;
wire n_1590;
wire n_5072;
wire n_7241;
wire n_10419;
wire n_7172;
wire n_3106;
wire n_15427;
wire n_17364;
wire n_10333;
wire n_12430;
wire n_18330;
wire n_7235;
wire n_6239;
wire n_2340;
wire n_13407;
wire n_5896;
wire n_13676;
wire n_18391;
wire n_16694;
wire n_12557;
wire n_13788;
wire n_6974;
wire n_16537;
wire n_18227;
wire n_18666;
wire n_8939;
wire n_13584;
wire n_428;
wire n_15471;
wire n_12139;
wire n_9030;
wire n_7657;
wire n_822;
wire n_2791;
wire n_19433;
wire n_9665;
wire n_5044;
wire n_5134;
wire n_7096;
wire n_3063;
wire n_13327;
wire n_1550;
wire n_19098;
wire n_11197;
wire n_491;
wire n_7442;
wire n_1591;
wire n_3632;
wire n_10093;
wire n_15428;
wire n_15014;
wire n_1344;
wire n_6174;
wire n_2730;
wire n_7999;
wire n_10675;
wire n_6087;
wire n_16311;
wire n_538;
wire n_4164;
wire n_10107;
wire n_3225;
wire n_15536;
wire n_13224;
wire n_11469;
wire n_5022;
wire n_14046;
wire n_7041;
wire n_10742;
wire n_10829;
wire n_19115;
wire n_12389;
wire n_9309;
wire n_19632;
wire n_10620;
wire n_13971;
wire n_16750;
wire n_7672;
wire n_2551;
wire n_5047;
wire n_7318;
wire n_19325;
wire n_12995;
wire n_18261;
wire n_14406;
wire n_13209;
wire n_11883;
wire n_14959;
wire n_3269;
wire n_15387;
wire n_11901;
wire n_6352;
wire n_15973;
wire n_8542;
wire n_10859;
wire n_18446;
wire n_8576;
wire n_14807;
wire n_8038;
wire n_11572;
wire n_5141;
wire n_3603;
wire n_14493;
wire n_18306;
wire n_13113;
wire n_13387;
wire n_8716;
wire n_3822;
wire n_5535;
wire n_19411;
wire n_3812;
wire n_16807;
wire n_18538;
wire n_2696;
wire n_17576;
wire n_4080;
wire n_6002;
wire n_541;
wire n_18665;
wire n_15538;
wire n_2073;
wire n_2273;
wire n_4941;
wire n_5506;
wire n_11399;
wire n_17578;
wire n_8768;
wire n_10884;
wire n_1162;
wire n_15870;
wire n_12035;
wire n_13006;
wire n_12791;
wire n_7600;
wire n_14742;
wire n_2831;
wire n_4158;
wire n_6644;
wire n_17878;
wire n_4795;
wire n_19528;
wire n_12810;
wire n_16930;
wire n_3824;
wire n_13947;
wire n_11322;
wire n_17562;
wire n_4544;
wire n_5841;
wire n_12241;
wire n_9343;
wire n_15895;
wire n_16554;
wire n_17779;
wire n_5108;
wire n_7347;
wire n_11057;
wire n_2355;
wire n_10969;
wire n_14474;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_8863;
wire n_18501;
wire n_7759;
wire n_11551;
wire n_18049;
wire n_7479;
wire n_2866;
wire n_10598;
wire n_8947;
wire n_15494;
wire n_10717;
wire n_11118;
wire n_18579;
wire n_3649;
wire n_2821;
wire n_6067;
wire n_12674;
wire n_17727;
wire n_17839;
wire n_8510;
wire n_11410;
wire n_12230;
wire n_19282;
wire n_1563;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_17122;
wire n_1359;
wire n_5367;
wire n_16778;
wire n_3794;
wire n_12220;
wire n_6868;
wire n_1335;
wire n_5970;
wire n_16133;
wire n_12283;
wire n_7174;
wire n_9421;
wire n_5202;
wire n_19055;
wire n_13383;
wire n_18787;
wire n_17079;
wire n_8021;
wire n_3346;
wire n_7803;
wire n_15124;
wire n_12595;
wire n_11429;
wire n_15802;
wire n_15163;
wire n_13983;
wire n_9416;
wire n_6225;
wire n_5502;
wire n_3428;
wire n_4552;
wire n_6218;
wire n_17489;
wire n_9929;
wire n_13317;
wire n_12920;
wire n_2519;
wire n_9953;
wire n_1063;
wire n_6648;
wire n_15578;
wire n_10955;
wire n_7927;
wire n_11011;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_4837;
wire n_9850;
wire n_12141;
wire n_9346;
wire n_7920;
wire n_437;
wire n_12774;
wire n_4169;
wire n_14687;
wire n_11904;
wire n_8480;
wire n_697;
wire n_17399;
wire n_388;
wire n_7025;
wire n_15886;
wire n_17022;
wire n_15856;
wire n_1757;
wire n_8484;
wire n_9472;
wire n_14304;
wire n_14357;
wire n_13044;
wire n_13228;
wire n_13518;
wire n_4070;
wire n_3885;
wire n_1369;
wire n_14008;
wire n_17069;
wire n_12746;
wire n_4031;
wire n_16162;
wire n_10970;
wire n_16285;
wire n_14927;
wire n_13881;
wire n_3209;
wire n_17205;
wire n_5547;
wire n_13747;
wire n_1391;
wire n_12532;
wire n_10238;
wire n_8931;
wire n_5596;
wire n_4653;
wire n_4435;
wire n_8334;
wire n_4019;
wire n_1071;
wire n_11681;
wire n_10890;
wire n_11202;
wire n_19513;
wire n_10552;
wire n_5815;
wire n_15254;
wire n_6595;
wire n_8539;
wire n_10205;
wire n_16947;
wire n_15747;
wire n_3727;
wire n_13899;
wire n_6306;
wire n_19386;
wire n_1714;
wire n_16235;
wire n_11663;
wire n_542;
wire n_11331;
wire n_305;
wire n_19472;
wire n_9528;
wire n_14348;
wire n_12201;
wire n_7583;
wire n_19334;
wire n_14086;
wire n_12499;
wire n_19173;
wire n_12448;
wire n_10610;
wire n_11187;
wire n_12761;
wire n_16455;
wire n_15004;
wire n_16625;
wire n_16025;
wire n_5520;
wire n_2638;
wire n_14552;
wire n_7353;
wire n_9490;
wire n_5669;
wire n_14575;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_5772;
wire n_7571;
wire n_145;
wire n_4775;
wire n_16249;
wire n_16435;
wire n_4674;
wire n_16723;
wire n_11446;
wire n_10910;
wire n_294;
wire n_8242;
wire n_11540;
wire n_13248;
wire n_17296;
wire n_19237;
wire n_9819;
wire n_15338;
wire n_8184;
wire n_425;
wire n_6525;
wire n_4286;
wire n_13119;
wire n_2958;
wire n_12642;
wire n_3731;
wire n_1822;
wire n_12484;
wire n_6128;
wire n_13549;
wire n_2489;
wire n_17361;
wire n_16080;
wire n_4525;
wire n_9992;
wire n_15180;
wire n_15692;
wire n_5712;
wire n_12669;
wire n_14296;
wire n_6702;
wire n_19490;
wire n_11179;
wire n_17074;
wire n_2520;
wire n_446;
wire n_7749;
wire n_10078;
wire n_11321;
wire n_14313;
wire n_9500;
wire n_18496;
wire n_8705;
wire n_19107;
wire n_11779;
wire n_7508;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_14211;
wire n_7574;
wire n_4306;
wire n_13516;
wire n_14273;
wire n_12462;
wire n_4453;
wire n_16462;
wire n_18648;
wire n_4005;
wire n_6169;
wire n_18775;
wire n_15230;
wire n_3546;
wire n_3661;
wire n_12735;
wire n_10709;
wire n_12646;
wire n_15875;
wire n_7352;
wire n_10244;
wire n_755;
wire n_18512;
wire n_12999;
wire n_12682;
wire n_14802;
wire n_6848;
wire n_17415;
wire n_3509;
wire n_10043;
wire n_14834;
wire n_5919;
wire n_8159;
wire n_14346;
wire n_16955;
wire n_7439;
wire n_17653;
wire n_2504;
wire n_14506;
wire n_2623;
wire n_18822;
wire n_16018;
wire n_14615;
wire n_15222;
wire n_6850;
wire n_18991;
wire n_15285;
wire n_5005;
wire n_13294;
wire n_6098;
wire n_7112;
wire n_11307;
wire n_19021;
wire n_17860;
wire n_18274;
wire n_9545;
wire n_596;
wire n_9603;
wire n_9629;
wire n_18003;
wire n_12719;
wire n_10342;
wire n_15361;
wire n_3322;
wire n_19037;
wire n_16244;
wire n_17862;
wire n_4654;
wire n_13438;
wire n_3640;
wire n_1159;
wire n_995;
wire n_15850;
wire n_9930;
wire n_14371;
wire n_12925;
wire n_5775;
wire n_14988;
wire n_9659;
wire n_3226;
wire n_2780;
wire n_16293;
wire n_9897;
wire n_9241;
wire n_14590;
wire n_14603;
wire n_8185;
wire n_11466;
wire n_5061;
wire n_15265;
wire n_15040;
wire n_6775;
wire n_9291;
wire n_4063;
wire n_11982;
wire n_2601;
wire n_773;
wire n_11873;
wire n_15821;
wire n_920;
wire n_10185;
wire n_11182;
wire n_3212;
wire n_16250;
wire n_15768;
wire n_8220;
wire n_18807;
wire n_4721;
wire n_14145;
wire n_11991;
wire n_848;
wire n_12875;
wire n_15064;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_13918;
wire n_13775;
wire n_9851;
wire n_11799;
wire n_8009;
wire n_7852;
wire n_1881;
wire n_10983;
wire n_9987;
wire n_7984;
wire n_18307;
wire n_2720;
wire n_18110;
wire n_14973;
wire n_16751;
wire n_7220;
wire n_18015;
wire n_1323;
wire n_2627;
wire n_18242;
wire n_6550;
wire n_3004;
wire n_8841;
wire n_12196;
wire n_5483;
wire n_3625;
wire n_15136;
wire n_1764;
wire n_10354;
wire n_7465;
wire n_13177;
wire n_4546;
wire n_12724;
wire n_14958;
wire n_6672;
wire n_16744;
wire n_17876;
wire n_1551;
wire n_15992;
wire n_7738;
wire n_17406;
wire n_19079;
wire n_8395;
wire n_6634;
wire n_14758;
wire n_18392;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_4635;
wire n_16802;
wire n_17909;
wire n_18439;
wire n_5735;
wire n_19022;
wire n_13311;
wire n_2278;
wire n_16020;
wire n_11513;
wire n_7464;
wire n_8937;
wire n_7115;
wire n_2924;
wire n_12087;
wire n_13675;
wire n_15022;
wire n_18693;
wire n_3595;
wire n_6104;
wire n_10537;
wire n_421;
wire n_6082;
wire n_18305;
wire n_1270;
wire n_10426;
wire n_1852;
wire n_9167;
wire n_12082;
wire n_9655;
wire n_11436;
wire n_11729;
wire n_3230;
wire n_19276;
wire n_1499;
wire n_12989;
wire n_504;
wire n_5877;
wire n_8845;
wire n_15198;
wire n_6018;
wire n_17902;
wire n_13620;
wire n_1503;
wire n_7702;
wire n_6676;
wire n_2819;
wire n_9976;
wire n_2423;
wire n_8042;
wire n_17144;
wire n_12464;
wire n_9560;
wire n_18362;
wire n_18886;
wire n_1182;
wire n_15007;
wire n_15197;
wire n_167;
wire n_8519;
wire n_5582;
wire n_5886;
wire n_1216;
wire n_6032;
wire n_18982;
wire n_9319;
wire n_5446;
wire n_3010;
wire n_12450;
wire n_5224;
wire n_14648;
wire n_11767;
wire n_2486;
wire n_3560;
wire n_10985;
wire n_9401;
wire n_11586;
wire n_12149;
wire n_12002;
wire n_12836;
wire n_19506;
wire n_17084;
wire n_13548;
wire n_15710;
wire n_2232;
wire n_11195;
wire n_4038;
wire n_16240;
wire n_2790;
wire n_9747;
wire n_5414;
wire n_14526;
wire n_13487;
wire n_17190;
wire n_3784;
wire n_17973;
wire n_220;
wire n_8586;
wire n_9058;
wire n_18707;
wire n_1472;
wire n_18547;
wire n_16700;
wire n_5454;
wire n_800;
wire n_10780;
wire n_17940;
wire n_8756;
wire n_1840;
wire n_4434;
wire n_13406;
wire n_16371;
wire n_7923;
wire n_14040;
wire n_8602;
wire n_14054;
wire n_1346;
wire n_13469;
wire n_10411;
wire n_13249;
wire n_12984;
wire n_18840;
wire n_13587;
wire n_5913;
wire n_10090;
wire n_14872;
wire n_1102;
wire n_8112;
wire n_18959;
wire n_258;
wire n_11567;
wire n_2766;
wire n_19428;
wire n_9292;
wire n_18771;
wire n_12197;
wire n_356;
wire n_17753;
wire n_19134;
wire n_4833;
wire n_11580;
wire n_13326;
wire n_6474;
wire n_13082;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_152;
wire n_18518;
wire n_12403;
wire n_10856;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_2782;
wire n_13692;
wire n_9584;
wire n_8194;
wire n_8055;
wire n_8579;
wire n_10914;
wire n_8360;
wire n_4279;
wire n_6425;
wire n_1456;
wire n_6493;
wire n_14382;
wire n_13396;
wire n_10071;
wire n_8755;
wire n_2099;
wire n_11565;
wire n_3388;
wire n_14911;
wire n_15405;
wire n_5810;
wire n_4461;
wire n_3245;
wire n_4007;
wire n_15643;
wire n_15420;
wire n_13052;
wire n_11013;
wire n_5991;
wire n_1676;
wire n_1319;
wire n_16762;
wire n_16634;
wire n_10035;
wire n_5702;
wire n_18094;
wire n_18673;
wire n_18980;
wire n_14962;
wire n_1633;
wire n_17435;
wire n_8108;
wire n_2820;
wire n_17065;
wire n_12068;
wire n_5250;
wire n_3074;
wire n_17285;
wire n_10041;
wire n_15499;
wire n_5590;
wire n_14514;
wire n_17612;
wire n_8498;
wire n_14256;
wire n_17073;
wire n_16773;
wire n_2727;
wire n_2533;
wire n_5349;
wire n_19320;
wire n_2759;
wire n_2361;
wire n_2266;
wire n_14082;
wire n_7280;
wire n_5833;
wire n_7886;
wire n_15728;
wire n_6884;
wire n_7664;
wire n_18292;
wire n_7012;
wire n_299;
wire n_1248;
wire n_17354;
wire n_12486;
wire n_902;
wire n_2189;
wire n_7376;
wire n_5816;
wire n_15347;
wire n_10137;
wire n_12084;
wire n_16517;
wire n_706;
wire n_1794;
wire n_1236;
wire n_11863;
wire n_17868;
wire n_17033;
wire n_17234;
wire n_430;
wire n_16174;
wire n_18059;
wire n_19015;
wire n_10794;
wire n_14703;
wire n_13533;
wire n_6274;
wire n_8838;
wire n_12109;
wire n_16283;
wire n_9562;
wire n_3097;
wire n_7007;
wire n_2975;
wire n_16088;
wire n_2856;
wire n_4498;
wire n_12320;
wire n_19245;
wire n_9759;
wire n_6992;
wire n_15226;
wire n_646;
wire n_528;
wire n_10206;
wire n_1329;
wire n_17736;
wire n_6322;
wire n_5167;
wire n_15425;
wire n_5661;
wire n_16878;
wire n_3589;
wire n_262;
wire n_897;
wire n_7616;
wire n_1800;
wire n_18294;
wire n_9733;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_8481;
wire n_13011;
wire n_9981;
wire n_18514;
wire n_5558;
wire n_5687;
wire n_16513;
wire n_6378;
wire n_14495;
wire n_1759;
wire n_16879;
wire n_12269;
wire n_853;
wire n_13486;
wire n_11463;
wire n_3585;
wire n_17541;
wire n_5954;
wire n_5025;
wire n_933;
wire n_17394;
wire n_7587;
wire n_3135;
wire n_17496;
wire n_6930;
wire n_17472;
wire n_19121;
wire n_12802;
wire n_11569;
wire n_10064;
wire n_7197;
wire n_9676;
wire n_7393;
wire n_11332;
wire n_13629;
wire n_13207;
wire n_310;
wire n_5766;
wire n_18025;
wire n_7358;
wire n_2796;
wire n_9950;
wire n_18088;
wire n_13589;
wire n_15730;
wire n_18089;
wire n_4534;
wire n_17967;
wire n_6929;
wire n_16706;
wire n_11309;
wire n_955;
wire n_8045;
wire n_16032;
wire n_18910;
wire n_2969;
wire n_2395;
wire n_16959;
wire n_8209;
wire n_14477;
wire n_9213;
wire n_7291;
wire n_14522;
wire n_669;
wire n_16971;
wire n_2290;
wire n_2005;
wire n_13561;
wire n_14720;
wire n_7437;
wire n_16873;
wire n_1408;
wire n_7618;
wire n_8575;
wire n_5733;
wire n_6620;
wire n_6597;
wire n_11105;
wire n_13698;
wire n_13894;
wire n_452;
wire n_6586;
wire n_10474;
wire n_12689;
wire n_18939;
wire n_8789;
wire n_7953;
wire n_13540;
wire n_6428;
wire n_5328;
wire n_14642;
wire n_12042;
wire n_14827;
wire n_15481;
wire n_5657;
wire n_174;
wire n_1173;
wire n_13465;
wire n_11130;
wire n_16149;
wire n_11664;
wire n_18705;
wire n_17430;
wire n_15388;
wire n_19242;
wire n_10652;
wire n_13733;
wire n_13098;
wire n_3334;
wire n_9388;
wire n_12654;
wire n_4985;
wire n_10869;
wire n_3823;
wire n_18708;
wire n_19112;
wire n_11783;
wire n_2255;
wire n_17837;
wire n_4678;
wire n_2649;
wire n_9911;
wire n_19603;
wire n_5579;
wire n_414;
wire n_16317;
wire n_1922;
wire n_15187;
wire n_17897;
wire n_10346;
wire n_12419;
wire n_13763;
wire n_4363;
wire n_10473;
wire n_15712;
wire n_5107;
wire n_16985;
wire n_5095;
wire n_8493;
wire n_10957;
wire n_13517;
wire n_11188;
wire n_3404;
wire n_10442;
wire n_1509;
wire n_3290;
wire n_13973;
wire n_7150;
wire n_8252;
wire n_11774;
wire n_3671;
wire n_7015;
wire n_2015;
wire n_3982;
wire n_13206;
wire n_7249;
wire n_1161;
wire n_15939;
wire n_3840;
wire n_3461;
wire n_7985;
wire n_13637;
wire n_3513;
wire n_16705;
wire n_18163;
wire n_8893;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_15904;
wire n_592;
wire n_12768;
wire n_1156;
wire n_18369;
wire n_16047;
wire n_3508;
wire n_10165;
wire n_8156;
wire n_868;
wire n_14923;
wire n_13031;
wire n_19029;
wire n_19316;
wire n_17912;
wire n_13155;
wire n_469;
wire n_1218;
wire n_13410;
wire n_19581;
wire n_7814;
wire n_8660;
wire n_985;
wire n_2440;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_19546;
wire n_561;
wire n_8606;
wire n_9663;
wire n_16584;
wire n_18340;
wire n_1244;
wire n_9743;
wire n_19048;
wire n_11584;
wire n_2285;
wire n_5280;
wire n_14169;
wire n_7700;
wire n_4451;
wire n_10158;
wire n_10582;
wire n_16151;
wire n_10427;
wire n_11816;
wire n_18808;
wire n_3563;
wire n_16420;
wire n_201;
wire n_11693;
wire n_3495;
wire n_15429;
wire n_9248;
wire n_6138;
wire n_5369;
wire n_10835;
wire n_975;
wire n_11411;
wire n_5576;
wire n_13823;
wire n_11386;
wire n_11604;
wire n_13323;
wire n_3359;
wire n_12164;
wire n_16919;
wire n_12824;
wire n_13434;
wire n_16680;
wire n_16938;
wire n_3187;
wire n_10844;
wire n_17793;
wire n_14153;
wire n_6802;
wire n_10654;
wire n_6909;
wire n_13445;
wire n_17177;
wire n_19074;
wire n_18182;
wire n_4336;
wire n_15760;
wire n_16712;
wire n_14746;
wire n_11097;
wire n_4981;
wire n_14606;
wire n_12052;
wire n_9746;
wire n_8073;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_8821;
wire n_9440;
wire n_3955;
wire n_17253;
wire n_2280;
wire n_203;
wire n_1868;
wire n_17264;
wire n_2079;
wire n_15475;
wire n_8663;
wire n_2185;
wire n_5861;
wire n_1836;
wire n_10553;
wire n_8309;
wire n_1486;
wire n_5258;
wire n_8945;
wire n_15121;
wire n_10988;
wire n_19209;
wire n_784;
wire n_6112;
wire n_16192;
wire n_18030;
wire n_9041;
wire n_862;
wire n_8166;
wire n_2098;
wire n_5606;
wire n_1935;
wire n_10108;
wire n_13865;
wire n_5920;
wire n_10307;
wire n_1449;
wire n_361;
wire n_8215;
wire n_19538;
wire n_17497;
wire n_6180;
wire n_8809;
wire n_12382;
wire n_5527;
wire n_6476;
wire n_14428;
wire n_6566;
wire n_5172;
wire n_11173;
wire n_16218;
wire n_6872;
wire n_13998;
wire n_5254;
wire n_17825;
wire n_10587;
wire n_8713;
wire n_15450;
wire n_7111;
wire n_13522;
wire n_7967;
wire n_15609;
wire n_16423;
wire n_9002;
wire n_14670;
wire n_9130;
wire n_19016;
wire n_7180;
wire n_13530;
wire n_16362;
wire n_8604;
wire n_7263;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_677;
wire n_14318;
wire n_4686;
wire n_17673;
wire n_17004;
wire n_11802;
wire n_3706;
wire n_8005;
wire n_2179;
wire n_13942;
wire n_18230;
wire n_1547;
wire n_12570;
wire n_11905;
wire n_19326;
wire n_893;
wire n_3801;
wire n_5267;
wire n_10202;
wire n_3564;
wire n_9104;
wire n_15295;
wire n_17050;
wire n_17408;
wire n_15445;
wire n_8272;
wire n_13997;
wire n_14402;
wire n_14882;
wire n_11051;
wire n_11214;
wire n_2628;
wire n_7000;
wire n_7398;
wire n_18335;
wire n_1078;
wire n_14232;
wire n_12882;
wire n_19300;
wire n_18057;
wire n_12617;
wire n_8236;
wire n_13137;
wire n_3345;
wire n_19612;
wire n_15933;
wire n_17188;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_10348;
wire n_12495;
wire n_9581;
wire n_8070;
wire n_4696;
wire n_18468;
wire n_16786;
wire n_7802;
wire n_17118;
wire n_3877;
wire n_15353;
wire n_19623;
wire n_1455;
wire n_6629;
wire n_15993;
wire n_5279;
wire n_5894;
wire n_17699;
wire n_19605;
wire n_8175;
wire n_567;
wire n_8953;
wire n_17546;
wire n_17279;
wire n_19111;
wire n_4814;
wire n_10373;
wire n_3979;
wire n_3077;
wire n_9525;
wire n_10816;
wire n_9725;
wire n_19511;
wire n_6914;
wire n_14121;
wire n_10381;
wire n_713;
wire n_1400;
wire n_10947;
wire n_16984;
wire n_6015;
wire n_11261;
wire n_16012;
wire n_1560;
wire n_734;
wire n_13929;
wire n_17739;
wire n_10767;
wire n_14646;
wire n_14095;
wire n_15069;
wire n_14520;
wire n_14780;
wire n_4950;
wire n_4729;
wire n_4268;
wire n_11447;
wire n_12652;
wire n_15507;
wire n_8142;
wire n_11627;
wire n_6404;
wire n_12209;
wire n_6674;
wire n_5680;
wire n_17883;
wire n_13606;
wire n_11659;
wire n_13501;
wire n_4102;
wire n_9106;
wire n_4662;
wire n_8869;
wire n_3959;
wire n_2268;
wire n_8381;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_17149;
wire n_9520;
wire n_2080;
wire n_14931;
wire n_18774;
wire n_7770;
wire n_6968;
wire n_16268;
wire n_12371;
wire n_4507;
wire n_11497;
wire n_14900;
wire n_792;
wire n_15846;
wire n_13454;
wire n_5306;
wire n_16662;
wire n_9042;
wire n_17329;
wire n_3488;
wire n_8987;
wire n_11805;
wire n_1910;
wire n_14935;
wire n_2998;
wire n_237;
wire n_6282;
wire n_12770;
wire n_4294;
wire n_19551;
wire n_11635;
wire n_15434;
wire n_16530;
wire n_12951;
wire n_9453;
wire n_8118;
wire n_12393;
wire n_16442;
wire n_9718;
wire n_10281;
wire n_3927;
wire n_3888;
wire n_764;
wire n_12831;
wire n_2895;
wire n_6431;
wire n_733;
wire n_19620;
wire n_15767;
wire n_1290;
wire n_12427;
wire n_1354;
wire n_7533;
wire n_7221;
wire n_16026;
wire n_15159;
wire n_1701;
wire n_10656;
wire n_6575;
wire n_6055;
wire n_8246;
wire n_8952;
wire n_3875;
wire n_5609;
wire n_4717;
wire n_871;
wire n_15154;
wire n_9680;
wire n_12172;
wire n_5658;
wire n_4731;
wire n_12923;
wire n_12147;
wire n_3052;
wire n_19624;
wire n_13227;
wire n_8848;
wire n_12825;
wire n_5667;
wire n_8259;
wire n_2624;
wire n_5865;
wire n_15182;
wire n_8349;
wire n_6836;
wire n_11998;
wire n_8776;
wire n_19391;
wire n_7753;
wire n_6771;
wire n_14732;
wire n_9947;
wire n_16659;
wire n_1750;
wire n_1462;
wire n_10138;
wire n_12117;
wire n_10375;
wire n_14535;
wire n_6795;
wire n_5314;
wire n_12960;
wire n_18972;
wire n_14094;
wire n_13033;
wire n_15703;
wire n_19353;
wire n_7648;
wire n_515;
wire n_4418;
wire n_12131;
wire n_12851;
wire n_7452;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_514;
wire n_15518;
wire n_14217;
wire n_10903;
wire n_17596;
wire n_15574;
wire n_14062;
wire n_8453;
wire n_12740;
wire n_2393;
wire n_2921;
wire n_3237;
wire n_8949;
wire n_10831;
wire n_9131;
wire n_17580;
wire n_10517;
wire n_16889;
wire n_10323;
wire n_10842;
wire n_17620;
wire n_3542;
wire n_16465;
wire n_2763;
wire n_2762;
wire n_11146;
wire n_10883;
wire n_17785;
wire n_1296;
wire n_19249;
wire n_3073;
wire n_5343;
wire n_1294;
wire n_3696;
wire n_12278;
wire n_18918;
wire n_19018;
wire n_1779;
wire n_524;
wire n_17672;
wire n_4329;
wire n_18036;
wire n_5135;
wire n_17414;
wire n_10123;
wire n_10651;
wire n_4697;
wire n_3763;
wire n_17483;
wire n_17689;
wire n_18975;
wire n_14785;
wire n_8500;
wire n_17857;
wire n_2145;
wire n_4964;
wire n_12804;
wire n_12116;
wire n_17438;
wire n_1932;
wire n_13755;
wire n_1101;
wire n_10468;
wire n_4636;
wire n_14126;
wire n_14105;
wire n_8285;
wire n_8483;
wire n_4946;
wire n_4767;
wire n_4287;
wire n_19145;
wire n_17696;
wire n_1451;
wire n_639;
wire n_11370;
wire n_16731;
wire n_4576;
wire n_9020;
wire n_4615;
wire n_1018;
wire n_9895;
wire n_16452;
wire n_11585;
wire n_13140;
wire n_13962;
wire n_4389;
wire n_13753;
wire n_1376;
wire n_15365;
wire n_17141;
wire n_948;
wire n_12560;
wire n_19295;
wire n_18171;
wire n_977;
wire n_13610;
wire n_536;
wire n_8851;
wire n_13332;
wire n_15293;
wire n_19405;
wire n_6097;
wire n_19214;
wire n_7093;
wire n_4098;
wire n_5026;
wire n_4476;
wire n_432;
wire n_3700;
wire n_3104;
wire n_2239;
wire n_7840;
wire n_18797;
wire n_10024;
wire n_16386;
wire n_17101;
wire n_15695;
wire n_7080;
wire n_17984;
wire n_2191;
wire n_14156;
wire n_10711;
wire n_7624;
wire n_1426;
wire n_16185;
wire n_9186;
wire n_10818;
wire n_1529;
wire n_4634;
wire n_2069;
wire n_18851;
wire n_2362;
wire n_4096;
wire n_15178;
wire n_2698;
wire n_12222;
wire n_11951;
wire n_7003;
wire n_13604;
wire n_5427;
wire n_10788;
wire n_17163;
wire n_10563;
wire n_8810;
wire n_3631;
wire n_2772;
wire n_14518;
wire n_16310;
wire n_16477;
wire n_13397;
wire n_10178;
wire n_5052;
wire n_4541;
wire n_17731;
wire n_15360;
wire n_929;
wire n_4551;
wire n_2857;
wire n_13132;
wire n_6609;
wire n_10115;
wire n_17157;
wire n_5326;
wire n_16927;
wire n_12793;
wire n_11778;
wire n_1183;
wire n_2494;
wire n_12406;
wire n_998;
wire n_717;
wire n_1383;
wire n_7484;
wire n_16639;
wire n_6414;
wire n_1000;
wire n_9470;
wire n_3810;
wire n_552;
wire n_15516;
wire n_3006;
wire n_216;
wire n_13792;
wire n_5010;
wire n_1201;
wire n_4592;
wire n_18229;
wire n_9405;
wire n_1395;
wire n_6264;
wire n_2199;
wire n_17426;
wire n_13480;
wire n_1955;
wire n_19583;
wire n_312;
wire n_13571;
wire n_10984;
wire n_5104;
wire n_18742;
wire n_12001;
wire n_7883;
wire n_589;
wire n_1310;
wire n_13715;
wire n_3591;
wire n_16675;
wire n_2797;
wire n_7458;
wire n_4746;
wire n_15186;
wire n_16935;
wire n_18576;
wire n_13810;
wire n_14403;
wire n_7435;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_3964;
wire n_19292;
wire n_13473;
wire n_18267;
wire n_5985;
wire n_556;
wire n_15963;
wire n_14353;
wire n_16589;
wire n_1602;
wire n_19213;
wire n_11742;
wire n_6891;
wire n_10031;
wire n_276;
wire n_19163;
wire n_12235;
wire n_5232;
wire n_7663;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_14386;
wire n_18784;
wire n_16472;
wire n_17830;
wire n_12098;
wire n_4428;
wire n_1533;
wire n_7917;
wire n_12579;
wire n_2274;
wire n_9203;
wire n_15073;
wire n_7532;
wire n_9613;
wire n_5761;
wire n_13982;
wire n_18703;
wire n_12611;
wire n_13269;
wire n_7375;
wire n_13369;
wire n_7968;
wire n_6382;
wire n_317;
wire n_18542;
wire n_1679;
wire n_9141;
wire n_15867;
wire n_5760;
wire n_2146;
wire n_11027;
wire n_11852;
wire n_5472;
wire n_8377;
wire n_9913;
wire n_2575;
wire n_9286;
wire n_19646;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_10819;
wire n_1179;
wire n_324;
wire n_14521;
wire n_9704;
wire n_19468;
wire n_19025;
wire n_9046;
wire n_16576;
wire n_6339;
wire n_8814;
wire n_8530;
wire n_9193;
wire n_16882;
wire n_7711;
wire n_16181;
wire n_15948;
wire n_8984;
wire n_17123;
wire n_3663;
wire n_3299;
wire n_9290;
wire n_351;
wire n_259;
wire n_14580;
wire n_5745;
wire n_1645;
wire n_14028;
wire n_19131;
wire n_14772;
wire n_956;
wire n_13827;
wire n_14542;
wire n_18632;
wire n_3845;
wire n_664;
wire n_1869;
wire n_7230;
wire n_17552;
wire n_7989;
wire n_9778;
wire n_18986;
wire n_2016;
wire n_5171;
wire n_18280;
wire n_15003;
wire n_13200;
wire n_1937;
wire n_16783;
wire n_12848;
wire n_18963;
wire n_341;
wire n_1744;
wire n_828;
wire n_10315;
wire n_18321;
wire n_607;
wire n_19104;
wire n_17187;
wire n_4028;
wire n_17031;
wire n_11455;
wire n_12368;
wire n_5255;
wire n_3756;
wire n_17240;
wire n_3406;
wire n_13193;
wire n_951;
wire n_952;
wire n_8462;
wire n_18953;
wire n_9380;
wire n_10062;
wire n_18235;
wire n_19476;
wire n_2375;
wire n_1934;
wire n_10514;
wire n_8429;
wire n_1434;
wire n_12785;
wire n_3981;
wire n_15312;
wire n_14155;
wire n_1275;
wire n_1510;
wire n_7620;
wire n_5783;
wire n_3120;
wire n_5821;
wire n_15818;
wire n_6079;
wire n_16481;
wire n_16430;
wire n_19313;
wire n_3864;
wire n_16715;
wire n_8492;
wire n_16565;
wire n_248;
wire n_2302;
wire n_8135;
wire n_16620;
wire n_8445;
wire n_1037;
wire n_6427;
wire n_3592;
wire n_468;
wire n_4230;
wire n_14978;
wire n_2637;
wire n_18353;
wire n_12639;
wire n_991;
wire n_8895;
wire n_3817;
wire n_7811;
wire n_340;
wire n_14649;
wire n_15940;
wire n_12175;
wire n_5003;
wire n_13536;
wire n_10512;
wire n_14714;
wire n_11384;
wire n_4827;
wire n_8273;
wire n_12353;
wire n_14129;
wire n_6065;
wire n_9761;
wire n_16962;
wire n_4610;
wire n_9087;
wire n_4472;
wire n_17832;
wire n_3081;
wire n_17316;
wire n_15333;
wire n_10434;
wire n_12869;
wire n_8312;
wire n_6781;
wire n_18585;
wire n_13830;
wire n_6133;
wire n_14184;
wire n_11889;
wire n_14183;
wire n_6127;
wire n_4990;
wire n_19172;
wire n_17751;
wire n_2498;
wire n_11362;
wire n_19256;
wire n_8078;
wire n_4515;
wire n_14200;
wire n_6006;
wire n_16558;
wire n_7926;
wire n_19118;
wire n_6598;
wire n_172;
wire n_15568;
wire n_12502;
wire n_2392;
wire n_4131;
wire n_16859;
wire n_1043;
wire n_18800;
wire n_16703;
wire n_2305;
wire n_13191;
wire n_10131;
wire n_15464;
wire n_17741;
wire n_6867;
wire n_12600;
wire n_14536;
wire n_16338;
wire n_6139;
wire n_12133;
wire n_7965;
wire n_12919;
wire n_3356;
wire n_10273;
wire n_11416;
wire n_3210;
wire n_937;
wire n_17485;
wire n_14321;
wire n_1682;
wire n_7474;
wire n_11169;
wire n_8650;
wire n_17843;
wire n_14654;
wire n_10503;
wire n_4905;
wire n_14664;
wire n_13215;
wire n_4601;
wire n_16834;
wire n_962;
wire n_10465;
wire n_16073;
wire n_10590;
wire n_3647;
wire n_13782;
wire n_15476;
wire n_8526;
wire n_1186;
wire n_13751;
wire n_17150;
wire n_14019;
wire n_19140;
wire n_19418;
wire n_6759;
wire n_10786;
wire n_3988;
wire n_7028;
wire n_9890;
wire n_11492;
wire n_19653;
wire n_394;
wire n_18904;
wire n_6535;
wire n_18801;
wire n_16644;
wire n_9817;
wire n_1524;
wire n_11160;
wire n_18899;
wire n_9782;
wire n_1920;
wire n_3292;
wire n_1225;
wire n_12319;
wire n_10805;
wire n_17214;
wire n_6643;
wire n_17982;
wire n_9471;
wire n_3712;
wire n_4608;
wire n_2506;
wire n_17012;
wire n_14896;
wire n_17440;
wire n_12930;
wire n_17181;
wire n_1567;
wire n_4037;
wire n_8351;
wire n_9069;
wire n_17371;
wire n_3562;
wire n_14030;
wire n_8603;
wire n_17274;
wire n_16660;
wire n_11343;
wire n_3007;
wire n_19143;
wire n_12575;
wire n_11451;
wire n_4571;
wire n_16853;
wire n_3698;
wire n_13384;
wire n_3355;
wire n_2114;
wire n_16048;
wire n_16262;
wire n_17127;
wire n_15422;
wire n_9003;
wire n_2154;
wire n_18874;
wire n_12418;
wire n_5290;
wire n_4185;
wire n_14837;
wire n_7312;
wire n_4219;
wire n_11269;
wire n_16849;
wire n_3985;
wire n_1447;
wire n_14103;
wire n_4774;
wire n_6689;
wire n_7632;
wire n_9172;
wire n_14653;
wire n_4232;
wire n_3000;
wire n_19464;
wire n_17275;
wire n_8980;
wire n_5571;
wire n_17573;
wire n_11311;
wire n_6698;
wire n_18553;
wire n_17345;
wire n_17770;
wire n_13242;
wire n_7707;
wire n_13282;
wire n_14436;
wire n_12113;
wire n_14599;
wire n_16087;
wire n_4736;
wire n_1725;
wire n_3743;
wire n_13352;
wire n_17648;
wire n_18116;
wire n_17853;
wire n_14812;
wire n_17871;
wire n_11293;
wire n_14728;
wire n_19184;
wire n_545;
wire n_2671;
wire n_6363;
wire n_2715;
wire n_8619;
wire n_3511;
wire n_19224;
wire n_18217;
wire n_18812;
wire n_15122;
wire n_10134;
wire n_11603;
wire n_1477;
wire n_7277;
wire n_11271;
wire n_14778;
wire n_15714;
wire n_17270;
wire n_12015;
wire n_8146;
wire n_13690;
wire n_2833;
wire n_11562;
wire n_10194;
wire n_17085;
wire n_8910;
wire n_1001;
wire n_6408;
wire n_6150;
wire n_10077;
wire n_4708;
wire n_13619;
wire n_4657;
wire n_18508;
wire n_12031;
wire n_1191;
wire n_9278;
wire n_855;
wire n_10889;
wire n_10010;
wire n_14996;
wire n_12126;
wire n_14543;
wire n_8550;
wire n_11094;
wire n_14747;
wire n_10599;
wire n_9667;
wire n_6401;
wire n_9739;
wire n_14358;
wire n_4536;
wire n_9480;
wire n_17886;
wire n_1976;
wire n_12195;
wire n_19369;
wire n_6679;
wire n_19294;
wire n_1824;
wire n_13289;
wire n_13182;
wire n_16265;
wire n_16466;
wire n_13324;
wire n_9541;
wire n_11286;
wire n_15215;
wire n_18947;
wire n_17748;
wire n_16379;
wire n_16728;
wire n_823;
wire n_1074;
wire n_7097;
wire n_8140;
wire n_15111;
wire n_1097;
wire n_781;
wire n_18563;
wire n_1810;
wire n_5915;
wire n_8527;
wire n_12899;
wire n_18917;
wire n_1583;
wire n_17621;
wire n_2295;
wire n_1643;
wire n_19570;
wire n_7909;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_15759;
wire n_10734;
wire n_16441;
wire n_15383;
wire n_11560;
wire n_10395;
wire n_3617;
wire n_14966;
wire n_11435;
wire n_1598;
wire n_15255;
wire n_6214;
wire n_9370;
wire n_918;
wire n_13136;
wire n_763;
wire n_6692;
wire n_2485;
wire n_14322;
wire n_12331;
wire n_8093;
wire n_6036;
wire n_13349;
wire n_9956;
wire n_17007;
wire n_6552;
wire n_17096;
wire n_8327;
wire n_13096;
wire n_15314;
wire n_10991;
wire n_14173;
wire n_17005;
wire n_1702;
wire n_4947;
wire n_9487;
wire n_16791;
wire n_14608;
wire n_7306;
wire n_16153;
wire n_10118;
wire n_795;
wire n_18791;
wire n_7470;
wire n_13800;
wire n_19593;
wire n_1245;
wire n_7693;
wire n_3215;
wire n_4740;
wire n_15662;
wire n_1112;
wire n_10002;
wire n_2081;
wire n_911;
wire n_11242;
wire n_17974;
wire n_2862;
wire n_472;
wire n_15923;
wire n_2474;
wire n_3703;
wire n_13694;
wire n_4863;
wire n_17494;
wire n_2267;
wire n_668;
wire n_1821;
wire n_9660;
wire n_16233;
wire n_17344;
wire n_13093;
wire n_9328;
wire n_16511;
wire n_15274;
wire n_16410;
wire n_7653;
wire n_8354;
wire n_14276;
wire n_6959;
wire n_8353;
wire n_6388;
wire n_5045;
wire n_13185;
wire n_11053;
wire n_18635;
wire n_12159;
wire n_9434;
wire n_18450;
wire n_13855;
wire n_10902;
wire n_19596;
wire n_8348;
wire n_7032;
wire n_19086;
wire n_18806;
wire n_8211;
wire n_1816;
wire n_11304;
wire n_9681;
wire n_5848;
wire n_10485;
wire n_7475;
wire n_18448;
wire n_4612;
wire n_6435;
wire n_10536;
wire n_2531;
wire n_9079;
wire n_15544;
wire n_18738;
wire n_19564;
wire n_16145;
wire n_19424;
wire n_17512;
wire n_18931;
wire n_18988;
wire n_714;
wire n_8653;
wire n_8920;
wire n_17521;
wire n_10950;
wire n_5485;
wire n_17477;
wire n_6682;
wire n_6823;
wire n_14550;
wire n_9089;
wire n_4390;
wire n_15346;
wire n_13477;
wire n_18200;
wire n_2095;
wire n_8942;
wire n_10978;
wire n_8222;
wire n_13808;
wire n_6822;
wire n_3295;
wire n_8553;
wire n_1998;
wire n_240;
wire n_19608;
wire n_17068;
wire n_10187;
wire n_11014;
wire n_17508;
wire n_15033;
wire n_2640;
wire n_3288;
wire n_583;
wire n_17789;
wire n_3876;
wire n_9564;
wire n_7391;
wire n_9230;
wire n_19301;
wire n_941;
wire n_19297;
wire n_10768;
wire n_14067;
wire n_6389;
wire n_15903;
wire n_2471;
wire n_6983;
wire n_10494;
wire n_8398;
wire n_13970;
wire n_15247;
wire n_16656;
wire n_4580;
wire n_1055;
wire n_2197;
wire n_10065;
wire n_8700;
wire n_4148;
wire n_2461;
wire n_271;
wire n_13408;
wire n_17585;
wire n_15248;
wire n_13727;
wire n_17500;
wire n_13025;
wire n_10268;
wire n_18728;
wire n_14801;
wire n_12601;
wire n_15399;
wire n_17549;
wire n_13641;
wire n_2634;
wire n_1761;
wire n_19588;
wire n_19493;
wire n_8750;
wire n_17473;
wire n_17746;
wire n_5868;
wire n_10305;
wire n_2308;
wire n_16862;
wire n_3001;
wire n_12807;
wire n_15669;
wire n_18018;
wire n_3795;
wire n_7321;
wire n_5289;
wire n_8200;
wire n_4138;
wire n_16055;
wire n_19053;
wire n_18179;
wire n_18564;
wire n_3815;
wire n_12981;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_339;
wire n_434;
wire n_13542;
wire n_288;
wire n_8212;
wire n_5612;
wire n_14426;
wire n_9016;
wire n_15456;
wire n_11545;
wire n_8846;
wire n_4834;
wire n_12665;
wire n_19469;
wire n_16526;
wire n_16397;
wire n_11850;
wire n_9194;
wire n_8760;
wire n_12592;
wire n_17467;
wire n_9029;
wire n_6837;
wire n_3813;
wire n_18860;
wire n_1613;
wire n_11043;
wire n_9414;
wire n_18539;
wire n_7023;
wire n_9615;
wire n_14205;
wire n_1189;
wire n_18532;
wire n_5034;
wire n_726;
wire n_10779;
wire n_11061;
wire n_16495;
wire n_17922;
wire n_5375;
wire n_15742;
wire n_16686;
wire n_16347;
wire n_5370;
wire n_9811;
wire n_5784;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_16385;
wire n_19141;
wire n_1708;
wire n_805;
wire n_14723;
wire n_2051;
wire n_5112;
wire n_19205;
wire n_1402;
wire n_1691;
wire n_10520;
wire n_17437;
wire n_13531;
wire n_7797;
wire n_3668;
wire n_18641;
wire n_13880;
wire n_7687;
wire n_2491;
wire n_1264;
wire n_18251;
wire n_4087;
wire n_7582;
wire n_10541;
wire n_14587;
wire n_8959;
wire n_17326;
wire n_10614;
wire n_18834;
wire n_7809;
wire n_461;
wire n_16877;
wire n_18169;
wire n_8425;
wire n_11257;
wire n_15176;
wire n_9910;
wire n_16790;
wire n_10217;
wire n_17255;
wire n_2513;
wire n_10743;
wire n_2247;
wire n_13424;
wire n_14658;
wire n_15066;
wire n_1579;
wire n_9651;
wire n_3275;
wire n_836;
wire n_15474;
wire n_15316;
wire n_10270;
wire n_11115;
wire n_8001;
wire n_2094;
wire n_1511;
wire n_17417;
wire n_7529;
wire n_14233;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_1313;
wire n_3607;
wire n_3316;
wire n_2418;
wire n_6881;
wire n_3371;
wire n_19269;
wire n_9544;
wire n_3261;
wire n_17324;
wire n_666;
wire n_7520;
wire n_9831;
wire n_4187;
wire n_940;
wire n_18245;
wire n_9697;
wire n_18878;
wire n_5317;
wire n_18414;
wire n_494;
wire n_8362;
wire n_2394;
wire n_5540;
wire n_6300;
wire n_8256;
wire n_5716;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_12091;
wire n_8704;
wire n_17589;
wire n_6132;
wire n_5211;
wire n_17493;
wire n_9294;
wire n_11747;
wire n_6395;
wire n_976;
wire n_7054;
wire n_2686;
wire n_5327;
wire n_4392;
wire n_11858;
wire n_14027;
wire n_7433;
wire n_16316;
wire n_10075;
wire n_10423;
wire n_17762;
wire n_4334;
wire n_3351;
wire n_6171;
wire n_17291;
wire n_17895;
wire n_5519;
wire n_11895;
wire n_13458;
wire n_4047;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_10886;
wire n_18720;
wire n_13003;
wire n_3791;
wire n_13091;
wire n_6387;
wire n_10192;
wire n_9465;
wire n_13811;
wire n_5139;
wire n_757;
wire n_19459;
wire n_14011;
wire n_166;
wire n_10436;
wire n_19026;
wire n_12794;
wire n_15496;
wire n_6342;
wire n_17744;
wire n_15260;
wire n_15104;
wire n_12483;
wire n_16374;
wire n_18173;
wire n_17251;
wire n_3883;
wire n_18945;
wire n_261;
wire n_5866;
wire n_3728;
wire n_2925;
wire n_5822;
wire n_17381;
wire n_9959;
wire n_15055;
wire n_3949;
wire n_11015;
wire n_18712;
wire n_5364;
wire n_3315;
wire n_9631;
wire n_14751;
wire n_6194;
wire n_4893;
wire n_18313;
wire n_12815;
wire n_15913;
wire n_10431;
wire n_9945;
wire n_1413;
wire n_2228;
wire n_17694;
wire n_5039;
wire n_16314;
wire n_2455;
wire n_4772;
wire n_15115;
wire n_8746;
wire n_11183;
wire n_10019;
wire n_8531;
wire n_12093;
wire n_19296;
wire n_11581;
wire n_4468;
wire n_4161;
wire n_6459;
wire n_8379;
wire n_13100;
wire n_4961;
wire n_4454;
wire n_16154;
wire n_12334;
wire n_18397;
wire n_9209;
wire n_7311;
wire n_3686;
wire n_18234;
wire n_7669;
wire n_8793;
wire n_12355;
wire n_19340;
wire n_15052;
wire n_9838;
wire n_9767;
wire n_1713;
wire n_4277;
wire n_9300;
wire n_11500;
wire n_12943;
wire n_17598;
wire n_530;
wire n_17956;
wire n_618;
wire n_11021;
wire n_8543;
wire n_16502;
wire n_3069;
wire n_7189;
wire n_13067;
wire n_6258;
wire n_16688;
wire n_10243;
wire n_9700;
wire n_18114;
wire n_18802;
wire n_3725;
wire n_8533;
wire n_15483;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_5554;
wire n_1175;
wire n_10596;
wire n_903;
wire n_12140;
wire n_1802;
wire n_286;
wire n_254;
wire n_8063;
wire n_3961;
wire n_12599;
wire n_2347;
wire n_19419;
wire n_816;
wire n_8032;
wire n_7427;
wire n_2967;
wire n_13250;
wire n_11190;
wire n_11794;
wire n_10519;
wire n_2467;
wire n_17630;
wire n_10163;
wire n_17409;
wire n_3983;
wire n_3538;
wire n_16544;
wire n_2824;
wire n_17529;
wire n_18979;
wire n_12330;
wire n_950;
wire n_15871;
wire n_14819;
wire n_14890;
wire n_8129;
wire n_13906;
wire n_3009;
wire n_5824;
wire n_6760;
wire n_14265;
wire n_13664;
wire n_13566;
wire n_12591;
wire n_12466;
wire n_9509;
wire n_3526;
wire n_4367;
wire n_10874;
wire n_6825;
wire n_19558;
wire n_11831;
wire n_16213;
wire n_14399;
wire n_9628;
wire n_18940;
wire n_19348;
wire n_2583;
wire n_18279;
wire n_19655;
wire n_10250;
wire n_1033;
wire n_1052;
wire n_2794;
wire n_18658;
wire n_14063;
wire n_16657;
wire n_2078;
wire n_2932;
wire n_3431;
wire n_3450;
wire n_17584;
wire n_12041;
wire n_449;
wire n_16734;
wire n_17783;
wire n_2728;
wire n_15157;
wire n_13074;
wire n_3183;
wire n_1067;
wire n_14716;
wire n_255;
wire n_1952;
wire n_12876;
wire n_15286;
wire n_14698;
wire n_19152;
wire n_18633;
wire n_6468;
wire n_3937;
wire n_3159;
wire n_14323;
wire n_18565;
wire n_13071;
wire n_6857;
wire n_3576;
wire n_1863;
wire n_12536;
wire n_10795;
wire n_16333;
wire n_872;
wire n_15116;
wire n_8049;
wire n_7762;
wire n_9467;
wire n_7186;
wire n_13739;
wire n_11157;
wire n_9097;
wire n_1513;
wire n_14364;
wire n_15472;
wire n_837;
wire n_5087;
wire n_13234;
wire n_9314;
wire n_7017;
wire n_16718;
wire n_2060;
wire n_7830;
wire n_5131;
wire n_19217;
wire n_17380;
wire n_8084;
wire n_14113;
wire n_8289;
wire n_11178;
wire n_5887;
wire n_16428;
wire n_19010;
wire n_14938;
wire n_14784;
wire n_2816;
wire n_11432;
wire n_14179;
wire n_17755;
wire n_7191;
wire n_14979;
wire n_10412;
wire n_12650;
wire n_4443;
wire n_14324;
wire n_614;
wire n_5460;
wire n_1615;
wire n_4114;
wire n_12859;
wire n_2119;
wire n_17763;
wire n_7961;
wire n_5899;
wire n_17176;
wire n_10617;
wire n_3185;
wire n_2605;
wire n_16524;
wire n_10544;
wire n_13030;
wire n_2848;
wire n_919;
wire n_17819;
wire n_18475;
wire n_15094;
wire n_16880;
wire n_11952;
wire n_6422;
wire n_1299;
wire n_13896;
wire n_5339;
wire n_3837;
wire n_16473;
wire n_1436;
wire n_9873;
wire n_13299;
wire n_13042;
wire n_4818;
wire n_15658;
wire n_10095;
wire n_15873;
wire n_8268;
wire n_6160;
wire n_7066;
wire n_18128;
wire n_796;
wire n_7789;
wire n_184;
wire n_6192;
wire n_10056;
wire n_16597;
wire n_17627;
wire n_18815;
wire n_6039;
wire n_2144;
wire n_11919;
wire n_1142;
wire n_11414;
wire n_17705;
wire n_5719;
wire n_17728;
wire n_19457;
wire n_17618;
wire n_7344;
wire n_9888;
wire n_10037;
wire n_2259;
wire n_18029;
wire n_6707;
wire n_12744;
wire n_19601;
wire n_11136;
wire n_3142;
wire n_19527;
wire n_6787;
wire n_11620;
wire n_15480;
wire n_10179;
wire n_4709;
wire n_2132;
wire n_14038;
wire n_18726;
wire n_11215;
wire n_2860;
wire n_2330;
wire n_11890;
wire n_9366;
wire n_14253;
wire n_7915;
wire n_5893;
wire n_9077;
wire n_2281;
wire n_8406;
wire n_15919;
wire n_16652;
wire n_12443;
wire n_6463;
wire n_11683;
wire n_8554;
wire n_386;
wire n_6051;
wire n_2301;
wire n_7538;
wire n_12934;
wire n_3270;
wire n_19547;
wire n_18981;
wire n_970;
wire n_6799;
wire n_19368;
wire n_444;
wire n_3311;
wire n_3913;
wire n_6487;
wire n_8818;
wire n_16648;
wire n_4348;
wire n_16724;
wire n_10466;
wire n_11953;
wire n_4404;
wire n_439;
wire n_6563;
wire n_2828;
wire n_7554;
wire n_2384;
wire n_4204;
wire n_19005;
wire n_759;
wire n_18881;
wire n_2724;
wire n_15926;
wire n_4513;
wire n_16943;
wire n_11089;
wire n_6341;
wire n_13422;
wire n_7421;
wire n_10166;
wire n_7489;
wire n_1647;
wire n_14702;
wire n_13179;
wire n_15844;
wire n_2306;
wire n_11839;
wire n_18039;
wire n_3683;
wire n_4801;
wire n_13834;
wire n_401;
wire n_18277;
wire n_2550;
wire n_8341;
wire n_11193;
wire n_17800;
wire n_17613;
wire n_7188;
wire n_3736;
wire n_11217;
wire n_15651;
wire n_17759;
wire n_6923;
wire n_9287;
wire n_7991;
wire n_10877;
wire n_16737;
wire n_14686;
wire n_3284;
wire n_12214;
wire n_427;
wire n_16259;
wire n_8926;
wire n_2995;
wire n_10766;
wire n_4438;
wire n_4844;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_13924;
wire n_4149;
wire n_9608;
wire n_501;
wire n_19539;
wire n_8817;
wire n_8190;
wire n_1668;
wire n_2777;
wire n_11488;
wire n_13671;
wire n_14876;
wire n_18571;
wire n_1129;
wire n_6987;
wire n_18265;
wire n_11037;
wire n_16925;
wire n_18740;
wire n_14319;
wire n_2911;
wire n_1429;
wire n_5706;
wire n_16763;
wire n_3429;
wire n_17462;
wire n_1593;
wire n_15287;
wire n_1202;
wire n_7671;
wire n_13150;
wire n_5431;
wire n_15103;
wire n_12541;
wire n_8649;
wire n_14818;
wire n_19508;
wire n_8303;
wire n_6153;
wire n_16512;
wire n_13809;
wire n_8059;
wire n_18364;
wire n_11665;
wire n_6579;
wire n_13590;
wire n_16747;
wire n_11138;
wire n_5798;
wire n_575;
wire n_11731;
wire n_5875;
wire n_16257;
wire n_5621;
wire n_16200;
wire n_16041;
wire n_732;
wire n_2983;
wire n_16023;
wire n_6789;
wire n_12100;
wire n_1042;
wire n_15327;
wire n_17718;
wire n_1728;
wire n_13471;
wire n_17615;
wire n_845;
wire n_19063;
wire n_140;
wire n_8862;
wire n_16161;
wire n_10580;
wire n_17287;
wire n_4870;
wire n_6164;
wire n_13261;
wire n_768;
wire n_9675;
wire n_7786;
wire n_16923;
wire n_11454;
wire n_7609;
wire n_3449;
wire n_2598;
wire n_8900;
wire n_597;
wire n_12523;
wire n_6934;
wire n_1403;
wire n_6737;
wire n_18388;
wire n_4488;
wire n_3767;
wire n_8478;
wire n_16988;
wire n_6695;
wire n_12395;
wire n_4211;
wire n_5867;
wire n_17475;
wire n_17363;
wire n_4656;
wire n_3839;
wire n_8497;
wire n_10770;
wire n_6410;
wire n_17873;
wire n_4915;
wire n_15592;
wire n_16064;
wire n_18524;
wire n_15319;
wire n_235;
wire n_5662;
wire n_3730;
wire n_14452;
wire n_17894;
wire n_13464;
wire n_12670;
wire n_16817;
wire n_18336;
wire n_7667;
wire n_10203;
wire n_10980;
wire n_9174;
wire n_17835;
wire n_2737;
wire n_17459;
wire n_10082;
wire n_7182;
wire n_7365;
wire n_10467;
wire n_9849;
wire n_1622;
wire n_17476;
wire n_9856;
wire n_18449;
wire n_17591;
wire n_18672;
wire n_18848;
wire n_11668;
wire n_7885;
wire n_15684;
wire n_2171;
wire n_16720;
wire n_9349;
wire n_17423;
wire n_3136;
wire n_11091;
wire n_4192;
wire n_10940;
wire n_16463;
wire n_15976;
wire n_2808;
wire n_18100;
wire n_17723;
wire n_8839;
wire n_4174;
wire n_12891;
wire n_11615;
wire n_1171;
wire n_11059;
wire n_16403;
wire n_1827;
wire n_14616;
wire n_16799;
wire n_2187;
wire n_6058;
wire n_17965;
wire n_7745;
wire n_12941;
wire n_2872;
wire n_14258;
wire n_12200;
wire n_14024;
wire n_2046;
wire n_17212;
wire n_8684;
wire n_13682;
wire n_6249;
wire n_11060;
wire n_5480;
wire n_18943;
wire n_4831;
wire n_11461;
wire n_10714;
wire n_6969;
wire n_7459;
wire n_6161;
wire n_2970;
wire n_8206;
wire n_18070;
wire n_2882;
wire n_4260;
wire n_18338;
wire n_6607;
wire n_9335;
wire n_1974;
wire n_4122;
wire n_9452;
wire n_11427;
wire n_19293;
wire n_934;
wire n_5284;
wire n_12673;
wire n_14694;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_19208;
wire n_9427;
wire n_17817;
wire n_6294;
wire n_543;
wire n_9611;
wire n_18371;
wire n_9021;
wire n_16269;
wire n_9250;
wire n_11212;
wire n_13145;
wire n_804;
wire n_9550;
wire n_16591;
wire n_11263;
wire n_10641;
wire n_959;
wire n_4312;
wire n_18805;
wire n_16566;
wire n_13195;
wire n_8694;
wire n_13965;
wire n_5048;
wire n_11994;
wire n_13358;
wire n_2195;
wire n_3208;
wire n_18759;
wire n_16693;
wire n_14519;
wire n_6123;
wire n_11000;
wire n_16125;
wire n_4935;
wire n_19403;
wire n_8191;
wire n_10325;
wire n_16354;
wire n_10298;
wire n_6922;
wire n_16701;
wire n_7698;
wire n_12854;
wire n_16427;
wire n_16336;
wire n_8431;
wire n_19631;
wire n_2945;
wire n_3061;
wire n_16248;
wire n_3932;
wire n_3469;
wire n_2960;
wire n_10400;
wire n_19081;
wire n_9177;
wire n_9060;
wire n_11947;
wire n_14496;
wire n_9096;
wire n_13952;
wire n_11697;
wire n_16963;
wire n_18074;
wire n_7891;
wire n_14413;
wire n_8517;
wire n_3008;
wire n_4776;
wire n_4153;
wire n_11034;
wire n_10901;
wire n_10549;
wire n_12115;
wire n_1962;
wire n_11499;
wire n_10825;
wire n_4723;
wire n_17292;
wire n_4269;
wire n_18023;
wire n_14777;
wire n_14057;
wire n_5459;
wire n_17788;
wire n_4143;
wire n_876;
wire n_16406;
wire n_12558;
wire n_11984;
wire n_11948;
wire n_4719;
wire n_7477;
wire n_17028;
wire n_15654;
wire n_1904;
wire n_17289;
wire n_2588;
wire n_11402;
wire n_1353;
wire n_11401;
wire n_17828;
wire n_17820;
wire n_2366;
wire n_10581;
wire n_14949;
wire n_17487;
wire n_4423;
wire n_2210;
wire n_3602;
wire n_18372;
wire n_12086;
wire n_1411;
wire n_16952;
wire n_566;
wire n_16449;
wire n_2951;
wire n_11589;
wire n_11246;
wire n_1807;
wire n_18266;
wire n_16606;
wire n_14460;
wire n_13216;
wire n_209;
wire n_12849;
wire n_11312;
wire n_13786;
wire n_5909;
wire n_9344;
wire n_671;
wire n_10865;
wire n_740;
wire n_10738;
wire n_7378;
wire n_9798;
wire n_15491;
wire n_14925;
wire n_11612;
wire n_4229;
wire n_12447;
wire n_13417;
wire n_12296;
wire n_13414;
wire n_3865;
wire n_4073;
wire n_5400;
wire n_7498;
wire n_3846;
wire n_11916;
wire n_180;
wire n_3512;
wire n_7501;
wire n_5201;
wire n_10421;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_12764;
wire n_15325;
wire n_1326;
wire n_4783;
wire n_18987;
wire n_19091;
wire n_14238;
wire n_16918;
wire n_12409;
wire n_11625;
wire n_1130;
wire n_17054;
wire n_6592;
wire n_9712;
wire n_8585;
wire n_6626;
wire n_14042;
wire n_9220;
wire n_17312;
wire n_12763;
wire n_378;
wire n_18460;
wire n_17272;
wire n_16394;
wire n_18869;
wire n_15310;
wire n_17989;
wire n_1283;
wire n_4917;
wire n_8698;
wire n_12584;
wire n_14435;
wire n_4432;
wire n_10376;
wire n_15510;
wire n_7515;
wire n_17567;
wire n_344;
wire n_9994;
wire n_14226;
wire n_7309;
wire n_15811;
wire n_5114;
wire n_1392;
wire n_8559;
wire n_5693;
wire n_17670;
wire n_15618;
wire n_2463;
wire n_10224;
wire n_15849;
wire n_611;
wire n_18758;
wire n_3062;
wire n_2679;
wire n_9391;
wire n_16105;
wire n_8514;
wire n_9134;
wire n_14159;
wire n_14515;
wire n_12268;
wire n_18990;
wire n_12077;
wire n_15321;
wire n_14757;
wire n_1017;
wire n_5396;
wire n_12534;
wire n_6846;
wire n_13271;
wire n_11481;
wire n_10175;
wire n_15812;
wire n_16292;
wire n_18458;
wire n_6886;
wire n_17019;
wire n_5365;
wire n_8405;
wire n_15223;
wire n_11350;
wire n_626;
wire n_11925;
wire n_16033;
wire n_8672;
wire n_1104;
wire n_4920;
wire n_1253;
wire n_6446;
wire n_3256;
wire n_7218;
wire n_19279;
wire n_9430;
wire n_11407;
wire n_2118;
wire n_19548;
wire n_12710;
wire n_19331;
wire n_2188;
wire n_8440;
wire n_7005;
wire n_9776;
wire n_16736;
wire n_6777;
wire n_18156;
wire n_11987;
wire n_18208;
wire n_19206;
wire n_8475;
wire n_8029;
wire n_18845;
wire n_18527;
wire n_4861;
wire n_4064;
wire n_1829;
wire n_13089;
wire n_15459;
wire n_15192;
wire n_5266;
wire n_4828;
wire n_1638;
wire n_18360;
wire n_16836;
wire n_13167;
wire n_12329;
wire n_519;
wire n_15013;
wire n_6953;
wire n_3669;
wire n_16710;
wire n_14945;
wire n_4316;
wire n_5122;
wire n_5390;
wire n_18660;
wire n_18348;
wire n_19658;
wire n_18487;
wire n_9834;
wire n_16353;
wire n_2047;
wire n_12318;
wire n_5385;
wire n_13278;
wire n_13597;
wire n_5322;
wire n_3989;
wire n_7089;
wire n_2490;
wire n_18232;
wire n_3841;
wire n_1996;
wire n_6332;
wire n_1442;
wire n_7403;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_4909;
wire n_13938;
wire n_13251;
wire n_8566;
wire n_7343;
wire n_12766;
wire n_18913;
wire n_8317;
wire n_12229;
wire n_269;
wire n_6116;
wire n_7492;
wire n_13319;
wire n_9071;
wire n_10415;
wire n_7694;
wire n_11711;
wire n_18637;
wire n_15666;
wire n_11931;
wire n_8109;
wire n_2055;
wire n_18971;
wire n_12780;
wire n_13267;
wire n_14017;
wire n_7987;
wire n_9133;
wire n_16054;
wire n_12664;
wire n_14942;
wire n_7434;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_15359;
wire n_9063;
wire n_7787;
wire n_1494;
wire n_2325;
wire n_1850;
wire n_5304;
wire n_15035;
wire n_18500;
wire n_19085;
wire n_18536;
wire n_6261;
wire n_4281;
wire n_4648;
wire n_10096;
wire n_13617;
wire n_10025;
wire n_412;
wire n_18779;
wire n_6299;
wire n_11753;
wire n_7425;
wire n_19061;
wire n_1059;
wire n_11150;
wire n_18199;
wire n_4360;
wire n_16111;
wire n_3263;
wire n_6316;
wire n_6292;
wire n_9726;
wire n_1748;
wire n_13884;
wire n_17125;
wire n_7719;
wire n_5615;
wire n_6220;
wire n_12783;
wire n_1885;
wire n_1240;
wire n_17671;
wire n_1234;
wire n_14195;
wire n_18363;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_3152;
wire n_7935;
wire n_8458;
wire n_6772;
wire n_16902;
wire n_16646;
wire n_14300;
wire n_6077;
wire n_1003;
wire n_11512;
wire n_17090;
wire n_14678;
wire n_13599;
wire n_17282;
wire n_15008;
wire n_5188;
wire n_13647;
wire n_4490;
wire n_13683;
wire n_1575;
wire n_19094;
wire n_10147;
wire n_17921;
wire n_17197;
wire n_18503;
wire n_9298;
wire n_18058;
wire n_16939;
wire n_14497;
wire n_1991;
wire n_5161;
wire n_14280;
wire n_4078;
wire n_13724;
wire n_9301;
wire n_3046;
wire n_5382;
wire n_12054;
wire n_15827;
wire n_5659;
wire n_17256;
wire n_8099;
wire n_11595;
wire n_17806;
wire n_13768;
wire n_1415;
wire n_16707;
wire n_8578;
wire n_1370;
wire n_7222;
wire n_13838;
wire n_10046;
wire n_2291;
wire n_2184;
wire n_10397;
wire n_2982;
wire n_19379;
wire n_10936;
wire n_12442;
wire n_8611;
wire n_1517;
wire n_8819;
wire n_17927;
wire n_2630;
wire n_15123;
wire n_9835;
wire n_15021;
wire n_12839;
wire n_6697;
wire n_13153;
wire n_7875;
wire n_7643;
wire n_13441;
wire n_16082;
wire n_13857;
wire n_10207;
wire n_18872;
wire n_1143;
wire n_10401;
wire n_19352;
wire n_7242;
wire n_17737;
wire n_19240;
wire n_13816;
wire n_18355;
wire n_2013;
wire n_17215;
wire n_14736;
wire n_10139;
wire n_13246;
wire n_14061;
wire n_12986;
wire n_11381;
wire n_16378;
wire n_16109;
wire n_7224;
wire n_12441;
wire n_15789;
wire n_16611;
wire n_16172;
wire n_7746;
wire n_3662;
wire n_2981;
wire n_18108;
wire n_16277;
wire n_16598;
wire n_17588;
wire n_12516;
wire n_8414;
wire n_13921;
wire n_6297;
wire n_16806;
wire n_6653;
wire n_15512;
wire n_18836;
wire n_12377;
wire n_638;
wire n_18486;
wire n_5492;
wire n_9965;
wire n_13650;
wire n_16789;
wire n_887;
wire n_15636;
wire n_15946;
wire n_6501;
wire n_18063;
wire n_9990;
wire n_10005;
wire n_12905;
wire n_11426;
wire n_2599;
wire n_15311;
wire n_8505;
wire n_3368;
wire n_17667;
wire n_7884;
wire n_11258;
wire n_15498;
wire n_7417;
wire n_18097;
wire n_4881;
wire n_12513;
wire n_5734;
wire n_13395;
wire n_4255;
wire n_4071;
wire n_7388;
wire n_3568;
wire n_11657;
wire n_8717;
wire n_5770;
wire n_5705;
wire n_3313;
wire n_9064;
wire n_17420;
wire n_2725;
wire n_14135;
wire n_16482;
wire n_8571;
wire n_4305;
wire n_12514;
wire n_10048;
wire n_16809;
wire n_14194;
wire n_619;
wire n_13825;
wire n_18942;
wire n_8243;
wire n_6347;
wire n_9593;
wire n_606;
wire n_13398;
wire n_8449;
wire n_17605;
wire n_630;
wire n_13204;
wire n_4094;
wire n_14331;
wire n_18994;
wire n_4765;
wire n_2522;
wire n_4364;
wire n_9406;
wire n_8967;
wire n_9322;
wire n_15017;
wire n_5959;
wire n_3720;
wire n_8031;
wire n_15591;
wire n_264;
wire n_12188;
wire n_16609;
wire n_4745;
wire n_5642;
wire n_9232;
wire n_15167;
wire n_12299;
wire n_16739;
wire n_15706;
wire n_1680;
wire n_3842;
wire n_993;
wire n_1605;
wire n_11327;
wire n_4979;
wire n_1988;
wire n_15900;
wire n_12000;
wire n_17281;
wire n_19004;
wire n_1233;
wire n_14182;
wire n_241;
wire n_10279;
wire n_15853;
wire n_4520;
wire n_5299;
wire n_3455;
wire n_14352;
wire n_13889;
wire n_17864;
wire n_7081;
wire n_13015;
wire n_7319;
wire n_15831;
wire n_7644;
wire n_11176;
wire n_9883;
wire n_11135;
wire n_5668;
wire n_11275;
wire n_268;
wire n_18850;
wire n_5463;
wire n_12700;
wire n_12904;
wire n_5489;
wire n_1165;
wire n_14623;
wire n_4773;
wire n_7910;
wire n_6009;
wire n_3281;
wire n_9034;
wire n_7084;
wire n_5923;
wire n_14073;
wire n_8074;
wire n_13639;
wire n_15989;
wire n_8860;
wire n_2676;
wire n_3940;
wire n_1214;
wire n_15514;
wire n_9266;
wire n_3453;
wire n_3410;
wire n_16210;
wire n_10027;
wire n_12784;
wire n_1813;
wire n_18639;
wire n_825;
wire n_12877;
wire n_14261;
wire n_14677;
wire n_18020;
wire n_10616;
wire n_8587;
wire n_5366;
wire n_16016;
wire n_15550;
wire n_15528;
wire n_6925;
wire n_6878;
wire n_9078;
wire n_16297;
wire n_16896;
wire n_13198;
wire n_15914;
wire n_3289;
wire n_13741;
wire n_12610;
wire n_14416;
wire n_11251;
wire n_12293;
wire n_2036;
wire n_6470;
wire n_11598;
wire n_8368;
wire n_15691;
wire n_17560;
wire n_8322;
wire n_16127;
wire n_6187;
wire n_8300;
wire n_9378;
wire n_678;
wire n_12206;
wire n_18112;
wire n_17488;
wire n_17427;
wire n_11400;
wire n_19532;
wire n_6693;
wire n_15848;
wire n_11563;
wire n_362;
wire n_12444;
wire n_18586;
wire n_16409;
wire n_5419;
wire n_14513;
wire n_2943;
wire n_12778;
wire n_12485;
wire n_3253;
wire n_15995;
wire n_14602;
wire n_11468;
wire n_16150;
wire n_4603;
wire n_9683;
wire n_17403;
wire n_15132;
wire n_1527;
wire n_495;
wire n_5732;
wire n_11878;
wire n_15843;
wire n_16666;
wire n_4471;
wire n_15749;
wire n_7449;
wire n_15638;
wire n_16547;
wire n_14289;
wire n_1493;
wire n_16479;
wire n_10751;
wire n_16967;
wire n_10240;
wire n_10691;
wire n_2535;
wire n_9561;
wire n_19351;
wire n_16104;
wire n_9773;
wire n_2436;
wire n_3838;
wire n_9745;
wire n_3941;
wire n_15413;
wire n_10216;
wire n_15628;
wire n_17733;
wire n_1514;
wire n_10150;
wire n_12581;
wire n_17395;
wire n_4994;
wire n_6652;
wire n_10971;
wire n_5168;
wire n_4661;
wire n_18506;
wire n_7674;
wire n_14516;
wire n_18484;
wire n_12305;
wire n_12170;
wire n_2853;
wire n_9630;
wire n_13927;
wire n_13313;
wire n_15308;
wire n_17025;
wire n_9255;
wire n_10231;
wire n_8310;
wire n_16500;
wire n_9758;
wire n_15175;
wire n_8936;
wire n_18413;
wire n_7126;
wire n_15206;
wire n_9691;
wire n_12997;
wire n_14005;
wire n_14293;
wire n_14334;
wire n_7690;
wire n_15245;
wire n_15225;
wire n_3229;
wire n_11223;
wire n_13562;
wire n_14537;
wire n_6950;
wire n_10038;
wire n_17794;
wire n_15614;
wire n_2012;
wire n_5066;
wire n_18101;
wire n_2842;
wire n_19087;
wire n_11221;
wire n_15772;
wire n_14245;
wire n_17659;
wire n_11448;
wire n_17321;
wire n_18272;
wire n_1809;
wire n_8328;
wire n_15502;
wire n_15076;
wire n_12576;
wire n_7258;
wire n_10579;
wire n_13345;
wire n_3677;
wire n_8336;
wire n_3996;
wire n_17492;
wire n_19324;
wire n_4218;
wire n_11445;
wire n_13151;
wire n_3685;
wire n_11552;
wire n_15102;
wire n_14733;
wire n_417;
wire n_14317;
wire n_4459;
wire n_16220;
wire n_9852;
wire n_11623;
wire n_3019;
wire n_3471;
wire n_5295;
wire n_2368;
wire n_18599;
wire n_14131;
wire n_10676;
wire n_8041;
wire n_17931;
wire n_4175;
wire n_10299;
wire n_10540;
wire n_16993;
wire n_12845;
wire n_11645;
wire n_10200;
wire n_3259;
wire n_2524;
wire n_13164;
wire n_2460;
wire n_13662;
wire n_3867;
wire n_3593;
wire n_1073;
wire n_16275;
wire n_17062;
wire n_13340;
wire n_17887;
wire n_17192;
wire n_4140;
wire n_2481;
wire n_9939;
wire n_7766;
wire n_19397;
wire n_12797;
wire n_6758;
wire n_5160;
wire n_9481;
wire n_17081;
wire n_7955;
wire n_1207;
wire n_12012;
wire n_7287;
wire n_10076;
wire n_880;
wire n_6464;
wire n_18675;
wire n_3540;
wire n_11554;
wire n_150;
wire n_1478;
wire n_3777;
wire n_4203;
wire n_767;
wire n_1837;
wire n_4533;
wire n_9635;
wire n_19619;
wire n_1410;
wire n_14308;
wire n_5408;
wire n_1736;
wire n_3848;
wire n_319;
wire n_8181;
wire n_2511;
wire n_8254;
wire n_13452;
wire n_8071;
wire n_5271;
wire n_17480;
wire n_562;
wire n_5964;
wire n_6004;
wire n_11628;
wire n_1136;
wire n_11549;
wire n_17162;
wire n_12286;
wire n_9001;
wire n_19517;
wire n_2329;
wire n_16107;
wire n_14545;
wire n_18031;
wire n_8013;
wire n_146;
wire n_193;
wire n_16683;
wire n_17804;
wire n_12347;
wire n_19346;
wire n_17424;
wire n_296;
wire n_651;
wire n_3407;
wire n_5992;
wire n_217;
wire n_1185;
wire n_19394;
wire n_215;
wire n_17818;
wire n_12698;
wire n_2621;
wire n_6540;
wire n_16086;
wire n_5513;
wire n_5614;
wire n_497;
wire n_17383;
wire n_11871;
wire n_16857;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_15326;
wire n_17555;
wire n_18957;
wire n_7722;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_4056;
wire n_9240;
wire n_8293;
wire n_14726;
wire n_14180;
wire n_18697;
wire n_10548;
wire n_12957;
wire n_11616;
wire n_8791;
wire n_8288;
wire n_1091;
wire n_1425;
wire n_12786;
wire n_983;
wire n_10678;
wire n_6757;
wire n_17752;
wire n_18045;
wire n_1390;
wire n_2289;
wire n_8323;
wire n_10391;
wire n_13176;
wire n_9784;
wire n_19647;
wire n_7990;
wire n_18368;
wire n_10036;
wire n_17631;
wire n_5278;
wire n_14905;
wire n_15128;
wire n_3688;
wire n_8720;
wire n_12205;
wire n_11989;
wire n_16912;
wire n_16215;
wire n_1905;
wire n_14009;
wire n_3466;
wire n_5704;
wire n_15787;
wire n_7148;
wire n_5956;
wire n_9417;
wire n_2139;
wire n_12020;
wire n_18875;
wire n_6835;
wire n_1203;
wire n_11624;
wire n_8826;
wire n_15083;
wire n_11352;
wire n_19290;
wire n_5516;
wire n_2841;
wire n_6247;
wire n_11234;
wire n_10919;
wire n_12099;
wire n_12858;
wire n_4399;
wire n_15351;
wire n_2487;
wire n_18170;
wire n_19159;
wire n_7544;
wire n_9336;
wire n_3572;
wire n_8854;
wire n_6645;
wire n_16177;
wire n_10727;
wire n_10885;
wire n_443;
wire n_13201;
wire n_14759;
wire n_13274;
wire n_18621;
wire n_9312;
wire n_5174;
wire n_7469;
wire n_5538;
wire n_5017;
wire n_10895;
wire n_198;
wire n_11977;
wire n_15576;
wire n_11696;
wire n_11734;
wire n_9533;
wire n_9494;
wire n_5241;
wire n_11507;
wire n_17290;
wire n_15337;
wire n_17276;
wire n_14749;
wire n_7082;
wire n_18731;
wire n_3108;
wire n_19306;
wire n_11320;
wire n_11837;
wire n_19458;
wire n_8260;
wire n_3417;
wire n_13898;
wire n_16507;
wire n_4124;
wire n_16543;
wire n_11938;
wire n_6418;
wire n_17003;
wire n_5153;
wire n_18814;
wire n_609;
wire n_10571;
wire n_19202;
wire n_19664;
wire n_9807;
wire n_9057;
wire n_8706;
wire n_2607;
wire n_7945;
wire n_8894;
wire n_19244;
wire n_2890;
wire n_12053;
wire n_15947;
wire n_17738;
wire n_12619;
wire n_1320;
wire n_11289;
wire n_13555;
wire n_2499;
wire n_12582;
wire n_5487;
wire n_18919;
wire n_12423;
wire n_15426;
wire n_14137;
wire n_16905;
wire n_17765;
wire n_14163;
wire n_15523;
wire n_2472;
wire n_7328;
wire n_19298;
wire n_10958;
wire n_15682;
wire n_9479;
wire n_15556;
wire n_3957;
wire n_14041;
wire n_18622;
wire n_9181;
wire n_19338;
wire n_19385;
wire n_6578;
wire n_3040;
wire n_14763;
wire n_19319;
wire n_17686;
wire n_18381;
wire n_10879;
wire n_19481;
wire n_5951;
wire n_6589;
wire n_1864;
wire n_10639;
wire n_16359;
wire n_3475;
wire n_17448;
wire n_18657;
wire n_16037;
wire n_13351;
wire n_9276;
wire n_579;
wire n_5152;
wire n_16805;
wire n_15937;
wire n_16141;
wire n_5574;
wire n_4927;
wire n_9821;
wire n_11112;
wire n_4258;
wire n_2699;
wire n_11723;
wire n_650;
wire n_16647;
wire n_1940;
wire n_1405;
wire n_5469;
wire n_14393;
wire n_456;
wire n_12364;
wire n_3878;
wire n_12420;
wire n_6567;
wire n_313;
wire n_5895;
wire n_5804;
wire n_9508;
wire n_3134;
wire n_16231;
wire n_896;
wire n_4553;
wire n_3278;
wire n_17805;
wire n_17318;
wire n_11906;
wire n_2673;
wire n_2456;
wire n_14298;
wire n_9741;
wire n_1637;
wire n_3307;
wire n_1407;
wire n_2871;
wire n_420;
wire n_10180;
wire n_4183;
wire n_14112;
wire n_10650;
wire n_12120;
wire n_12021;
wire n_10157;
wire n_7423;
wire n_10402;
wire n_12515;
wire n_17283;
wire n_9166;
wire n_1640;
wire n_12895;
wire n_12045;
wire n_2141;
wire n_6940;
wire n_12726;
wire n_12668;
wire n_7835;
wire n_15437;
wire n_6320;
wire n_799;
wire n_3044;
wire n_9969;
wire n_11437;
wire n_14068;
wire n_14853;
wire n_16735;
wire n_11869;
wire n_5620;
wire n_10836;
wire n_159;
wire n_16375;
wire n_2125;
wire n_8072;
wire n_13117;
wire n_7130;
wire n_2992;
wire n_1241;
wire n_3221;
wire n_11282;
wire n_17720;
wire n_14700;
wire n_16382;
wire n_7491;
wire n_1706;
wire n_18944;
wire n_18474;
wire n_4052;
wire n_9636;
wire n_7559;
wire n_13175;
wire n_2441;
wire n_9833;
wire n_9095;
wire n_15757;
wire n_18465;
wire n_5907;
wire n_15979;
wire n_19076;
wire n_1559;
wire n_6731;
wire n_4315;
wire n_2888;
wire n_6154;
wire n_6943;
wire n_4301;
wire n_3744;
wire n_12038;
wire n_8210;
wire n_12644;
wire n_1360;
wire n_11826;
wire n_18241;
wire n_3781;
wire n_10888;
wire n_2484;
wire n_10116;
wire n_16764;
wire n_14808;
wire n_2126;
wire n_18135;
wire n_3843;
wire n_11764;
wire n_6600;
wire n_817;
wire n_14140;
wire n_5402;
wire n_10696;
wire n_7355;
wire n_18688;
wire n_9331;
wire n_10170;
wire n_6031;
wire n_14479;
wire n_8331;
wire n_3216;
wire n_332;
wire n_1882;
wire n_18109;
wire n_14172;
wire n_7270;
wire n_591;
wire n_18721;
wire n_5417;
wire n_6967;
wire n_19241;
wire n_6742;
wire n_18117;
wire n_13525;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_14997;
wire n_15931;
wire n_6691;
wire n_14799;
wire n_10689;
wire n_13909;
wire n_6172;
wire n_19062;
wire n_12634;
wire n_14774;
wire n_12680;
wire n_11613;
wire n_10233;
wire n_751;
wire n_15492;
wire n_18443;
wire n_17343;
wire n_4652;
wire n_10810;
wire n_12176;
wire n_10311;
wire n_9140;
wire n_2163;
wire n_18533;
wire n_2815;
wire n_19427;
wire n_4577;
wire n_4748;
wire n_337;
wire n_5814;
wire n_12094;
wire n_3231;
wire n_9736;
wire n_2979;
wire n_5531;
wire n_12517;
wire n_6517;
wire n_18431;
wire n_15441;
wire n_9225;
wire n_17353;
wire n_2946;
wire n_12071;
wire n_11923;
wire n_13832;
wire n_3430;
wire n_2269;
wire n_8105;
wire n_9031;
wire n_4225;
wire n_19406;
wire n_13087;
wire n_13972;
wire n_15436;
wire n_17920;
wire n_15633;
wire n_2565;
wire n_12339;
wire n_10602;
wire n_16630;
wire n_14632;
wire n_5655;
wire n_15969;
wire n_6393;
wire n_8154;
wire n_2175;
wire n_2182;
wire n_13849;
wire n_11131;
wire n_10778;
wire n_17961;
wire n_13258;
wire n_1506;
wire n_3473;
wire n_957;
wire n_1994;
wire n_9014;
wire n_13166;
wire n_8509;
wire n_6364;
wire n_16754;
wire n_15482;
wire n_16217;
wire n_19467;
wire n_11003;
wire n_6061;
wire n_18132;
wire n_12723;
wire n_14097;
wire n_18741;
wire n_2685;
wire n_8372;
wire n_17042;
wire n_10088;
wire n_14887;
wire n_7225;
wire n_8077;
wire n_18530;
wire n_16948;
wire n_6755;
wire n_18934;
wire n_2265;
wire n_13762;
wire n_13037;
wire n_11573;
wire n_4409;
wire n_7509;
wire n_10145;
wire n_14225;
wire n_11005;
wire n_4629;
wire n_6255;
wire n_18611;
wire n_4638;
wire n_6840;
wire n_17675;
wire n_8423;
wire n_9577;
wire n_19149;
wire n_12589;
wire n_14143;
wire n_6488;
wire n_904;
wire n_8337;
wire n_709;
wire n_7164;
wire n_14044;
wire n_17431;
wire n_3868;
wire n_18249;
wire n_18561;
wire n_18134;
wire n_17000;
wire n_12699;
wire n_1085;
wire n_12927;
wire n_2042;
wire n_16588;
wire n_771;
wire n_8199;
wire n_17456;
wire n_1149;
wire n_8656;
wire n_265;
wire n_14909;
wire n_10918;
wire n_13122;
wire n_2592;
wire n_15553;
wire n_2666;
wire n_1585;
wire n_12663;
wire n_1799;
wire n_2564;
wire n_16349;
wire n_17165;
wire n_15841;
wire n_17623;
wire n_4259;
wire n_2035;
wire n_11127;
wire n_18083;
wire n_7134;
wire n_4572;
wire n_9547;
wire n_4104;
wire n_16350;
wire n_8346;
wire n_8761;
wire n_15458;
wire n_9085;
wire n_13734;
wire n_8226;
wire n_17532;
wire n_7079;
wire n_9084;
wire n_5928;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_3219;
wire n_14051;
wire n_17680;
wire n_9889;
wire n_12375;
wire n_12556;
wire n_2010;
wire n_1198;
wire n_13723;
wire n_10168;
wire n_2174;
wire n_12156;
wire n_13128;
wire n_13490;
wire n_4727;
wire n_4594;
wire n_17663;
wire n_14913;
wire n_10621;
wire n_9731;
wire n_6572;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_15382;
wire n_4051;
wire n_7755;
wire n_16031;
wire n_6080;
wire n_4865;
wire n_8387;
wire n_12076;
wire n_10613;
wire n_6717;
wire n_7473;
wire n_11359;
wire n_19404;
wire n_19064;
wire n_15997;
wire n_19562;
wire n_10561;
wire n_19335;
wire n_14695;
wire n_16251;
wire n_13212;
wire n_16978;
wire n_15166;
wire n_18304;
wire n_15138;
wire n_16516;
wire n_18517;
wire n_2879;
wire n_17533;
wire n_14405;
wire n_967;
wire n_7038;
wire n_14081;
wire n_4341;
wire n_1819;
wire n_8177;
wire n_17616;
wire n_12025;
wire n_8962;
wire n_9538;
wire n_14254;
wire n_16137;
wire n_6145;
wire n_6539;
wire n_6926;
wire n_13421;
wire n_1632;
wire n_13495;
wire n_13474;
wire n_14903;
wire n_13949;
wire n_12383;
wire n_11912;
wire n_4973;
wire n_14967;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3950;
wire n_9423;
wire n_16619;
wire n_2927;
wire n_4750;
wire n_12962;
wire n_18823;
wire n_16263;
wire n_11666;
wire n_12459;
wire n_2166;
wire n_2899;
wire n_7105;
wire n_14500;
wire n_13568;
wire n_10140;
wire n_12612;
wire n_16369;
wire n_5903;
wire n_17213;
wire n_5986;
wire n_3065;
wire n_6710;
wire n_1423;
wire n_18326;
wire n_19402;
wire n_17664;
wire n_4959;
wire n_9056;
wire n_4426;
wire n_12496;
wire n_12814;
wire n_3002;
wire n_649;
wire n_15943;
wire n_18714;
wire n_11921;
wire n_8495;
wire n_14532;
wire n_8783;
wire n_14557;
wire n_1199;
wire n_12603;
wire n_15392;
wire n_14340;
wire n_18444;
wire n_14032;
wire n_16944;
wire n_15702;
wire n_7262;
wire n_212;
wire n_3773;
wire n_12967;
wire n_14899;
wire n_12232;
wire n_18115;
wire n_18847;
wire n_11859;
wire n_15773;
wire n_798;
wire n_15307;
wire n_14111;
wire n_6719;
wire n_13580;
wire n_7178;
wire n_9553;
wire n_11633;
wire n_7506;
wire n_8551;
wire n_14361;
wire n_12760;
wire n_18291;
wire n_2647;
wire n_19633;
wire n_14943;
wire n_4578;
wire n_4777;
wire n_2672;
wire n_12590;
wire n_2299;
wire n_15605;
wire n_5871;
wire n_18951;
wire n_7142;
wire n_12577;
wire n_17711;
wire n_10182;
wire n_16813;
wire n_13928;
wire n_19342;
wire n_7125;
wire n_1172;
wire n_11655;
wire n_3626;
wire n_2313;
wire n_12069;
wire n_16899;
wire n_15656;
wire n_18455;
wire n_16957;
wire n_10317;
wire n_4029;
wire n_375;
wire n_12270;
wire n_4617;
wire n_16021;
wire n_9196;
wire n_4010;
wire n_1649;
wire n_5882;
wire n_5650;
wire n_6057;
wire n_14555;
wire n_10893;
wire n_1572;
wire n_5021;
wire n_9251;
wire n_9973;
wire n_11117;
wire n_8064;
wire n_8468;
wire n_4325;
wire n_3251;
wire n_10201;
wire n_2212;
wire n_12210;
wire n_8778;
wire n_17106;
wire n_14168;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_15342;
wire n_15534;
wire n_10539;
wire n_14080;
wire n_5625;
wire n_11777;
wire n_17402;
wire n_4919;
wire n_3737;
wire n_13975;
wire n_5969;
wire n_10121;
wire n_8198;
wire n_19054;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_12189;
wire n_1211;
wire n_9270;
wire n_14142;
wire n_6041;
wire n_9099;
wire n_7350;
wire n_10814;
wire n_5276;
wire n_16034;
wire n_9627;
wire n_17008;
wire n_16563;
wire n_6664;
wire n_196;
wire n_17575;
wire n_2985;
wire n_13131;
wire n_14941;
wire n_1446;
wire n_3938;
wire n_11154;
wire n_3507;
wire n_11700;
wire n_5855;
wire n_3531;
wire n_16128;
wire n_10975;
wire n_1054;
wire n_9460;
wire n_17698;
wire n_11652;
wire n_14320;
wire n_11056;
wire n_19229;
wire n_6238;
wire n_13932;
wire n_2397;
wire n_16804;
wire n_3931;
wire n_15606;
wire n_10459;
wire n_2113;
wire n_1918;
wire n_5429;
wire n_6545;
wire n_11583;
wire n_15866;
wire n_9766;
wire n_4163;
wire n_10463;
wire n_14764;
wire n_645;
wire n_7074;
wire n_8734;
wire n_2633;
wire n_12564;
wire n_19443;
wire n_13433;
wire n_15505;
wire n_10403;
wire n_7037;
wire n_13697;
wire n_11784;
wire n_5298;
wire n_9025;
wire n_3396;
wire n_14244;
wire n_7928;
wire n_12886;
wire n_6532;
wire n_821;
wire n_4372;
wire n_7293;
wire n_18638;
wire n_13000;
wire n_14362;
wire n_5640;
wire n_15996;
wire n_408;
wire n_4318;
wire n_6721;
wire n_18825;
wire n_2123;
wire n_3716;
wire n_6108;
wire n_8258;
wire n_10370;
wire n_18537;
wire n_9597;
wire n_11892;
wire n_5744;
wire n_5384;
wire n_3248;
wire n_15731;
wire n_8299;
wire n_12473;
wire n_4032;
wire n_1064;
wire n_11421;
wire n_1396;
wire n_18704;
wire n_11966;
wire n_19530;
wire n_17450;
wire n_18011;
wire n_12748;
wire n_4337;
wire n_16829;
wire n_3092;
wire n_9692;
wire n_7395;
wire n_13402;
wire n_3734;
wire n_17305;
wire n_18047;
wire n_7078;
wire n_8188;
wire n_2580;
wire n_13831;
wire n_16792;
wire n_18572;
wire n_11423;
wire n_1875;
wire n_1865;
wire n_5701;
wire n_18378;
wire n_9567;
wire n_9061;
wire n_3419;
wire n_1297;
wire n_17154;
wire n_16922;
wire n_8664;
wire n_922;
wire n_16552;
wire n_16867;
wire n_16638;
wire n_14783;
wire n_13268;
wire n_10740;
wire n_10457;
wire n_19042;
wire n_17968;
wire n_1896;
wire n_3058;
wire n_14158;
wire n_9701;
wire n_675;
wire n_19247;
wire n_14236;
wire n_1540;
wire n_18849;
wire n_13510;
wire n_14640;
wire n_6659;
wire n_9709;
wire n_242;
wire n_9295;
wire n_4371;
wire n_2994;
wire n_3689;
wire n_16678;
wire n_10264;
wire n_5850;
wire n_15029;
wire n_14286;
wire n_12528;
wire n_17640;
wire n_6182;
wire n_12717;
wire n_6520;
wire n_12660;
wire n_3918;
wire n_1965;
wire n_2476;
wire n_17662;
wire n_17651;
wire n_598;
wire n_11547;
wire n_13520;
wire n_8501;
wire n_10301;
wire n_3271;
wire n_295;
wire n_4248;
wire n_13018;
wire n_18240;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_15139;
wire n_8076;
wire n_6826;
wire n_1792;
wire n_11395;
wire n_9107;
wire n_19630;
wire n_3809;
wire n_11279;
wire n_18370;
wire n_11724;
wire n_11789;
wire n_14152;
wire n_3139;
wire n_14869;
wire n_19354;
wire n_881;
wire n_8014;
wire n_19030;
wire n_7768;
wire n_8638;
wire n_16294;
wire n_4018;
wire n_14651;
wire n_694;
wire n_7982;
wire n_8804;
wire n_297;
wire n_3337;
wire n_11383;
wire n_1044;
wire n_2165;
wire n_15882;
wire n_17740;
wire n_6879;
wire n_17059;
wire n_7567;
wire n_8433;
wire n_6074;
wire n_4588;
wire n_585;
wire n_10932;
wire n_10619;
wire n_1756;
wire n_5411;
wire n_17263;
wire n_9156;
wire n_16113;
wire n_16848;
wire n_1968;
wire n_4728;
wire n_4385;
wire n_18749;
wire n_10248;
wire n_9748;
wire n_3616;
wire n_13365;
wire n_7771;
wire n_11780;
wire n_6027;
wire n_5695;
wire n_2870;
wire n_16289;
wire n_2151;
wire n_7701;
wire n_16342;
wire n_1839;
wire n_17278;
wire n_5235;
wire n_6720;
wire n_11930;
wire n_6888;
wire n_826;
wire n_3747;
wire n_12628;
wire n_8122;
wire n_17095;
wire n_13444;
wire n_16504;
wire n_8432;
wire n_4330;
wire n_7592;
wire n_14209;
wire n_19462;
wire n_18651;
wire n_5311;
wire n_6590;
wire n_3522;
wire n_2747;
wire n_18243;
wire n_791;
wire n_11876;
wire n_5572;
wire n_19110;
wire n_7151;
wire n_8950;
wire n_18683;
wire n_10758;
wire n_2861;
wire n_13431;
wire n_3975;
wire n_1838;
wire n_4683;
wire n_12538;
wire n_14025;
wire n_7758;
wire n_13779;
wire n_12446;
wire n_2316;
wire n_15954;
wire n_9355;
wire n_5060;
wire n_15386;
wire n_4986;
wire n_14620;
wire n_5888;
wire n_15349;
wire n_9582;
wire n_2208;
wire n_5884;
wire n_11009;
wire n_9288;
wire n_6308;
wire n_7897;
wire n_17701;
wire n_7118;
wire n_2134;
wire n_8284;
wire n_9702;
wire n_18767;
wire n_15378;
wire n_7422;
wire n_1431;
wire n_17881;
wire n_3835;
wire n_6738;
wire n_12307;
wire n_8703;
wire n_15839;
wire n_16135;
wire n_17661;
wire n_14999;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_19377;
wire n_3557;
wire n_2610;
wire n_3620;
wire n_13720;
wire n_478;
wire n_7339;
wire n_3832;
wire n_13706;
wire n_13903;
wire n_9051;
wire n_3693;
wire n_8545;
wire n_10385;
wire n_10105;
wire n_2372;
wire n_1490;
wire n_15785;
wire n_19056;
wire n_3674;
wire n_2959;
wire n_17114;
wire n_10251;
wire n_15234;
wire n_293;
wire n_18796;
wire n_1070;
wire n_2403;
wire n_4700;
wire n_17524;
wire n_9980;
wire n_14394;
wire n_4224;
wire n_18679;
wire n_6005;
wire n_17261;
wire n_9555;
wire n_14845;
wire n_1358;
wire n_7713;
wire n_4564;
wire n_15372;
wire n_13560;
wire n_15700;
wire n_16182;
wire n_2424;
wire n_3201;
wire n_19239;
wire n_1475;
wire n_10304;
wire n_3103;
wire n_5860;
wire n_6936;
wire n_15934;
wire n_16827;
wire n_16121;
wire n_7487;
wire n_9986;
wire n_527;
wire n_13794;
wire n_3627;
wire n_13537;
wire n_9397;
wire n_18616;
wire n_1137;
wire n_3612;
wire n_17574;
wire n_4695;
wire n_9855;
wire n_10568;
wire n_2966;
wire n_2294;
wire n_13463;
wire n_600;
wire n_9496;
wire n_16241;
wire n_10796;
wire n_10016;
wire n_10030;
wire n_12864;
wire n_9653;
wire n_10272;
wire n_8989;
wire n_9640;
wire n_1339;
wire n_13936;
wire n_13933;
wire n_7815;
wire n_403;
wire n_7934;
wire n_3244;
wire n_11578;
wire n_6865;
wire n_1141;
wire n_7276;
wire n_18595;
wire n_1755;
wire n_5043;
wire n_8739;
wire n_17078;
wire n_6747;
wire n_13714;
wire n_2025;
wire n_12725;
wire n_6640;
wire n_16030;
wire n_2250;
wire n_3033;
wire n_16079;
wire n_11908;
wire n_18166;
wire n_6462;
wire n_17372;
wire n_6034;
wire n_13159;
wire n_9781;
wire n_418;
wire n_14788;
wire n_13287;
wire n_11913;
wire n_7034;
wire n_1618;
wire n_4867;
wire n_13389;
wire n_17726;
wire n_1653;
wire n_9906;
wire n_4237;
wire n_5029;
wire n_12317;
wire n_13302;
wire n_10092;
wire n_6833;
wire n_6793;
wire n_16766;
wire n_17834;
wire n_11815;
wire n_6295;
wire n_3386;
wire n_11231;
wire n_463;
wire n_13740;
wire n_17966;
wire n_19278;
wire n_8137;
wire n_12027;
wire n_3205;
wire n_15218;
wire n_17366;
wire n_19114;
wire n_17514;
wire n_7014;
wire n_17975;
wire n_10430;
wire n_16697;
wire n_8305;
wire n_18147;
wire n_1636;
wire n_4001;
wire n_18751;
wire n_6709;
wire n_17525;
wire n_960;
wire n_6712;
wire n_7416;
wire n_778;
wire n_14553;
wire n_5177;
wire n_9657;
wire n_16594;
wire n_16370;
wire n_6743;
wire n_16223;
wire n_1610;
wire n_12412;
wire n_11880;
wire n_5785;
wire n_14528;
wire n_4583;
wire n_9485;
wire n_13940;
wire n_2515;
wire n_11249;
wire n_15449;
wire n_4054;
wire n_10119;
wire n_11986;
wire n_14798;
wire n_5966;
wire n_3349;
wire n_17579;
wire n_368;
wire n_12118;
wire n_14409;
wire n_14724;
wire n_18451;
wire n_14291;
wire n_1020;
wire n_8625;
wire n_4214;
wire n_6919;
wire n_13756;
wire n_7805;
wire n_10995;
wire n_9192;
wire n_1138;
wire n_5752;
wire n_11618;
wire n_14266;
wire n_12594;
wire n_8179;
wire n_19360;
wire n_11861;
wire n_8511;
wire n_6973;
wire n_12081;
wire n_4413;
wire n_7453;
wire n_10684;
wire n_2381;
wire n_18095;
wire n_2052;
wire n_5081;
wire n_15039;
wire n_17929;
wire n_17027;
wire n_8806;
wire n_17400;
wire n_19234;
wire n_6619;
wire n_16434;
wire n_5189;
wire n_13930;
wire n_8149;
wire n_3041;
wire n_603;
wire n_10390;
wire n_1657;
wire n_7210;
wire n_5869;
wire n_2439;
wire n_2404;
wire n_6718;
wire n_4238;
wire n_3011;
wire n_15400;
wire n_2061;
wire n_17411;
wire n_16866;
wire n_15485;
wire n_18499;
wire n_18789;
wire n_14841;
wire n_16726;
wire n_13624;
wire n_5632;
wire n_5425;
wire n_18603;
wire n_19480;
wire n_8269;
wire n_13805;
wire n_18786;
wire n_3650;
wire n_8968;
wire n_16243;
wire n_7855;
wire n_14029;
wire n_4590;
wire n_3137;
wire n_14056;
wire n_5678;
wire n_13695;
wire n_6981;
wire n_13288;
wire n_19465;
wire n_16917;
wire n_3238;
wire n_218;
wire n_11519;
wire n_13065;
wire n_11229;
wire n_18655;
wire n_16159;
wire n_17570;
wire n_11397;
wire n_12840;
wire n_5437;
wire n_12846;
wire n_14705;
wire n_17660;
wire n_8401;
wire n_7854;
wire n_10577;
wire n_11324;
wire n_12945;
wire n_5307;
wire n_17385;
wire n_10151;
wire n_6439;
wire n_2446;
wire n_8240;
wire n_12850;
wire n_7714;
wire n_16193;
wire n_2017;
wire n_3029;
wire n_3597;
wire n_9305;
wire n_9999;
wire n_17495;
wire n_1121;
wire n_11361;
wire n_1963;
wire n_6945;
wire n_18617;
wire n_3790;
wire n_7029;
wire n_19009;
wire n_10186;
wire n_17236;
wire n_11841;
wire n_6618;
wire n_14453;
wire n_17545;
wire n_13094;
wire n_7317;
wire n_17558;
wire n_3977;
wire n_227;
wire n_9461;
wire n_6816;
wire n_10928;
wire n_5008;
wire n_6502;
wire n_6250;
wire n_6288;
wire n_5974;
wire n_7522;
wire n_4133;
wire n_9618;
wire n_6118;
wire n_18961;
wire n_4561;
wire n_464;
wire n_11808;
wire n_17970;
wire n_13257;
wire n_17160;
wire n_18778;
wire n_4239;
wire n_18509;
wire n_4184;
wire n_17636;
wire n_1830;
wire n_13393;
wire n_6251;
wire n_9828;
wire n_3915;
wire n_13922;
wire n_13423;
wire n_18149;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_2293;
wire n_10252;
wire n_16641;
wire n_11555;
wire n_6869;
wire n_3102;
wire n_14625;
wire n_10345;
wire n_2026;
wire n_10059;
wire n_8325;
wire n_7621;
wire n_7359;
wire n_550;
wire n_3321;
wire n_2322;
wire n_12394;
wire n_4782;
wire n_13578;
wire n_19540;
wire n_14204;
wire n_9005;
wire n_4378;
wire n_8274;
wire n_12954;
wire n_4876;
wire n_6146;
wire n_8504;
wire n_10464;
wire n_14688;
wire n_10644;
wire n_12801;
wire n_18594;
wire n_13708;
wire n_10365;
wire n_11781;
wire n_9648;
wire n_2653;
wire n_12965;
wire n_12788;
wire n_9498;
wire n_15707;
wire n_16328;
wire n_3156;
wire n_15396;
wire n_15909;
wire n_672;
wire n_3483;
wire n_11884;
wire n_19516;
wire n_13371;
wire n_4493;
wire n_7971;
wire n_743;
wire n_12264;
wire n_8232;
wire n_9649;
wire n_8904;
wire n_16977;
wire n_19287;
wire n_10629;
wire n_660;
wire n_7070;
wire n_8382;
wire n_4421;
wire n_18950;
wire n_2839;
wire n_4793;
wire n_13856;
wire n_15607;
wire n_15879;
wire n_7259;
wire n_12274;
wire n_14588;
wire n_2944;
wire n_8128;
wire n_15746;
wire n_3831;
wire n_15921;
wire n_19545;
wire n_5932;
wire n_5830;
wire n_11345;
wire n_12380;
wire n_13245;
wire n_12586;
wire n_3391;
wire n_8794;
wire n_11760;
wire n_19203;
wire n_1463;
wire n_4505;
wire n_17222;
wire n_1826;
wire n_5126;
wire n_8205;
wire n_9907;
wire n_13088;
wire n_6976;
wire n_13538;
wire n_11024;
wire n_18437;
wire n_6304;
wire n_5236;
wire n_7640;
wire n_13701;
wire n_10498;
wire n_11424;
wire n_12585;
wire n_5012;
wire n_14021;
wire n_1256;
wire n_10635;
wire n_13626;
wire n_19218;
wire n_12832;
wire n_8067;
wire n_12301;
wire n_9643;
wire n_4630;
wire n_18973;
wire n_18402;
wire n_15822;
wire n_11881;
wire n_14980;
wire n_2109;
wire n_7727;
wire n_18968;
wire n_11935;
wire n_17561;
wire n_18766;
wire n_1204;
wire n_18901;
wire n_233;
wire n_8719;
wire n_16140;
wire n_19223;
wire n_18046;
wire n_2787;
wire n_15493;
wire n_12615;
wire n_13357;
wire n_10802;
wire n_17148;
wire n_769;
wire n_4786;
wire n_7565;
wire n_16624;
wire n_7631;
wire n_13869;
wire n_16903;
wire n_7387;
wire n_9212;
wire n_12167;
wire n_9473;
wire n_13026;
wire n_10490;
wire n_15019;
wire n_13499;
wire n_17107;
wire n_14843;
wire n_2736;
wire n_10647;
wire n_3493;
wire n_9320;
wire n_10523;
wire n_16781;
wire n_12298;
wire n_10081;
wire n_3774;
wire n_12569;
wire n_2910;
wire n_14929;
wire n_18497;
wire n_5148;
wire n_2584;
wire n_866;
wire n_12456;
wire n_8655;
wire n_17039;
wire n_10808;
wire n_6333;
wire n_8745;
wire n_5791;
wire n_18504;
wire n_8086;
wire n_15466;
wire n_13943;
wire n_17124;
wire n_7379;
wire n_17530;
wire n_8901;
wire n_11078;
wire n_8695;
wire n_4911;
wire n_8173;
wire n_12072;
wire n_4436;
wire n_10545;
wire n_1174;
wire n_17945;
wire n_16557;
wire n_14141;
wire n_5602;
wire n_647;
wire n_9379;
wire n_11992;
wire n_15790;
wire n_844;
wire n_17061;
wire n_14880;
wire n_13142;
wire n_13180;
wire n_3584;
wire n_10453;
wire n_16975;
wire n_3556;
wire n_16716;
wire n_13785;
wire n_5831;
wire n_7742;
wire n_9274;
wire n_3456;
wire n_10331;
wire n_11439;
wire n_14655;
wire n_17230;
wire n_12863;
wire n_10352;
wire n_19449;
wire n_1122;
wire n_4059;
wire n_16830;
wire n_1109;
wire n_17851;
wire n_3309;
wire n_8507;
wire n_8415;
wire n_2609;
wire n_10713;
wire n_6680;
wire n_10954;
wire n_7432;
wire n_16036;
wire n_13978;
wire n_13941;
wire n_15339;
wire n_13439;
wire n_228;
wire n_16152;
wire n_14133;
wire n_14433;
wire n_13187;
wire n_13162;
wire n_2600;
wire n_7505;
wire n_18521;
wire n_15059;
wire n_8244;
wire n_7494;
wire n_18380;
wire n_4353;
wire n_735;
wire n_17071;
wire n_13661;
wire n_9546;
wire n_7589;
wire n_17764;
wire n_4346;
wire n_4351;
wire n_11296;
wire n_13770;
wire n_18636;
wire n_8723;
wire n_13511;
wire n_18016;
wire n_11019;
wire n_980;
wire n_7843;
wire n_1651;
wire n_19544;
wire n_4784;
wire n_19258;
wire n_14569;
wire n_7902;
wire n_1685;
wire n_6496;
wire n_3066;
wire n_15744;
wire n_7756;
wire n_2844;
wire n_15557;
wire n_18244;
wire n_8342;
wire n_8940;
wire n_14154;
wire n_8472;
wire n_4332;
wire n_810;
wire n_10000;
wire n_12812;
wire n_7988;
wire n_14174;
wire n_7500;
wire n_10246;
wire n_3198;
wire n_18236;
wire n_14269;
wire n_9822;
wire n_13991;
wire n_17523;
wire n_14821;
wire n_17330;
wire n_15096;
wire n_5272;
wire n_14992;
wire n_10125;
wire n_9065;
wire n_16637;
wire n_3218;
wire n_18627;
wire n_9086;
wire n_9153;
wire n_10505;
wire n_582;
wire n_861;
wire n_11064;
wire n_6908;
wire n_8237;
wire n_9093;
wire n_2968;
wire n_4201;
wire n_7266;
wire n_19046;
wire n_17928;
wire n_8046;
wire n_5646;
wire n_13284;
wire n_4852;
wire n_4210;
wire n_16521;
wire n_2709;
wire n_9198;
wire n_8335;
wire n_9142;
wire n_17697;
wire n_15820;
wire n_18239;
wire n_5214;
wire n_15486;
wire n_9493;
wire n_19371;
wire n_11330;
wire n_12720;
wire n_7794;
wire n_19139;
wire n_13318;
wire n_15917;
wire n_1274;
wire n_3333;
wire n_6605;
wire n_12687;
wire n_18278;
wire n_17510;
wire n_19106;
wire n_13208;
wire n_13867;
wire n_15594;
wire n_17807;
wire n_17841;
wire n_5380;
wire n_5776;
wire n_11796;
wire n_18339;
wire n_16881;
wire n_12789;
wire n_2677;
wire n_12127;
wire n_17232;
wire n_3283;
wire n_16976;
wire n_14119;
wire n_13673;
wire n_8037;
wire n_1742;
wire n_16775;
wire n_12573;
wire n_2542;
wire n_1671;
wire n_19400;
wire n_15214;
wire n_13045;
wire n_741;
wire n_1351;
wire n_17347;
wire n_18684;
wire n_6806;
wire n_13146;
wire n_13235;
wire n_15125;
wire n_5019;
wire n_2332;
wire n_5138;
wire n_4388;
wire n_6960;
wire n_3089;
wire n_8169;
wire n_12265;
wire n_783;
wire n_5409;
wire n_5301;
wire n_17777;
wire n_188;
wire n_1854;
wire n_3222;
wire n_7504;
wire n_15971;
wire n_442;
wire n_11678;
wire n_8023;
wire n_12251;
wire n_1975;
wire n_16307;
wire n_8130;
wire n_16911;
wire n_15294;
wire n_5055;
wire n_18676;
wire n_16288;
wire n_7116;
wire n_4249;
wire n_17992;
wire n_6999;
wire n_14741;
wire n_11046;
wire n_11079;
wire n_5548;
wire n_15581;
wire n_11065;
wire n_8339;
wire n_19058;
wire n_14215;
wire n_17368;
wire n_852;
wire n_544;
wire n_5900;
wire n_4273;
wire n_18104;
wire n_8499;
wire n_15356;
wire n_18525;
wire n_6882;
wire n_10775;
wire n_2129;
wire n_9526;
wire n_17511;
wire n_18762;
wire n_15571;
wire n_7983;
wire n_10863;
wire n_4997;
wire n_2399;
wire n_4843;
wire n_1232;
wire n_17138;
wire n_17700;
wire n_13993;
wire n_10986;
wire n_8366;
wire n_8102;
wire n_19126;
wire n_18087;
wire n_8022;
wire n_17226;
wire n_19212;
wire n_10262;
wire n_5239;
wire n_1781;
wire n_10239;
wire n_14577;
wire n_5332;
wire n_14984;
wire n_2004;
wire n_1106;
wire n_18183;
wire n_8913;
wire n_155;
wire n_4956;
wire n_16772;
wire n_14699;
wire n_454;
wire n_10335;
wire n_15362;
wire n_5129;
wire n_11301;
wire n_15101;
wire n_5070;
wire n_18154;
wire n_11703;
wire n_6374;
wire n_17013;
wire n_6628;
wire n_13483;
wire n_18923;
wire n_4262;
wire n_16551;
wire n_17803;
wire n_1894;
wire n_6570;
wire n_8556;
wire n_8040;
wire n_11821;
wire n_13121;
wire n_13989;
wire n_10755;
wire n_16998;
wire n_15200;
wire n_17349;
wire n_10682;
wire n_3928;
wire n_6371;
wire n_8079;
wire n_2613;
wire n_3535;
wire n_8595;
wire n_2708;
wire n_1648;
wire n_2011;
wire n_5684;
wire n_15887;
wire n_10022;
wire n_5729;
wire n_13803;
wire n_14066;
wire n_7856;
wire n_564;
wire n_6148;
wire n_7625;
wire n_686;
wire n_1641;
wire n_3871;
wire n_12775;
wire n_6989;
wire n_7863;
wire n_8958;
wire n_12833;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_13687;
wire n_7623;
wire n_7217;
wire n_1699;
wire n_14540;
wire n_16784;
wire n_8115;
wire n_608;
wire n_2101;
wire n_9398;
wire n_15320;
wire n_3484;
wire n_4677;
wire n_12915;
wire n_6196;
wire n_13149;
wire n_18748;
wire n_2616;
wire n_5275;
wire n_14091;
wire n_15755;
wire n_8412;
wire n_2811;
wire n_6485;
wire n_14478;
wire n_17848;
wire n_10177;
wire n_6107;
wire n_16689;
wire n_11944;
wire n_1075;
wire n_7796;
wire n_6994;
wire n_15986;
wire n_14570;
wire n_16068;
wire n_13797;
wire n_13013;
wire n_13238;
wire n_4810;
wire n_175;
wire n_9446;
wire n_11129;
wire n_7234;
wire n_3914;
wire n_8119;
wire n_10296;
wire n_8641;
wire n_12988;
wire n_17136;
wire n_13344;
wire n_11139;
wire n_17766;
wire n_12685;
wire n_8436;
wire n_14239;
wire n_8659;
wire n_14045;
wire n_19575;
wire n_4369;
wire n_7849;
wire n_12667;
wire n_18747;
wire n_15635;
wire n_4331;
wire n_7297;
wire n_10018;
wire n_15183;
wire n_4972;
wire n_4993;
wire n_15118;
wire n_7298;
wire n_5536;
wire n_9129;
wire n_10141;
wire n_14162;
wire n_8224;
wire n_2678;
wire n_15679;
wire n_4613;
wire n_13014;
wire n_1167;
wire n_2428;
wire n_10897;
wire n_210;
wire n_10449;
wire n_7861;
wire n_14303;
wire n_7039;
wire n_11349;
wire n_5046;
wire n_2749;
wire n_3273;
wire n_7077;
wire n_12540;
wire n_19160;
wire n_5305;
wire n_4681;
wire n_13239;
wire n_15942;
wire n_17583;
wire n_4752;
wire n_18552;
wire n_9143;
wire n_8287;
wire n_2092;
wire n_7950;
wire n_8607;
wire n_2514;
wire n_604;
wire n_17032;
wire n_6248;
wire n_16768;
wire n_16134;
wire n_10452;
wire n_7806;
wire n_3942;
wire n_15928;
wire n_16092;
wire n_7595;
wire n_8066;
wire n_5795;
wire n_12349;
wire n_14282;
wire n_5552;
wire n_6715;
wire n_6714;
wire n_11308;
wire n_890;
wire n_16266;
wire n_8416;
wire n_4518;
wire n_14167;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_10363;
wire n_2252;
wire n_13623;
wire n_11511;
wire n_15833;
wire n_16046;
wire n_760;
wire n_15974;
wire n_9393;
wire n_13845;
wire n_12709;
wire n_13432;
wire n_12771;
wire n_17760;
wire n_1858;
wire n_14787;
wire n_19502;
wire n_7303;
wire n_3021;
wire n_17100;
wire n_6616;
wire n_10781;
wire n_7315;
wire n_9886;
wire n_1164;
wire n_13244;
wire n_4288;
wire n_18969;
wire n_6185;
wire n_5529;
wire n_3733;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_13843;
wire n_17191;
wire n_13404;
wire n_3614;
wire n_874;
wire n_382;
wire n_5183;
wire n_18689;
wire n_7268;
wire n_4228;
wire n_3423;
wire n_10094;
wire n_16295;
wire n_10084;
wire n_19259;
wire n_13870;
wire n_13791;
wire n_3644;
wire n_6955;
wire n_2706;
wire n_1127;
wire n_1512;
wire n_9932;
wire n_16745;
wire n_320;
wire n_13900;
wire n_16224;
wire n_14652;
wire n_1139;
wire n_3179;
wire n_8741;
wire n_4000;
wire n_2897;
wire n_3970;
wire n_7232;
wire n_7377;
wire n_19461;
wire n_996;
wire n_16132;
wire n_19425;
wire n_6646;
wire n_15149;
wire n_14844;
wire n_16907;
wire n_14391;
wire n_6033;
wire n_11541;
wire n_15495;
wire n_4873;
wire n_9801;
wire n_19312;
wire n_3782;
wire n_8773;
wire n_6369;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_581;
wire n_7542;
wire n_5636;
wire n_13213;
wire n_12231;
wire n_989;
wire n_17643;
wire n_8410;
wire n_14756;
wire n_18144;
wire n_7739;
wire n_4939;
wire n_19474;
wire n_14384;
wire n_15905;
wire n_5530;
wire n_2473;
wire n_12552;
wire n_11069;
wire n_2539;
wire n_4123;
wire n_5595;
wire n_9941;
wire n_16795;
wire n_17131;
wire n_3119;
wire n_3735;
wire n_11369;
wire n_4379;
wire n_14210;
wire n_486;
wire n_5388;
wire n_4718;
wire n_15788;
wire n_13362;
wire n_5962;
wire n_7010;
wire n_648;
wire n_9728;
wire n_16690;
wire n_2057;
wire n_7219;
wire n_9662;
wire n_12896;
wire n_15694;
wire n_8774;
wire n_18690;
wire n_19494;
wire n_7299;
wire n_4872;
wire n_9936;
wire n_6195;
wire n_9530;
wire n_14692;
wire n_7471;
wire n_10455;
wire n_15488;
wire n_5300;
wire n_11393;
wire n_7741;
wire n_5035;
wire n_9466;
wire n_16525;
wire n_7790;
wire n_16315;
wire n_19283;
wire n_6149;
wire n_17918;
wire n_7002;
wire n_12428;
wire n_3025;
wire n_1626;
wire n_15814;
wire n_1388;
wire n_10265;
wire n_16676;
wire n_18736;
wire n_15756;
wire n_19495;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_11995;
wire n_14378;
wire n_18299;
wire n_11371;
wire n_5394;
wire n_14191;
wire n_19267;
wire n_16546;
wire n_18252;
wire n_17454;
wire n_16144;
wire n_16669;
wire n_474;
wire n_6902;
wire n_3331;
wire n_10100;
wire n_18607;
wire n_5741;
wire n_15743;
wire n_2773;
wire n_7478;
wire n_19587;
wire n_19130;
wire n_5405;
wire n_7456;
wire n_13600;
wire n_964;
wire n_8503;
wire n_4756;
wire n_8196;
wire n_16062;
wire n_17712;
wire n_10846;
wire n_9787;
wire n_13363;
wire n_19648;
wire n_4970;
wire n_211;
wire n_9786;
wire n_18681;
wire n_14908;
wire n_2292;
wire n_12908;
wire n_18692;
wire n_3441;
wire n_17168;
wire n_2416;
wire n_311;
wire n_14201;
wire n_8923;
wire n_13315;
wire n_18900;
wire n_6736;
wire n_19231;
wire n_1769;
wire n_14597;
wire n_15663;
wire n_3605;
wire n_4633;
wire n_3306;
wire n_9115;
wire n_4584;
wire n_3090;
wire n_11833;
wire n_3724;
wire n_4276;
wire n_11897;
wire n_2990;
wire n_1773;
wire n_5001;
wire n_5176;
wire n_7443;
wire n_11285;
wire n_3323;
wire n_9977;
wire n_8051;
wire n_16719;
wire n_518;
wire n_9242;
wire n_4618;
wire n_4679;
wire n_914;
wire n_11262;
wire n_4496;
wire n_12880;
wire n_4805;
wire n_8651;
wire n_13959;
wire n_3454;
wire n_10732;
wire n_6885;
wire n_10851;
wire n_10221;
wire n_3547;
wire n_9299;
wire n_11162;
wire n_13685;
wire n_3816;
wire n_14693;
wire n_8842;
wire n_3214;
wire n_16915;
wire n_1917;
wire n_14486;
wire n_1580;
wire n_7730;
wire n_11592;
wire n_15090;
wire n_8467;
wire n_17043;
wire n_15385;
wire n_3109;
wire n_16094;
wire n_2863;
wire n_6417;
wire n_13281;
wire n_1731;
wire n_5648;
wire n_15627;
wire n_2135;
wire n_4707;
wire n_1832;
wire n_10996;
wire n_858;
wire n_8676;
wire n_9853;
wire n_13192;
wire n_7448;
wire n_17170;
wire n_19045;
wire n_410;
wire n_17351;
wire n_18060;
wire n_1594;
wire n_15048;
wire n_16393;
wire n_17135;
wire n_6199;
wire n_9823;
wire n_15739;
wire n_12937;
wire n_10698;
wire n_16891;
wire n_18118;
wire n_14665;
wire n_6726;
wire n_580;
wire n_7011;
wire n_5261;
wire n_10870;
wire n_11066;
wire n_17327;
wire n_4252;
wire n_13886;
wire n_16887;
wire n_6576;
wire n_2448;
wire n_8906;
wire n_17117;
wire n_8482;
wire n_7952;
wire n_16242;
wire n_14489;
wire n_13774;
wire n_13847;
wire n_6915;
wire n_19645;
wire n_12529;
wire n_12103;
wire n_7834;
wire n_17072;
wire n_5185;
wire n_8409;
wire n_17889;
wire n_974;
wire n_14053;
wire n_5023;
wire n_2656;
wire n_4952;
wire n_19321;
wire n_5906;
wire n_8930;
wire n_16564;
wire n_14581;
wire n_628;
wire n_18811;
wire n_1573;
wire n_7890;
wire n_3973;
wire n_11950;
wire n_6024;
wire n_12461;
wire n_485;
wire n_11415;
wire n_7265;
wire n_7986;
wire n_17809;
wire n_2024;
wire n_17900;
wire n_202;
wire n_9879;
wire n_1749;
wire n_18744;
wire n_3474;
wire n_11390;
wire n_17238;
wire n_11669;
wire n_1669;
wire n_1024;
wire n_14712;
wire n_15717;
wire n_5556;
wire n_8250;
wire n_10601;
wire n_9158;
wire n_18591;
wire n_1667;
wire n_16945;
wire n_7717;
wire n_9518;
wire n_18187;
wire n_18462;
wire n_18260;
wire n_5143;
wire n_11739;
wire n_10497;
wire n_14561;
wire n_18405;
wire n_1639;
wire n_13301;
wire n_8298;
wire n_466;
wire n_5215;
wire n_7860;
wire n_14212;
wire n_2548;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_13158;
wire n_1108;
wire n_11044;
wire n_15967;
wire n_15530;
wire n_1601;
wire n_11679;
wire n_8450;
wire n_17665;
wire n_3648;
wire n_17799;
wire n_7499;
wire n_3042;
wire n_7292;
wire n_12398;
wire n_17089;
wire n_5433;
wire n_9043;
wire n_6075;
wire n_7397;
wire n_10789;
wire n_17020;
wire n_12705;
wire n_1430;
wire n_1316;
wire n_7977;
wire n_12847;
wire n_13047;
wire n_6861;
wire n_14470;
wire n_15497;
wire n_7847;
wire n_15952;
wire n_13178;
wire n_3723;
wire n_18609;
wire n_1190;
wire n_12404;
wire n_397;
wire n_11606;
wire n_5978;
wire n_11452;
wire n_15734;
wire n_6217;
wire n_5031;
wire n_10797;
wire n_7289;
wire n_17656;
wire n_14110;
wire n_14806;
wire n_1673;
wire n_7354;
wire n_18312;
wire n_13824;
wire n_3424;
wire n_239;
wire n_7960;
wire n_15620;
wire n_2326;
wire n_18053;
wire n_12912;
wire n_12211;
wire n_6115;
wire n_13377;
wire n_2120;
wire n_16493;
wire n_6048;
wire n_6416;
wire n_2964;
wire n_352;
wire n_6838;
wire n_10068;
wire n_11988;
wire n_3485;
wire n_4077;
wire n_1361;
wire n_19034;
wire n_6256;
wire n_15645;
wire n_6613;
wire n_11438;
wire n_15965;
wire n_5221;
wire n_5641;
wire n_18877;
wire n_6361;
wire n_14981;
wire n_11348;
wire n_9685;
wire n_11685;
wire n_5731;
wire n_6678;
wire n_8662;
wire n_15058;
wire n_16539;
wire n_14971;
wire n_12429;
wire n_14734;
wire n_14494;
wire n_14956;
wire n_4623;
wire n_7325;
wire n_14866;
wire n_19123;
wire n_5007;
wire n_3320;
wire n_6370;
wire n_9923;
wire n_13743;
wire n_7166;
wire n_7356;
wire n_13378;
wire n_11319;
wire n_3476;
wire n_16981;
wire n_5629;
wire n_3439;
wire n_7873;
wire n_2688;
wire n_1489;
wire n_16418;
wire n_19363;
wire n_17795;
wire n_12640;
wire n_10063;
wire n_13092;
wire n_2852;
wire n_14292;
wire n_8419;
wire n_1496;
wire n_19497;
wire n_9862;
wire n_11385;
wire n_1485;
wire n_11355;
wire n_18659;
wire n_11674;
wire n_1846;
wire n_12535;
wire n_19031;
wire n_12327;
wire n_879;
wire n_2310;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_8430;
wire n_15719;
wire n_12058;
wire n_14879;
wire n_16143;
wire n_18387;
wire n_5852;
wire n_15164;
wire n_7052;
wire n_16755;
wire n_10496;
wire n_5960;
wire n_14149;
wire n_2454;
wire n_18225;
wire n_5321;
wire n_9960;
wire n_157;
wire n_4215;
wire n_10998;
wire n_19180;
wire n_7502;
wire n_1484;
wire n_14216;
wire n_16380;
wire n_3752;
wire n_7919;
wire n_10800;
wire n_17962;
wire n_7085;
wire n_1373;
wire n_12065;
wire n_3958;
wire n_13950;
wire n_18952;
wire n_5210;
wire n_13732;
wire n_16422;
wire n_14968;
wire n_10993;
wire n_15542;
wire n_14985;
wire n_15910;
wire n_17734;
wire n_14443;
wire n_1047;
wire n_3899;
wire n_16136;
wire n_14285;
wire n_1385;
wire n_9734;
wire n_7288;
wire n_16325;
wire n_16842;
wire n_17355;
wire n_4987;
wire n_10495;
wire n_9004;
wire n_834;
wire n_3818;
wire n_6610;
wire n_3124;
wire n_10612;
wire n_1741;
wire n_10260;
wire n_12285;
wire n_6750;
wire n_9150;
wire n_14508;
wire n_15092;
wire n_12683;
wire n_18535;
wire n_2614;
wire n_18457;
wire n_3694;
wire n_14566;
wire n_2937;
wire n_7869;
wire n_7165;
wire n_13386;
wire n_13846;
wire n_4376;
wire n_7683;
wire n_16437;
wire n_9587;
wire n_1076;
wire n_10671;
wire n_10193;
wire n_1377;
wire n_11718;
wire n_19333;
wire n_695;
wire n_14383;
wire n_16695;
wire n_4081;
wire n_11680;
wire n_14683;
wire n_18685;
wire n_17052;
wire n_7322;
wire n_17378;
wire n_11658;
wire n_12226;
wire n_13492;
wire n_14001;
wire n_5562;
wire n_15397;
wire n_978;
wire n_15840;
wire n_7880;
wire n_4382;
wire n_749;
wire n_16855;
wire n_19120;
wire n_16937;
wire n_2140;
wire n_9919;
wire n_12135;
wire n_19485;
wire n_5577;
wire n_568;
wire n_17092;
wire n_8829;
wire n_19308;
wire n_13381;
wire n_739;
wire n_5413;
wire n_8971;
wire n_18076;
wire n_16667;
wire n_1338;
wire n_16897;
wire n_10558;
wire n_9579;
wire n_9475;
wire n_17603;
wire n_15273;
wire n_573;
wire n_9049;
wire n_13718;
wire n_18701;
wire n_4480;
wire n_14775;
wire n_18809;
wire n_11045;
wire n_16756;
wire n_222;
wire n_11340;
wire n_16965;
wire n_7675;
wire n_11903;
wire n_13279;
wire n_13644;
wire n_13291;
wire n_742;
wire n_691;
wire n_10174;
wire n_377;
wire n_7524;
wire n_2935;
wire n_15897;
wire n_4046;
wire n_11564;
wire n_14015;
wire n_8925;
wire n_12946;
wire n_16729;
wire n_18406;
wire n_13513;
wire n_4027;
wire n_12916;
wire n_1227;
wire n_3520;
wire n_8471;
wire n_12521;
wire n_18925;
wire n_9800;
wire n_11382;
wire n_19578;
wire n_10098;
wire n_11745;
wire n_1570;
wire n_15240;
wire n_1780;
wire n_15564;
wire n_1347;
wire n_17002;
wire n_14350;
wire n_7733;
wire n_17405;
wire n_18711;
wire n_4631;
wire n_19090;
wire n_1561;
wire n_13773;
wire n_14109;
wire n_6982;
wire n_2168;
wire n_5847;
wire n_7345;
wire n_17526;
wire n_14136;
wire n_10923;
wire n_7385;
wire n_5159;
wire n_2615;
wire n_14176;
wire n_4625;
wire n_11149;
wire n_12635;
wire n_3962;
wire n_8488;
wire n_9543;
wire n_11443;
wire n_15765;
wire n_6855;
wire n_18176;
wire n_3362;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_4188;
wire n_13467;
wire n_3667;
wire n_712;
wire n_18374;
wire n_18700;
wire n_7907;
wire n_5568;
wire n_6312;
wire n_11532;
wire n_2505;
wire n_9415;
wire n_4115;
wire n_14343;
wire n_18619;
wire n_9147;
wire n_470;
wire n_11209;
wire n_3680;
wire n_15918;
wire n_5723;
wire n_5918;
wire n_16212;
wire n_11790;
wire n_1972;
wire n_19189;
wire n_4491;
wire n_19444;
wire n_363;
wire n_18148;
wire n_16313;
wire n_10420;
wire n_17058;
wire n_18309;
wire n_16363;
wire n_503;
wire n_6131;
wire n_15232;
wire n_12105;
wire n_14329;
wire n_19392;
wire n_15721;
wire n_5163;
wire n_307;
wire n_10444;
wire n_3361;
wire n_11377;
wire n_3478;
wire n_8018;
wire n_18557;
wire n_7937;
wire n_9176;
wire n_7819;
wire n_10631;
wire n_7305;
wire n_6334;
wire n_16780;
wire n_3096;
wire n_2651;
wire n_8884;
wire n_5537;
wire n_19222;
wire n_1574;
wire n_253;
wire n_2918;
wire n_8751;
wire n_4307;
wire n_11864;
wire n_11006;
wire n_15018;
wire n_6617;
wire n_3552;
wire n_7511;
wire n_6533;
wire n_849;
wire n_4091;
wire n_14108;
wire n_1753;
wire n_3095;
wire n_15439;
wire n_16049;
wire n_2807;
wire n_8178;
wire n_14000;
wire n_14372;
wire n_3618;
wire n_4758;
wire n_17911;
wire n_12046;
wire n_10212;
wire n_18566;
wire n_5335;
wire n_12917;
wire n_14629;
wire n_9425;
wire n_11172;
wire n_10089;
wire n_14947;
wire n_5505;
wire n_8560;
wire n_14748;
wire n_18895;
wire n_18466;
wire n_10004;
wire n_12488;
wire n_3852;
wire n_1365;
wire n_11110;
wire n_17338;
wire n_16211;
wire n_15001;
wire n_3896;
wire n_8674;
wire n_5274;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_13328;
wire n_4093;
wire n_10892;
wire n_18556;
wire n_10493;
wire n_19195;
wire n_10405;
wire n_15037;
wire n_4794;
wire n_17386;
wire n_7964;
wire n_17091;
wire n_629;
wire n_14349;
wire n_6278;
wire n_7022;
wire n_12691;
wire n_11033;
wire n_19072;
wire n_18203;
wire n_14356;
wire n_19028;
wire n_5581;
wire n_16926;
wire n_16006;
wire n_992;
wire n_12651;
wire n_19194;
wire n_16476;
wire n_7486;
wire n_6756;
wire n_16373;
wire n_18792;
wire n_14190;
wire n_8563;
wire n_17223;
wire n_15546;
wire n_11534;
wire n_14157;
wire n_14344;
wire n_9221;
wire n_509;
wire n_1209;
wire n_7906;
wire n_5248;
wire n_6411;
wire n_350;
wire n_10285;
wire n_4370;
wire n_14488;
wire n_11032;
wire n_2359;
wire n_13582;
wire n_142;
wire n_17950;
wire n_7302;
wire n_18162;
wire n_11174;
wire n_18574;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_18544;
wire n_10294;
wire n_4359;
wire n_10106;
wire n_17865;
wire n_9934;
wire n_3487;
wire n_287;
wire n_9234;
wire n_10674;
wire n_6534;
wire n_3340;
wire n_230;
wire n_5227;
wire n_16011;
wire n_6265;
wire n_2989;
wire n_5778;
wire n_18185;
wire n_8087;
wire n_7607;
wire n_14458;
wire n_17540;
wire n_12073;
wire n_13655;
wire n_6898;
wire n_6596;
wire n_13565;
wire n_14643;
wire n_10249;
wire n_8361;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_522;
wire n_18965;
wire n_3440;
wire n_13784;
wire n_13468;
wire n_2356;
wire n_12363;
wire n_18201;
wire n_7553;
wire n_1772;
wire n_1119;
wire n_6824;
wire n_19625;
wire n_5788;
wire n_11788;
wire n_2739;
wire n_12544;
wire n_13036;
wire n_14146;
wire n_13199;
wire n_6903;
wire n_2864;
wire n_13009;
wire n_1180;
wire n_10908;
wire n_10339;
wire n_9908;
wire n_9486;
wire n_13002;
wire n_13868;
wire n_7903;
wire n_18596;
wire n_11877;
wire n_8864;
wire n_7384;
wire n_18674;
wire n_13285;
wire n_8610;
wire n_19075;
wire n_7894;
wire n_11750;
wire n_3532;
wire n_7055;
wire n_18722;
wire n_8520;
wire n_16458;
wire n_13374;
wire n_12055;
wire n_381;
wire n_7639;
wire n_16520;
wire n_4327;
wire n_3765;
wire n_4125;
wire n_12811;
wire n_12186;
wire n_13032;
wire n_3067;
wire n_2155;
wire n_11001;
wire n_9512;
wire n_14199;
wire n_17858;
wire n_13684;
wire n_2364;
wire n_9170;
wire n_15108;
wire n_9616;
wire n_3803;
wire n_2085;
wire n_917;
wire n_16898;
wire n_3639;
wire n_9073;
wire n_12897;
wire n_5192;
wire n_18325;
wire n_12272;
wire n_9302;
wire n_19068;
wire n_13948;
wire n_11798;
wire n_9062;
wire n_3413;
wire n_9171;
wire n_3412;
wire n_8279;
wire n_12191;
wire n_17432;
wire n_9580;
wire n_8019;
wire n_13963;
wire n_17707;
wire n_4575;
wire n_699;
wire n_4320;
wire n_18842;
wire n_7832;
wire n_9540;
wire n_17242;
wire n_11137;
wire n_451;
wire n_8390;
wire n_8898;
wire n_14316;
wire n_5231;
wire n_2190;
wire n_8613;
wire n_3438;
wire n_18300;
wire n_8464;
wire n_15701;
wire n_6423;
wire n_1441;
wire n_15612;
wire n_3373;
wire n_18804;
wire n_7441;
wire n_513;
wire n_12112;
wire n_13060;
wire n_16187;
wire n_9449;
wire n_14817;
wire n_9050;
wire n_433;
wire n_6121;
wire n_5726;
wire n_14087;
wire n_2792;
wire n_15980;
wire n_3798;
wire n_788;
wire n_329;
wire n_14438;
wire n_2674;
wire n_4641;
wire n_16253;
wire n_7133;
wire n_12202;
wire n_13836;
wire n_1866;
wire n_8661;
wire n_2130;
wire n_7424;
wire n_3714;
wire n_16671;
wire n_12870;
wire n_11156;
wire n_10611;
wire n_10715;
wire n_12333;
wire n_8609;
wire n_17666;
wire n_17219;
wire n_13576;
wire n_7626;
wire n_2714;
wire n_2245;
wire n_7310;
wire n_17451;
wire n_12119;
wire n_12618;
wire n_16093;
wire n_1265;
wire n_17266;
wire n_15129;
wire n_17146;
wire n_16209;
wire n_14306;
wire n_8873;
wire n_11891;
wire n_16276;
wire n_199;
wire n_18427;
wire n_12401;
wire n_13055;
wire n_7323;
wire n_7301;
wire n_3715;
wire n_18600;
wire n_612;
wire n_17633;
wire n_13829;
wire n_16533;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_14657;
wire n_3933;
wire n_17815;
wire n_7244;
wire n_10745;
wire n_2311;
wire n_1012;
wire n_3691;
wire n_7633;
wire n_18760;
wire n_13937;
wire n_4146;
wire n_5711;
wire n_9437;
wire n_18724;
wire n_8640;
wire n_14359;
wire n_4855;
wire n_6186;
wire n_16933;
wire n_6803;
wire n_8437;
wire n_8427;
wire n_1188;
wire n_10605;
wire n_14013;
wire n_14419;
wire n_9933;
wire n_11449;
wire n_2916;
wire n_15251;
wire n_9892;
wire n_18976;
wire n_16727;
wire n_9462;
wire n_5972;
wire n_19447;
wire n_15854;
wire n_3145;
wire n_19438;
wire n_5444;
wire n_12501;
wire n_961;
wire n_4356;
wire n_17518;
wire n_8843;
wire n_9891;
wire n_15810;
wire n_2377;
wire n_701;
wire n_10643;
wire n_16974;
wire n_3719;
wire n_4361;
wire n_10872;
wire n_13987;
wire n_15626;
wire n_1630;
wire n_4136;
wire n_13416;
wire n_12798;
wire n_14885;
wire n_2619;
wire n_5329;
wire n_9925;
wire n_16066;
wire n_9757;
wire n_10008;
wire n_13726;
wire n_507;
wire n_14412;
wire n_17587;
wire n_2271;
wire n_12243;
wire n_8562;
wire n_12614;
wire n_11378;
wire n_2606;
wire n_14631;
wire n_5728;
wire n_10032;
wire n_462;
wire n_304;
wire n_13425;
wire n_9806;
wire n_17105;
wire n_17233;
wire n_7021;
wire n_13591;
wire n_18296;
wire n_11713;
wire n_16972;
wire n_15586;
wire n_6355;
wire n_2954;
wire n_17821;
wire n_12931;
wire n_15525;
wire n_7215;
wire n_17790;
wire n_2493;
wire n_4802;
wire n_17566;
wire n_2705;
wire n_5523;
wire n_14332;
wire n_18379;
wire n_3405;
wire n_8016;
wire n_5423;
wire n_10645;
wire n_11096;
wire n_10604;
wire n_5074;
wire n_17398;
wire n_4044;
wire n_6564;
wire n_11161;
wire n_8709;
wire n_2631;
wire n_12491;
wire n_11216;
wire n_14368;
wire n_1293;
wire n_18390;
wire n_4701;
wire n_10966;
wire n_794;
wire n_727;
wire n_19310;
wire n_3385;
wire n_19650;
wire n_4851;
wire n_6442;
wire n_18359;
wire n_3293;
wire n_5204;
wire n_7925;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_15126;
wire n_4991;
wire n_19289;
wire n_5422;
wire n_6871;
wire n_16846;
wire n_9389;
wire n_1913;
wire n_12074;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5292;
wire n_12745;
wire n_9752;
wire n_14473;
wire n_12887;
wire n_18997;
wire n_10341;
wire n_19521;
wire n_4011;
wire n_15816;
wire n_18314;
wire n_7138;
wire n_17341;
wire n_4753;
wire n_8712;
wire n_631;
wire n_2262;
wire n_3611;
wire n_19254;
wire n_5059;
wire n_8837;
wire n_843;
wire n_17652;
wire n_2604;
wire n_14641;
wire n_16506;
wire n_17543;
wire n_15433;
wire n_15953;
wire n_5219;
wire n_9721;
wire n_11344;
wire n_3537;
wire n_12658;
wire n_1022;
wire n_9197;
wire n_19167;
wire n_1474;
wire n_14740;
wire n_9210;
wire n_6893;
wire n_5686;
wire n_8905;
wire n_13008;
wire n_18832;
wire n_18691;
wire n_7807;
wire n_18126;
wire n_14198;
wire n_14846;
wire n_3654;
wire n_1849;
wire n_9917;
wire n_12056;
wire n_14539;
wire n_8106;
wire n_4264;
wire n_12238;
wire n_5937;
wire n_19226;
wire n_12976;
wire n_14420;
wire n_18562;
wire n_6040;
wire n_11888;
wire n_13243;
wire n_14314;
wire n_16642;
wire n_14227;
wire n_10309;
wire n_11099;
wire n_5465;
wire n_8974;
wire n_4339;
wire n_14164;
wire n_3324;
wire n_10050;
wire n_9871;
wire n_19652;
wire n_1195;
wire n_10306;
wire n_7606;
wire n_1811;
wire n_7193;
wire n_3987;
wire n_1519;
wire n_18180;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_5721;
wire n_1048;
wire n_18142;
wire n_13632;
wire n_13020;
wire n_6012;
wire n_13148;
wire n_1418;
wire n_10429;
wire n_292;
wire n_11470;
wire n_3072;
wire n_13871;
wire n_4874;
wire n_4401;
wire n_889;
wire n_9903;
wire n_17208;
wire n_11102;
wire n_1110;
wire n_9228;
wire n_11539;
wire n_7710;
wire n_17792;
wire n_16166;
wire n_11899;
wire n_7892;
wire n_13168;
wire n_9522;
wire n_15617;
wire n_15463;
wire n_4658;
wire n_11076;
wire n_14339;
wire n_505;
wire n_1787;
wire n_16005;
wire n_6769;
wire n_9148;
wire n_11054;
wire n_2776;
wire n_10754;
wire n_5742;
wire n_3909;
wire n_9275;
wire n_10223;
wire n_1220;
wire n_8896;
wire n_7206;
wire n_5539;
wire n_6895;
wire n_13598;
wire n_2488;
wire n_17979;
wire n_10228;
wire n_1252;
wire n_511;
wire n_8758;
wire n_6026;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_17953;
wire n_13966;
wire n_12530;
wire n_1597;
wire n_9463;
wire n_4839;
wire n_2596;
wire n_1153;
wire n_13077;
wire n_16309;
wire n_10425;
wire n_8069;
wire n_6481;
wire n_19144;
wire n_4006;
wire n_15201;
wire n_9997;
wire n_6384;
wire n_13828;
wire n_7541;
wire n_6906;
wire n_14562;
wire n_9844;
wire n_12826;
wire n_8318;
wire n_10366;
wire n_15015;
wire n_19122;
wire n_7334;
wire n_5807;
wire n_16376;
wire n_2227;
wire n_5216;
wire n_14991;
wire n_10225;
wire n_4869;
wire n_6257;
wire n_4386;
wire n_8383;
wire n_12621;
wire n_4955;
wire n_11290;
wire n_17080;
wire n_12518;
wire n_19033;
wire n_3234;
wire n_14047;
wire n_9052;
wire n_856;
wire n_17447;
wire n_2830;
wire n_17678;
wire n_6587;
wire n_7781;
wire n_7360;
wire n_14568;
wire n_2181;
wire n_11702;
wire n_19395;
wire n_16970;
wire n_11372;
wire n_2826;
wire n_10817;
wire n_15324;
wire n_326;
wire n_8355;
wire n_19501;
wire n_17098;
wire n_12741;
wire n_18041;
wire n_7101;
wire n_1635;
wire n_7530;
wire n_15006;
wire n_15619;
wire n_18911;
wire n_9860;
wire n_12510;
wire n_11756;
wire n_2851;
wire n_8369;
wire n_9022;
wire n_160;
wire n_9103;
wire n_17142;
wire n_8831;
wire n_1508;
wire n_5608;
wire n_2240;
wire n_392;
wire n_12233;
wire n_8853;
wire n_4582;
wire n_6252;
wire n_18403;
wire n_6211;
wire n_15716;
wire n_5844;
wire n_17499;
wire n_1549;
wire n_17898;
wire n_17172;
wire n_8081;
wire n_16608;
wire n_17310;
wire n_13442;
wire n_1916;
wire n_14444;
wire n_18531;
wire n_10484;
wire n_11744;
wire n_17247;
wire n_10288;
wire n_18838;
wire n_10388;
wire n_6189;
wire n_15299;
wire n_4016;
wire n_11072;
wire n_621;
wire n_750;
wire n_2823;
wire n_5597;
wire n_13944;
wire n_9492;
wire n_6413;
wire n_7419;
wire n_6506;
wire n_18476;
wire n_1997;
wire n_710;
wire n_1818;
wire n_17086;
wire n_9727;
wire n_6935;
wire n_13019;
wire n_12703;
wire n_13079;
wire n_4397;
wire n_18343;
wire n_5050;
wire n_746;
wire n_3416;
wire n_3498;
wire n_15369;
wire n_15134;
wire n_16110;
wire n_2957;
wire n_1740;
wire n_19420;
wire n_9375;
wire n_17715;
wire n_5980;
wire n_8770;
wire n_3672;
wire n_15453;
wire n_5318;
wire n_6105;
wire n_6022;
wire n_10964;
wire n_3382;
wire n_12493;
wire n_13135;
wire n_8075;
wire n_5053;
wire n_7841;
wire n_9458;
wire n_8466;
wire n_6527;
wire n_15275;
wire n_19092;
wire n_8094;
wire n_4824;
wire n_2037;
wire n_4567;
wire n_6430;
wire n_782;
wire n_18268;
wire n_809;
wire n_10987;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_1797;
wire n_4595;
wire n_402;
wire n_1870;
wire n_11965;
wire n_4904;
wire n_1152;
wire n_14696;
wire n_5988;
wire n_5585;
wire n_15093;
wire n_12324;
wire n_711;
wire n_3105;
wire n_14006;
wire n_6666;
wire n_3692;
wire n_8321;
wire n_19116;
wire n_9954;
wire n_8735;
wire n_1695;
wire n_11722;
wire n_2272;
wire n_2760;
wire n_972;
wire n_12310;
wire n_5348;
wire n_6594;
wire n_624;
wire n_19471;
wire n_7095;
wire n_3045;
wire n_16672;
wire n_11701;
wire n_885;
wire n_3666;
wire n_4916;
wire n_18010;
wire n_13917;
wire n_7184;
wire n_9617;
wire n_13546;
wire n_14595;
wire n_17001;
wire n_7908;
wire n_7974;
wire n_7551;
wire n_11980;
wire n_11255;
wire n_13592;
wire n_3858;
wire n_17224;
wire n_11720;
wire n_3502;
wire n_5461;
wire n_13874;
wire n_6482;
wire n_5147;
wire n_15506;
wire n_1355;
wire n_9810;
wire n_14469;
wire n_16201;
wire n_2562;
wire n_17690;
wire n_1522;
wire n_5755;
wire n_8043;
wire n_16377;
wire n_14492;
wire n_1548;
wire n_1155;
wire n_14134;
wire n_4944;
wire n_11990;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_15457;
wire n_14345;
wire n_16847;
wire n_6841;
wire n_10153;
wire n_17622;
wire n_17952;
wire n_5054;
wire n_2962;
wire n_8171;
wire n_9006;
wire n_19641;
wire n_6774;
wire n_16964;
wire n_8600;
wire n_1925;
wire n_4407;
wire n_14816;
wire n_8710;
wire n_12806;
wire n_4045;
wire n_14302;
wire n_8549;
wire n_10172;
wire n_8054;
wire n_13904;
wire n_16614;
wire n_3258;
wire n_18694;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_17045;
wire n_15784;
wire n_18613;
wire n_3149;
wire n_11969;
wire n_7914;
wire n_16388;
wire n_3365;
wire n_6521;
wire n_3379;
wire n_8857;
wire n_14243;
wire n_9040;
wire n_6162;
wire n_8010;
wire n_3939;
wire n_6432;
wire n_1375;
wire n_3972;
wire n_1650;
wire n_13574;
wire n_12762;
wire n_16740;
wire n_9830;
wire n_18870;
wire n_10761;
wire n_2761;
wire n_3776;
wire n_18781;
wire n_11579;
wire n_1019;
wire n_15303;
wire n_8291;
wire n_18017;
wire n_4170;
wire n_11535;
wire n_2845;
wire n_18400;
wire n_5173;
wire n_12975;
wire n_16291;
wire n_13850;
wire n_6740;
wire n_1113;
wire n_11510;
wire n_6315;
wire n_17866;
wire n_12736;
wire n_5283;
wire n_9111;
wire n_7156;
wire n_9163;
wire n_15461;
wire n_6910;
wire n_6262;
wire n_14800;
wire n_2827;
wire n_7703;
wire n_6319;
wire n_17352;
wire n_14888;
wire n_12350;
wire n_12542;
wire n_13860;
wire n_1879;
wire n_6536;
wire n_256;
wire n_6175;
wire n_7040;
wire n_8280;
wire n_12390;
wire n_367;
wire n_18898;
wire n_2569;
wire n_10235;
wire n_6978;
wire n_5351;
wire n_12805;
wire n_6093;
wire n_11649;
wire n_16306;
wire n_703;
wire n_18485;
wire n_9190;
wire n_6947;
wire n_14918;
wire n_5293;
wire n_8203;
wire n_6099;
wire n_1324;
wire n_1435;
wire n_3920;
wire n_4892;
wire n_6140;
wire n_15489;
wire n_12914;
wire n_17721;
wire n_17159;
wire n_9506;
wire n_18440;
wire n_6415;
wire n_4439;
wire n_18883;
wire n_16542;
wire n_15158;
wire n_10828;
wire n_18866;
wire n_12300;
wire n_15389;
wire n_7549;
wire n_17308;
wire n_17425;
wire n_11281;
wire n_13056;
wire n_16019;
wire n_17732;
wire n_12337;
wire n_18520;
wire n_13466;
wire n_15082;
wire n_8871;
wire n_11114;
wire n_19442;
wire n_8418;
wire n_7740;
wire n_3679;
wire n_5891;
wire n_13050;
wire n_10860;
wire n_18259;
wire n_17517;
wire n_4930;
wire n_16208;
wire n_19327;
wire n_15209;
wire n_12273;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_12712;
wire n_360;
wire n_2149;
wire n_15078;
wire n_4557;
wire n_13012;
wire n_895;
wire n_8924;
wire n_12752;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_15511;
wire n_4593;
wire n_4465;
wire n_3622;
wire n_19600;
wire n_18204;
wire n_4495;
wire n_14278;
wire n_5117;
wire n_12777;
wire n_14706;
wire n_8214;
wire n_5990;
wire n_7043;
wire n_11462;
wire n_11732;
wire n_5024;
wire n_4559;
wire n_18137;
wire n_12819;
wire n_10214;
wire n_8241;
wire n_838;
wire n_3336;
wire n_8442;
wire n_2952;
wire n_9572;
wire n_15282;
wire n_9229;
wire n_19505;
wire n_16812;
wire n_16038;
wire n_12237;
wire n_18350;
wire n_6134;
wire n_1656;
wire n_5803;
wire n_2112;
wire n_13372;
wire n_2430;
wire n_653;
wire n_11375;
wire n_11267;
wire n_9602;
wire n_9311;
wire n_4335;
wire n_19482;
wire n_2034;
wire n_576;
wire n_6593;
wire n_8630;
wire n_2683;
wire n_19432;
wire n_9884;
wire n_9876;
wire n_9260;
wire n_14534;
wire n_13630;
wire n_16535;
wire n_13700;
wire n_10406;
wire n_3204;
wire n_17859;
wire n_6746;
wire n_11985;
wire n_8447;
wire n_6443;
wire n_14290;
wire n_7980;
wire n_348;
wire n_8828;
wire n_18631;
wire n_17687;
wire n_390;
wire n_1148;
wire n_6749;
wire n_10965;
wire n_10798;
wire n_19657;
wire n_7732;
wire n_13325;
wire n_15135;
wire n_14850;
wire n_16196;
wire n_11911;
wire n_4265;
wire n_11442;
wire n_2950;
wire n_5634;
wire n_719;
wire n_18862;
wire n_14064;
wire n_14524;
wire n_1090;
wire n_8859;
wire n_16883;
wire n_11388;
wire n_11651;
wire n_1362;
wire n_17946;
wire n_10154;
wire n_18663;
wire n_7922;
wire n_17469;
wire n_15826;
wire n_5580;
wire n_1450;
wire n_19101;
wire n_10033;
wire n_1789;
wire n_17877;
wire n_8311;
wire n_12253;
wire n_15005;
wire n_11147;
wire n_12928;
wire n_9877;
wire n_8764;
wire n_19361;
wire n_16167;
wire n_2161;
wire n_19452;
wire n_12990;
wire n_14246;
wire n_5764;
wire n_6920;
wire n_11817;
wire n_8729;
wire n_10359;
wire n_3344;
wire n_2334;
wire n_14957;
wire n_5133;
wire n_1763;
wire n_6907;
wire n_13447;
wire n_7144;
wire n_16579;
wire n_11479;
wire n_11737;
wire n_8048;
wire n_635;
wire n_12028;
wire n_3786;
wire n_7072;
wire n_13095;
wire n_4254;
wire n_8253;
wire n_4303;
wire n_18592;
wire n_15032;
wire n_1158;
wire n_11600;
wire n_2248;
wire n_16607;
wire n_15085;
wire n_16390;
wire n_10722;
wire n_8088;
wire n_17855;
wire n_10666;
wire n_3147;
wire n_15440;
wire n_753;
wire n_3925;
wire n_3180;
wire n_8516;
wire n_8302;
wire n_17717;
wire n_15610;
wire n_359;
wire n_15329;
wire n_8167;
wire n_7859;
wire n_14315;
wire n_7872;
wire n_1479;
wire n_4768;
wire n_13858;
wire n_17913;
wire n_3717;
wire n_7480;
wire n_5410;
wire n_571;
wire n_2215;
wire n_16255;
wire n_8944;
wire n_1884;
wire n_10023;
wire n_10999;
wire n_665;
wire n_5156;
wire n_18716;
wire n_10410;
wire n_4447;
wire n_3445;
wire n_373;
wire n_16983;
wire n_8975;
wire n_1833;
wire n_17009;
wire n_11305;
wire n_17668;
wire n_9101;
wire n_15631;
wire n_14755;
wire n_8825;
wire n_12969;
wire n_1856;
wire n_12260;
wire n_12016;
wire n_8266;
wire n_5691;
wire n_8981;
wire n_4957;
wire n_17082;
wire n_165;
wire n_8771;
wire n_15750;
wire n_4039;
wire n_457;
wire n_3800;
wire n_4566;
wire n_12939;
wire n_15038;
wire n_17925;
wire n_10404;
wire n_8138;
wire n_6638;
wire n_12779;
wire n_17505;
wire n_17199;
wire n_2930;
wire n_15531;
wire n_13547;
wire n_12816;
wire n_9211;
wire n_8124;
wire n_7366;
wire n_9395;
wire n_5269;
wire n_17348;
wire n_1538;
wire n_8147;
wire n_5468;
wire n_4730;
wire n_8127;
wire n_9402;
wire n_14014;
wire n_10700;
wire n_17743;
wire n_10968;
wire n_3579;
wire n_14247;
wire n_3335;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_700;
wire n_3178;
wire n_16155;
wire n_15418;
wire n_5256;
wire n_11970;
wire n_7918;
wire n_4168;
wire n_6651;
wire n_12308;
wire n_1923;
wire n_10783;
wire n_12163;
wire n_3952;
wire n_11523;
wire n_12944;
wire n_3911;
wire n_7472;
wire n_9737;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_14709;
wire n_10812;
wire n_12297;
wire n_13848;
wire n_6366;
wire n_2997;
wire n_10001;
wire n_13280;
wire n_12145;
wire n_11088;
wire n_5939;
wire n_5509;
wire n_8160;
wire n_3619;
wire n_11405;
wire n_19274;
wire n_1786;
wire n_13103;
wire n_18385;
wire n_15630;
wire n_4198;
wire n_1371;
wire n_10977;
wire n_2886;
wire n_11299;
wire n_10615;
wire n_1803;
wire n_11542;
wire n_4065;
wire n_229;
wire n_7647;
wire n_12426;
wire n_16222;
wire n_15068;
wire n_15442;
wire n_9054;
wire n_2470;
wire n_4446;
wire n_10532;
wire n_17776;
wire n_4417;
wire n_13995;
wire n_13073;
wire n_6728;
wire n_2286;
wire n_4743;
wire n_16029;
wire n_2018;
wire n_1903;
wire n_13556;
wire n_13367;
wire n_10771;
wire n_11441;
wire n_14203;
wire n_17269;
wire n_693;
wire n_1056;
wire n_12844;
wire n_5851;
wire n_7073;
wire n_9755;
wire n_5110;
wire n_10104;
wire n_772;
wire n_2806;
wire n_9117;
wire n_19426;
wire n_3028;
wire n_9381;
wire n_3076;
wire n_12049;
wire n_14498;
wire n_886;
wire n_343;
wire n_3624;
wire n_1820;
wire n_6549;
wire n_539;
wire n_6096;
wire n_7853;
wire n_12526;
wire n_2836;
wire n_8890;
wire n_16575;
wire n_7721;
wire n_7192;
wire n_19602;
wire n_11206;
wire n_11593;
wire n_15807;
wire n_3906;
wire n_11786;
wire n_12737;
wire n_4954;
wire n_17258;
wire n_15113;
wire n_9273;
wire n_2612;
wire n_8970;
wire n_16910;
wire n_2591;
wire n_1815;
wire n_10640;
wire n_2593;
wire n_10729;
wire n_14656;
wire n_16052;
wire n_14745;
wire n_19243;
wire n_4605;
wire n_7635;
wire n_11268;
wire n_17121;
wire n_14760;
wire n_3943;
wire n_11501;
wire n_7227;
wire n_13390;
wire n_8030;
wire n_6052;
wire n_13264;
wire n_8687;
wire n_5374;
wire n_12010;
wire n_1843;
wire n_9738;
wire n_12026;
wire n_4227;
wire n_521;
wire n_17481;
wire n_8633;
wire n_17645;
wire n_7689;
wire n_6511;
wire n_18470;
wire n_1309;
wire n_916;
wire n_4415;
wire n_7099;
wire n_1970;
wire n_14676;
wire n_6358;
wire n_2059;
wire n_2669;
wire n_18880;
wire n_11313;
wire n_10438;
wire n_6986;
wire n_8801;
wire n_3912;
wire n_3118;
wire n_1907;
wire n_2529;
wire n_16438;
wire n_860;
wire n_8219;
wire n_15373;
wire n_18580;
wire n_1302;
wire n_10575;
wire n_11028;
wire n_12171;
wire n_14193;
wire n_12935;
wire n_14906;
wire n_7827;
wire n_15211;
wire n_10760;
wire n_4792;
wire n_15334;
wire n_7731;
wire n_11527;
wire n_18404;
wire n_3514;
wire n_16486;
wire n_9535;
wire n_2654;
wire n_5302;
wire n_966;
wire n_12490;
wire n_3357;
wire n_692;
wire n_5781;
wire n_3895;
wire n_8486;
wire n_12829;
wire n_4118;
wire n_2176;
wire n_2459;
wire n_18662;
wire n_1111;
wire n_1251;
wire n_11610;
wire n_12739;
wire n_7132;
wire n_2711;
wire n_17021;
wire n_17710;
wire n_6663;
wire n_12609;
wire n_4441;
wire n_18248;
wire n_8155;
wire n_11360;
wire n_11868;
wire n_1664;
wire n_3022;
wire n_8098;
wire n_9191;
wire n_17791;
wire n_5654;
wire n_2345;
wire n_18202;
wire n_6376;
wire n_18141;
wire n_5113;
wire n_12888;
wire n_5479;
wire n_19407;
wire n_8485;
wire n_14852;
wire n_7001;
wire n_13070;
wire n_4822;
wire n_9650;
wire n_850;
wire n_5692;
wire n_8473;
wire n_13640;
wire n_14147;
wire n_14491;
wire n_15011;
wire n_17607;
wire n_3768;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_9664;
wire n_3785;
wire n_14928;
wire n_2602;
wire n_2980;
wire n_13778;
wire n_696;
wire n_9931;
wire n_16419;
wire n_16470;
wire n_1082;
wire n_1317;
wire n_16956;
wire n_3227;
wire n_4055;
wire n_14634;
wire n_2178;
wire n_10753;
wire n_13174;
wire n_7108;
wire n_14455;
wire n_1796;
wire n_17164;
wire n_11879;
wire n_2082;
wire n_7876;
wire n_17175;
wire n_9656;
wire n_3707;
wire n_8148;
wire n_8150;
wire n_3578;
wire n_909;
wire n_12596;
wire n_15398;
wire n_15593;
wire n_18175;
wire n_4925;
wire n_16424;
wire n_5415;
wire n_13945;
wire n_8986;
wire n_19367;
wire n_12697;
wire n_7260;
wire n_6409;
wire n_11939;
wire n_1634;
wire n_3252;
wire n_627;
wire n_14347;
wire n_7552;
wire n_19052;
wire n_17969;
wire n_12166;
wire n_2133;
wire n_1712;
wire n_1523;
wire n_10646;
wire n_15725;
wire n_1627;
wire n_11704;
wire n_17506;
wire n_18050;
wire n_8763;
wire n_5208;
wire n_8679;
wire n_7239;
wire n_15582;
wire n_16415;
wire n_9848;
wire n_14447;
wire n_11962;
wire n_5690;
wire n_9227;
wire n_7050;
wire n_17137;
wire n_2573;
wire n_2646;
wire n_6623;
wire n_13951;
wire n_13968;
wire n_10378;
wire n_16924;
wire n_1364;
wire n_13316;
wire n_10313;
wire n_13689;
wire n_8139;
wire n_17268;
wire n_18000;
wire n_19384;
wire n_3037;
wire n_19288;
wire n_3729;
wire n_19431;
wire n_10773;
wire n_18210;
wire n_2537;
wire n_8830;
wire n_4483;
wire n_5347;
wire n_14836;
wire n_12867;
wire n_4988;
wire n_15960;
wire n_15343;
wire n_7568;
wire n_6354;
wire n_6344;
wire n_12123;
wire n_9772;
wire n_18885;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_15370;
wire n_7949;
wire n_7724;
wire n_18001;
wire n_4284;
wire n_6305;
wire n_1947;
wire n_12547;
wire n_16148;
wire n_15577;
wire n_3426;
wire n_16550;
wire n_4971;
wire n_19066;
wire n_5857;
wire n_8646;
wire n_13415;
wire n_10259;
wire n_7107;
wire n_17111;
wire n_6457;
wire n_8597;
wire n_17951;
wire n_17379;
wire n_987;
wire n_7123;
wire n_5499;
wire n_720;
wire n_8117;
wire n_15169;
wire n_1707;
wire n_10213;
wire n_13888;
wire n_16592;
wire n_8208;
wire n_797;
wire n_2933;
wire n_19373;
wire n_1878;
wire n_8536;
wire n_17252;
wire n_9435;
wire n_7229;
wire n_8350;
wire n_16475;
wire n_5190;
wire n_13892;
wire n_16361;
wire n_14559;
wire n_16831;
wire n_4097;
wire n_1666;
wire n_5392;
wire n_17110;
wire n_14052;
wire n_14311;
wire n_13765;
wire n_10332;
wire n_7709;
wire n_15290;
wire n_11874;
wire n_13926;
wire n_10171;
wire n_15184;
wire n_1228;
wire n_5455;
wire n_18131;
wire n_5442;
wire n_6386;
wire n_12803;
wire n_5948;
wire n_19518;
wire n_5511;
wire n_2898;
wire n_6208;
wire n_6739;
wire n_15779;
wire n_8202;
wire n_15366;
wire n_3200;
wire n_12734;
wire n_3167;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_10269;
wire n_19504;
wire n_12262;
wire n_14910;
wire n_14385;
wire n_14499;
wire n_8738;
wire n_9126;
wire n_15368;
wire n_19077;
wire n_11376;
wire n_9438;
wire n_18433;
wire n_7808;
wire n_6544;
wire n_9122;
wire n_14731;
wire n_683;
wire n_5140;
wire n_4992;
wire n_5197;
wire n_16337;
wire n_17691;
wire n_8721;
wire n_12820;
wire n_9912;
wire n_6356;
wire n_13558;
wire n_3577;
wire n_2432;
wire n_10148;
wire n_19491;
wire n_1363;
wire n_3641;
wire n_2218;
wire n_16890;
wire n_13890;
wire n_5481;
wire n_9264;
wire n_14483;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_5184;
wire n_5794;
wire n_15179;
wire n_7638;
wire n_15724;
wire n_19303;
wire n_4053;
wire n_10234;
wire n_8836;
wire n_7019;
wire n_11325;
wire n_14838;
wire n_15207;
wire n_13521;
wire n_4167;
wire n_14926;
wire n_10731;
wire n_9878;
wire n_14591;
wire n_14363;
wire n_14576;
wire n_4431;
wire n_17797;
wire n_1125;
wire n_11498;
wire n_10513;
wire n_441;
wire n_7296;
wire n_4299;
wire n_7575;
wire n_3571;
wire n_7083;
wire n_1775;
wire n_7720;
wire n_11643;
wire n_1093;
wire n_6268;
wire n_5827;
wire n_5199;
wire n_6456;
wire n_11103;
wire n_16823;
wire n_16966;
wire n_14088;
wire n_5313;
wire n_17926;
wire n_13817;
wire n_3856;
wire n_9971;
wire n_19579;
wire n_3425;
wire n_10894;
wire n_14118;
wire n_18082;
wire n_9524;
wire n_6467;
wire n_9243;
wire n_9282;
wire n_1453;
wire n_6796;
wire n_18821;
wire n_12417;
wire n_4830;
wire n_13225;
wire n_17006;
wire n_1224;
wire n_10208;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_10804;
wire n_6486;
wire n_3960;
wire n_17246;
wire n_17167;
wire n_18357;
wire n_8438;
wire n_13355;
wire n_18160;
wire n_4693;
wire n_18614;
wire n_10793;
wire n_2000;
wire n_14672;
wire n_4267;
wire n_15127;
wire n_6732;
wire n_2270;
wire n_12711;
wire n_12219;
wire n_906;
wire n_10440;
wire n_1733;
wire n_9695;
wire n_11306;
wire n_19169;
wire n_4609;
wire n_1687;
wire n_8757;
wire n_2328;
wire n_13035;
wire n_7020;
wire n_13021;
wire n_613;
wire n_12893;
wire n_8596;
wire n_3314;
wire n_3016;
wire n_11292;
wire n_554;
wire n_13502;
wire n_5223;
wire n_6298;
wire n_5474;
wire n_12289;
wire n_10813;
wire n_1889;
wire n_10757;
wire n_13046;
wire n_13935;
wire n_435;
wire n_16670;
wire n_762;
wire n_11431;
wire n_1778;
wire n_5287;
wire n_13646;
wire n_1079;
wire n_5083;
wire n_6007;
wire n_3338;
wire n_18186;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_8834;
wire n_3636;
wire n_2327;
wire n_16429;
wire n_15262;
wire n_10822;
wire n_18773;
wire n_7104;
wire n_7467;
wire n_14609;
wire n_2597;
wire n_9534;
wire n_3194;
wire n_13380;
wire n_5771;
wire n_17369;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_11836;
wire n_349;
wire n_6602;
wire n_10924;
wire n_17421;
wire n_11186;
wire n_9742;
wire n_6484;
wire n_19642;
wire n_3637;
wire n_12527;
wire n_4574;
wire n_1859;
wire n_9019;
wire n_13891;
wire n_1718;
wire n_8985;
wire n_7692;
wire n_19463;
wire n_12477;
wire n_4234;
wire n_14325;
wire n_15503;
wire n_10418;
wire n_1768;
wire n_19589;
wire n_3974;
wire n_10875;
wire n_1847;
wire n_3634;
wire n_11736;
wire n_7560;
wire n_16270;
wire n_14729;
wire n_11846;
wire n_1397;
wire n_12400;
wire n_901;
wire n_2755;
wire n_4660;
wire n_1623;
wire n_16861;
wire n_9145;
wire n_12092;
wire n_3112;
wire n_12295;
wire n_9754;
wire n_19549;
wire n_9315;
wire n_18483;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_6734;
wire n_7476;
wire n_5570;
wire n_18096;
wire n_785;
wire n_7392;
wire n_7495;
wire n_5435;
wire n_9765;
wire n_3213;
wire n_3820;
wire n_5200;
wire n_6941;
wire n_1168;
wire n_5115;
wire n_1943;
wire n_5566;
wire n_7829;
wire n_3249;
wire n_8680;
wire n_2722;
wire n_4152;
wire n_16522;
wire n_10394;
wire n_11391;
wire n_15462;
wire n_5244;
wire n_12714;
wire n_16779;
wire n_5889;
wire n_19024;
wire n_5391;
wire n_1938;
wire n_9763;
wire n_11070;
wire n_13337;
wire n_15112;
wire n_18146;
wire n_3394;
wire n_9162;
wire n_1715;
wire n_14849;
wire n_1443;
wire n_1272;
wire n_16661;
wire n_5849;
wire n_11648;
wire n_4554;
wire n_19044;
wire n_10322;
wire n_7135;
wire n_8555;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_15912;
wire n_16206;
wire n_8508;
wire n_19509;
wire n_18827;
wire n_16529;
wire n_1705;
wire n_3905;
wire n_8207;
wire n_11653;
wire n_4680;
wire n_3013;
wire n_11717;
wire n_15246;
wire n_14940;
wire n_6165;
wire n_19153;
wire n_17553;
wire n_15395;
wire n_12838;
wire n_2670;
wire n_18813;
wire n_13505;
wire n_5910;
wire n_12776;
wire n_1569;
wire n_7033;
wire n_13156;
wire n_15529;
wire n_10710;
wire n_5557;
wire n_411;
wire n_8850;
wire n_14647;
wire n_18384;
wire n_8002;
wire n_19610;
wire n_1795;
wire n_16722;
wire n_9090;
wire n_16412;
wire n_12008;
wire n_6119;
wire n_1545;
wire n_4145;
wire n_4821;
wire n_3121;
wire n_9261;
wire n_8301;
wire n_17453;
wire n_12223;
wire n_18706;
wire n_16758;
wire n_548;
wire n_10942;
wire n_11430;
wire n_13010;
wire n_19073;
wire n_345;
wire n_11239;
wire n_4943;
wire n_10953;
wire n_7842;
wire n_2629;
wire n_2172;
wire n_6202;
wire n_17831;
wire n_12898;
wire n_4682;
wire n_19523;
wire n_15540;
wire n_10343;
wire n_4942;
wire n_9258;
wire n_1086;
wire n_10286;
wire n_10371;
wire n_14990;
wire n_2561;
wire n_16691;
wire n_7236;
wire n_10257;
wire n_3305;
wire n_11219;
wire n_10047;
wire n_14541;
wire n_3267;
wire n_16186;
wire n_1914;
wire n_1318;
wire n_13766;
wire n_11226;
wire n_3005;
wire n_16989;
wire n_11413;
wire n_4840;
wire n_1029;
wire n_16617;
wire n_5320;
wire n_5353;
wire n_13710;
wire n_11232;
wire n_2417;
wire n_9105;
wire n_12080;
wire n_16261;
wire n_5093;
wire n_1556;
wire n_19512;
wire n_5979;
wire n_9668;
wire n_13335;
wire n_14022;
wire n_2083;
wire n_5517;
wire n_3207;
wire n_11276;
wire n_5605;
wire n_3401;
wire n_10744;
wire n_3242;
wire n_9870;
wire n_3613;
wire n_11334;
wire n_7678;
wire n_1045;
wire n_13075;
wire n_13736;
wire n_13129;
wire n_9178;
wire n_6063;
wire n_16118;
wire n_1325;
wire n_6504;
wire n_2923;
wire n_1727;
wire n_13586;
wire n_15813;
wire n_10597;
wire n_17382;
wire n_16281;
wire n_11827;
wire n_13049;
wire n_13961;
wire n_17413;
wire n_15745;
wire n_3814;
wire n_6003;
wire n_6684;
wire n_19084;
wire n_13063;
wire n_5451;
wire n_9323;
wire n_6961;
wire n_3543;
wire n_13252;
wire n_9922;
wire n_12024;
wire n_13084;
wire n_2903;
wire n_16622;
wire n_15374;
wire n_3808;
wire n_4365;
wire n_18123;
wire n_16440;
wire n_7929;
wire n_16821;
wire n_10572;
wire n_16431;
wire n_1007;
wire n_1929;
wire n_19272;
wire n_1592;
wire n_19455;
wire n_13985;
wire n_3758;
wire n_17594;
wire n_14124;
wire n_19119;
wire n_17658;
wire n_13552;
wire n_18086;
wire n_12681;
wire n_3343;
wire n_18419;
wire n_13022;
wire n_18583;
wire n_2752;
wire n_17047;
wire n_9513;
wire n_16447;
wire n_16124;
wire n_4885;
wire n_15446;
wire n_10555;
wire n_19179;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_13656;
wire n_18967;
wire n_3658;
wire n_6834;
wire n_6817;
wire n_6927;
wire n_5209;
wire n_16841;
wire n_15470;
wire n_6215;
wire n_4212;
wire n_5699;
wire n_181;
wire n_5765;
wire n_15754;
wire n_17375;
wire n_7862;
wire n_16708;
wire n_17439;
wire n_10630;
wire n_17955;
wire n_8808;
wire n_10061;
wire n_300;
wire n_15599;
wire n_11865;
wire n_13024;
wire n_10694;
wire n_11041;
wire n_14490;
wire n_9708;
wire n_5064;
wire n_15479;
wire n_7119;
wire n_8889;
wire n_601;
wire n_13986;
wire n_9790;
wire n_11973;
wire n_5759;
wire n_13329;
wire n_7874;
wire n_8490;
wire n_10329;
wire n_9979;
wire n_8767;
wire n_13946;
wire n_9505;
wire n_2566;
wire n_15028;
wire n_2702;
wire n_7102;
wire n_7420;
wire n_13618;
wire n_4568;
wire n_10662;
wire n_5559;
wire n_18653;
wire n_17534;
wire n_14993;
wire n_14327;
wire n_8624;
wire n_11022;
wire n_10247;
wire n_5377;
wire n_1016;
wire n_8796;
wire n_4106;
wire n_1501;
wire n_17829;
wire n_10733;
wire n_10472;
wire n_12597;
wire n_13744;
wire n_12834;
wire n_10066;
wire n_17239;
wire n_14335;
wire n_6419;
wire n_3553;
wire n_18989;
wire n_2275;
wire n_15087;
wire n_2568;
wire n_2022;
wire n_3494;
wire n_6244;
wire n_6900;
wire n_9337;
wire n_15219;
wire n_908;
wire n_9432;
wire n_17295;
wire n_19563;
wire n_7705;
wire n_2106;
wire n_5350;
wire n_5470;
wire n_7932;
wire n_18331;
wire n_7058;
wire n_15009;
wire n_8262;
wire n_5700;
wire n_7981;
wire n_9874;
wire n_12588;
wire n_17203;
wire n_15648;
wire n_17548;
wire n_5874;
wire n_9231;
wire n_3328;
wire n_18612;
wire n_7973;
wire n_6815;
wire n_15634;
wire n_9569;
wire n_14823;
wire n_14691;
wire n_2530;
wire n_16908;
wire n_16508;
wire n_9719;
wire n_8358;
wire n_9552;
wire n_13822;
wire n_14948;
wire n_6317;
wire n_475;
wire n_492;
wire n_4012;
wire n_10756;
wire n_3645;
wire n_17099;
wire n_14387;
wire n_16572;
wire n_11797;
wire n_18889;
wire n_18933;
wire n_14106;
wire n_18788;
wire n_13616;
wire n_18667;
wire n_7820;
wire n_8881;
wire n_7844;
wire n_14301;
wire n_15468;
wire n_9633;
wire n_3422;
wire n_4845;
wire n_3086;
wire n_2033;
wire n_13627;
wire n_878;
wire n_19040;
wire n_5120;
wire n_13112;
wire n_10042;
wire n_10478;
wire n_16581;
wire n_981;
wire n_18597;
wire n_13163;
wire n_3702;
wire n_8754;
wire n_9847;
wire n_16968;
wire n_2233;
wire n_18098;
wire n_10367;
wire n_3233;
wire n_10867;
wire n_3310;
wire n_4061;
wire n_7460;
wire n_9519;
wire n_14814;
wire n_6367;
wire n_13564;
wire n_12671;
wire n_8714;
wire n_13260;
wire n_17302;
wire n_10085;
wire n_1051;
wire n_8182;
wire n_16165;
wire n_14090;
wire n_6056;
wire n_7200;
wire n_3206;
wire n_2363;
wire n_553;
wire n_15424;
wire n_4903;
wire n_17301;
wire n_15554;
wire n_15836;
wire n_15966;
wire n_16009;
wire n_15309;
wire n_14463;
wire n_2540;
wire n_973;
wire n_5743;
wire n_13503;
wire n_11152;
wire n_16318;
wire n_14166;
wire n_4522;
wire n_10122;
wire n_679;
wire n_9327;
wire n_16175;
wire n_5368;
wire n_4263;
wire n_14271;
wire n_7059;
wire n_915;
wire n_14425;
wire n_5971;
wire n_6327;
wire n_11964;
wire n_3155;
wire n_7826;
wire n_19078;
wire n_5933;
wire n_7076;
wire n_4780;
wire n_11403;
wire n_2697;
wire n_6866;
wire n_17108;
wire n_2512;
wire n_9387;
wire n_3039;
wire n_14596;
wire n_6514;
wire n_9794;
wire n_1322;
wire n_16387;
wire n_11142;
wire n_1958;
wire n_17434;
wire n_1197;
wire n_17509;
wire n_4984;
wire n_3420;
wire n_10862;
wire n_4283;
wire n_8911;
wire n_900;
wire n_8248;
wire n_11476;
wire n_2659;
wire n_13633;
wire n_14538;
wire n_2116;
wire n_19534;
wire n_1013;
wire n_17999;
wire n_11367;
wire n_15478;
wire n_2183;
wire n_16797;
wire n_12676;
wire n_18755;
wire n_3392;
wire n_13913;
wire n_19166;
wire n_8733;
wire n_6050;
wire n_7976;
wire n_13080;
wire n_13403;
wire n_17444;
wire n_1581;
wire n_1357;
wire n_14952;
wire n_1853;
wire n_10386;
wire n_12128;
wire n_14060;
wire n_14018;
wire n_15959;
wire n_5563;
wire n_1348;
wire n_11026;
wire n_13309;
wire n_15292;
wire n_11467;
wire n_12672;
wire n_12063;
wire n_8330;
wire n_1009;
wire n_15560;
wire n_1160;
wire n_15065;
wire n_5717;
wire n_1247;
wire n_6017;
wire n_9696;
wire n_15771;
wire n_15508;
wire n_471;
wire n_17990;
wire n_14148;
wire n_5720;
wire n_4702;
wire n_4895;
wire n_12924;
wire n_16331;
wire n_12732;
wire n_17171;
wire n_12649;
wire n_5898;
wire n_17458;
wire n_6858;
wire n_9464;
wire n_9252;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_12843;
wire n_14279;
wire n_1140;
wire n_1670;
wire n_2344;
wire n_17856;
wire n_2365;
wire n_19573;
wire n_15687;
wire n_11248;
wire n_2447;
wire n_8540;
wire n_9915;
wire n_5940;
wire n_6089;
wire n_7588;
wire n_18480;
wire n_4969;
wire n_10017;
wire n_11141;
wire n_5105;
wire n_11093;
wire n_19556;
wire n_17716;
wire n_5263;
wire n_2510;
wire n_6713;
wire n_18750;
wire n_15968;
wire n_17893;
wire n_4602;
wire n_13181;
wire n_18303;
wire n_1163;
wire n_16487;
wire n_17592;
wire n_15047;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_7593;
wire n_17156;
wire n_17908;
wire n_14085;
wire n_8068;
wire n_19599;
wire n_2173;
wire n_7764;
wire n_19634;
wire n_10196;
wire n_493;
wire n_14573;
wire n_17433;
wire n_19453;
wire n_2108;
wire n_8693;
wire n_6454;
wire n_12625;
wire n_12177;
wire n_7307;
wire n_14512;
wire n_1280;
wire n_6918;
wire n_16214;
wire n_13761;
wire n_19576;
wire n_3296;
wire n_19065;
wire n_16219;
wire n_17017;
wire n_14456;
wire n_13364;
wire n_11494;
wire n_14743;
wire n_10218;
wire n_18492;
wire n_3792;
wire n_4791;
wire n_19127;
wire n_14859;
wire n_8062;
wire n_11832;
wire n_6375;
wire n_12974;
wire n_13078;
wire n_1956;
wire n_7047;
wire n_6632;
wire n_4549;
wire n_17241;
wire n_15795;
wire n_10542;
wire n_16814;
wire n_4349;
wire n_10681;
wire n_15162;
wire n_9732;
wire n_16494;
wire n_13370;
wire n_11894;
wire n_10222;
wire n_10524;
wire n_6705;
wire n_17988;
wire n_8629;
wire n_818;
wire n_9517;
wire n_15237;
wire n_15862;
wire n_6591;
wire n_2207;
wire n_13643;
wire n_9780;
wire n_3482;
wire n_2198;
wire n_13607;
wire n_6289;
wire n_3272;
wire n_8524;
wire n_19355;
wire n_18907;
wire n_4393;
wire n_14114;
wire n_1068;
wire n_932;
wire n_14904;
wire n_3317;
wire n_3978;
wire n_5560;
wire n_6512;
wire n_4074;
wire n_4918;
wire n_13820;
wire n_4013;
wire n_6703;
wire n_12122;
wire n_13428;
wire n_354;
wire n_17958;
wire n_2941;
wire n_547;
wire n_17194;
wire n_6086;
wire n_16668;
wire n_4147;
wire n_4477;
wire n_18139;
wire n_3168;
wire n_12184;
wire n_10210;
wire n_1793;
wire n_5611;
wire n_12571;
wire n_6219;
wire n_11853;
wire n_19626;
wire n_16770;
wire n_4742;
wire n_9609;
wire n_10029;
wire n_1703;
wire n_6761;
wire n_8972;
wire n_11725;
wire n_13635;
wire n_10801;
wire n_9206;
wire n_3384;
wire n_18488;
wire n_15698;
wire n_1950;
wire n_6811;
wire n_16865;
wire n_18642;
wire n_11622;
wire n_4838;
wire n_12336;
wire n_18345;
wire n_12543;
wire n_16129;
wire n_347;
wire n_9705;
wire n_16585;
wire n_17490;
wire n_2965;
wire n_9624;
wire n_3861;
wire n_1977;
wire n_10389;
wire n_3891;
wire n_15688;
wire n_1655;
wire n_13677;
wire n_1886;
wire n_14036;
wire n_13757;
wire n_12463;
wire n_10990;
wire n_11640;
wire n_12263;
wire n_8982;
wire n_17899;
wire n_13910;
wire n_4673;
wire n_7086;
wire n_3415;
wire n_2947;
wire n_9532;
wire n_18195;
wire n_6601;
wire n_16247;
wire n_13196;
wire n_17482;
wire n_5088;
wire n_19261;
wire n_8034;
wire n_484;
wire n_15824;
wire n_5856;
wire n_9836;
wire n_2497;
wire n_11525;
wire n_11999;
wire n_10837;
wire n_3545;
wire n_18921;
wire n_10554;
wire n_3993;
wire n_8994;
wire n_17827;
wire n_8413;
wire n_4685;
wire n_10149;
wire n_19473;
wire n_19393;
wire n_2663;
wire n_5825;
wire n_2938;
wire n_3780;
wire n_15791;
wire n_12190;
wire n_15484;
wire n_15152;
wire n_11847;
wire n_11976;
wire n_12511;
wire n_2750;
wire n_11167;
wire n_2775;
wire n_8765;
wire n_3477;
wire n_2349;
wire n_2684;
wire n_8213;
wire n_1495;
wire n_14472;
wire n_10534;
wire n_11049;
wire n_14974;
wire n_8451;
wire n_19410;
wire n_1128;
wire n_12743;
wire n_16523;
wire n_8731;
wire n_8385;
wire n_4999;
wire n_15587;
wire n_4922;
wire n_7370;
wire n_15322;
wire n_13539;
wire n_9350;
wire n_18324;
wire n_19383;
wire n_17917;
wire n_7026;
wire n_7053;
wire n_14618;
wire n_9226;
wire n_1765;
wire n_2707;
wire n_18810;
wire n_10608;
wire n_16355;
wire n_7173;
wire n_7042;
wire n_17314;
wire n_718;
wire n_17915;
wire n_5331;
wire n_19225;
wire n_19011;
wire n_16774;
wire n_16436;
wire n_2089;
wire n_10638;
wire n_17923;
wire n_9112;
wire n_18582;
wire n_18970;
wire n_4216;
wire n_19284;
wire n_5797;
wire n_9235;
wire n_16570;
wire n_19124;
wire n_4240;
wire n_3491;
wire n_13852;
wire n_9333;
wire n_704;
wire n_4162;
wire n_17813;
wire n_14089;
wire n_15758;
wire n_1999;
wire n_2731;
wire n_622;
wire n_147;
wire n_3353;
wire n_11804;
wire n_14234;
wire n_3018;
wire n_14125;
wire n_5800;
wire n_6562;
wire n_12809;
wire n_18770;
wire n_4785;
wire n_2002;
wire n_2138;
wire n_2414;
wire n_1771;
wire n_11052;
wire n_3148;
wire n_17350;
wire n_18598;
wire n_6671;
wire n_13470;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_19151;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_13068;
wire n_19158;
wire n_3775;
wire n_18795;
wire n_1176;
wire n_7792;
wire n_15985;
wire n_8161;
wire n_18798;
wire n_5763;
wire n_10014;
wire n_15723;
wire n_16840;
wire n_6029;
wire n_18698;
wire n_10677;
wire n_18269;
wire n_5751;
wire n_15852;
wire n_18857;
wire n_19216;
wire n_12321;
wire n_5924;
wire n_11247;
wire n_290;
wire n_18581;
wire n_8384;
wire n_6445;
wire n_18079;
wire n_13106;
wire n_14294;
wire n_17609;
wire n_6701;
wire n_14862;
wire n_7380;
wire n_8736;
wire n_11514;
wire n_4497;
wire n_1568;
wire n_12470;
wire n_12994;
wire n_18604;
wire n_10215;
wire n_18768;
wire n_14059;
wire n_4871;
wire n_10834;
wire n_17632;
wire n_17611;
wire n_1665;
wire n_19341;
wire n_154;
wire n_12064;
wire n_2127;
wire n_12696;
wire n_18024;
wire n_15735;
wire n_11133;
wire n_5449;
wire n_17143;
wire n_18341;
wire n_10871;
wire n_16405;
wire n_5926;
wire n_2354;
wire n_5398;
wire n_4573;
wire n_14624;
wire n_16600;
wire n_15036;
wire n_17695;
wire n_18193;
wire n_19489;
wire n_11571;
wire n_14120;
wire n_8844;
wire n_13147;
wire n_7641;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_14407;
wire n_14260;
wire n_16845;
wire n_18924;
wire n_17307;
wire n_7169;
wire n_10407;
wire n_19330;
wire n_14175;
wire n_11941;
wire n_4368;
wire n_15780;
wire n_18085;
wire n_1942;
wire n_3196;
wire n_15189;
wire n_8110;
wire n_5319;
wire n_9008;
wire n_12079;
wire n_15335;
wire n_399;
wire n_1440;
wire n_19147;
wire n_2063;
wire n_15227;
wire n_8805;
wire n_6014;
wire n_7209;
wire n_18908;
wire n_15026;
wire n_13895;
wire n_2475;
wire n_5181;
wire n_6979;
wire n_13222;
wire n_3144;
wire n_1268;
wire n_17284;
wire n_5583;
wire n_15987;
wire n_10462;
wire n_642;
wire n_3481;
wire n_11769;
wire n_8856;
wire n_19362;
wire n_303;
wire n_6142;
wire n_14901;
wire n_7769;
wire n_2374;
wire n_416;
wire n_17034;
wire n_10291;
wire n_4597;
wire n_18575;
wire n_18764;
wire n_3364;
wire n_17502;
wire n_14333;
wire n_8732;
wire n_7233;
wire n_13506;
wire n_7602;
wire n_9296;
wire n_18587;
wire n_7390;
wire n_10669;
wire n_19515;
wire n_8231;
wire n_13717;
wire n_5127;
wire n_2920;
wire n_7598;
wire n_12440;
wire n_19032;
wire n_8908;
wire n_1374;
wire n_2648;
wire n_16085;
wire n_1169;
wire n_6767;
wire n_12782;
wire n_3093;
wire n_10111;
wire n_19186;
wire n_19629;
wire n_15300;
wire n_6385;
wire n_11354;
wire n_17796;
wire n_7045;
wire n_3169;
wire n_8740;
wire n_11727;
wire n_6788;
wire n_12192;
wire n_2204;
wire n_177;
wire n_2087;
wire n_17342;
wire n_14465;
wire n_13412;
wire n_4422;
wire n_11749;
wire n_11300;
wire n_6143;
wire n_13457;
wire n_12551;
wire n_18066;
wire n_12497;
wire n_15043;
wire n_4632;
wire n_3084;
wire n_16602;
wire n_2343;
wire n_5967;
wire n_4963;
wire n_16864;
wire n_16761;
wire n_2942;
wire n_4966;
wire n_4714;
wire n_7679;
wire n_18133;
wire n_7936;
wire n_8966;
wire n_4847;
wire n_10287;
wire n_8538;
wire n_12101;
wire n_11145;
wire n_3586;
wire n_3653;
wire n_16684;
wire n_19594;
wire n_725;
wire n_10349;
wire n_4668;
wire n_5213;
wire n_16340;
wire n_7490;
wire n_7545;
wire n_1273;
wire n_7160;
wire n_9809;
wire n_10750;
wire n_617;
wire n_7295;
wire n_14338;
wire n_7348;
wire n_19071;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_17554;
wire n_16071;
wire n_3991;
wire n_15394;
wire n_3516;
wire n_16875;
wire n_15941;
wire n_610;
wire n_9558;
wire n_11594;
wire n_8715;
wire n_12474;
wire n_4036;
wire n_4759;
wire n_2153;
wire n_7162;
wire n_16655;
wire n_12346;
wire n_517;
wire n_18167;
wire n_4182;
wire n_667;
wire n_8371;
wire n_13916;
wire n_15195;
wire n_1279;
wire n_11458;
wire n_17056;
wire n_12244;
wire n_18753;
wire n_16188;
wire n_15644;
wire n_14255;
wire n_11670;
wire n_7681;
wire n_11504;
wire n_16850;
wire n_13981;
wire n_4637;
wire n_11516;
wire n_2412;
wire n_8392;
wire n_14659;
wire n_8095;
wire n_10830;
wire n_16868;
wire n_17644;
wire n_5118;
wire n_7503;
wire n_6854;
wire n_17254;
wire n_2757;
wire n_18733;
wire n_4977;
wire n_2716;
wire n_12953;
wire n_2452;
wire n_15224;
wire n_9215;
wire n_11406;
wire n_3043;
wire n_14963;
wire n_11047;
wire n_8050;
wire n_12817;
wire n_8399;
wire n_2543;
wire n_5090;
wire n_16916;
wire n_13866;
wire n_3177;
wire n_12435;
wire n_10946;
wire n_18106;
wire n_7065;
wire n_9216;
wire n_1262;
wire n_4835;
wire n_11961;
wire n_6122;
wire n_7911;
wire n_17486;
wire n_17504;
wire n_7330;
wire n_14605;
wire n_9202;
wire n_2373;
wire n_13543;
wire n_10351;
wire n_13772;
wire n_4734;
wire n_7493;
wire n_12940;
wire n_10460;
wire n_15487;
wire n_19221;
wire n_10334;
wire n_2244;
wire n_11614;
wire n_4290;
wire n_1684;
wire n_1352;
wire n_5407;
wire n_15242;
wire n_8422;
wire n_12224;
wire n_7088;
wire n_9394;
wire n_2704;
wire n_8878;
wire n_7440;
wire n_17681;
wire n_260;
wire n_17676;
wire n_14797;
wire n_9622;
wire n_14177;
wire n_14093;
wire n_3318;
wire n_14607;
wire n_10191;
wire n_4888;
wire n_17919;
wire n_776;
wire n_6000;
wire n_12679;
wire n_14921;
wire n_11168;
wire n_10911;
wire n_12756;
wire n_5004;
wire n_5294;
wire n_16097;
wire n_9845;
wire n_16147;
wire n_7374;
wire n_14389;
wire n_19514;
wire n_11937;
wire n_17277;
wire n_2229;
wire n_4527;
wire n_6046;
wire n_8251;
wire n_5323;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_14621;
wire n_3184;
wire n_18864;
wire n_3075;
wire n_17875;
wire n_11192;
wire n_4949;
wire n_6852;
wire n_8677;
wire n_9091;
wire n_17206;
wire n_13914;
wire n_14663;
wire n_16921;
wire n_17559;
wire n_2536;
wire n_9699;
wire n_13277;
wire n_12340;
wire n_18143;
wire n_16742;
wire n_18464;
wire n_13494;
wire n_5260;
wire n_9751;
wire n_5809;
wire n_10543;
wire n_7924;
wire n_17225;
wire n_560;
wire n_1321;
wire n_7659;
wire n_569;
wire n_3530;
wire n_16203;
wire n_8875;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_1235;
wire n_12662;
wire n_1292;
wire n_15697;
wire n_17879;
wire n_18140;
wire n_9293;
wire n_12503;
wire n_18510;
wire n_15202;
wire n_18218;
wire n_12871;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_18224;
wire n_16400;
wire n_2246;
wire n_4469;
wire n_431;
wire n_10809;
wire n_16934;
wire n_10899;
wire n_9639;
wire n_11898;
wire n_15250;
wire n_17193;
wire n_6711;
wire n_1941;
wire n_11997;
wire n_8946;
wire n_13090;
wire n_18984;
wire n_13541;
wire n_16958;
wire n_4924;
wire n_13908;
wire n_9646;
wire n_8017;
wire n_17396;
wire n_766;
wire n_1746;
wire n_7275;
wire n_8795;
wire n_7195;
wire n_11199;
wire n_17642;
wire n_11264;
wire n_2062;
wire n_4539;
wire n_7610;
wire n_6072;
wire n_12303;
wire n_9501;
wire n_11896;
wire n_16229;
wire n_10006;
wire n_11757;
wire n_2070;
wire n_18447;
wire n_12622;
wire n_6353;
wire n_4953;
wire n_12659;
wire n_2348;
wire n_6818;
wire n_391;
wire n_2066;
wire n_7539;
wire n_1476;
wire n_12629;
wire n_12868;
wire n_19263;
wire n_10275;
wire n_3458;
wire n_7775;
wire n_11392;
wire n_3190;
wire n_7930;
wire n_7661;
wire n_5383;
wire n_16498;
wire n_14165;
wire n_17309;
wire n_19413;
wire n_13787;
wire n_875;
wire n_1678;
wire n_13674;
wire n_18311;
wire n_13912;
wire n_10292;
wire n_7969;
wire n_6864;
wire n_14445;
wire n_11278;
wire n_3787;
wire n_7548;
wire n_16732;
wire n_4450;
wire n_6156;
wire n_12913;
wire n_7064;
wire n_19285;
wire n_16839;
wire n_16798;
wire n_12154;
wire n_8000;
wire n_14427;
wire n_5645;
wire n_3990;
wire n_18327;
wire n_6917;
wire n_6937;
wire n_1628;
wire n_9963;
wire n_988;
wire n_17211;
wire n_7324;
wire n_2507;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_17568;
wire n_1536;
wire n_6301;
wire n_18061;
wire n_16815;
wire n_18022;
wire n_1132;
wire n_15570;
wire n_15562;
wire n_17207;
wire n_1327;
wire n_19000;
wire n_7729;
wire n_246;
wire n_19622;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_16987;
wire n_18337;
wire n_2380;
wire n_6699;
wire n_12926;
wire n_14809;
wire n_4579;
wire n_14725;
wire n_16892;
wire n_4811;
wire n_6874;
wire n_6259;
wire n_9340;
wire n_16527;
wire n_17963;
wire n_6677;
wire n_12161;
wire n_3432;
wire n_11735;
wire n_4282;
wire n_1196;
wire n_8769;
wire n_6764;
wire n_10324;
wire n_11189;
wire n_8815;
wire n_12044;
wire n_748;
wire n_9303;
wire n_1785;
wire n_3057;
wire n_8261;
wire n_13104;
wire n_2287;
wire n_7139;
wire n_5727;
wire n_16819;
wire n_16612;
wire n_761;
wire n_5946;
wire n_3778;
wire n_9722;
wire n_12155;
wire n_15664;
wire n_4974;
wire n_12373;
wire n_5975;
wire n_19376;
wire n_14579;
wire n_17930;
wire n_4569;
wire n_8665;
wire n_15847;
wire n_5097;
wire n_7751;
wire n_2234;
wire n_18763;
wire n_14718;
wire n_4384;
wire n_19253;
wire n_2741;
wire n_3114;
wire n_18298;
wire n_888;
wire n_13116;
wire n_2203;
wire n_14589;
wire n_5246;
wire n_236;
wire n_12386;
wire n_14257;
wire n_16492;
wire n_16811;
wire n_3836;
wire n_8835;
wire n_18645;
wire n_10688;
wire n_16771;
wire n_1215;
wire n_12964;
wire n_16404;
wire n_15099;
wire n_779;
wire n_2205;
wire n_7579;
wire n_16874;
wire n_4025;
wire n_11687;
wire n_4121;
wire n_8870;
wire n_7155;
wire n_4313;
wire n_6475;
wire n_7699;
wire n_15951;
wire n_6103;
wire n_5546;
wire n_232;
wire n_6394;
wire n_8781;
wire n_18618;
wire n_14102;
wire n_17196;
wire n_4246;
wire n_12267;
wire n_15803;
wire n_8365;
wire n_3690;
wire n_2483;
wire n_4532;
wire n_13780;
wire n_16699;
wire n_7194;
wire n_4049;
wire n_6752;
wire n_6426;
wire n_984;
wire n_5626;
wire n_8025;
wire n_8502;
wire n_7612;
wire n_16999;
wire n_18843;
wire n_11120;
wire n_6350;
wire n_7736;
wire n_16040;
wire n_14259;
wire n_5921;
wire n_3596;
wire n_4537;
wire n_6159;
wire n_13360;
wire n_2429;
wire n_8479;
wire n_14214;
wire n_15558;
wire n_3521;
wire n_802;
wire n_17306;
wire n_6235;
wire n_17996;
wire n_2360;
wire n_12647;
wire n_7662;
wire n_15340;
wire n_16061;
wire n_7773;
wire n_5340;
wire n_3947;
wire n_16776;
wire n_13048;
wire n_13563;
wire n_17905;
wire n_7555;
wire n_1194;
wire n_4506;
wire n_2742;
wire n_3695;
wire n_12060;
wire n_3976;
wire n_18254;
wire n_10199;
wire n_8658;
wire n_11910;
wire n_15377;
wire n_15583;
wire n_13347;
wire n_5925;
wire n_2909;
wire n_8866;
wire n_8061;
wire n_5730;
wire n_16623;
wire n_17186;
wire n_13111;
wire n_15563;
wire n_10117;
wire n_12716;
wire n_467;
wire n_16341;
wire n_16679;
wire n_13456;
wire n_10198;
wire n_7157;
wire n_13237;
wire n_15448;
wire n_857;
wire n_7411;
wire n_16851;
wire n_2221;
wire n_588;
wire n_7871;
wire n_12051;
wire n_1010;
wire n_6477;
wire n_15298;
wire n_11533;
wire n_8652;
wire n_534;
wire n_7198;
wire n_1578;
wire n_9904;
wire n_17891;
wire n_19182;
wire n_1557;
wire n_3945;
wire n_6184;
wire n_730;
wire n_5817;
wire n_10973;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_4278;
wire n_5586;
wire n_11036;
wire n_3433;
wire n_17362;
wire n_4463;
wire n_10267;
wire n_10551;
wire n_18589;
wire n_17029;
wire n_3833;
wire n_2774;
wire n_17924;
wire n_18323;
wire n_13127;
wire n_18004;
wire n_4129;
wire n_11002;
wire n_19637;
wire n_5032;
wire n_14075;
wire n_9032;
wire n_6313;
wire n_18884;
wire n_16184;
wire n_3965;
wire n_7145;
wire n_12325;
wire n_9245;
wire n_5065;
wire n_9357;
wire n_3085;
wire n_19060;
wire n_5826;
wire n_15766;
wire n_18121;
wire n_2991;
wire n_16759;
wire n_14530;
wire n_17724;
wire n_7994;
wire n_14206;
wire n_17328;
wire n_4703;
wire n_7349;
wire n_9598;
wire n_14481;
wire n_17993;
wire n_15044;
wire n_12504;
wire n_12602;
wire n_12062;
wire n_15375;
wire n_16100;
wire n_12335;
wire n_12949;
wire n_13611;
wire n_801;
wire n_4452;
wire n_15268;
wire n_4649;
wire n_5315;
wire n_10487;
wire n_5362;
wire n_2157;
wire n_10960;
wire n_6141;
wire n_18540;
wire n_3849;
wire n_10931;
wire n_11574;
wire n_15049;
wire n_15181;
wire n_8168;
wire n_3257;
wire n_14870;
wire n_7190;
wire n_1387;
wire n_12322;
wire n_1151;
wire n_14196;
wire n_2317;
wire n_5524;
wire n_10236;
wire n_11205;
wire n_11776;
wire n_11650;
wire n_5818;
wire n_5963;
wire n_19197;
wire n_12179;
wire n_14439;
wire n_9896;
wire n_11856;
wire n_14825;
wire n_11536;
wire n_5950;
wire n_1192;
wire n_14914;
wire n_1844;
wire n_10283;
wire n_5057;
wire n_3030;
wire n_5838;
wire n_6324;
wire n_13437;
wire n_15623;
wire n_2838;
wire n_5325;
wire n_16696;
wire n_18865;
wire n_2926;
wire n_8411;
wire n_2019;
wire n_5102;
wire n_16733;
wire n_18799;
wire n_13221;
wire n_2074;
wire n_2919;
wire n_11163;
wire n_13657;
wire n_945;
wire n_14099;
wire n_15632;
wire n_16245;
wire n_11419;
wire n_12095;
wire n_13990;
wire n_16302;
wire n_9018;
wire n_13663;
wire n_6660;
wire n_13298;
wire n_9055;
wire n_4347;
wire n_14939;
wire n_11740;
wire n_17471;
wire n_8444;
wire n_17227;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_12392;
wire n_11979;
wire n_7596;
wire n_6280;
wire n_18090;
wire n_18626;
wire n_2786;
wire n_10759;
wire n_9036;
wire n_9551;
wire n_13210;
wire n_18211;
wire n_8977;
wire n_15797;
wire n_9962;
wire n_2873;
wire n_11104;
wire n_3452;
wire n_3107;
wire n_11537;
wire n_13814;
wire n_18993;
wire n_12707;
wire n_15194;
wire n_7686;
wire n_1421;
wire n_14861;
wire n_1936;
wire n_5337;
wire n_18894;
wire n_15572;
wire n_12424;
wire n_1660;
wire n_3047;
wire n_11699;
wire n_8125;
wire n_14811;
wire n_17608;
wire n_10226;
wire n_6526;
wire n_1088;
wire n_17401;
wire n_7196;
wire n_3347;
wire n_907;
wire n_14864;
wire n_4110;
wire n_17936;
wire n_16643;
wire n_1658;
wire n_12107;
wire n_10161;
wire n_9842;
wire n_9614;
wire n_3999;
wire n_16024;
wire n_10699;
wire n_4751;
wire n_7846;
wire n_5151;
wire n_8598;
wire n_7256;
wire n_281;
wire n_16078;
wire n_7331;
wire n_13509;
wire n_17637;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_14791;
wire n_14485;
wire n_10606;
wire n_11164;
wire n_4296;
wire n_12203;
wire n_7147;
wire n_5902;
wire n_512;
wire n_12359;
wire n_19175;
wire n_5063;
wire n_9037;
wire n_1328;
wire n_15983;
wire n_12548;
wire n_15874;
wire n_3900;
wire n_3732;
wire n_14461;
wire n_2832;
wire n_4226;
wire n_1762;
wire n_13958;
wire n_17619;
wire n_3980;
wire n_4366;
wire n_6863;
wire n_10012;
wire n_13754;
wire n_12985;
wire n_4445;
wire n_2692;
wire n_16191;
wire n_14171;
wire n_6768;
wire n_4456;
wire n_15212;
wire n_15977;
wire n_9128;
wire n_9872;
wire n_14380;
wire n_10310;
wire n_15896;
wire n_6151;
wire n_16843;
wire n_7110;
wire n_5476;
wire n_17273;
wire n_13920;
wire n_18119;
wire n_2922;
wire n_10097;
wire n_3882;
wire n_2068;
wire n_8915;
wire n_16509;
wire n_9866;
wire n_9858;
wire n_2072;
wire n_586;
wire n_423;
wire n_4375;
wire n_13977;
wire n_8727;
wire n_18494;
wire n_3935;
wire n_5130;
wire n_16538;
wire n_11662;
wire n_1726;
wire n_16992;
wire n_2878;
wire n_18065;
wire n_3012;
wire n_10266;
wire n_17949;
wire n_4877;
wire n_2641;
wire n_8955;
wire n_7734;
wire n_178;
wire n_17781;
wire n_12384;
wire n_15438;
wire n_11260;
wire n_3298;
wire n_11351;
wire n_4467;
wire n_195;
wire n_780;
wire n_15611;
wire n_14388;
wire n_12249;
wire n_2350;
wire n_14977;
wire n_10628;
wire n_13429;
wire n_4220;
wire n_7905;
wire n_5281;
wire n_11775;
wire n_10769;
wire n_10256;
wire n_1654;
wire n_13999;
wire n_14037;
wire n_11706;
wire n_11800;
wire n_18382;
wire n_1588;
wire n_11642;
wire n_4381;
wire n_11143;
wire n_17103;
wire n_11074;
wire n_6831;
wire n_16352;
wire n_18713;
wire n_18032;
wire n_11934;
wire n_4473;
wire n_6043;
wire n_687;
wire n_7677;
wire n_5457;
wire n_10396;
wire n_13919;
wire n_19357;
wire n_190;
wire n_13642;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_1709;
wire n_10693;
wire n_2657;
wire n_15872;
wire n_13240;
wire n_949;
wire n_3500;
wire n_12578;
wire n_4589;
wire n_12194;
wire n_2972;
wire n_7519;
wire n_7400;
wire n_15649;
wire n_9724;
wire n_9281;
wire n_10101;
wire n_15863;
wire n_6581;
wire n_2279;
wire n_161;
wire n_7013;
wire n_14150;
wire n_12125;
wire n_7290;
wire n_18830;
wire n_595;
wire n_4921;
wire n_9687;
wire n_18052;
wire n_19108;
wire n_9426;
wire n_2712;
wire n_7889;
wire n_9102;
wire n_11526;
wire n_16115;
wire n_14128;
wire n_11851;
wire n_898;
wire n_18983;
wire n_17323;
wire n_6965;
wire n_9144;
wire n_18191;
wire n_7461;
wire n_15133;
wire n_16885;
wire n_4137;
wire n_9521;
wire n_15288;
wire n_16900;
wire n_13040;
wire n_963;
wire n_7278;
wire n_6509;
wire n_7454;
wire n_11253;
wire n_17102;
wire n_15527;
wire n_12861;
wire n_17443;
wire n_16146;
wire n_16654;
wire n_3400;
wire n_1521;
wire n_12918;
wire n_1366;
wire n_18332;
wire n_5501;
wire n_5342;
wire n_4345;
wire n_18145;
wire n_13353;
wire n_8648;
wire n_12388;
wire n_12102;
wire n_16991;
wire n_18051;
wire n_19051;
wire n_4664;
wire n_13716;
wire n_7069;
wire n_7904;
wire n_11691;
wire n_14408;
wire n_9410;
wire n_2643;
wire n_5748;
wire n_12865;
wire n_10712;
wire n_4713;
wire n_7168;
wire n_17604;
wire n_18765;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_3435;
wire n_842;
wire n_10972;
wire n_6359;
wire n_1432;
wire n_10945;
wire n_8800;
wire n_10845;
wire n_8229;
wire n_18743;
wire n_14863;
wire n_5811;
wire n_6766;
wire n_1035;
wire n_7629;
wire n_9735;
wire n_18831;
wire n_5397;
wire n_14711;
wire n_9802;
wire n_1448;
wire n_14373;
wire n_8107;
wire n_12992;
wire n_11108;
wire n_11004;
wire n_2445;
wire n_6519;
wire n_15752;
wire n_11686;
wire n_6530;
wire n_4440;
wire n_10566;
wire n_17798;
wire n_19592;
wire n_16568;
wire n_17581;
wire n_18906;
wire n_12104;
wire n_17954;
wire n_6402;
wire n_12469;
wire n_19554;
wire n_15829;
wire n_19568;
wire n_7326;
wire n_17522;
wire n_7067;
wire n_14835;
wire n_15391;
wire n_16226;
wire n_14871;
wire n_8691;
wire n_14907;
wire n_3342;
wire n_6748;
wire n_11719;
wire n_19307;
wire n_16685;
wire n_19498;
wire n_3656;
wire n_16979;
wire n_1424;
wire n_18282;
wire n_15358;
wire n_14636;
wire n_1507;
wire n_2482;
wire n_7528;
wire n_8026;
wire n_9638;
wire n_16069;
wire n_8174;
wire n_13524;
wire n_912;
wire n_11175;
wire n_10040;
wire n_2661;
wire n_8861;
wire n_5359;
wire n_8644;
wire n_931;
wire n_1791;
wire n_12304;
wire n_15156;
wire n_1897;
wire n_2064;
wire n_13138;
wire n_7117;
wire n_18490;
wire n_6205;
wire n_7136;
wire n_6754;
wire n_12692;
wire n_1334;
wire n_7939;
wire n_13602;
wire n_17436;
wire n_16785;
wire n_9612;
wire n_10790;
wire n_14919;
wire n_16653;
wire n_6723;
wire n_9108;
wire n_16692;
wire n_6440;
wire n_7436;
wire n_14101;
wire n_9376;
wire n_8446;
wire n_17654;
wire n_3534;
wire n_12996;
wire n_15171;
wire n_13625;
wire n_12643;
wire n_3944;
wire n_6124;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_19265;
wire n_1939;
wire n_8197;
wire n_2209;
wire n_6622;
wire n_11521;
wire n_12827;
wire n_12678;
wire n_15868;
wire n_1053;
wire n_17249;
wire n_7747;
wire n_9779;
wire n_8082;
wire n_8730;
wire n_15533;
wire n_266;
wire n_6528;
wire n_15165;
wire n_13475;
wire n_15079;
wire n_13859;
wire n_18640;
wire n_1745;
wire n_3479;
wire n_12713;
wire n_13144;
wire n_18129;
wire n_488;
wire n_19488;
wire n_10660;
wire n_7430;
wire n_18560;
wire n_9937;
wire n_5679;
wire n_7912;
wire n_5100;
wire n_16749;
wire n_5973;
wire n_8281;
wire n_4807;
wire n_1243;
wire n_301;
wire n_2928;
wire n_5166;
wire n_19437;
wire n_18876;
wire n_19430;
wire n_11428;
wire n_2822;
wire n_17626;
wire n_1281;
wire n_11677;
wire n_7281;
wire n_9717;
wire n_13577;
wire n_2572;
wire n_1520;
wire n_3126;
wire n_18523;
wire n_1419;
wire n_19176;
wire n_5688;
wire n_13769;
wire n_18044;
wire n_4676;
wire n_13672;
wire n_19036;
wire n_17600;
wire n_6763;
wire n_8956;
wire n_7858;
wire n_663;
wire n_4880;
wire n_6542;
wire n_15681;
wire n_2781;
wire n_4126;
wire n_17262;
wire n_1696;
wire n_6556;
wire n_12374;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_8998;
wire n_10538;
wire n_1790;
wire n_4014;
wire n_13342;
wire n_18856;
wire n_9123;
wire n_17374;
wire n_6471;
wire n_5949;
wire n_15545;
wire n_4048;
wire n_14924;
wire n_4444;
wire n_11867;
wire n_12796;
wire n_3919;
wire n_16053;
wire n_19185;
wire n_15708;
wire n_19441;
wire n_11716;
wire n_8979;
wire n_7245;
wire n_18858;
wire n_6675;
wire n_6270;
wire n_18111;
wire n_6808;
wire n_2884;
wire n_16091;
wire n_11886;
wire n_7006;
wire n_16264;
wire n_14160;
wire n_6245;
wire n_14932;
wire n_17231;
wire n_3797;
wire n_10925;
wire n_4770;
wire n_11158;
wire n_9861;
wire n_15878;
wire n_2549;
wire n_4690;
wire n_14390;
wire n_18678;
wire n_8264;
wire n_7381;
wire n_16160;
wire n_12078;
wire n_15647;
wire n_9832;
wire n_6580;
wire n_18790;
wire n_9898;
wire n_5500;
wire n_6412;
wire n_18410;
wire n_183;
wire n_13293;
wire n_3967;
wire n_6437;
wire n_14381;
wire n_2526;
wire n_15709;
wire n_18590;
wire n_8408;
wire n_3277;
wire n_10661;
wire n_9495;
wire n_10028;
wire n_13878;
wire n_15000;
wire n_11771;
wire n_16870;
wire n_19082;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_13833;
wire n_16518;
wire n_1960;
wire n_2694;
wire n_1686;
wire n_9867;
wire n_6059;
wire n_14441;
wire n_9688;
wire n_5094;
wire n_10967;
wire n_7870;
wire n_3228;
wire n_18377;
wire n_3657;
wire n_1287;
wire n_6117;
wire n_11828;
wire n_12326;
wire n_1586;
wire n_14264;
wire n_19317;
wire n_14115;
wire n_16635;
wire n_3464;
wire n_380;
wire n_8963;
wire n_4380;
wire n_5247;
wire n_4996;
wire n_4398;
wire n_4193;
wire n_3570;
wire n_12309;
wire n_7399;
wire n_3828;
wire n_1539;
wire n_13953;
wire n_7482;
wire n_14847;
wire n_10312;
wire n_4090;
wire n_18308;
wire n_9223;
wire n_17465;
wire n_15930;
wire n_13226;
wire n_5931;
wire n_19416;
wire n_2371;
wire n_17943;
wire n_662;
wire n_16433;
wire n_3262;
wire n_11244;
wire n_4008;
wire n_18577;
wire n_14432;
wire n_1642;
wire n_10209;
wire n_13253;
wire n_4689;
wire n_8183;
wire n_16098;
wire n_4547;
wire n_11245;
wire n_13354;
wire n_6085;
wire n_12422;
wire n_15616;
wire n_17614;
wire n_3329;
wire n_14422;
wire n_9694;
wire n_3826;
wire n_16636;
wire n_9948;
wire n_14630;
wire n_17048;
wire n_3681;
wire n_18966;
wire n_19390;
wire n_10887;
wire n_16876;
wire n_5883;
wire n_6554;
wire n_12146;
wire n_5754;
wire n_6560;
wire n_14055;
wire n_1720;
wire n_12136;
wire n_17046;
wire n_16138;
wire n_12399;
wire n_942;
wire n_12342;
wire n_7414;
wire n_9744;
wire n_9548;
wire n_8973;
wire n_6448;
wire n_1964;
wire n_12378;
wire n_19155;
wire n_12533;
wire n_5434;
wire n_5934;
wire n_7431;
wire n_12178;
wire n_18871;
wire n_11346;
wire n_17210;
wire n_2626;
wire n_5880;
wire n_18206;
wire n_14810;
wire n_8249;
wire n_12257;
wire n_3528;
wire n_15770;
wire n_13394;
wire n_13391;
wire n_14680;
wire n_8234;
wire n_16835;
wire n_1066;
wire n_18438;
wire n_16863;
wire n_9280;
wire n_18285;
wire n_13263;
wire n_14877;
wire n_5145;
wire n_15203;
wire n_1229;
wire n_11491;
wire n_14048;
wire n_2427;
wire n_11772;
wire n_16063;
wire n_16237;
wire n_16112;
wire n_15891;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_12769;
wire n_4190;
wire n_5149;
wire n_12641;
wire n_10765;
wire n_3375;
wire n_15263;
wire n_11792;
wire n_18776;
wire n_2668;
wire n_8558;
wire n_10489;
wire n_12421;
wire n_2128;
wire n_7274;
wire n_10159;
wire n_14351;
wire n_7466;
wire n_1002;
wire n_13310;
wire n_2508;
wire n_11568;
wire n_2054;
wire n_7429;
wire n_11766;
wire n_11038;
wire n_13798;
wire n_16894;
wire n_18890;
wire n_17294;
wire n_16932;
wire n_15842;
wire n_14822;
wire n_2758;
wire n_8813;
wire n_10356;
wire n_17461;
wire n_18216;
wire n_10173;
wire n_4789;
wire n_19162;
wire n_12311;
wire n_14374;
wire n_2241;
wire n_6555;
wire n_14815;
wire n_9448;
wire n_10739;
wire n_8470;
wire n_1690;
wire n_5341;
wire n_16480;
wire n_4512;
wire n_1378;
wire n_17657;
wire n_14831;
wire n_11170;
wire n_17683;
wire n_11758;
wire n_1542;
wire n_9396;
wire n_19486;
wire n_14450;
wire n_7061;
wire n_12480;
wire n_14192;
wire n_1716;
wire n_278;
wire n_9053;
wire n_15504;
wire n_11893;
wire n_10573;
wire n_3303;
wire n_4324;
wire n_10850;
wire n_384;
wire n_9185;
wire n_13376;
wire n_2905;
wire n_8092;
wire n_13864;
wire n_3954;
wire n_15279;
wire n_11456;
wire n_10546;
wire n_5622;
wire n_3160;
wire n_6574;
wire n_6571;
wire n_17484;
wire n_143;
wire n_9151;
wire n_7824;
wire n_17202;
wire n_18080;
wire n_698;
wire n_13236;
wire n_3569;
wire n_14299;
wire n_7094;
wire n_2528;
wire n_16320;
wire n_4639;
wire n_7036;
wire n_13777;
wire n_19359;
wire n_1730;
wire n_814;
wire n_5779;
wire n_2020;
wire n_6260;
wire n_7413;
wire n_16803;
wire n_17229;
wire n_6286;
wire n_8267;
wire n_4023;
wire n_18929;
wire n_721;
wire n_7175;
wire n_6019;
wire n_4344;
wire n_9978;
wire n_11914;
wire n_9670;
wire n_3154;
wire n_9334;
wire n_15131;
wire n_3898;
wire n_12531;
wire n_4391;
wire n_11302;
wire n_946;
wire n_1303;
wire n_19006;
wire n_4095;
wire n_9413;
wire n_12727;
wire n_15509;
wire n_3551;
wire n_3064;
wire n_11707;
wire n_1689;
wire n_7697;
wire n_1944;
wire n_13835;
wire n_16260;
wire n_7547;
wire n_6013;
wire n_13815;
wire n_9557;
wire n_15957;
wire n_16319;
wire n_448;
wire n_3853;
wire n_17259;
wire n_14039;
wire n_6348;
wire n_6744;
wire n_18578;
wire n_8582;
wire n_5068;
wire n_6293;
wire n_234;
wire n_6049;
wire n_1460;
wire n_9762;
wire n_8957;
wire n_18646;
wire n_15793;
wire n_6558;
wire n_12227;
wire n_12258;
wire n_14117;
wire n_18209;
wire n_2437;
wire n_2444;
wire n_9271;
wire n_17747;
wire n_3035;
wire n_13688;
wire n_4166;
wire n_11396;
wire n_15196;
wire n_16176;
wire n_9483;
wire n_19649;
wire n_1058;
wire n_19435;
wire n_14754;
wire n_15020;
wire n_2934;
wire n_6091;
wire n_14252;
wire n_15830;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_8747;
wire n_9539;
wire n_4817;
wire n_2014;
wire n_9385;
wire n_1584;
wire n_13462;
wire n_5381;
wire n_9785;
wire n_3468;
wire n_8922;
wire n_9027;
wire n_12750;
wire n_4383;
wire n_6995;
wire n_5696;
wire n_455;
wire n_4486;
wire n_19315;
wire n_9233;
wire n_3024;
wire n_16895;
wire n_10282;
wire n_17602;
wire n_4529;
wire n_500;
wire n_15142;
wire n_291;
wire n_10913;
wire n_18803;
wire n_18409;
wire n_17838;
wire n_15991;
wire n_5823;
wire n_13388;
wire n_2800;
wire n_13731;
wire n_10703;
wire n_9666;
wire n_14503;
wire n_12248;
wire n_8678;
wire n_10565;
wire n_10011;
wire n_17754;
wire n_14886;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_3161;
wire n_2799;
wire n_14644;
wire n_11715;
wire n_7071;
wire n_15454;
wire n_10642;
wire n_15213;
wire n_756;
wire n_18859;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_18428;
wire n_12181;
wire n_18670;
wire n_14560;
wire n_17257;
wire n_3992;
wire n_14829;
wire n_15473;
wire n_11007;
wire n_249;
wire n_15584;
wire n_3125;
wire n_10316;
wire n_9795;
wire n_18386;
wire n_4684;
wire n_3116;
wire n_6429;
wire n_6407;
wire n_16515;
wire n_5027;
wire n_17914;
wire n_10479;
wire n_13660;
wire n_19280;
wire n_6801;
wire n_1921;
wire n_18099;
wire n_5630;
wire n_12738;
wire n_4057;
wire n_15062;
wire n_1170;
wire n_5379;
wire n_11599;
wire n_308;
wire n_3444;
wire n_6113;
wire n_10070;
wire n_16178;
wire n_1890;
wire n_18841;
wire n_2477;
wire n_17304;
wire n_18393;
wire n_14983;
wire n_2333;
wire n_8439;
wire n_18434;
wire n_9641;
wire n_1089;
wire n_12755;
wire n_18522;
wire n_12059;
wire n_18541;
wire n_18257;
wire n_15845;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_9138;
wire n_18072;
wire n_18048;
wire n_7537;
wire n_10516;
wire n_8675;
wire n_1616;
wire n_15924;
wire n_17906;
wire n_12567;
wire n_9367;
wire n_15130;
wire n_4197;
wire n_4482;
wire n_2547;
wire n_2415;
wire n_11887;
wire n_17852;
wire n_17442;
wire n_10026;
wire n_9729;
wire n_5073;
wire n_827;
wire n_12471;
wire n_12451;
wire n_17243;
wire n_15740;
wire n_9411;
wire n_3660;
wire n_3766;
wire n_12507;
wire n_1027;
wire n_3266;
wire n_3574;
wire n_14564;
wire n_11277;
wire n_4907;
wire n_5077;
wire n_18416;
wire n_17606;
wire n_7410;
wire n_365;
wire n_8777;
wire n_2534;
wire n_4975;
wire n_13581;
wire n_2451;
wire n_12972;
wire n_13789;
wire n_4815;
wire n_14511;
wire n_13286;
wire n_9951;
wire n_396;
wire n_19023;
wire n_9424;
wire n_480;
wire n_4134;
wire n_10507;
wire n_11968;
wire n_19003;
wire n_1238;
wire n_4092;
wire n_10045;
wire n_11335;
wire n_18606;
wire n_13988;
wire n_4755;
wire n_4960;
wire n_1700;
wire n_15272;
wire n_4933;
wire n_17169;
wire n_13609;
wire n_4591;
wire n_5528;
wire n_16886;
wire n_5111;
wire n_13679;
wire n_11785;
wire n_873;
wire n_10417;
wire n_3946;
wire n_12841;
wire n_12855;
wire n_17370;
wire n_15834;
wire n_13276;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_16058;
wire n_2509;
wire n_11801;
wire n_16994;
wire n_16519;
wire n_3757;
wire n_17810;
wire n_1704;
wire n_250;
wire n_4884;
wire n_14830;
wire n_7867;
wire n_14281;
wire n_14594;
wire n_18213;
wire n_6135;
wire n_17303;
wire n_3678;
wire n_6814;
wire n_10557;
wire n_8669;
wire n_7525;
wire n_19219;
wire n_7257;
wire n_9372;
wire n_4692;
wire n_6791;
wire n_616;
wire n_3165;
wire n_11915;
wire n_13704;
wire n_11016;
wire n_9326;
wire n_14976;
wire n_1902;
wire n_1735;
wire n_3890;
wire n_641;
wire n_3750;
wire n_7650;
wire n_17297;
wire n_13043;
wire n_4311;
wire n_4722;
wire n_17260;
wire n_12620;
wire n_12632;
wire n_6309;
wire n_19618;
wire n_11303;
wire n_405;
wire n_213;
wire n_6733;
wire n_19047;
wire n_1094;
wire n_5430;
wire n_5942;
wire n_9902;
wire n_4820;
wire n_9900;
wire n_17367;
wire n_18937;
wire n_15521;
wire n_18415;
wire n_7202;
wire n_12416;
wire n_8265;
wire n_4619;
wire n_5762;
wire n_11609;
wire n_1961;
wire n_18287;
wire n_16464;
wire n_5036;
wire n_4221;
wire n_19597;
wire n_3297;
wire n_12494;
wire n_10327;
wire n_13826;
wire n_7605;
wire n_11556;
wire n_15140;
wire n_11529;
wire n_10437;
wire n_10021;
wire n_16673;
wire n_9146;
wire n_15753;
wire n_2996;
wire n_8131;
wire n_8941;
wire n_5014;
wire n_17093;
wire n_17685;
wire n_16357;
wire n_12623;
wire n_11444;
wire n_659;
wire n_6269;
wire n_5233;
wire n_12213;
wire n_6654;
wire n_9358;
wire n_3164;
wire n_9565;
wire n_8257;
wire n_13072;
wire n_18120;
wire n_7726;
wire n_5436;
wire n_17026;
wire n_13839;
wire n_594;
wire n_6120;
wire n_6068;
wire n_4141;
wire n_13954;
wire n_8799;
wire n_2850;
wire n_572;
wire n_6641;
wire n_5789;
wire n_2104;
wire n_19215;
wire n_10124;
wire n_19595;
wire n_14689;
wire n_10245;
wire n_14132;
wire n_10905;
wire n_11235;
wire n_19020;
wire n_6399;
wire n_4499;
wire n_5195;
wire n_9563;
wire n_17077;
wire n_17702;
wire n_11166;
wire n_7031;
wire n_9285;
wire n_263;
wire n_18093;
wire n_16595;
wire n_7763;
wire n_1543;
wire n_8033;
wire n_1599;
wire n_15172;
wire n_4458;
wire n_19470;
wire n_5103;
wire n_8393;
wire n_16561;
wire n_10784;
wire n_1876;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_10944;
wire n_10211;
wire n_18554;
wire n_18077;
wire n_12431;
wire n_11855;
wire n_6790;
wire n_3099;
wire n_17628;
wire n_13799;
wire n_16084;
wire n_13854;
wire n_18250;
wire n_15380;
wire n_2457;
wire n_6686;
wire n_15956;
wire n_4119;
wire n_18835;
wire n_11787;
wire n_5958;
wire n_16059;
wire n_8103;
wire n_2971;
wire n_715;
wire n_4526;
wire n_14752;
wire n_5792;
wire n_6183;
wire n_11544;
wire n_15447;
wire n_10730;
wire n_2028;
wire n_1069;
wire n_10564;
wire n_8682;
wire n_7655;
wire n_18276;
wire n_4485;
wire n_1504;
wire n_11509;
wire n_19191;
wire n_11960;
wire n_1801;
wire n_3917;
wire n_7878;
wire n_9514;
wire n_6210;
wire n_6500;
wire n_12465;
wire n_2206;
wire n_13532;
wire n_11029;
wire n_13118;
wire n_17390;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_19415;
wire n_6785;
wire n_10454;
wire n_15401;
wire n_13339;
wire n_4940;
wire n_8039;
wire n_5757;
wire n_19323;
wire n_8916;
wire n_10087;
wire n_3510;
wire n_10146;
wire n_12959;
wire n_9946;
wire n_9885;
wire n_6849;
wire n_8162;
wire n_18263;
wire n_7457;
wire n_8744;
wire n_5488;
wire n_10701;
wire n_3827;
wire n_891;
wire n_2067;
wire n_7752;
wire n_15775;
wire n_4245;
wire n_17346;
wire n_8286;
wire n_9015;
wire n_6452;
wire n_16408;
wire n_1008;
wire n_6611;
wire n_4560;
wire n_18828;
wire n_4899;
wire n_18297;
wire n_5471;
wire n_11433;
wire n_10592;
wire n_5164;
wire n_18130;
wire n_7207;
wire n_8218;
wire n_17978;
wire n_1767;
wire n_8537;
wire n_10126;
wire n_14421;
wire n_15890;
wire n_4663;
wire n_2893;
wire n_13653;
wire n_5484;
wire n_12566;
wire n_6227;
wire n_13680;
wire n_3421;
wire n_16077;
wire n_9066;
wire n_10302;
wire n_12546;
wire n_13058;
wire n_18342;
wire n_12036;
wire n_17650;
wire n_8782;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_12911;
wire n_15715;
wire n_9857;
wire n_12781;
wire n_10057;
wire n_10882;
wire n_894;
wire n_9338;
wire n_353;
wire n_8144;
wire n_10435;
wire n_9542;
wire n_10921;
wire n_7171;
wire n_12061;
wire n_3922;
wire n_14585;
wire n_11085;
wire n_16541;
wire n_7068;
wire n_13649;
wire n_10609;
wire n_14804;
wire n_2554;
wire n_9783;
wire n_13806;
wire n_19542;
wire n_4934;
wire n_9404;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_18351;
wire n_16198;
wire n_14466;
wire n_7777;
wire n_12138;
wire n_2765;
wire n_5403;
wire n_2590;
wire n_7652;
wire n_10220;
wire n_3150;
wire n_11347;
wire n_17635;
wire n_4479;
wire n_2608;
wire n_10550;
wire n_14673;
wire n_12365;
wire n_1959;
wire n_3133;
wire n_13738;
wire n_14972;
wire n_765;
wire n_1492;
wire n_16996;
wire n_9306;
wire n_14138;
wire n_1340;
wire n_10232;
wire n_10461;
wire n_14586;
wire n_7966;
wire n_8591;
wire n_8811;
wire n_19188;
wire n_1277;
wire n_14031;
wire n_5242;
wire n_10326;
wire n_8417;
wire n_2675;
wire n_5631;
wire n_6008;
wire n_3887;
wire n_12487;
wire n_7997;
wire n_6420;
wire n_4587;
wire n_1577;
wire n_12288;
wire n_17300;
wire n_1117;
wire n_12130;
wire n_13120;
wire n_3223;
wire n_16299;
wire n_12271;
wire n_12704;
wire n_7680;
wire n_15190;
wire n_16909;
wire n_12958;
wire n_8172;
wire n_19559;
wire n_9502;
wire n_6447;
wire n_5981;
wire n_3788;
wire n_4891;
wire n_14761;
wire n_6751;
wire n_2718;
wire n_15243;
wire n_1384;
wire n_11087;
wire n_11477;
wire n_3325;
wire n_2238;
wire n_8375;
wire n_8612;
wire n_4624;
wire n_8345;
wire n_13725;
wire n_3600;
wire n_6741;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_5015;
wire n_1178;
wire n_2338;
wire n_19414;
wire n_17551;
wire n_19417;
wire n_9164;
wire n_7183;
wire n_13197;
wire n_10878;
wire n_18408;
wire n_7140;
wire n_14860;
wire n_10450;
wire n_623;
wire n_19609;
wire n_11472;
wire n_9114;
wire n_11978;
wire n_8515;
wire n_10529;
wire n_1502;
wire n_14685;
wire n_5773;
wire n_5482;
wire n_14892;
wire n_8812;
wire n_14505;
wire n_12254;
wire n_9392;
wire n_1250;
wire n_14531;
wire n_3615;
wire n_11538;
wire n_3087;
wire n_2121;
wire n_9698;
wire n_13435;
wire n_15408;
wire n_15173;
wire n_4015;
wire n_477;
wire n_9644;
wire n_11353;
wire n_18745;
wire n_2213;
wire n_2389;
wire n_9499;
wire n_2892;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_14771;
wire n_1564;
wire n_5296;
wire n_3718;
wire n_7750;
wire n_11597;
wire n_537;
wire n_15902;
wire n_6277;
wire n_1919;
wire n_3705;
wire n_3211;
wire n_546;
wire n_10920;
wire n_14398;
wire n_3582;
wire n_11126;
wire n_4223;
wire n_5674;
wire n_18453;
wire n_5282;
wire n_9409;
wire n_18629;
wire n_1060;
wire n_1951;
wire n_17814;
wire n_12555;
wire n_11646;
wire n_1223;
wire n_5121;
wire n_9768;
wire n_6070;
wire n_1286;
wire n_12980;
wire n_9881;
wire n_5013;
wire n_6807;
wire n_7251;
wire n_4489;
wire n_7254;
wire n_18178;
wire n_12973;
wire n_3163;
wire n_17313;
wire n_13123;
wire n_14669;
wire n_5589;
wire n_12234;
wire n_10776;
wire n_7882;
wire n_16348;
wire n_16514;
wire n_17704;
wire n_10848;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_11482;
wire n_1625;
wire n_5006;
wire n_7816;
wire n_2226;
wire n_2801;
wire n_10164;
wire n_15809;
wire n_1901;
wire n_3869;
wire n_15579;
wire n_18549;
wire n_18084;
wire n_15585;
wire n_3753;
wire n_12033;
wire n_1892;
wire n_1614;
wire n_3742;
wire n_14376;
wire n_3260;
wire n_9595;
wire n_18978;
wire n_15555;
wire n_13923;
wire n_13051;
wire n_11524;
wire n_17220;
wire n_9265;
wire n_8239;
wire n_16114;
wire n_13330;
wire n_2159;
wire n_2315;
wire n_11228;
wire n_5273;
wire n_7898;
wire n_18286;
wire n_9789;
wire n_5936;
wire n_7646;
wire n_17537;
wire n_3220;
wire n_14627;
wire n_13699;
wire n_6069;
wire n_171;
wire n_169;
wire n_7665;
wire n_9354;
wire n_10501;
wire n_14026;
wire n_2379;
wire n_17782;
wire n_9436;
wire n_18157;
wire n_8489;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_12730;
wire n_6887;
wire n_18926;
wire n_16123;
wire n_13152;
wire n_17221;
wire n_4374;
wire n_6637;
wire n_9238;
wire n_358;
wire n_6633;
wire n_2420;
wire n_11031;
wire n_3722;
wire n_186;
wire n_4400;
wire n_17365;
wire n_9839;
wire n_18479;
wire n_15704;
wire n_7900;
wire n_6569;
wire n_10807;
wire n_12478;
wire n_2538;
wire n_724;
wire n_3250;
wire n_17265;
wire n_13545;
wire n_557;
wire n_13760;
wire n_1871;
wire n_13883;
wire n_10511;
wire n_7576;
wire n_19499;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_2102;
wire n_10873;
wire n_14484;
wire n_7676;
wire n_18956;
wire n_9017;
wire n_4304;
wire n_15726;
wire n_14307;
wire n_2544;
wire n_15302;
wire n_8865;
wire n_10337;
wire n_7779;
wire n_8999;
wire n_1206;
wire n_11626;
wire n_12148;
wire n_16872;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_16312;
wire n_16204;
wire n_8820;
wire n_16793;
wire n_16443;
wire n_6090;
wire n_18456;
wire n_5515;
wire n_3131;
wire n_18281;
wire n_12132;
wire n_1298;
wire n_10593;
wire n_5862;
wire n_16801;
wire n_2088;
wire n_12182;
wire n_12043;
wire n_10636;
wire n_16478;
wire n_18489;
wire n_5697;
wire n_2401;
wire n_18723;
wire n_8992;
wire n_8880;
wire n_8690;
wire n_2900;
wire n_6234;
wire n_3994;
wire n_1497;
wire n_7818;
wire n_11721;
wire n_13573;
wire n_19019;
wire n_6608;
wire n_9109;
wire n_5498;
wire n_2571;
wire n_3138;
wire n_7896;
wire n_12482;
wire n_18839;
wire n_15208;
wire n_6860;
wire n_12137;
wire n_12306;
wire n_11328;
wire n_2988;
wire n_1350;
wire n_11200;
wire n_14442;
wire n_15210;
wire n_4109;
wire n_16536;
wire n_13418;
wire n_5175;
wire n_7996;
wire n_986;
wire n_10533;
wire n_460;
wire n_5987;
wire n_16681;
wire n_10176;
wire n_7517;
wire n_8080;
wire n_450;
wire n_4150;
wire n_12345;
wire n_13551;
wire n_19135;
wire n_19178;
wire n_16060;
wire n_8772;
wire n_8786;
wire n_15597;
wire n_4643;
wire n_12694;
wire n_8083;
wire n_10155;
wire n_1332;
wire n_9805;
wire n_13593;
wire n_8157;
wire n_2346;
wire n_19660;
wire n_936;
wire n_3821;
wire n_13902;
wire n_3676;
wire n_4896;
wire n_3675;
wire n_9110;
wire n_18358;
wire n_5904;
wire n_599;
wire n_14468;
wire n_6062;
wire n_12550;
wire n_13861;
wire n_13350;
wire n_10051;
wire n_4209;
wire n_10414;
wire n_8344;
wire n_17597;
wire n_1341;
wire n_8120;
wire n_3003;
wire n_9075;
wire n_12961;
wire n_18882;
wire n_11496;
wire n_4128;
wire n_12225;
wire n_4271;
wire n_2258;
wire n_8621;
wire n_12884;
wire n_325;
wire n_5845;
wire n_19171;
wire n_6246;
wire n_8868;
wire n_8134;
wire n_4716;
wire n_12207;
wire n_9975;
wire n_1782;
wire n_5600;
wire n_12011;
wire n_707;
wire n_6053;
wire n_7252;
wire n_3246;
wire n_6843;
wire n_4715;
wire n_10626;
wire n_6901;
wire n_19014;
wire n_13273;
wire n_4694;
wire n_18855;
wire n_8101;
wire n_5448;
wire n_6489;
wire n_7402;
wire n_737;
wire n_3517;
wire n_3893;
wire n_19552;
wire n_11273;
wire n_138;
wire n_19089;
wire n_16954;
wire n_12472;
wire n_19526;
wire n_14035;
wire n_13218;
wire n_9081;
wire n_333;
wire n_4084;
wire n_9236;
wire n_6844;
wire n_11762;
wire n_459;
wire n_4850;
wire n_10156;
wire n_9607;
wire n_2840;
wire n_6779;
wire n_10774;
wire n_12332;
wire n_7216;
wire n_3855;
wire n_15990;
wire n_15364;
wire n_3091;
wire n_6543;
wire n_19585;
wire n_6178;
wire n_9621;
wire n_3398;
wire n_5685;
wire n_18075;
wire n_2793;
wire n_4235;
wire n_16117;
wire n_10398;
wire n_17947;
wire n_16459;
wire n_774;
wire n_17987;
wire n_18165;
wire n_15661;
wire n_17932;
wire n_7706;
wire n_1860;
wire n_5016;
wire n_479;
wire n_6458;
wire n_7642;
wire n_1777;
wire n_12506;
wire n_18356;
wire n_3308;
wire n_12718;
wire n_1600;
wire n_2253;
wire n_12638;
wire n_14116;
wire n_4799;
wire n_2261;
wire n_18710;
wire n_2516;
wire n_16453;
wire n_16645;
wire n_1177;
wire n_10470;
wire n_15034;
wire n_14240;
wire n_14504;
wire n_13449;
wire n_12747;
wire n_10625;
wire n_12561;
wire n_18420;
wire n_5514;
wire n_8388;
wire n_18469;
wire n_14730;
wire n_18732;
wire n_9589;
wire n_4543;
wire n_10445;
wire n_15110;
wire n_8988;
wire n_15025;
wire n_19329;
wire n_18161;
wire n_12900;
wire n_18761;
wire n_8569;
wire n_14598;
wire n_3255;
wire n_1401;
wire n_10679;
wire n_1516;
wire n_11323;
wire n_10799;
wire n_2029;
wire n_5890;
wire n_17228;
wire n_1394;
wire n_10585;
wire n_18519;
wire n_13696;
wire n_12948;
wire n_7931;
wire n_13322;
wire n_9092;
wire n_10034;
wire n_935;
wire n_11148;
wire n_9451;
wire n_18729;
wire n_13934;
wire n_6899;
wire n_7373;
wire n_7895;
wire n_676;
wire n_15331;
wire n_17109;
wire n_832;
wire n_13254;
wire n_3049;
wire n_15191;
wire n_17617;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_18783;
wire n_15676;
wire n_17044;
wire n_9011;
wire n_7613;
wire n_3541;
wire n_6101;
wire n_14440;
wire n_7556;
wire n_5935;
wire n_10528;
wire n_372;
wire n_314;
wire n_13875;
wire n_17319;
wire n_17774;
wire n_338;
wire n_19255;
wire n_14076;
wire n_506;
wire n_11220;
wire n_17709;
wire n_9012;
wire n_2396;
wire n_18150;
wire n_2450;
wire n_14638;
wire n_2284;
wire n_7238;
wire n_2769;
wire n_14936;
wire n_16469;
wire n_8047;
wire n_11596;
wire n_6273;
wire n_5663;
wire n_525;
wire n_7572;
wire n_11955;
wire n_1677;
wire n_18818;
wire n_16156;
wire n_11654;
wire n_18361;
wire n_12982;
wire n_4160;
wire n_4231;
wire n_11619;
wire n_10649;
wire n_2779;
wire n_5203;
wire n_19638;
wire n_6311;
wire n_7590;
wire n_5162;
wire n_1464;
wire n_5285;
wire n_2721;
wire n_12275;
wire n_13742;
wire n_270;
wire n_15177;
wire n_12376;
wire n_563;
wire n_13114;
wire n_8583;
wire n_4521;
wire n_10447;
wire n_15063;
wire n_7176;
wire n_9353;
wire n_13054;
wire n_8948;
wire n_5715;
wire n_8295;
wire n_498;
wire n_5395;
wire n_10522;
wire n_13793;
wire n_11782;
wire n_16532;
wire n_1693;
wire n_16618;
wire n_10278;
wire n_15384;
wire n_13882;
wire n_9750;
wire n_14139;
wire n_9749;
wire n_2915;
wire n_15686;
wire n_9263;
wire n_11082;
wire n_1989;
wire n_15950;
wire n_2802;
wire n_6181;
wire n_7447;
wire n_17998;
wire n_19156;
wire n_18928;
wire n_12721;
wire n_18301;
wire n_5672;
wire n_16008;
wire n_11730;
wire n_3098;
wire n_6924;
wire n_9804;
wire n_1851;
wire n_9304;
wire n_5799;
wire n_8380;
wire n_12039;
wire n_3123;
wire n_3380;
wire n_5617;
wire n_10377;
wire n_9926;
wire n_570;
wire n_15161;
wire n_620;
wire n_2523;
wire n_10858;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_1482;
wire n_16303;
wire n_9843;
wire n_3130;
wire n_16559;
wire n_1710;
wire n_13320;
wire n_1301;
wire n_6683;
wire n_10683;
wire n_2282;
wire n_9921;
wire n_19606;
wire n_6229;
wire n_1609;
wire n_13488;
wire n_15907;
wire n_7286;
wire n_13668;
wire n_13016;
wire n_6177;
wire n_16961;
wire n_14708;
wire n_2867;
wire n_2726;
wire n_17293;
wire n_12048;
wire n_5982;
wire n_10930;
wire n_17972;
wire n_8749;
wire n_18264;
wire n_2662;
wire n_12057;
wire n_6696;
wire n_17590;
wire n_9527;
wire n_16450;
wire n_19651;
wire n_2795;
wire n_18352;
wire n_14875;
wire n_3472;
wire n_15056;
wire n_15860;
wire n_19460;
wire n_17288;
wire n_5376;
wire n_16197;
wire n_14003;
wire n_5106;
wire n_9511;
wire n_6730;
wire n_17822;
wire n_13670;
wire n_11254;
wire n_15023;
wire n_11617;
wire n_18184;
wire n_5561;
wire n_404;
wire n_158;
wire n_18436;
wire n_6170;
wire n_9459;
wire n_14185;
wire n_6094;
wire n_9098;
wire n_14953;
wire n_15604;
wire n_4826;
wire n_16000;
wire n_3903;
wire n_12360;
wire n_9268;
wire n_17116;
wire n_15431;
wire n_3854;
wire n_3235;
wire n_8673;
wire n_18702;
wire n_19174;
wire n_5378;
wire n_10456;
wire n_3673;
wire n_13186;
wire n_18824;
wire n_5916;
wire n_15655;
wire n_11907;
wire n_3094;
wire n_10627;
wire n_10475;
wire n_965;
wire n_1428;
wire n_15430;
wire n_1576;
wire n_2077;
wire n_8581;
wire n_15732;
wire n_12457;
wire n_16070;
wire n_16045;
wire n_4951;
wire n_17772;
wire n_540;
wire n_14170;
wire n_3070;
wire n_13496;
wire n_8058;
wire n_9308;
wire n_3504;
wire n_11838;
wire n_10508;
wire n_18008;
wire n_10811;
wire n_18696;
wire n_8333;
wire n_17152;
wire n_7619;
wire n_6985;
wire n_18551;
wire n_7170;
wire n_13853;
wire n_8823;
wire n_11457;
wire n_12751;
wire n_15284;
wire n_3054;
wire n_5399;
wire n_4620;
wire n_5421;
wire n_4127;
wire n_17901;
wire n_15443;
wire n_5206;
wire n_18228;
wire n_17833;
wire n_18471;
wire n_4517;
wire n_16852;
wire n_18817;
wire n_6916;
wire n_15524;
wire n_2260;
wire n_10725;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_18354;
wire n_8290;
wire n_7536;
wire n_1743;
wire n_18152;
wire n_6230;
wire n_16108;
wire n_11107;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_12757;
wire n_14379;
wire n_8840;
wire n_16284;
wire n_16001;
wire n_18873;
wire n_13189;
wire n_5881;
wire n_18915;
wire n_2382;
wire n_3754;
wire n_19492;
wire n_12328;
wire n_415;
wire n_9083;
wire n_17271;
wire n_383;
wire n_2974;
wire n_4213;
wire n_200;
wire n_6483;
wire n_10994;
wire n_14004;
wire n_17023;
wire n_5863;
wire n_2645;
wire n_16221;
wire n_3904;
wire n_8036;
wire n_11485;
wire n_1444;
wire n_7300;
wire n_6975;
wire n_14666;
wire n_1263;
wire n_13605;
wire n_17387;
wire n_11048;
wire n_4733;
wire n_14237;
wire n_6729;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_11240;
wire n_13841;
wire n_3080;
wire n_11634;
wire n_12580;
wire n_10013;
wire n_17166;
wire n_2865;
wire n_16119;
wire n_6076;
wire n_8933;
wire n_19344;
wire n_15876;
wire n_18819;
wire n_15231;
wire n_11287;
wire n_943;
wire n_9774;
wire n_4879;
wire n_6390;
wire n_13409;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_9720;
wire n_15727;
wire n_10169;
wire n_12690;
wire n_7563;
wire n_12475;
wire n_1345;
wire n_4556;
wire n_11765;
wire n_8434;
wire n_13405;
wire n_12302;
wire n_10477;
wire n_19510;
wire n_4117;
wire n_14414;
wire n_15565;
wire n_5995;
wire n_17823;
wire n_2378;
wire n_5905;
wire n_9149;
wire n_2655;
wire n_7035;
wire n_6193;
wire n_1467;
wire n_4250;
wire n_16858;
wire n_16980;
wire n_224;
wire n_3963;
wire n_9345;
wire n_11550;
wire n_17315;
wire n_7527;
wire n_13061;
wire n_9682;
wire n_2214;
wire n_17719;
wire n_6582;
wire n_18432;
wire n_12545;
wire n_18320;
wire n_1230;
wire n_3850;
wire n_18078;
wire n_9924;
wire n_14744;
wire n_15091;
wire n_5525;
wire n_17527;
wire n_163;
wire n_1644;
wire n_12753;
wire n_2277;
wire n_7090;
wire n_9254;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_11641;
wire n_7415;
wire n_11211;
wire n_13375;
wire n_13691;
wire n_824;
wire n_6745;
wire n_6972;
wire n_18526;
wire n_16913;
wire n_16663;
wire n_11857;
wire n_395;
wire n_6240;
wire n_13482;
wire n_18069;
wire n_5297;
wire n_15778;
wire n_7121;
wire n_9469;
wire n_15869;
wire n_2961;
wire n_15598;
wire n_15988;
wire n_16593;
wire n_6515;
wire n_483;
wire n_16604;
wire n_2546;
wire n_13873;
wire n_15805;
wire n_476;
wire n_1957;
wire n_17836;
wire n_4732;
wire n_18769;
wire n_11201;
wire n_10531;
wire n_14964;
wire n_8918;
wire n_12878;
wire n_19273;
wire n_8932;
wire n_17756;
wire n_4581;
wire n_16603;
wire n_9249;
wire n_2143;
wire n_8180;
wire n_15580;
wire n_9444;
wire n_10772;
wire n_2031;
wire n_7114;
wire n_4878;
wire n_15984;
wire n_6770;
wire n_17730;
wire n_15151;
wire n_16626;
wire n_5639;
wire n_487;
wire n_8943;
wire n_14767;
wire n_18463;
wire n_4503;
wire n_14773;
wire n_10127;
wire n_13654;
wire n_5361;
wire n_11814;
wire n_12255;
wire n_4199;
wire n_1912;
wire n_9723;
wire n_19446;
wire n_1982;
wire n_3872;
wire n_1312;
wire n_19577;
wire n_5330;
wire n_7199;
wire n_10039;
wire n_10854;
wire n_11358;
wire n_13366;
wire n_247;
wire n_5892;
wire n_7940;
wire n_16467;
wire n_6782;
wire n_18746;
wire n_2008;
wire n_2192;
wire n_328;
wire n_17669;
wire n_1386;
wire n_6503;
wire n_19423;
wire n_12017;
wire n_17357;
wire n_15381;
wire n_18477;
wire n_11958;
wire n_6621;
wire n_15624;
wire n_16103;
wire n_19041;
wire n_16460;
wire n_690;
wire n_8271;
wire n_4800;
wire n_1157;
wire n_12728;
wire n_1752;
wire n_16651;
wire n_4958;
wire n_6783;
wire n_12259;
wire n_8699;
wire n_16305;
wire n_19409;
wire n_2963;
wire n_15861;
wire n_3873;
wire n_8225;
wire n_9536;
wire n_14250;
wire n_16818;
wire n_16573;
wire n_18671;
wire n_16562;
wire n_6296;
wire n_7708;
wire n_11671;
wire n_10328;
wire n_5968;
wire n_2644;
wire n_3326;
wire n_6497;
wire n_15705;
wire n_2411;
wire n_16816;
wire n_7333;
wire n_15376;
wire n_8546;
wire n_10963;
wire n_16358;
wire n_18035;
wire n_7371;
wire n_17547;
wire n_15050;
wire n_8152;
wire n_10826;
wire n_7463;
wire n_8525;
wire n_17767;
wire n_18680;
wire n_283;
wire n_12160;
wire n_590;
wire n_9620;
wire n_1990;
wire n_3805;
wire n_5205;
wire n_17145;
wire n_11119;
wire n_7954;
wire n_1465;
wire n_2622;
wire n_7951;
wire n_8096;
wire n_13901;
wire n_7231;
wire n_5080;
wire n_3128;
wire n_15252;
wire n_18043;
wire n_16238;
wire n_5372;
wire n_14050;
wire n_15763;
wire n_17983;
wire n_2691;
wire n_15317;
wire n_7772;
wire n_2690;
wire n_14197;
wire n_18159;
wire n_19364;
wire n_8996;
wire n_12070;
wire n_9714;
wire n_3078;
wire n_14898;
wire n_15672;
wire n_3793;
wire n_15920;
wire n_11928;
wire n_5071;
wire n_14395;
wire n_5801;
wire n_13528;
wire n_6047;
wire n_8292;
wire n_8601;
wire n_9377;
wire n_11932;
wire n_6970;
wire n_19328;
wire n_1308;
wire n_13027;
wire n_12607;
wire n_7272;
wire n_15782;
wire n_19553;
wire n_12075;
wire n_4540;
wire n_13489;
wire n_2097;
wire n_18887;
wire n_3499;
wire n_13877;
wire n_1005;
wire n_6209;
wire n_11922;
wire n_14020;
wire n_1469;
wire n_12358;
wire n_7408;
wire n_2650;
wire n_10488;
wire n_8969;
wire n_14187;
wire n_11577;
wire n_17840;
wire n_16914;
wire n_18513;
wire n_153;
wire n_3348;
wire n_19165;
wire n_17907;
wire n_11475;
wire n_9048;
wire n_5228;
wire n_10274;
wire n_1723;
wire n_189;
wire n_6694;
wire n_15318;
wire n_9168;
wire n_14220;
wire n_13837;
wire n_2335;
wire n_18570;
wire n_529;
wire n_5507;
wire n_5569;
wire n_15559;
wire n_16871;
wire n_14221;
wire n_13964;
wire n_10832;
wire n_3173;
wire n_18829;
wire n_6856;
wire n_1049;
wire n_6466;
wire n_16039;
wire n_7864;
wire n_18295;
wire n_6727;
wire n_14360;
wire n_10584;
wire n_1717;
wire n_2449;
wire n_3880;
wire n_13601;
wire n_17457;
wire n_17115;
wire n_19281;
wire n_18155;
wire n_4545;
wire n_272;
wire n_6820;
wire n_2896;
wire n_2639;
wire n_17083;
wire n_458;
wire n_5490;
wire n_19007;
wire n_4771;
wire n_13392;
wire n_5836;
wire n_17563;
wire n_9169;
wire n_252;
wire n_5834;
wire n_3191;
wire n_10229;
wire n_5584;
wire n_7512;
wire n_3561;
wire n_19008;
wire n_18401;
wire n_6469;
wire n_6700;
wire n_3032;
wire n_6223;
wire n_11398;
wire n_8798;
wire n_9600;
wire n_2877;
wire n_8085;
wire n_11274;
wire n_1021;
wire n_8123;
wire n_811;
wire n_17997;
wire n_12512;
wire n_9927;
wire n_5497;
wire n_16973;
wire n_15657;
wire n_17571;
wire n_3598;
wire n_7127;
wire n_831;
wire n_15513;
wire n_8666;
wire n_2435;
wire n_12284;
wire n_18322;
wire n_1382;
wire n_7801;
wire n_9155;
wire n_1483;
wire n_10416;
wire n_15837;
wire n_1372;
wire n_14370;
wire n_1719;
wire n_13430;
wire n_7959;
wire n_1427;
wire n_2745;
wire n_14525;
wire n_7735;
wire n_8004;
wire n_6667;
wire n_10583;
wire n_10806;
wire n_2323;
wire n_162;
wire n_5234;
wire n_7546;
wire n_6272;
wire n_14274;
wire n_6588;
wire n_3265;
wire n_3755;
wire n_4042;
wire n_18125;
wire n_15403;
wire n_13081;
wire n_15602;
wire n_12252;
wire n_16743;
wire n_10439;
wire n_12627;
wire n_19378;
wire n_16730;
wire n_15637;
wire n_14272;
wire n_11237;
wire n_2410;
wire n_18868;
wire n_6222;
wire n_15012;
wire n_1783;
wire n_4176;
wire n_14551;
wire n_15720;
wire n_11181;
wire n_13651;
wire n_7521;
wire n_12968;
wire n_10663;
wire n_15517;
wire n_3894;
wire n_13974;
wire n_12277;
wire n_14917;
wire n_3127;
wire n_3623;
wire n_5312;
wire n_16075;
wire n_6625;
wire n_15680;
wire n_2502;
wire n_3646;
wire n_17441;
wire n_14855;
wire n_16757;
wire n_2783;
wire n_8487;
wire n_4034;
wire n_18601;
wire n_1470;
wire n_8141;
wire n_4887;
wire n_14058;
wire n_11020;
wire n_13141;
wire n_16461;
wire n_14065;
wire n_11920;
wire n_17299;
wire n_3862;
wire n_14366;
wire n_10481;
wire n_19250;
wire n_6876;
wire n_16022;
wire n_5049;
wire n_19001;
wire n_19627;
wire n_9573;
wire n_5846;
wire n_7636;
wire n_9799;
wire n_17235;
wire n_5592;
wire n_6954;
wire n_6938;
wire n_1855;
wire n_3051;
wire n_15143;
wire n_11198;
wire n_18932;
wire n_18346;
wire n_18238;
wire n_385;
wire n_1439;
wire n_2859;
wire n_1331;
wire n_3525;
wire n_5157;
wire n_2100;
wire n_11840;
wire n_13157;
wire n_1134;
wire n_10261;
wire n_4003;
wire n_5708;
wire n_3751;
wire n_4894;
wire n_14084;
wire n_4113;
wire n_5649;
wire n_9827;
wire n_13334;
wire n_10907;
wire n_4983;
wire n_14002;
wire n_419;
wire n_7214;
wire n_3907;
wire n_16205;
wire n_13399;
wire n_1254;
wire n_7075;
wire n_19503;
wire n_14697;
wire n_7124;
wire n_13967;
wire n_3291;
wire n_2304;
wire n_7799;
wire n_5698;
wire n_11092;
wire n_14310;
wire n_5084;
wire n_15792;
wire n_15281;
wire n_15675;
wire n_8917;
wire n_15515;
wire n_9647;
wire n_15106;
wire n_4710;
wire n_12067;
wire n_9214;
wire n_17030;
wire n_19537;
wire n_4101;
wire n_7776;
wire n_19621;
wire n_14309;
wire n_9864;
wire n_16256;
wire n_3236;
wire n_17416;
wire n_16741;
wire n_923;
wire n_11770;
wire n_19201;
wire n_13996;
wire n_17944;
wire n_17679;
wire n_9000;
wire n_18442;
wire n_18505;
wire n_10864;
wire n_18412;
wire n_14704;
wire n_8307;
wire n_9383;
wire n_17692;
wire n_4611;
wire n_15258;
wire n_2337;
wire n_12174;
wire n_16322;
wire n_15220;
wire n_6400;
wire n_19611;
wire n_16304;
wire n_18417;
wire n_7543;
wire n_13504;
wire n_16787;
wire n_13169;
wire n_7877;
wire n_9672;
wire n_15291;
wire n_8855;
wire n_18375;
wire n_8885;
wire n_5486;
wire n_15345;
wire n_137;
wire n_1596;
wire n_5092;
wire n_14721;
wire n_1734;
wire n_3172;
wire n_13265;
wire n_4832;
wire n_2902;
wire n_12153;
wire n_7284;
wire n_7264;
wire n_13666;
wire n_19192;
wire n_6537;
wire n_10702;
wire n_13730;
wire n_3536;
wire n_12405;
wire n_2894;
wire n_3710;
wire n_4195;
wire n_10319;
wire n_9654;
wire n_8802;
wire n_9859;
wire n_5240;
wire n_2225;
wire n_6092;
wire n_6241;
wire n_1692;
wire n_8667;
wire n_18996;
wire n_2006;
wire n_3402;
wire n_8121;
wire n_9645;
wire n_7754;
wire n_15549;
wire n_18777;
wire n_2789;
wire n_12792;
wire n_1828;
wire n_19661;
wire n_8320;
wire n_9796;
wire n_18219;
wire n_18231;
wire n_4862;
wire n_15889;
wire n_2376;
wire n_11830;
wire n_12438;
wire n_16173;
wire n_16665;
wire n_8766;
wire n_9165;
wire n_2700;
wire n_19555;
wire n_1041;
wire n_12539;
wire n_565;
wire n_5965;
wire n_9596;
wire n_13652;
wire n_13703;
wire n_18461;
wire n_14369;
wire n_1062;
wire n_7240;
wire n_15354;
wire n_10476;
wire n_9966;
wire n_16794;
wire n_1222;
wire n_2635;
wire n_11486;
wire n_15999;
wire n_15280;
wire n_12677;
wire n_4321;
wire n_7237;
wire n_17867;
wire n_16456;
wire n_6877;
wire n_12873;
wire n_16364;
wire n_6949;
wire n_19356;
wire n_17036;
wire n_806;
wire n_13401;
wire n_584;
wire n_12276;
wire n_9893;
wire n_14122;
wire n_17565;
wire n_8126;
wire n_15819;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4757;
wire n_15603;
wire n_12352;
wire n_17267;
wire n_2809;
wire n_18528;
wire n_787;
wire n_10099;
wire n_9961;
wire n_16833;
wire n_14895;
wire n_7163;
wire n_1528;
wire n_1146;
wire n_16582;
wire n_18028;
wire n_2021;
wire n_15270;
wire n_17964;
wire n_10181;
wire n_15670;
wire n_4604;
wire n_5724;
wire n_7201;
wire n_3157;
wire n_16825;
wire n_2422;
wire n_10949;
wire n_3457;
wire n_3762;
wire n_18197;
wire n_3411;
wire n_4519;
wire n_5355;
wire n_13969;
wire n_16548;
wire n_5186;
wire n_1498;
wire n_12693;
wire n_6792;
wire n_1210;
wire n_9316;
wire n_5438;
wire n_13259;
wire n_1269;
wire n_19164;
wire n_14954;
wire n_12648;
wire n_655;
wire n_4726;
wire n_6045;
wire n_1872;
wire n_9914;
wire n_8132;
wire n_19541;
wire n_10917;
wire n_16050;
wire n_3761;
wire n_18006;
wire n_7821;
wire n_12407;
wire n_11284;
wire n_14668;
wire n_14776;
wire n_10458;
wire n_2041;
wire n_11656;
wire n_13134;
wire n_10271;
wire n_15415;
wire n_16808;
wire n_18902;
wire n_1098;
wire n_5746;
wire n_6673;
wire n_18207;
wire n_11909;
wire n_12637;
wire n_7887;
wire n_398;
wire n_6060;
wire n_15414;
wire n_15783;
wire n_3726;
wire n_12009;
wire n_2369;
wire n_13612;
wire n_19388;
wire n_10648;
wire n_2587;
wire n_7550;
wire n_17498;
wire n_15077;
wire n_3199;
wire n_12414;
wire n_9760;
wire n_10690;
wire n_15733;
wire n_15864;
wire n_14207;
wire n_1953;
wire n_19080;
wire n_13863;
wire n_14305;
wire n_9863;
wire n_15330;
wire n_10500;
wire n_5432;
wire n_15261;
wire n_11929;
wire n_11075;
wire n_7851;
wire n_16605;
wire n_9791;
wire n_19228;
wire n_5453;
wire n_4900;
wire n_11177;
wire n_13667;
wire n_18056;
wire n_5842;
wire n_13126;
wire n_7798;
wire n_5253;
wire n_10857;
wire n_18491;
wire n_11310;
wire n_13275;
wire n_11165;
wire n_14411;
wire n_12823;
wire n_2953;
wire n_15412;
wire n_4295;
wire n_5943;
wire n_12193;
wire n_2500;
wire n_1729;
wire n_6088;
wire n_5777;
wire n_15257;
wire n_8528;
wire n_8204;
wire n_11733;
wire n_15646;
wire n_1389;
wire n_18214;
wire n_7100;
wire n_3583;
wire n_3860;
wire n_18347;
wire n_14738;
wire n_12242;
wire n_5610;
wire n_3015;
wire n_13796;
wire n_10502;
wire n_15522;
wire n_17577;
wire n_17874;
wire n_6722;
wire n_17892;
wire n_7622;
wire n_11123;
wire n_8512;
wire n_14464;
wire n_387;
wire n_744;
wire n_971;
wire n_8635;
wire n_3241;
wire n_2906;
wire n_4342;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_1205;
wire n_15535;
wire n_16633;
wire n_7831;
wire n_10227;
wire n_10574;
wire n_19271;
wire n_2180;
wire n_16323;
wire n_2858;
wire n_18624;
wire n_6201;
wire n_12218;
wire n_5737;
wire n_3604;
wire n_12343;
wire n_4373;
wire n_8919;
wire n_17014;
wire n_12316;
wire n_14937;
wire n_14454;
wire n_4711;
wire n_11478;
wire n_16067;
wire n_3068;
wire n_15650;
wire n_12236;
wire n_12902;
wire n_16230;
wire n_7784;
wire n_9272;
wire n_5768;
wire n_13038;
wire n_2465;
wire n_12892;
wire n_17768;
wire n_3811;
wire n_11294;
wire n_910;
wire n_15667;
wire n_3486;
wire n_4086;
wire n_10289;
wire n_6565;
wire n_6942;
wire n_11819;
wire n_19389;
wire n_2032;
wire n_4812;
wire n_13420;
wire n_6862;
wire n_5858;
wire n_17200;
wire n_15053;
wire n_13005;
wire n_708;
wire n_14805;
wire n_6037;
wire n_2312;
wire n_11844;
wire n_1266;
wire n_15390;
wire n_6635;
wire n_185;
wire n_13184;
wire n_1276;
wire n_13535;
wire n_14982;
wire n_12247;
wire n_14770;
wire n_11100;
wire n_298;
wire n_1582;
wire n_5588;
wire n_3286;
wire n_19350;
wire n_7167;
wire n_6480;
wire n_15105;
wire n_5075;
wire n_3682;
wire n_18927;
wire n_3771;
wire n_18383;
wire n_12765;
wire n_7865;
wire n_15690;
wire n_9289;
wire n_11315;
wire n_6561;
wire n_12706;
wire n_11153;
wire n_17128;
wire n_859;
wire n_406;
wire n_6875;
wire n_10934;
wire n_1770;
wire n_10197;
wire n_18999;
wire n_3285;
wire n_19584;
wire n_11949;
wire n_8402;
wire n_9690;
wire n_2071;
wire n_11746;
wire n_9371;
wire n_16837;
wire n_7267;
wire n_4599;
wire n_12315;
wire n_18668;
wire n_5222;
wire n_7850;
wire n_14100;
wire n_12998;
wire n_7812;
wire n_13143;
wire n_9080;
wire n_14549;
wire n_8133;
wire n_6176;
wire n_14717;
wire n_3881;
wire n_16426;
wire n_14459;
wire n_4508;
wire n_11530;
wire n_13411;
wire n_7056;
wire n_8193;
wire n_12445;
wire n_12856;
wire n_19520;
wire n_7813;
wire n_7514;
wire n_7649;
wire n_18734;
wire n_12525;
wire n_16116;
wire n_1039;
wire n_6078;
wire n_2043;
wire n_1480;
wire n_15823;
wire n_5832;
wire n_13758;
wire n_1305;
wire n_7688;
wire n_4562;
wire n_16820;
wire n_3383;
wire n_8707;
wire n_12357;
wire n_9208;
wire n_11791;
wire n_19525;
wire n_7611;
wire n_17218;
wire n_15216;
wire n_11848;
wire n_3610;
wire n_11632;
wire n_15352;
wire n_7795;
wire n_12180;
wire n_2065;
wire n_15608;
wire n_10935;
wire n_2001;
wire n_7723;
wire n_11621;
wire n_19448;
wire n_225;
wire n_16171;
wire n_3555;
wire n_11667;
wire n_7450;
wire n_17311;
wire n_7362;
wire n_17455;
wire n_12208;
wire n_1131;
wire n_3110;
wire n_14565;
wire n_17248;
wire n_11298;
wire n_15796;
wire n_1888;
wire n_8993;
wire n_6204;
wire n_13314;
wire n_670;
wire n_11741;
wire n_3908;
wire n_15537;
wire n_3467;
wire n_12773;
wire n_9044;
wire n_12381;
wire n_19302;
wire n_18174;
wire n_14883;
wire n_17024;
wire n_6451;
wire n_9813;
wire n_1226;
wire n_3740;
wire n_18482;
wire n_3186;
wire n_640;
wire n_17322;
wire n_9244;
wire n_15304;
wire n_7049;
wire n_15271;
wire n_2632;
wire n_14865;
wire n_8278;
wire n_11644;
wire n_6345;
wire n_15893;
wire n_9094;
wire n_15432;
wire n_13108;
wire n_364;
wire n_5782;
wire n_5041;
wire n_13170;
wire n_1915;
wire n_4275;
wire n_14471;
wire n_11357;
wire n_19387;
wire n_4425;
wire n_9985;
wire n_4449;
wire n_12089;
wire n_7057;
wire n_17888;
wire n_11959;
wire n_19586;
wire n_1612;
wire n_4809;
wire n_12987;
wire n_8529;
wire n_625;
wire n_10254;
wire n_18625;
wire n_14715;
wire n_15970;
wire n_11208;
wire n_15978;
wire n_12452;
wire n_15961;
wire n_8574;
wire n_1038;
wire n_12292;
wire n_4241;
wire n_12818;
wire n_11420;
wire n_12500;
wire n_8044;
wire n_16330;
wire n_9439;
wire n_1380;
wire n_15239;
wire n_2557;
wire n_11630;
wire n_2405;
wire n_15444;
wire n_15289;
wire n_13172;
wire n_2336;
wire n_16234;
wire n_2521;
wire n_9120;
wire n_17335;
wire n_17610;
wire n_19522;
wire n_424;
wire n_12168;
wire n_16496;
wire n_8903;
wire n_141;
wire n_1985;
wire n_16057;
wire n_16401;
wire n_4531;
wire n_3282;
wire n_15781;
wire n_14448;
wire n_1532;
wire n_11017;
wire n_7247;
wire n_14622;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_3031;
wire n_14739;
wire n_16649;
wire n_12613;
wire n_14365;
wire n_9325;
wire n_16448;
wire n_4555;
wire n_17173;
wire n_9384;
wire n_6216;
wire n_7340;
wire n_12695;
wire n_15467;
wire n_4308;
wire n_14219;
wire n_3463;
wire n_11576;
wire n_1954;
wire n_2729;
wire n_2582;
wire n_1798;
wire n_3998;
wire n_12006;
wire n_2495;
wire n_10128;
wire n_371;
wire n_18319;
wire n_12246;
wire n_18220;
wire n_9955;
wire n_19477;
wire n_3829;
wire n_9007;
wire n_10143;
wire n_1471;
wire n_18715;
wire n_3655;
wire n_17884;
wire n_3825;
wire n_2880;
wire n_13085;
wire n_19260;
wire n_7780;
wire n_8452;
wire n_11518;
wire n_5670;
wire n_8557;
wire n_10303;
wire n_16189;
wire n_15097;
wire n_18892;
wire n_11252;
wire n_8012;
wire n_1445;
wire n_1526;
wire n_17055;
wire n_1978;
wire n_6472;
wire n_18067;
wire n_574;
wire n_8114;
wire n_4202;
wire n_16227;
wire n_5879;
wire n_14563;
wire n_4403;
wire n_5238;
wire n_16329;
wire n_11256;
wire n_6166;
wire n_12370;
wire n_9136;
wire n_12860;
wire n_16278;
wire n_473;
wire n_17404;
wire n_559;
wire n_19635;
wire n_7063;
wire n_14768;
wire n_4139;
wire n_13885;
wire n_1986;
wire n_13631;
wire n_18103;
wire n_6081;
wire n_16746;
wire n_15929;
wire n_6724;
wire n_813;
wire n_11336;
wire n_12758;
wire n_17410;
wire n_19248;
wire n_11849;
wire n_3910;
wire n_9204;
wire n_12142;
wire n_9476;
wire n_9689;
wire n_16711;
wire n_10659;
wire n_7585;
wire n_4948;
wire n_5268;
wire n_6946;
wire n_3319;
wire n_12983;
wire n_3748;
wire n_6424;
wire n_11210;
wire n_7599;
wire n_16271;
wire n_15541;
wire n_13980;
wire n_16366;
wire n_982;
wire n_11191;
wire n_10547;
wire n_6778;
wire n_17359;
wire n_13205;
wire n_1697;
wire n_979;
wire n_5544;
wire n_5067;
wire n_15283;
wire n_12396;
wire n_15407;
wire n_7614;
wire n_19381;
wire n_1278;
wire n_7839;
wire n_9837;
wire n_634;
wire n_10896;
wire n_136;
wire n_17761;
wire n_4130;
wire n_10562;
wire n_16042;
wire n_5941;
wire n_2009;
wire n_14417;
wire n_3601;
wire n_6340;
wire n_10054;
wire n_10355;
wire n_1289;
wire n_16893;
wire n_3055;
wire n_6706;
wire n_3966;
wire n_13034;
wire n_1014;
wire n_16828;
wire n_10007;
wire n_882;
wire n_11751;
wire n_17550;
wire n_3746;
wire n_17185;
wire n_14637;
wire n_11495;
wire n_4478;
wire n_1662;
wire n_17015;
wire n_7372;
wire n_19617;
wire n_2818;
wire n_17980;
wire n_674;
wire n_3921;
wire n_17535;
wire n_16822;
wire n_10704;
wire n_11520;
wire n_1927;
wire n_19614;
wire n_12169;
wire n_16788;
wire n_15088;
wire n_17976;
wire n_702;
wire n_4965;
wire n_16383;
wire n_17538;
wire n_11012;
wire n_6111;
wire n_11502;
wire n_15348;
wire n_11631;
wire n_13588;
wire n_13570;
wire n_2193;
wire n_4523;
wire n_6011;
wire n_11842;
wire n_14710;
wire n_3153;
wire n_877;
wire n_13737;
wire n_16590;
wire n_728;
wire n_18188;
wire n_4607;
wire n_16640;
wire n_11389;
wire n_7226;
wire n_9013;
wire n_18373;
wire n_4041;
wire n_9634;
wire n_17846;
wire n_5876;
wire n_10916;
wire n_8584;
wire n_11557;
wire n_17113;
wire n_16748;
wire n_15363;
wire n_7810;
wire n_14955;
wire n_9364;
wire n_8228;
wire n_1825;
wire n_16015;
wire n_170;
wire n_15642;
wire n_1412;
wire n_10929;
wire n_18854;
wire n_19372;
wire n_13862;
wire n_8100;
wire n_13446;
wire n_13086;
wire n_8091;
wire n_17155;
wire n_148;
wire n_4675;
wire n_5837;
wire n_5491;
wire n_2987;
wire n_5496;
wire n_5802;
wire n_14965;
wire n_13887;
wire n_12787;
wire n_12799;
wire n_4002;
wire n_5178;
wire n_9317;
wire n_12657;
wire n_9769;
wire n_15205;
wire n_8158;
wire n_1295;
wire n_8469;
wire n_18718;
wire n_18481;
wire n_10102;
wire n_5983;
wire n_3146;
wire n_1438;
wire n_3953;
wire n_11825;
wire n_1100;
wire n_14354;
wire n_7684;
wire n_15532;
wire n_5604;
wire n_673;
wire n_16083;
wire n_10589;
wire n_11611;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_865;
wire n_4191;
wire n_18221;
wire n_12408;
wire n_16287;
wire n_16169;
wire n_19314;
wire n_17556;
wire n_2341;
wire n_10110;
wire n_11230;
wire n_11688;
wire n_4350;
wire n_12715;
wire n_12434;
wire n_11709;
wire n_14328;
wire n_6095;
wire n_17049;
wire n_18938;
wire n_16540;
wire n_14429;
wire n_12979;
wire n_16901;
wire n_6559;
wire n_3924;
wire n_15799;
wire n_17195;
wire n_19050;
wire n_4621;
wire n_510;
wire n_1488;
wire n_2148;
wire n_5565;
wire n_14270;
wire n_15238;
wire n_2339;
wire n_10190;
wire n_19656;
wire n_5984;
wire n_6287;
wire n_13614;
wire n_17703;
wire n_8347;
wire n_19440;
wire n_1776;
wire n_1766;
wire n_14208;
wire n_9330;
wire n_4021;
wire n_3014;
wire n_15693;
wire n_12029;
wire n_4103;
wire n_9523;
wire n_14584;
wire n_4022;
wire n_19636;
wire n_10060;
wire n_18192;
wire n_9686;
wire n_4481;
wire n_17130;
wire n_19375;
wire n_1304;
wire n_10162;
wire n_4669;
wire n_15002;
wire n_9964;
wire n_17515;
wire n_13842;
wire n_7510;
wire n_6662;
wire n_11291;
wire n_13107;
wire n_5603;
wire n_9154;
wire n_14501;
wire n_3312;
wire n_7109;
wire n_2936;
wire n_3224;
wire n_14790;
wire n_8822;
wire n_1087;
wire n_17204;
wire n_12187;
wire n_657;
wire n_19662;
wire n_18772;
wire n_1505;
wire n_7253;
wire n_3129;
wire n_17201;
wire n_8476;
wire n_17745;
wire n_11927;
wire n_16674;
wire n_16326;
wire n_16571;
wire n_8359;
wire n_4484;
wire n_15808;
wire n_16497;
wire n_16752;
wire n_14574;
wire n_526;
wire n_14451;
wire n_2251;
wire n_9455;
wire n_8708;
wire n_14092;
wire n_2837;
wire n_4883;
wire n_14509;
wire n_11882;
wire n_17649;
wire n_11647;
wire n_15027;
wire n_15404;
wire n_10706;
wire n_3341;
wire n_19129;
wire n_8872;
wire n_3559;
wire n_8238;
wire n_15465;
wire n_11222;
wire n_9200;
wire n_16279;
wire n_5146;
wire n_3056;
wire n_745;
wire n_15858;
wire n_3447;
wire n_3971;
wire n_716;
wire n_1774;
wire n_18946;
wire n_2589;
wire n_4535;
wire n_14765;
wire n_7704;
wire n_18893;
wire n_16170;
wire n_14995;
wire n_6302;
wire n_2442;
wire n_17479;
wire n_7203;
wire n_11259;
wire n_7670;
wire n_18258;
wire n_16010;
wire n_14434;
wire n_9673;
wire n_2545;
wire n_8642;
wire n_11875;
wire n_18567;
wire n_12111;
wire n_8912;
wire n_19067;
wire n_1314;
wire n_864;
wire n_14275;
wire n_19309;
wire n_12903;
wire n_6343;
wire n_12593;
wire n_5270;
wire n_1534;
wire n_17849;
wire n_11602;
wire n_15689;
wire n_12413;
wire n_17474;
wire n_723;
wire n_13813;
wire n_16190;
wire n_18315;
wire n_8111;
wire n_10432;
wire n_19227;
wire n_16888;
wire n_18376;
wire n_8056;
wire n_3287;
wire n_9674;
wire n_2357;
wire n_6433;
wire n_18253;
wire n_15469;
wire n_17140;
wire n_18407;
wire n_1681;
wire n_520;
wire n_18816;
wire n_4020;
wire n_13636;
wire n_19332;
wire n_19456;
wire n_5220;
wire n_18920;
wire n_11341;
wire n_10787;
wire n_13256;
wire n_14567;
wire n_6870;
wire n_6221;
wire n_16308;
wire n_6279;
wire n_13905;
wire n_12290;
wire n_7881;
wire n_9369;
wire n_18896;
wire n_16986;
wire n_17872;
wire n_6071;
wire n_9583;
wire n_19422;
wire n_15119;
wire n_19117;
wire n_12150;
wire n_1617;
wire n_3370;
wire n_335;
wire n_15256;
wire n_18366;
wire n_8090;
wire n_8053;
wire n_10184;
wire n_15982;
wire n_274;
wire n_19643;
wire n_18647;
wire n_15452;
wire n_1267;
wire n_1806;
wire n_13615;
wire n_15625;
wire n_2023;
wire n_12633;
wire n_14779;
wire n_496;
wire n_15114;
wire n_4614;
wire n_3360;
wire n_10277;
wire n_17934;
wire n_3956;
wire n_8163;
wire n_16632;
wire n_16028;
wire n_10948;
wire n_10525;
wire n_14287;
wire n_9507;
wire n_11528;
wire n_15296;
wire n_15828;
wire n_18107;
wire n_19211;
wire n_3870;
wire n_16126;
wire n_18102;
wire n_18545;
wire n_16168;
wire n_15915;
wire n_793;
wire n_10049;
wire n_3749;
wire n_15551;
wire n_9457;
wire n_5780;
wire n_5037;
wire n_16738;
wire n_316;
wire n_6084;
wire n_11039;
wire n_14342;
wire n_2555;
wire n_13693;
wire n_18992;
wire n_12606;
wire n_10900;
wire n_2201;
wire n_14107;
wire n_14781;
wire n_13333;
wire n_13229;
wire n_994;
wire n_17336;
wire n_11380;
wire n_15737;
wire n_19567;
wire n_10792;
wire n_15573;
wire n_13296;
wire n_14611;
wire n_3448;
wire n_17863;
wire n_1036;
wire n_1661;
wire n_5360;
wire n_17088;
wire n_19100;
wire n_15051;
wire n_6548;
wire n_3926;
wire n_6993;
wire n_1095;
wire n_15916;
wire n_4405;
wire n_16468;
wire n_10241;
wire n_19598;
wire n_15639;
wire n_3670;
wire n_179;
wire n_4667;
wire n_8702;
wire n_17158;
wire n_8116;
wire n_1115;
wire n_8195;
wire n_7946;
wire n_14069;
wire n_18452;
wire n_1409;
wire n_9991;
wire n_11366;
wire n_11872;
wire n_10823;
wire n_14766;
wire n_11106;
wire n_1126;
wire n_14592;
wire n_15109;
wire n_11132;
wire n_17625;
wire n_18546;
wire n_18034;
wire n_3635;
wire n_18181;
wire n_17126;
wire n_10824;
wire n_4155;
wire n_19566;
wire n_16216;
wire n_19398;
wire n_14277;
wire n_19565;
wire n_13493;
wire n_16389;
wire n_9047;
wire n_12842;
wire n_18569;
wire n_12481;
wire n_18168;
wire n_11316;
wire n_9599;
wire n_11559;
wire n_9072;
wire n_4929;
wire n_9428;
wire n_10340;
wire n_17463;
wire n_15817;
wire n_15344;
wire n_2220;
wire n_2577;
wire n_13669;
wire n_17245;
wire n_3529;
wire n_17179;
wire n_11109;
wire n_13840;
wire n_16601;
wire n_11591;
wire n_14251;
wire n_11225;
wire n_6765;
wire n_4565;
wire n_4159;
wire n_8883;
wire n_10634;
wire n_4586;
wire n_11058;
wire n_15888;
wire n_1608;
wire n_7336;
wire n_11471;
wire n_7446;
wire n_3628;
wire n_14679;
wire n_10961;
wire n_7357;
wire n_1491;
wire n_17064;
wire n_8737;
wire n_13925;
wire n_18334;
wire n_10379;
wire n_16704;
wire n_2586;
wire n_18223;
wire n_13368;
wire n_14507;
wire n_9484;
wire n_10989;
wire n_17725;
wire n_10939;
wire n_19557;
wire n_1046;
wire n_2560;
wire n_1145;
wire n_11144;
wire n_14857;
wire n_6406;
wire n_14034;
wire n_10962;
wire n_11128;
wire n_15677;
wire n_10721;
wire n_8593;
wire n_11025;
wire n_12007;
wire n_5062;
wire n_15901;
wire n_321;
wire n_13481;
wire n_12018;
wire n_3588;
wire n_18040;
wire n_17393;
wire n_14457;
wire n_16931;
wire n_12872;
wire n_18189;
wire n_6492;
wire n_14517;
wire n_2288;
wire n_11460;
wire n_13713;
wire n_12372;
wire n_13608;
wire n_7046;
wire n_19059;
wire n_10956;
wire n_2642;
wire n_7468;
wire n_2383;
wire n_18785;
wire n_14934;
wire n_19663;
wire n_2351;
wire n_18844;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_2986;
wire n_17870;
wire n_139;
wire n_15652;
wire n_3489;
wire n_19466;
wire n_16713;
wire n_14578;
wire n_15653;
wire n_5914;
wire n_12955;
wire n_9321;
wire n_16856;
wire n_18555;
wire n_1282;
wire n_15016;
wire n_2567;
wire n_18493;
wire n_275;
wire n_3377;
wire n_9161;
wire n_2869;
wire n_7836;
wire n_10737;
wire n_17910;
wire n_17750;
wire n_346;
wire n_15865;
wire n_13448;
wire n_16928;
wire n_5813;
wire n_13767;
wire n_790;
wire n_2901;
wire n_2611;
wire n_11055;
wire n_4358;
wire n_16616;
wire n_14832;
wire n_10982;
wire n_5805;
wire n_5616;
wire n_17599;
wire n_14571;
wire n_6631;
wire n_12369;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_8927;
wire n_17985;
wire n_16396;
wire n_17531;
wire n_15155;
wire n_12686;
wire n_6228;
wire n_19336;
wire n_5416;
wire n_14881;
wire n_18588;
wire n_14527;
wire n_12822;
wire n_13307;
wire n_7279;
wire n_17460;
wire n_13312;
wire n_11761;
wire n_9984;
wire n_8474;
wire n_3524;
wire n_489;
wire n_2885;
wire n_10600;
wire n_6102;
wire n_636;
wire n_10833;
wire n_18329;
wire n_18649;
wire n_13023;
wire n_19343;
wire n_1607;
wire n_1454;
wire n_15315;
wire n_19210;
wire n_11185;
wire n_13440;
wire n_869;
wire n_1154;
wire n_13436;
wire n_19615;
wire n_19133;
wire n_16982;
wire n_846;
wire n_841;
wire n_508;
wire n_11081;
wire n_16687;
wire n_1562;
wire n_14858;
wire n_8787;
wire n_13911;
wire n_5051;
wire n_17544;
wire n_5587;
wire n_10941;
wire n_14617;
wire n_9816;
wire n_17132;
wire n_14263;
wire n_661;
wire n_8605;
wire n_10358;
wire n_3565;
wire n_17593;
wire n_9944;
wire n_6998;
wire n_16158;
wire n_4173;
wire n_12338;
wire n_7615;
wire n_5651;
wire n_9605;
wire n_1217;
wire n_7591;
wire n_11404;
wire n_16488;
wire n_15994;
wire n_15685;
wire n_9788;
wire n_16273;
wire n_10785;
wire n_18262;
wire n_13872;
wire n_17646;
wire n_12341;
wire n_18389;
wire n_5412;
wire n_14475;
wire n_10815;
wire n_1120;
wire n_555;
wire n_8784;
wire n_7382;
wire n_2048;
wire n_13955;
wire n_176;
wire n_17708;
wire n_14400;
wire n_4857;
wire n_16725;
wire n_16904;
wire n_16432;
wire n_12085;
wire n_2883;
wire n_18190;
wire n_13554;
wire n_18421;
wire n_863;
wire n_6780;
wire n_11582;
wire n_3268;
wire n_1147;
wire n_1754;
wire n_11705;
wire n_3701;
wire n_7673;
wire n_1812;
wire n_6830;
wire n_17391;
wire n_17682;
wire n_7282;
wire n_9968;
wire n_11474;
wire n_10657;
wire n_13595;
wire n_5997;
wire n_2492;
wire n_10687;
wire n_13283;
wire n_19543;
wire n_15615;
wire n_12110;
wire n_8363;
wire n_5119;
wire n_19445;
wire n_17802;
wire n_9669;
wire n_17775;
wire n_6510;
wire n_8282;
wire n_5938;
wire n_15972;
wire n_6237;
wire n_12040;
wire n_11752;
wire n_12216;
wire n_17446;
wire n_2117;
wire n_18573;
wire n_14975;
wire n_7581;
wire n_6360;
wire n_17960;
wire n_15217;
wire n_4858;
wire n_13308;
wire n_19049;
wire n_9952;
wire n_15323;
wire n_12183;
wire n_10668;
wire n_9256;
wire n_5750;
wire n_4823;
wire n_4309;
wire n_839;
wire n_14007;
wire n_7346;
wire n_1537;
wire n_13373;
wire n_4243;
wire n_7428;
wire n_12221;
wire n_5666;
wire n_9195;
wire n_16236;
wire n_17787;
wire n_7283;
wire n_4142;
wire n_6314;
wire n_10632;
wire n_18861;
wire n_9623;
wire n_3796;
wire n_6964;
wire n_3408;
wire n_19027;
wire n_19561;
wire n_1184;
wire n_18912;
wire n_19322;
wire n_16702;
wire n_1525;
wire n_2594;
wire n_11329;
wire n_6495;
wire n_5994;
wire n_17280;
wire n_9516;
wire n_4244;
wire n_2147;
wire n_13241;
wire n_16027;
wire n_2503;
wire n_8976;
wire n_17844;
wire n_18136;
wire n_10130;
wire n_11661;
wire n_9222;
wire n_8435;
wire n_8882;
wire n_16391;
wire n_4787;
wire n_15949;
wire n_10622;
wire n_5633;
wire n_5664;
wire n_6797;
wire n_15673;
wire n_14012;
wire n_8759;
wire n_16941;
wire n_7177;
wire n_357;
wire n_13066;
wire n_13665;
wire n_12993;
wire n_19604;
wire n_11314;
wire n_17784;
wire n_2681;
wire n_15678;
wire n_8235;
wire n_13083;
wire n_3764;
wire n_19093;
wire n_16164;
wire n_6152;
wire n_16444;
wire n_4075;
wire n_9820;
wire n_14071;
wire n_12749;
wire n_2303;
wire n_1619;
wire n_8448;
wire n_4538;
wire n_12066;
wire n_6513;
wire n_2367;
wire n_1034;
wire n_15908;
wire n_754;
wire n_11184;
wire n_11945;
wire n_11368;
wire n_6330;
wire n_17842;
wire n_19628;
wire n_8457;
wire n_19200;
wire n_18605;
wire n_18837;
wire n_9339;
wire n_14312;
wire n_9601;
wire n_15045;
wire n_11409;
wire n_18995;
wire n_2107;
wire n_2040;
wire n_18737;
wire n_12437;
wire n_5624;
wire n_10840;
wire n_6263;
wire n_10515;
wire n_15501;
wire n_6490;
wire n_15751;
wire n_11605;
wire n_1861;
wire n_10242;
wire n_10144;
wire n_9684;
wire n_15741;
wire n_16195;
wire n_14793;
wire n_18754;
wire n_13472;
wire n_2162;
wire n_15596;
wire n_207;
wire n_4763;
wire n_3587;
wire n_205;
wire n_18316;
wire n_6038;
wire n_15379;
wire n_16272;
wire n_14884;
wire n_3162;
wire n_8964;
wire n_16629;
wire n_1899;
wire n_9814;
wire n_4804;
wire n_5619;
wire n_5859;
wire n_14423;
wire n_16280;
wire n_16414;
wire n_4500;
wire n_13443;
wire n_4433;
wire n_5644;
wire n_2813;
wire n_14626;
wire n_2027;
wire n_2091;
wire n_8960;
wire n_5030;
wire n_15402;
wire n_4194;
wire n_18026;
wire n_8443;
wire n_7715;
wire n_2419;
wire n_8683;
wire n_18558;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_3182;
wire n_5756;
wire n_15306;
wire n_15981;
wire n_16367;

CKINVDCx5p33_ASAP7_75t_R g136 ( 
.A(n_78),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_60),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_44),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_70),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_0),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g146 ( 
.A(n_58),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_72),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_31),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_63),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_86),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_28),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_6),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_42),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_23),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_48),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_55),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_24),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_134),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_54),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_38),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_27),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_35),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_47),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_5),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_53),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_43),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_33),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_92),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_127),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_9),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_12),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_80),
.Y(n_180)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_122),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_111),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_57),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_81),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_56),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_4),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_19),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_101),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_71),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_51),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_93),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_36),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_82),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_41),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_67),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_95),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_100),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_116),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_132),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_124),
.Y(n_204)
);

BUFx8_ASAP7_75t_SL g205 ( 
.A(n_46),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_32),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_94),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_133),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_117),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_109),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_34),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_61),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_112),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_39),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_7),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_29),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_22),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_65),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_115),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_108),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_18),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_77),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_103),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_21),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_17),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_0),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_106),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_120),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_83),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_8),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_87),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_119),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_64),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_30),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

BUFx2_ASAP7_75t_SL g236 ( 
.A(n_131),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_128),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_84),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_98),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_79),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_37),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_14),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_97),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_11),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_129),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_130),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_110),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_52),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_15),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_91),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_13),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_74),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_121),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_25),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_123),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_75),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_66),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_126),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_3),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_113),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_40),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_85),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_45),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_69),
.Y(n_266)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_59),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_90),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_20),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_205),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_136),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_137),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_226),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_186),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_139),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_138),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_142),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_150),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_143),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_140),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_141),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_151),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_144),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_209),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_152),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_154),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_163),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_161),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_149),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_153),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_155),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_167),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_148),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_143),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_168),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_156),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_157),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_169),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_159),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_164),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_170),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_162),
.Y(n_303)
);

HB1xp67_ASAP7_75t_L g304 ( 
.A(n_171),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_166),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_174),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_178),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_173),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_176),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_165),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_267),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_179),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_278),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_271),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_279),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_177),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_276),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_281),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_282),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_287),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_288),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_293),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_290),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_294),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_291),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_292),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_285),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_297),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_300),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_296),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_303),
.Y(n_339)
);

BUFx6f_ASAP7_75t_SL g340 ( 
.A(n_273),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_305),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_302),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_308),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_289),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_301),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_216),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_309),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_274),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_275),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_270),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_280),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_295),
.B(n_181),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_271),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_277),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_310),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_321),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_353),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_313),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_240),
.Y(n_364)
);

CKINVDCx8_ASAP7_75t_R g365 ( 
.A(n_345),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_325),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_190),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_172),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_330),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_315),
.B(n_207),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_343),
.Y(n_378)
);

AOI22x1_ASAP7_75t_SL g379 ( 
.A1(n_355),
.A2(n_251),
.B1(n_220),
.B2(n_180),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_316),
.B(n_187),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_333),
.B(n_160),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_359),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_352),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_326),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_357),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_354),
.A2(n_199),
.B1(n_200),
.B2(n_213),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g388 ( 
.A1(n_344),
.A2(n_192),
.B(n_175),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_349),
.A2(n_219),
.B(n_257),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_348),
.A2(n_214),
.B1(n_215),
.B2(n_232),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_346),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_360),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_346),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_339),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_340),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_318),
.B(n_239),
.Y(n_397)
);

AND2x4_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_351),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_320),
.B(n_182),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

CKINVDCx6p67_ASAP7_75t_R g401 ( 
.A(n_341),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_329),
.B(n_244),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_331),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_342),
.Y(n_405)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_332),
.B(n_184),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_334),
.B(n_185),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_336),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_356),
.B(n_256),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_319),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_353),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_353),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_269),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_315),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_319),
.B(n_183),
.Y(n_416)
);

INVx4_ASAP7_75t_L g417 ( 
.A(n_315),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_315),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_321),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_353),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_319),
.A2(n_255),
.B1(n_266),
.B2(n_254),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_353),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

INVx6_ASAP7_75t_L g424 ( 
.A(n_321),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_321),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_319),
.A2(n_224),
.B1(n_250),
.B2(n_264),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_357),
.A2(n_249),
.B(n_265),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_356),
.B(n_222),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_330),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_353),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_319),
.A2(n_236),
.B1(n_263),
.B2(n_211),
.Y(n_431)
);

INVx5_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_356),
.B(n_246),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_353),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_353),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_319),
.A2(n_218),
.B1(n_248),
.B2(n_261),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g438 ( 
.A(n_333),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_321),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_353),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_319),
.A2(n_217),
.B1(n_241),
.B2(n_260),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g442 ( 
.A1(n_357),
.A2(n_235),
.B(n_262),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_353),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_319),
.A2(n_231),
.B1(n_259),
.B2(n_230),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_353),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_356),
.B(n_197),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g447 ( 
.A(n_321),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_321),
.Y(n_448)
);

AND2x6_ASAP7_75t_L g449 ( 
.A(n_352),
.B(n_245),
.Y(n_449)
);

OR2x6_ASAP7_75t_L g450 ( 
.A(n_321),
.B(n_206),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_353),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_356),
.B(n_198),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_319),
.B(n_191),
.Y(n_453)
);

OA21x2_ASAP7_75t_L g454 ( 
.A1(n_357),
.A2(n_201),
.B(n_258),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_319),
.B(n_210),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_347),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_321),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_353),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_319),
.B(n_195),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_353),
.Y(n_460)
);

AND2x2_ASAP7_75t_SL g461 ( 
.A(n_333),
.B(n_208),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_356),
.B(n_212),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_319),
.B(n_229),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_353),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_315),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_353),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_353),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_353),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_353),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_330),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_356),
.B(n_204),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_353),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_353),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_353),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_321),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_319),
.B(n_225),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_315),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_330),
.A2(n_189),
.B1(n_227),
.B2(n_221),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_315),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_353),
.Y(n_480)
);

OA21x2_ASAP7_75t_L g481 ( 
.A1(n_357),
.A2(n_234),
.B(n_233),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_321),
.B(n_196),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_321),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_353),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_330),
.A2(n_194),
.B1(n_193),
.B2(n_228),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_319),
.B(n_203),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_353),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_375),
.B(n_247),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_362),
.Y(n_489)
);

BUFx8_ASAP7_75t_L g490 ( 
.A(n_376),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_361),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_367),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_361),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_363),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_411),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_369),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_406),
.B(n_386),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_420),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_386),
.B(n_202),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_439),
.B(n_188),
.Y(n_501)
);

INVx5_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_419),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_456),
.B(n_223),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_368),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_419),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_371),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_391),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_393),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_416),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_374),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_385),
.A2(n_253),
.B1(n_252),
.B2(n_243),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_377),
.B(n_410),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_429),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_414),
.B(n_242),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_434),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_435),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_455),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_438),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_389),
.A2(n_238),
.B(n_237),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_422),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_460),
.Y(n_524)
);

NAND2x1_ASAP7_75t_L g525 ( 
.A(n_388),
.B(n_145),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_423),
.Y(n_526)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_425),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_433),
.B(n_146),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_446),
.B(n_146),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_430),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_466),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_364),
.B(n_146),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_462),
.B(n_145),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_459),
.B(n_145),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_463),
.B(n_476),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_486),
.B(n_268),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_425),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_440),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_443),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_398),
.B(n_146),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_445),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_451),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_469),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_470),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_458),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_464),
.B(n_146),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_447),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_467),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_468),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_473),
.B(n_143),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_474),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_370),
.B(n_245),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_472),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_415),
.B(n_2),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_402),
.B(n_143),
.Y(n_555)
);

INVxp33_ASAP7_75t_SL g556 ( 
.A(n_465),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_370),
.B(n_147),
.Y(n_558)
);

INVx6_ASAP7_75t_L g559 ( 
.A(n_437),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_480),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_457),
.B(n_147),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_484),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_487),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_402),
.B(n_143),
.Y(n_564)
);

OAI21x1_ASAP7_75t_L g565 ( 
.A1(n_392),
.A2(n_147),
.B(n_158),
.Y(n_565)
);

OA21x2_ASAP7_75t_L g566 ( 
.A1(n_373),
.A2(n_158),
.B(n_245),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_384),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_378),
.B(n_158),
.Y(n_568)
);

OA21x2_ASAP7_75t_L g569 ( 
.A1(n_428),
.A2(n_268),
.B(n_73),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_407),
.B(n_268),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_366),
.B(n_88),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_477),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_424),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_372),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_448),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_378),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_382),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_383),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_400),
.B(n_1),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_382),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_482),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_448),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_427),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_442),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_387),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_454),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_475),
.B(n_483),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_483),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_481),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_407),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_399),
.Y(n_592)
);

HB1xp67_ASAP7_75t_L g593 ( 
.A(n_432),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_R g594 ( 
.A(n_408),
.B(n_479),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_452),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_471),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_403),
.Y(n_597)
);

AND2x6_ASAP7_75t_L g598 ( 
.A(n_404),
.B(n_409),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_449),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_453),
.Y(n_600)
);

AND2x2_ASAP7_75t_SL g601 ( 
.A(n_381),
.B(n_461),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_449),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_426),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_441),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_444),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g606 ( 
.A(n_432),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_421),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_449),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_401),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_417),
.B(n_418),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_380),
.Y(n_611)
);

CKINVDCx8_ASAP7_75t_R g612 ( 
.A(n_394),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g613 ( 
.A(n_431),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_436),
.B(n_365),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_395),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_478),
.A2(n_485),
.B1(n_390),
.B2(n_405),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_379),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_362),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_367),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_362),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_367),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_367),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_361),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_411),
.B(n_397),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_362),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_362),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_362),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_362),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_411),
.B(n_397),
.Y(n_629)
);

AND2x4_ASAP7_75t_L g630 ( 
.A(n_439),
.B(n_457),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_362),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_361),
.Y(n_632)
);

AND2x4_ASAP7_75t_L g633 ( 
.A(n_439),
.B(n_457),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_362),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_367),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_411),
.B(n_390),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_361),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_362),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_390),
.A2(n_429),
.B1(n_330),
.B2(n_294),
.Y(n_639)
);

BUFx8_ASAP7_75t_L g640 ( 
.A(n_376),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_367),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_362),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_411),
.B(n_397),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_362),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_375),
.B(n_385),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_411),
.B(n_375),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_361),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_361),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_362),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_411),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_411),
.B(n_397),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_367),
.Y(n_652)
);

BUFx6f_ASAP7_75t_L g653 ( 
.A(n_361),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_362),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_397),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_362),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_367),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_362),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_367),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_411),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_424),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_361),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_375),
.B(n_385),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_375),
.B(n_385),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_367),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_375),
.B(n_385),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_362),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_375),
.B(n_385),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_362),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_367),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_362),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_367),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_375),
.B(n_385),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_375),
.B(n_385),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_362),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_362),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_362),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_367),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_362),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_362),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_362),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_361),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_361),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_364),
.B(n_400),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g685 ( 
.A(n_411),
.Y(n_685)
);

OA21x2_ASAP7_75t_L g686 ( 
.A1(n_389),
.A2(n_373),
.B(n_363),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_367),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_361),
.Y(n_688)
);

BUFx2_ASAP7_75t_L g689 ( 
.A(n_411),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_367),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_362),
.Y(n_691)
);

CKINVDCx6p67_ASAP7_75t_R g692 ( 
.A(n_432),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_367),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_362),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_411),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_362),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_367),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_362),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_411),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_361),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_362),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_411),
.B(n_375),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_362),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_362),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_362),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_362),
.Y(n_706)
);

AND3x1_ASAP7_75t_L g707 ( 
.A(n_375),
.B(n_397),
.C(n_364),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_375),
.B(n_385),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_375),
.B(n_385),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_367),
.Y(n_710)
);

AND2x4_ASAP7_75t_L g711 ( 
.A(n_439),
.B(n_457),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_361),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_362),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_362),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_411),
.B(n_375),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_361),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_367),
.Y(n_717)
);

BUFx2_ASAP7_75t_L g718 ( 
.A(n_411),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_361),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_411),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_361),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_362),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_361),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_424),
.Y(n_724)
);

OA21x2_ASAP7_75t_L g725 ( 
.A1(n_389),
.A2(n_373),
.B(n_363),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_367),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_375),
.B(n_385),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_411),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_367),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_411),
.B(n_375),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_411),
.B(n_397),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_362),
.Y(n_732)
);

HB1xp67_ASAP7_75t_L g733 ( 
.A(n_411),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_362),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_362),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_361),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_SL g737 ( 
.A1(n_390),
.A2(n_429),
.B1(n_330),
.B2(n_294),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_375),
.B(n_385),
.Y(n_738)
);

OAI21x1_ASAP7_75t_L g739 ( 
.A1(n_389),
.A2(n_388),
.B(n_385),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_375),
.A2(n_406),
.B1(n_411),
.B2(n_385),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_411),
.B(n_397),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_375),
.B(n_385),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_411),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_362),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_362),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_411),
.B(n_397),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_439),
.B(n_457),
.Y(n_747)
);

BUFx2_ASAP7_75t_L g748 ( 
.A(n_411),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_411),
.B(n_375),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_362),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_362),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_362),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_375),
.B(n_385),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_367),
.Y(n_754)
);

INVx4_ASAP7_75t_L g755 ( 
.A(n_424),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_367),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_362),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_362),
.Y(n_758)
);

CKINVDCx6p67_ASAP7_75t_R g759 ( 
.A(n_432),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_415),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_362),
.Y(n_761)
);

CKINVDCx16_ASAP7_75t_R g762 ( 
.A(n_438),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_362),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_456),
.B(n_375),
.Y(n_764)
);

HB1xp67_ASAP7_75t_L g765 ( 
.A(n_411),
.Y(n_765)
);

OA21x2_ASAP7_75t_L g766 ( 
.A1(n_389),
.A2(n_373),
.B(n_363),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_367),
.Y(n_767)
);

INVx3_ASAP7_75t_L g768 ( 
.A(n_361),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_SL g769 ( 
.A(n_417),
.B(n_418),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_362),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_362),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_SL g772 ( 
.A(n_417),
.B(n_418),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_367),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_362),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_415),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_362),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_362),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_362),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_367),
.Y(n_779)
);

BUFx8_ASAP7_75t_L g780 ( 
.A(n_376),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_362),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_367),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_397),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_411),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_SL g785 ( 
.A(n_411),
.B(n_390),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_367),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_456),
.A2(n_385),
.B1(n_411),
.B2(n_375),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_362),
.Y(n_788)
);

AND2x6_ASAP7_75t_L g789 ( 
.A(n_364),
.B(n_400),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_411),
.B(n_397),
.Y(n_790)
);

INVx3_ASAP7_75t_L g791 ( 
.A(n_361),
.Y(n_791)
);

NAND2xp33_ASAP7_75t_R g792 ( 
.A(n_614),
.B(n_535),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_567),
.Y(n_793)
);

BUFx10_ASAP7_75t_L g794 ( 
.A(n_590),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_489),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_494),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_505),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_764),
.B(n_514),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_508),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_645),
.B(n_663),
.Y(n_800)
);

INVx4_ASAP7_75t_L g801 ( 
.A(n_590),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_661),
.B(n_755),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_491),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_664),
.B(n_666),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_491),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_668),
.B(n_673),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_512),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_493),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_493),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_515),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_573),
.B(n_724),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_506),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_523),
.Y(n_813)
);

NAND2x1_ASAP7_75t_L g814 ( 
.A(n_583),
.B(n_584),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_596),
.B(n_595),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_526),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_SL g817 ( 
.A(n_556),
.B(n_572),
.Y(n_817)
);

AND2x6_ASAP7_75t_L g818 ( 
.A(n_597),
.B(n_586),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_674),
.B(n_708),
.Y(n_819)
);

INVx3_ASAP7_75t_L g820 ( 
.A(n_506),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_537),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_530),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_488),
.A2(n_709),
.B1(n_738),
.B2(n_727),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_742),
.B(n_753),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_740),
.B(n_655),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_538),
.Y(n_826)
);

BUFx2_ASAP7_75t_L g827 ( 
.A(n_510),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_539),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_541),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_760),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_707),
.B(n_769),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_542),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_603),
.A2(n_607),
.B1(n_604),
.B2(n_605),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_545),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_537),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_582),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_548),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_549),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_551),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_582),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_588),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_532),
.B(n_504),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_562),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_563),
.Y(n_844)
);

AOI22xp33_ASAP7_75t_L g845 ( 
.A1(n_585),
.A2(n_533),
.B1(n_620),
.B2(n_618),
.Y(n_845)
);

AOI21x1_ASAP7_75t_L g846 ( 
.A1(n_525),
.A2(n_529),
.B(n_528),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_624),
.B(n_629),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_643),
.B(n_651),
.Y(n_848)
);

BUFx4f_ASAP7_75t_L g849 ( 
.A(n_692),
.Y(n_849)
);

INVx2_ASAP7_75t_SL g850 ( 
.A(n_731),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_SL g851 ( 
.A(n_775),
.B(n_521),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_625),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_762),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_626),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_627),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_598),
.B(n_684),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_628),
.A2(n_631),
.B1(n_638),
.B2(n_634),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_642),
.Y(n_858)
);

INVx2_ASAP7_75t_SL g859 ( 
.A(n_741),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_644),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_SL g861 ( 
.A1(n_601),
.A2(n_616),
.B1(n_737),
.B2(n_639),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_746),
.B(n_790),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_588),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_507),
.B(n_783),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_649),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_654),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_656),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_658),
.B(n_667),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_772),
.B(n_787),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_623),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_669),
.B(n_671),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_509),
.B(n_646),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_623),
.Y(n_873)
);

AND3x4_ASAP7_75t_L g874 ( 
.A(n_575),
.B(n_615),
.C(n_591),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_675),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_676),
.B(n_677),
.Y(n_876)
);

INVx8_ASAP7_75t_L g877 ( 
.A(n_598),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_611),
.B(n_610),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_495),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_647),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_679),
.B(n_680),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_647),
.Y(n_882)
);

INVx4_ASAP7_75t_L g883 ( 
.A(n_648),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_681),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_691),
.Y(n_885)
);

BUFx10_ASAP7_75t_L g886 ( 
.A(n_559),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_650),
.B(n_689),
.Y(n_887)
);

NOR3xp33_ASAP7_75t_L g888 ( 
.A(n_498),
.B(n_785),
.C(n_636),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_694),
.B(n_696),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_698),
.A2(n_752),
.B1(n_751),
.B2(n_750),
.Y(n_890)
);

AO21x2_ASAP7_75t_L g891 ( 
.A1(n_589),
.A2(n_739),
.B(n_571),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_701),
.B(n_703),
.Y(n_892)
);

INVx5_ASAP7_75t_L g893 ( 
.A(n_579),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_660),
.Y(n_894)
);

AND2x6_ASAP7_75t_L g895 ( 
.A(n_600),
.B(n_555),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_704),
.Y(n_896)
);

INVx4_ASAP7_75t_L g897 ( 
.A(n_648),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_699),
.B(n_718),
.Y(n_898)
);

AND2x4_ASAP7_75t_L g899 ( 
.A(n_587),
.B(n_503),
.Y(n_899)
);

OR2x6_ASAP7_75t_L g900 ( 
.A(n_653),
.B(n_662),
.Y(n_900)
);

AND3x2_ASAP7_75t_L g901 ( 
.A(n_593),
.B(n_606),
.C(n_520),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_705),
.B(n_706),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_713),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_714),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_748),
.B(n_511),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_722),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_653),
.Y(n_907)
);

INVx4_ASAP7_75t_SL g908 ( 
.A(n_579),
.Y(n_908)
);

OAI22xp33_ASAP7_75t_L g909 ( 
.A1(n_613),
.A2(n_763),
.B1(n_734),
.B2(n_732),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_735),
.Y(n_910)
);

BUFx10_ASAP7_75t_L g911 ( 
.A(n_501),
.Y(n_911)
);

BUFx10_ASAP7_75t_L g912 ( 
.A(n_662),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_744),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_745),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_757),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_702),
.B(n_715),
.Y(n_916)
);

INVx6_ASAP7_75t_L g917 ( 
.A(n_490),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_682),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_758),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_544),
.B(n_516),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_791),
.B(n_527),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_761),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_770),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_682),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_L g925 ( 
.A1(n_771),
.A2(n_777),
.B1(n_788),
.B2(n_781),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_774),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_776),
.B(n_778),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_564),
.B(n_570),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_492),
.Y(n_929)
);

BUFx4f_ASAP7_75t_L g930 ( 
.A(n_759),
.Y(n_930)
);

HB1xp67_ASAP7_75t_L g931 ( 
.A(n_685),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_684),
.A2(n_789),
.B1(n_497),
.B2(n_499),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_684),
.A2(n_789),
.B1(n_496),
.B2(n_635),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_730),
.A2(n_749),
.B1(n_592),
.B2(n_765),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_594),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_683),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_695),
.B(n_720),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_518),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_728),
.B(n_733),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_789),
.B(n_574),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_743),
.B(n_784),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_519),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_578),
.B(n_524),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_513),
.B(n_540),
.C(n_517),
.Y(n_944)
);

AND3x2_ASAP7_75t_L g945 ( 
.A(n_617),
.B(n_581),
.C(n_630),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_531),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_543),
.B(n_553),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_633),
.B(n_711),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_576),
.B(n_577),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_683),
.Y(n_950)
);

INVx1_ASAP7_75t_SL g951 ( 
.A(n_700),
.Y(n_951)
);

INVx6_ASAP7_75t_L g952 ( 
.A(n_640),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_560),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_619),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_621),
.B(n_622),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_641),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_652),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_780),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_747),
.B(n_712),
.Y(n_959)
);

INVxp33_ASAP7_75t_L g960 ( 
.A(n_700),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_712),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_716),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_580),
.B(n_716),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_657),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_659),
.Y(n_965)
);

AO21x2_ASAP7_75t_L g966 ( 
.A1(n_546),
.A2(n_550),
.B(n_500),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_665),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_719),
.Y(n_968)
);

AND2x6_ASAP7_75t_L g969 ( 
.A(n_599),
.B(n_608),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_719),
.B(n_736),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_670),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_672),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_678),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_736),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_561),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_687),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_502),
.B(n_786),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_690),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_547),
.Y(n_979)
);

INVxp33_ASAP7_75t_L g980 ( 
.A(n_554),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_SL g981 ( 
.A(n_612),
.B(n_609),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_693),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_697),
.B(n_782),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_710),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_717),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_502),
.B(n_767),
.Y(n_986)
);

NAND2x1p5_ASAP7_75t_L g987 ( 
.A(n_557),
.B(n_637),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_726),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_632),
.B(n_688),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_721),
.B(n_723),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_729),
.B(n_779),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_754),
.B(n_773),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_756),
.B(n_534),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_686),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_768),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_766),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_536),
.A2(n_725),
.B1(n_602),
.B2(n_569),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_552),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_598),
.A2(n_579),
.B1(n_522),
.B2(n_568),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_558),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_565),
.B(n_566),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_655),
.B(n_624),
.Y(n_1002)
);

BUFx3_ASAP7_75t_L g1003 ( 
.A(n_573),
.Y(n_1003)
);

NAND3xp33_ASAP7_75t_L g1004 ( 
.A(n_764),
.B(n_375),
.C(n_377),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_567),
.Y(n_1005)
);

INVxp67_ASAP7_75t_SL g1006 ( 
.A(n_495),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_764),
.B(n_514),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_489),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_489),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_764),
.B(n_514),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_489),
.Y(n_1011)
);

INVxp67_ASAP7_75t_SL g1012 ( 
.A(n_495),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_567),
.Y(n_1013)
);

NAND3xp33_ASAP7_75t_L g1014 ( 
.A(n_764),
.B(n_375),
.C(n_377),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_514),
.B(n_645),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_489),
.Y(n_1016)
);

OR2x2_ASAP7_75t_L g1017 ( 
.A(n_655),
.B(n_294),
.Y(n_1017)
);

BUFx4f_ASAP7_75t_L g1018 ( 
.A(n_590),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_489),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_488),
.A2(n_604),
.B1(n_605),
.B2(n_406),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_567),
.Y(n_1021)
);

INVx1_ASAP7_75t_SL g1022 ( 
.A(n_655),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_590),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_514),
.B(n_764),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_764),
.B(n_514),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_489),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_SL g1027 ( 
.A(n_590),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_491),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_655),
.B(n_624),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_489),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_567),
.Y(n_1031)
);

INVx5_ASAP7_75t_L g1032 ( 
.A(n_590),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_567),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_567),
.Y(n_1034)
);

BUFx4f_ASAP7_75t_L g1035 ( 
.A(n_590),
.Y(n_1035)
);

INVx6_ASAP7_75t_L g1036 ( 
.A(n_490),
.Y(n_1036)
);

BUFx10_ASAP7_75t_L g1037 ( 
.A(n_590),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_514),
.B(n_645),
.Y(n_1038)
);

INVxp33_ASAP7_75t_SL g1039 ( 
.A(n_572),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_489),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_491),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_489),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_488),
.A2(n_604),
.B1(n_605),
.B2(n_406),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_489),
.Y(n_1044)
);

AND2x6_ASAP7_75t_L g1045 ( 
.A(n_596),
.B(n_595),
.Y(n_1045)
);

INVxp67_ASAP7_75t_SL g1046 ( 
.A(n_495),
.Y(n_1046)
);

INVx3_ASAP7_75t_L g1047 ( 
.A(n_491),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_572),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_489),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_567),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_573),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_590),
.B(n_661),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_514),
.B(n_764),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_514),
.B(n_645),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_567),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_489),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_SL g1057 ( 
.A(n_590),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_567),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_489),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_590),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_567),
.Y(n_1061)
);

XNOR2xp5_ASAP7_75t_L g1062 ( 
.A(n_639),
.B(n_429),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_489),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_655),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_489),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_590),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_573),
.Y(n_1067)
);

INVx2_ASAP7_75t_SL g1068 ( 
.A(n_624),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_489),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_567),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_590),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_572),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_590),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_514),
.B(n_645),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_764),
.B(n_375),
.C(n_377),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_764),
.B(n_514),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_514),
.B(n_764),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_590),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_567),
.Y(n_1079)
);

BUFx8_ASAP7_75t_SL g1080 ( 
.A(n_609),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_489),
.Y(n_1081)
);

INVx4_ASAP7_75t_SL g1082 ( 
.A(n_559),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_764),
.B(n_514),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_L g1084 ( 
.A(n_596),
.B(n_595),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_567),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_590),
.B(n_661),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_567),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_655),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_514),
.B(n_764),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_573),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_514),
.B(n_764),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_590),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_488),
.A2(n_604),
.B1(n_605),
.B2(n_406),
.Y(n_1093)
);

INVx8_ASAP7_75t_L g1094 ( 
.A(n_590),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_567),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_567),
.Y(n_1096)
);

INVx6_ASAP7_75t_L g1097 ( 
.A(n_490),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_567),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_489),
.Y(n_1099)
);

NAND2xp33_ASAP7_75t_L g1100 ( 
.A(n_596),
.B(n_595),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_514),
.B(n_645),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_567),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_764),
.B(n_514),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_567),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_567),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_510),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_489),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_567),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_514),
.B(n_645),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_624),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_489),
.Y(n_1111)
);

OAI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_514),
.A2(n_488),
.B1(n_663),
.B2(n_645),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_764),
.B(n_514),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_572),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_764),
.A2(n_603),
.B1(n_585),
.B2(n_514),
.Y(n_1115)
);

BUFx10_ASAP7_75t_L g1116 ( 
.A(n_590),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_567),
.Y(n_1117)
);

INVx4_ASAP7_75t_L g1118 ( 
.A(n_590),
.Y(n_1118)
);

BUFx4f_ASAP7_75t_L g1119 ( 
.A(n_590),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_624),
.Y(n_1120)
);

OR2x6_ASAP7_75t_L g1121 ( 
.A(n_590),
.B(n_661),
.Y(n_1121)
);

NOR2x1p5_ASAP7_75t_L g1122 ( 
.A(n_692),
.B(n_759),
.Y(n_1122)
);

BUFx3_ASAP7_75t_L g1123 ( 
.A(n_573),
.Y(n_1123)
);

OR2x6_ASAP7_75t_L g1124 ( 
.A(n_590),
.B(n_661),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_567),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_SL g1126 ( 
.A(n_514),
.B(n_645),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_489),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_514),
.B(n_764),
.Y(n_1128)
);

OAI22x1_ASAP7_75t_L g1129 ( 
.A1(n_764),
.A2(n_585),
.B1(n_740),
.B2(n_613),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_764),
.B(n_514),
.Y(n_1130)
);

CKINVDCx5p33_ASAP7_75t_R g1131 ( 
.A(n_572),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_514),
.B(n_764),
.Y(n_1132)
);

OR2x6_ASAP7_75t_L g1133 ( 
.A(n_590),
.B(n_661),
.Y(n_1133)
);

BUFx2_ASAP7_75t_L g1134 ( 
.A(n_510),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_567),
.Y(n_1135)
);

NOR2xp33_ASAP7_75t_L g1136 ( 
.A(n_764),
.B(n_514),
.Y(n_1136)
);

BUFx3_ASAP7_75t_L g1137 ( 
.A(n_573),
.Y(n_1137)
);

AND2x6_ASAP7_75t_L g1138 ( 
.A(n_596),
.B(n_595),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_764),
.B(n_514),
.Y(n_1139)
);

INVx5_ASAP7_75t_L g1140 ( 
.A(n_590),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_489),
.Y(n_1141)
);

NOR2x1p5_ASAP7_75t_L g1142 ( 
.A(n_692),
.B(n_759),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_491),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_567),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_567),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_489),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_764),
.B(n_514),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_489),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_489),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_491),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_655),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_514),
.B(n_764),
.Y(n_1152)
);

BUFx10_ASAP7_75t_L g1153 ( 
.A(n_590),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_573),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_590),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_514),
.B(n_764),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_489),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_489),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_567),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_567),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_491),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_590),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_567),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_514),
.B(n_645),
.Y(n_1164)
);

AO21x2_ASAP7_75t_L g1165 ( 
.A1(n_583),
.A2(n_586),
.B(n_584),
.Y(n_1165)
);

BUFx4f_ASAP7_75t_L g1166 ( 
.A(n_590),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_514),
.B(n_764),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_567),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_567),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_573),
.B(n_724),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_764),
.B(n_514),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_567),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_488),
.A2(n_604),
.B1(n_605),
.B2(n_406),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_489),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_514),
.B(n_764),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_489),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_514),
.B(n_764),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_SL g1178 ( 
.A(n_514),
.B(n_645),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_489),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_567),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_655),
.B(n_624),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_567),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_SL g1183 ( 
.A(n_514),
.B(n_645),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_491),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_567),
.Y(n_1185)
);

BUFx6f_ASAP7_75t_L g1186 ( 
.A(n_590),
.Y(n_1186)
);

INVx4_ASAP7_75t_L g1187 ( 
.A(n_590),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_567),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_764),
.B(n_514),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_489),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_596),
.A2(n_514),
.B1(n_595),
.B2(n_707),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_514),
.B(n_764),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_510),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_764),
.B(n_514),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_489),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_488),
.A2(n_604),
.B1(n_605),
.B2(n_406),
.Y(n_1196)
);

NAND2xp33_ASAP7_75t_L g1197 ( 
.A(n_596),
.B(n_595),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_489),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_567),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_590),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_573),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_514),
.B(n_764),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_514),
.B(n_764),
.Y(n_1203)
);

INVx3_ASAP7_75t_L g1204 ( 
.A(n_491),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_624),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_596),
.A2(n_514),
.B1(n_595),
.B2(n_707),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_590),
.Y(n_1207)
);

OR2x6_ASAP7_75t_L g1208 ( 
.A(n_590),
.B(n_661),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_491),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_596),
.A2(n_514),
.B1(n_595),
.B2(n_707),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_514),
.B(n_764),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_514),
.B(n_764),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_655),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_590),
.Y(n_1214)
);

INVx5_ASAP7_75t_L g1215 ( 
.A(n_590),
.Y(n_1215)
);

OAI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_514),
.A2(n_488),
.B1(n_663),
.B2(n_645),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_514),
.B(n_764),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_489),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_488),
.A2(n_604),
.B1(n_605),
.B2(n_406),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_489),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_572),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_SL g1222 ( 
.A(n_556),
.B(n_572),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_510),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_567),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_514),
.B(n_645),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_514),
.B(n_764),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_SL g1227 ( 
.A(n_514),
.B(n_645),
.Y(n_1227)
);

INVx3_ASAP7_75t_L g1228 ( 
.A(n_491),
.Y(n_1228)
);

INVx8_ASAP7_75t_L g1229 ( 
.A(n_590),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_567),
.Y(n_1230)
);

BUFx6f_ASAP7_75t_L g1231 ( 
.A(n_590),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_489),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_590),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_514),
.B(n_645),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_567),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_488),
.A2(n_604),
.B1(n_605),
.B2(n_406),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_514),
.B(n_764),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_514),
.B(n_764),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_590),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_514),
.B(n_764),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_514),
.B(n_764),
.Y(n_1241)
);

BUFx5_ASAP7_75t_L g1242 ( 
.A(n_969),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_798),
.B(n_1007),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1010),
.B(n_1025),
.Y(n_1245)
);

NOR2xp33_ASAP7_75t_L g1246 ( 
.A(n_1076),
.B(n_1083),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_795),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1032),
.B(n_1140),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1181),
.B(n_1103),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_810),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_SL g1252 ( 
.A(n_1039),
.B(n_830),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1113),
.B(n_1130),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1136),
.B(n_1139),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1147),
.B(n_1171),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1210),
.B(n_1112),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1216),
.B(n_1115),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1023),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1094),
.B(n_1229),
.Y(n_1259)
);

BUFx5_ASAP7_75t_L g1260 ( 
.A(n_969),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_796),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1189),
.B(n_1194),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1004),
.A2(n_1075),
.B(n_1014),
.C(n_819),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_797),
.Y(n_1264)
);

AND2x4_ASAP7_75t_L g1265 ( 
.A(n_1032),
.B(n_1140),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_799),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_807),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_813),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_816),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_828),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_832),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1024),
.B(n_1053),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_834),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_823),
.B(n_1077),
.Y(n_1274)
);

INVx2_ASAP7_75t_L g1275 ( 
.A(n_837),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1089),
.B(n_1241),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_1214),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1091),
.B(n_1240),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1128),
.B(n_1132),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1152),
.B(n_1156),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_822),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_794),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1167),
.B(n_1175),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_838),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1177),
.B(n_1192),
.Y(n_1285)
);

INVxp67_ASAP7_75t_L g1286 ( 
.A(n_1223),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_847),
.B(n_1202),
.Y(n_1287)
);

NOR2xp67_ASAP7_75t_L g1288 ( 
.A(n_1048),
.B(n_1072),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1203),
.B(n_1211),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1212),
.B(n_1217),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1226),
.B(n_1237),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_839),
.Y(n_1292)
);

NAND2xp33_ASAP7_75t_SL g1293 ( 
.A(n_1129),
.B(n_1023),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1238),
.B(n_800),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_826),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1020),
.A2(n_1093),
.B1(n_1173),
.B2(n_1043),
.Y(n_1296)
);

INVxp33_ASAP7_75t_L g1297 ( 
.A(n_920),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_829),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1015),
.B(n_1038),
.Y(n_1299)
);

INVx1_ASAP7_75t_SL g1300 ( 
.A(n_827),
.Y(n_1300)
);

BUFx5_ASAP7_75t_L g1301 ( 
.A(n_969),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1054),
.B(n_1074),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1101),
.B(n_1109),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1022),
.B(n_1064),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_844),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_843),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_SL g1307 ( 
.A(n_1114),
.B(n_1131),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1126),
.B(n_1164),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1178),
.B(n_1183),
.Y(n_1309)
);

INVx2_ASAP7_75t_SL g1310 ( 
.A(n_1214),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1225),
.B(n_1227),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_865),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_866),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1234),
.B(n_804),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_875),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_884),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_806),
.B(n_824),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_842),
.B(n_1196),
.Y(n_1318)
);

NAND3xp33_ASAP7_75t_L g1319 ( 
.A(n_1219),
.B(n_1236),
.C(n_1100),
.Y(n_1319)
);

AND2x4_ASAP7_75t_SL g1320 ( 
.A(n_1037),
.B(n_1116),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1106),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_833),
.B(n_815),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_815),
.B(n_1045),
.Y(n_1323)
);

INVx2_ASAP7_75t_L g1324 ( 
.A(n_903),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_848),
.B(n_862),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_906),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_852),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_815),
.B(n_1045),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_910),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_854),
.Y(n_1330)
);

BUFx5_ASAP7_75t_L g1331 ( 
.A(n_818),
.Y(n_1331)
);

BUFx5_ASAP7_75t_L g1332 ( 
.A(n_818),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1045),
.B(n_1138),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1134),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_913),
.Y(n_1335)
);

NOR2xp33_ASAP7_75t_L g1336 ( 
.A(n_1088),
.B(n_1151),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1215),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_914),
.Y(n_1338)
);

NAND2xp33_ASAP7_75t_L g1339 ( 
.A(n_1138),
.B(n_895),
.Y(n_1339)
);

NOR2xp67_ASAP7_75t_L g1340 ( 
.A(n_1221),
.B(n_1215),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_855),
.Y(n_1341)
);

INVxp67_ASAP7_75t_L g1342 ( 
.A(n_1193),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1138),
.B(n_1084),
.Y(n_1343)
);

INVx4_ASAP7_75t_L g1344 ( 
.A(n_1094),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_858),
.Y(n_1345)
);

NOR2xp67_ASAP7_75t_L g1346 ( 
.A(n_935),
.B(n_801),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1197),
.B(n_845),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_860),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_916),
.B(n_868),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_SL g1350 ( 
.A(n_817),
.B(n_1222),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_922),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_871),
.B(n_876),
.Y(n_1352)
);

BUFx5_ASAP7_75t_L g1353 ( 
.A(n_818),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_881),
.B(n_889),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_892),
.B(n_902),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_927),
.B(n_928),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1213),
.B(n_1017),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_867),
.B(n_885),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_872),
.B(n_1205),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_896),
.B(n_904),
.Y(n_1360)
);

AND2x2_ASAP7_75t_SL g1361 ( 
.A(n_851),
.B(n_981),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_915),
.B(n_919),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_850),
.B(n_859),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1080),
.Y(n_1364)
);

HB1xp67_ASAP7_75t_L g1365 ( 
.A(n_931),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_909),
.B(n_1068),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_923),
.B(n_926),
.Y(n_1367)
);

NOR2xp33_ASAP7_75t_L g1368 ( 
.A(n_825),
.B(n_939),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1008),
.B(n_1009),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1011),
.B(n_1016),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1019),
.B(n_1026),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_878),
.B(n_864),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1110),
.B(n_1120),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_938),
.Y(n_1374)
);

INVxp33_ASAP7_75t_L g1375 ( 
.A(n_1066),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_L g1376 ( 
.A(n_1066),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1030),
.B(n_1040),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1042),
.B(n_1044),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1049),
.B(n_1056),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1059),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1063),
.B(n_1065),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1069),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_942),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_SL g1384 ( 
.A(n_869),
.B(n_893),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1229),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1081),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1099),
.B(n_1107),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1111),
.B(n_1127),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1141),
.B(n_1146),
.Y(n_1389)
);

NAND2xp5_ASAP7_75t_SL g1390 ( 
.A(n_893),
.B(n_888),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1148),
.B(n_1149),
.Y(n_1391)
);

BUFx2_ASAP7_75t_R g1392 ( 
.A(n_853),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1071),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_879),
.B(n_894),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_962),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_954),
.Y(n_1396)
);

INVxp33_ASAP7_75t_L g1397 ( 
.A(n_1071),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1157),
.B(n_1158),
.Y(n_1398)
);

NAND3xp33_ASAP7_75t_L g1399 ( 
.A(n_861),
.B(n_792),
.C(n_857),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1174),
.B(n_1176),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_965),
.Y(n_1401)
);

NAND3xp33_ASAP7_75t_L g1402 ( 
.A(n_890),
.B(n_925),
.C(n_934),
.Y(n_1402)
);

NAND3xp33_ASAP7_75t_L g1403 ( 
.A(n_905),
.B(n_831),
.C(n_937),
.Y(n_1403)
);

INVxp33_ASAP7_75t_L g1404 ( 
.A(n_1073),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1179),
.B(n_1190),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_967),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1195),
.B(n_1198),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1218),
.B(n_1220),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_971),
.Y(n_1409)
);

NOR3xp33_ASAP7_75t_L g1410 ( 
.A(n_887),
.B(n_898),
.C(n_941),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1232),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1073),
.B(n_1078),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_973),
.Y(n_1413)
);

NOR2xp67_ASAP7_75t_L g1414 ( 
.A(n_1060),
.B(n_1118),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_895),
.B(n_793),
.Y(n_1415)
);

NAND2xp33_ASAP7_75t_L g1416 ( 
.A(n_895),
.B(n_877),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_947),
.Y(n_1417)
);

NOR2xp67_ASAP7_75t_L g1418 ( 
.A(n_1155),
.B(n_1162),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1005),
.B(n_1013),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1003),
.B(n_1051),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1021),
.B(n_1031),
.Y(n_1421)
);

NOR3xp33_ASAP7_75t_L g1422 ( 
.A(n_944),
.B(n_1233),
.C(n_1187),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_874),
.A2(n_856),
.B1(n_1050),
.B2(n_1235),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_984),
.Y(n_1424)
);

NOR2xp67_ASAP7_75t_L g1425 ( 
.A(n_1239),
.B(n_995),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1033),
.B(n_1034),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_955),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_SL g1428 ( 
.A(n_1078),
.B(n_1092),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1006),
.B(n_1012),
.Y(n_1429)
);

NOR3xp33_ASAP7_75t_L g1430 ( 
.A(n_948),
.B(n_1046),
.C(n_959),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1055),
.B(n_1058),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_988),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1061),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1070),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_SL g1435 ( 
.A(n_1092),
.B(n_1186),
.Y(n_1435)
);

NOR3xp33_ASAP7_75t_L g1436 ( 
.A(n_840),
.B(n_897),
.C(n_883),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_960),
.B(n_1186),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_932),
.A2(n_933),
.B1(n_940),
.B2(n_1224),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_943),
.B(n_946),
.C(n_929),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_983),
.Y(n_1440)
);

AO221x1_ASAP7_75t_L g1441 ( 
.A1(n_997),
.A2(n_1231),
.B1(n_1200),
.B2(n_880),
.C(n_936),
.Y(n_1441)
);

INVx8_ASAP7_75t_L g1442 ( 
.A(n_1027),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1079),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1085),
.B(n_1087),
.Y(n_1444)
);

NAND2x1_ASAP7_75t_L g1445 ( 
.A(n_900),
.B(n_970),
.Y(n_1445)
);

NOR2xp33_ASAP7_75t_L g1446 ( 
.A(n_1200),
.B(n_1231),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1095),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_950),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_991),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_992),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_951),
.B(n_1096),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1098),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1102),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1104),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1105),
.B(n_1108),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_SL g1456 ( 
.A(n_1018),
.B(n_1035),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1117),
.Y(n_1457)
);

INVxp67_ASAP7_75t_SL g1458 ( 
.A(n_805),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_989),
.B(n_990),
.Y(n_1459)
);

INVx4_ASAP7_75t_L g1460 ( 
.A(n_1052),
.Y(n_1460)
);

NAND2xp33_ASAP7_75t_L g1461 ( 
.A(n_877),
.B(n_805),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1119),
.B(n_1166),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_SL g1463 ( 
.A(n_1207),
.B(n_1125),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1135),
.B(n_1144),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1145),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_SL g1466 ( 
.A(n_849),
.B(n_930),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1159),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1160),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1163),
.B(n_1168),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1169),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1172),
.B(n_1180),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1182),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_SL g1473 ( 
.A(n_1185),
.B(n_1188),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_808),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1199),
.B(n_1230),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_953),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1153),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1062),
.A2(n_979),
.B1(n_899),
.B2(n_975),
.C(n_1057),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_L g1479 ( 
.A(n_956),
.B(n_957),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_964),
.B(n_972),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_976),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_978),
.Y(n_1482)
);

INVx5_ASAP7_75t_L g1483 ( 
.A(n_1052),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_982),
.Y(n_1484)
);

INVxp33_ASAP7_75t_L g1485 ( 
.A(n_811),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_985),
.B(n_998),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1165),
.Y(n_1487)
);

NOR2xp67_ASAP7_75t_L g1488 ( 
.A(n_961),
.B(n_1170),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_900),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_SL g1490 ( 
.A(n_886),
.B(n_958),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_L g1491 ( 
.A(n_808),
.B(n_809),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1000),
.B(n_949),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1086),
.B(n_1121),
.Y(n_1493)
);

NAND2xp33_ASAP7_75t_SL g1494 ( 
.A(n_809),
.B(n_821),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_814),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_963),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_993),
.B(n_1047),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_803),
.B(n_924),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_821),
.Y(n_1499)
);

NOR2xp67_ASAP7_75t_L g1500 ( 
.A(n_820),
.B(n_1228),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_994),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_968),
.B(n_1161),
.Y(n_1502)
);

NAND2xp33_ASAP7_75t_L g1503 ( 
.A(n_835),
.B(n_873),
.Y(n_1503)
);

INVx2_ASAP7_75t_SL g1504 ( 
.A(n_912),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_996),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_987),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1028),
.B(n_1209),
.Y(n_1507)
);

INVxp67_ASAP7_75t_L g1508 ( 
.A(n_970),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1041),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1143),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1150),
.Y(n_1511)
);

BUFx6f_ASAP7_75t_L g1512 ( 
.A(n_835),
.Y(n_1512)
);

NAND2xp33_ASAP7_75t_L g1513 ( 
.A(n_841),
.B(n_873),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_841),
.B(n_974),
.Y(n_1514)
);

NOR2x1_ASAP7_75t_L g1515 ( 
.A(n_1086),
.B(n_1208),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_863),
.B(n_974),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_863),
.B(n_870),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_870),
.B(n_882),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1184),
.B(n_1204),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_SL g1520 ( 
.A(n_882),
.B(n_908),
.Y(n_1520)
);

BUFx5_ASAP7_75t_L g1521 ( 
.A(n_812),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_836),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_921),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_907),
.B(n_918),
.Y(n_1524)
);

NOR2xp33_ASAP7_75t_L g1525 ( 
.A(n_1067),
.B(n_1123),
.Y(n_1525)
);

INVxp67_ASAP7_75t_L g1526 ( 
.A(n_1121),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_966),
.B(n_999),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_977),
.A2(n_986),
.B(n_1001),
.C(n_1090),
.Y(n_1528)
);

NAND2xp5_ASAP7_75t_L g1529 ( 
.A(n_1124),
.B(n_1208),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1124),
.B(n_1133),
.Y(n_1530)
);

NAND3xp33_ASAP7_75t_L g1531 ( 
.A(n_901),
.B(n_1133),
.C(n_1154),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_891),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1137),
.B(n_1201),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_945),
.B(n_802),
.Y(n_1534)
);

INVxp33_ASAP7_75t_L g1535 ( 
.A(n_980),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_802),
.B(n_846),
.Y(n_1536)
);

CKINVDCx20_ASAP7_75t_R g1537 ( 
.A(n_917),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_911),
.B(n_1082),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1142),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1122),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_952),
.B(n_1036),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1097),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1094),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_798),
.B(n_1007),
.Y(n_1546)
);

INVx2_ASAP7_75t_SL g1547 ( 
.A(n_1032),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_L g1548 ( 
.A(n_1023),
.Y(n_1548)
);

BUFx6f_ASAP7_75t_SL g1549 ( 
.A(n_886),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_798),
.B(n_1007),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_798),
.B(n_1007),
.Y(n_1551)
);

BUFx5_ASAP7_75t_L g1552 ( 
.A(n_969),
.Y(n_1552)
);

NOR2xp33_ASAP7_75t_L g1553 ( 
.A(n_798),
.B(n_1007),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1554)
);

AO221x1_ASAP7_75t_L g1555 ( 
.A1(n_1112),
.A2(n_616),
.B1(n_1216),
.B2(n_823),
.C(n_390),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_796),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_798),
.B(n_1007),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1023),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_798),
.B(n_1007),
.Y(n_1559)
);

AND2x2_ASAP7_75t_SL g1560 ( 
.A(n_851),
.B(n_601),
.Y(n_1560)
);

AO221x1_ASAP7_75t_L g1561 ( 
.A1(n_1112),
.A2(n_616),
.B1(n_1216),
.B2(n_823),
.C(n_390),
.Y(n_1561)
);

INVx4_ASAP7_75t_L g1562 ( 
.A(n_1032),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_796),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_798),
.B(n_1007),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_795),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_798),
.B(n_1007),
.Y(n_1566)
);

INVxp67_ASAP7_75t_L g1567 ( 
.A(n_1223),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_798),
.B(n_1007),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_798),
.B(n_1007),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1032),
.Y(n_1571)
);

NOR2xp67_ASAP7_75t_L g1572 ( 
.A(n_830),
.B(n_432),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_798),
.B(n_1007),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_796),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_796),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1032),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_SL g1577 ( 
.A(n_886),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1581)
);

NAND2xp33_ASAP7_75t_L g1582 ( 
.A(n_815),
.B(n_1045),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1032),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_796),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_798),
.B(n_1007),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_798),
.B(n_1007),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_798),
.B(n_1007),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_796),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_798),
.B(n_1007),
.Y(n_1591)
);

INVx2_ASAP7_75t_SL g1592 ( 
.A(n_1032),
.Y(n_1592)
);

AO221x1_ASAP7_75t_L g1593 ( 
.A1(n_1112),
.A2(n_616),
.B1(n_1216),
.B2(n_823),
.C(n_390),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_798),
.B(n_1007),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_798),
.B(n_1007),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_798),
.B(n_1007),
.Y(n_1596)
);

NAND3xp33_ASAP7_75t_L g1597 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_798),
.B(n_1007),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_798),
.B(n_1007),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_798),
.B(n_1007),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_798),
.B(n_1007),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_796),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_798),
.B(n_1007),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_798),
.B(n_1007),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_SL g1606 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1004),
.A2(n_1075),
.B1(n_1014),
.B2(n_798),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_796),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1094),
.B(n_1229),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_798),
.B(n_1007),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_796),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_827),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_795),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1024),
.B(n_1053),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_798),
.B(n_1007),
.Y(n_1618)
);

NOR3xp33_ASAP7_75t_L g1619 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_796),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_795),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_795),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_798),
.B(n_1007),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_L g1625 ( 
.A(n_815),
.B(n_1045),
.Y(n_1625)
);

INVxp67_ASAP7_75t_L g1626 ( 
.A(n_1223),
.Y(n_1626)
);

NAND2xp33_ASAP7_75t_L g1627 ( 
.A(n_815),
.B(n_1045),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_798),
.B(n_1007),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1629)
);

A2O1A1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_798),
.A2(n_1007),
.B(n_1025),
.C(n_1010),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_798),
.B(n_1007),
.Y(n_1632)
);

NOR3xp33_ASAP7_75t_L g1633 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1094),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_796),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_796),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_796),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_795),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_798),
.B(n_1007),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1032),
.B(n_1140),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_798),
.B(n_1007),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_798),
.B(n_1007),
.Y(n_1646)
);

BUFx6f_ASAP7_75t_L g1647 ( 
.A(n_1023),
.Y(n_1647)
);

A2O1A1Ixp33_ASAP7_75t_L g1648 ( 
.A1(n_798),
.A2(n_1007),
.B(n_1025),
.C(n_1010),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_796),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1032),
.B(n_1140),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_798),
.B(n_1007),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_795),
.Y(n_1652)
);

BUFx2_ASAP7_75t_R g1653 ( 
.A(n_1080),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_798),
.B(n_1007),
.Y(n_1654)
);

BUFx6f_ASAP7_75t_SL g1655 ( 
.A(n_886),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_827),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1094),
.Y(n_1657)
);

INVxp67_ASAP7_75t_L g1658 ( 
.A(n_1223),
.Y(n_1658)
);

INVx2_ASAP7_75t_L g1659 ( 
.A(n_796),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_798),
.B(n_1007),
.Y(n_1660)
);

NAND2xp33_ASAP7_75t_SL g1661 ( 
.A(n_1129),
.B(n_590),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_798),
.B(n_1007),
.Y(n_1663)
);

BUFx5_ASAP7_75t_L g1664 ( 
.A(n_969),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_798),
.B(n_1007),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_798),
.B(n_1007),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_798),
.B(n_1007),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_798),
.A2(n_1010),
.B1(n_1025),
.B2(n_1007),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_796),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_796),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_795),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1672)
);

NOR2xp33_ASAP7_75t_L g1673 ( 
.A(n_798),
.B(n_1007),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_SL g1674 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_798),
.B(n_1007),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_796),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1032),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_798),
.B(n_1007),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_796),
.Y(n_1681)
);

INVx2_ASAP7_75t_SL g1682 ( 
.A(n_1032),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_SL g1683 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_830),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_827),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1032),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_798),
.B(n_1007),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_795),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_796),
.Y(n_1689)
);

INVx2_ASAP7_75t_SL g1690 ( 
.A(n_1032),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_795),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_798),
.B(n_1007),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_796),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_798),
.B(n_1007),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_L g1697 ( 
.A(n_815),
.B(n_1045),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_798),
.B(n_1007),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_SL g1699 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1699)
);

AND2x4_ASAP7_75t_SL g1700 ( 
.A(n_794),
.B(n_1037),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_1032),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_798),
.B(n_1007),
.Y(n_1702)
);

NAND2xp33_ASAP7_75t_L g1703 ( 
.A(n_815),
.B(n_1045),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_798),
.B(n_1007),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_796),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_SL g1706 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_796),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1023),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_795),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_798),
.B(n_1007),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_795),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_798),
.B(n_1007),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_795),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_798),
.B(n_1007),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_796),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_798),
.B(n_1007),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_798),
.B(n_1007),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_SL g1719 ( 
.A(n_886),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1032),
.B(n_1140),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1024),
.B(n_1053),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_798),
.B(n_1007),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_795),
.Y(n_1724)
);

AO221x1_ASAP7_75t_L g1725 ( 
.A1(n_1112),
.A2(n_616),
.B1(n_1216),
.B2(n_823),
.C(n_390),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_798),
.B(n_1007),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_798),
.B(n_1007),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_SL g1729 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1729)
);

BUFx8_ASAP7_75t_L g1730 ( 
.A(n_1027),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_795),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_795),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_795),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_798),
.B(n_1007),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_795),
.Y(n_1738)
);

BUFx8_ASAP7_75t_L g1739 ( 
.A(n_1027),
.Y(n_1739)
);

INVx2_ASAP7_75t_SL g1740 ( 
.A(n_1032),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1023),
.Y(n_1741)
);

NOR2x1p5_ASAP7_75t_L g1742 ( 
.A(n_801),
.B(n_692),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1004),
.A2(n_1075),
.B1(n_1014),
.B2(n_798),
.Y(n_1743)
);

NOR2xp33_ASAP7_75t_L g1744 ( 
.A(n_798),
.B(n_1007),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_798),
.B(n_1007),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_798),
.B(n_1007),
.Y(n_1746)
);

NAND2x1_ASAP7_75t_L g1747 ( 
.A(n_969),
.B(n_818),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_SL g1748 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_798),
.B(n_1007),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_798),
.B(n_1007),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_798),
.B(n_1007),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_796),
.Y(n_1752)
);

NOR2xp33_ASAP7_75t_L g1753 ( 
.A(n_798),
.B(n_1007),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_798),
.B(n_1007),
.Y(n_1754)
);

AOI22xp33_ASAP7_75t_L g1755 ( 
.A1(n_1004),
.A2(n_1075),
.B1(n_1014),
.B2(n_798),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1223),
.Y(n_1756)
);

INVx1_ASAP7_75t_SL g1757 ( 
.A(n_827),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_795),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_795),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_798),
.B(n_1007),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_798),
.B(n_1007),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_795),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_798),
.B(n_1007),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_796),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_796),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_L g1766 ( 
.A(n_830),
.B(n_432),
.Y(n_1766)
);

NOR3xp33_ASAP7_75t_L g1767 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1768)
);

INVxp33_ASAP7_75t_SL g1769 ( 
.A(n_817),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_798),
.B(n_1007),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_795),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_798),
.B(n_1007),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_795),
.Y(n_1773)
);

BUFx3_ASAP7_75t_L g1774 ( 
.A(n_1094),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_795),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_795),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_795),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_798),
.B(n_1007),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_798),
.B(n_1007),
.Y(n_1780)
);

NOR3xp33_ASAP7_75t_L g1781 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_798),
.B(n_1007),
.Y(n_1782)
);

NOR3xp33_ASAP7_75t_L g1783 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_SL g1784 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1784)
);

BUFx5_ASAP7_75t_L g1785 ( 
.A(n_969),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_794),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_798),
.B(n_1007),
.Y(n_1787)
);

NOR3xp33_ASAP7_75t_L g1788 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_796),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_798),
.B(n_1007),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_798),
.B(n_1007),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_795),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_796),
.Y(n_1793)
);

NAND2xp33_ASAP7_75t_L g1794 ( 
.A(n_815),
.B(n_1045),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_796),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_794),
.Y(n_1796)
);

NAND2xp33_ASAP7_75t_L g1797 ( 
.A(n_815),
.B(n_1045),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_795),
.Y(n_1799)
);

BUFx6f_ASAP7_75t_L g1800 ( 
.A(n_1023),
.Y(n_1800)
);

INVx2_ASAP7_75t_SL g1801 ( 
.A(n_1032),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_798),
.B(n_1007),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_795),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_795),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_796),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_795),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_830),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_795),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_795),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_798),
.B(n_1007),
.Y(n_1810)
);

BUFx6f_ASAP7_75t_L g1811 ( 
.A(n_1023),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_796),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_798),
.B(n_1007),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_796),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_SL g1815 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1815)
);

BUFx6f_ASAP7_75t_L g1816 ( 
.A(n_1023),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_796),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_795),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_796),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1223),
.Y(n_1820)
);

BUFx6f_ASAP7_75t_L g1821 ( 
.A(n_1023),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_796),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_796),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_798),
.B(n_1007),
.Y(n_1825)
);

NOR3xp33_ASAP7_75t_L g1826 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1826)
);

NOR3xp33_ASAP7_75t_L g1827 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1827)
);

AND2x2_ASAP7_75t_SL g1828 ( 
.A(n_851),
.B(n_601),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_798),
.B(n_1007),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_795),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_798),
.B(n_1007),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_798),
.B(n_1007),
.Y(n_1832)
);

NOR2xp67_ASAP7_75t_L g1833 ( 
.A(n_830),
.B(n_432),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_SL g1834 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_SL g1835 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_798),
.B(n_1007),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_L g1837 ( 
.A(n_798),
.B(n_1007),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_798),
.B(n_1007),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_SL g1839 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1839)
);

BUFx6f_ASAP7_75t_L g1840 ( 
.A(n_1023),
.Y(n_1840)
);

NOR2xp67_ASAP7_75t_L g1841 ( 
.A(n_830),
.B(n_432),
.Y(n_1841)
);

AO221x1_ASAP7_75t_L g1842 ( 
.A1(n_1112),
.A2(n_616),
.B1(n_1216),
.B2(n_823),
.C(n_390),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_798),
.B(n_1007),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_798),
.B(n_1007),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_798),
.B(n_1007),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_796),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_795),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_795),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_798),
.B(n_1007),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1023),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_795),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_798),
.B(n_1007),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_SL g1853 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_830),
.Y(n_1855)
);

BUFx2_ASAP7_75t_L g1856 ( 
.A(n_827),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_SL g1858 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_795),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1032),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_795),
.Y(n_1861)
);

BUFx3_ASAP7_75t_L g1862 ( 
.A(n_1094),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_798),
.B(n_1007),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_796),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1094),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_SL g1867 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_798),
.B(n_1007),
.Y(n_1868)
);

NOR2xp67_ASAP7_75t_L g1869 ( 
.A(n_830),
.B(n_432),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_798),
.B(n_1007),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_798),
.B(n_1007),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1223),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_798),
.B(n_1007),
.Y(n_1873)
);

NOR2xp67_ASAP7_75t_L g1874 ( 
.A(n_830),
.B(n_432),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_796),
.Y(n_1875)
);

INVx8_ASAP7_75t_L g1876 ( 
.A(n_1094),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_795),
.Y(n_1877)
);

AOI22xp33_ASAP7_75t_L g1878 ( 
.A1(n_1004),
.A2(n_1075),
.B1(n_1014),
.B2(n_798),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_SL g1879 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_SL g1880 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_798),
.B(n_1007),
.Y(n_1881)
);

XOR2xp5_ASAP7_75t_L g1882 ( 
.A(n_853),
.B(n_429),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_795),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_795),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_795),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1094),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_798),
.B(n_1007),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_1023),
.Y(n_1888)
);

INVx8_ASAP7_75t_L g1889 ( 
.A(n_1094),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_798),
.B(n_1007),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_798),
.B(n_1007),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_798),
.B(n_1007),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_798),
.B(n_1007),
.Y(n_1893)
);

NOR3xp33_ASAP7_75t_L g1894 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_798),
.B(n_1007),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_798),
.B(n_1007),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_L g1897 ( 
.A(n_798),
.B(n_1007),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_795),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_798),
.B(n_1007),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_798),
.B(n_1007),
.Y(n_1900)
);

NAND3xp33_ASAP7_75t_L g1901 ( 
.A(n_1004),
.B(n_1075),
.C(n_1014),
.Y(n_1901)
);

INVx2_ASAP7_75t_SL g1902 ( 
.A(n_1032),
.Y(n_1902)
);

NAND2xp33_ASAP7_75t_L g1903 ( 
.A(n_815),
.B(n_1045),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_798),
.B(n_1007),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_798),
.B(n_1007),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_798),
.B(n_1007),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_796),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_SL g1909 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_798),
.B(n_1007),
.Y(n_1910)
);

NOR2xp33_ASAP7_75t_L g1911 ( 
.A(n_798),
.B(n_1007),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_798),
.B(n_1007),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_SL g1913 ( 
.A(n_1191),
.B(n_1206),
.Y(n_1913)
);

INVx2_ASAP7_75t_L g1914 ( 
.A(n_796),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1002),
.B(n_1029),
.Y(n_1915)
);

INVxp33_ASAP7_75t_L g1916 ( 
.A(n_1223),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_795),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_796),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_798),
.B(n_1007),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_795),
.Y(n_1920)
);

OA21x2_ASAP7_75t_L g1921 ( 
.A1(n_994),
.A2(n_996),
.B(n_739),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_798),
.B(n_1007),
.Y(n_1922)
);

NOR2xp33_ASAP7_75t_L g1923 ( 
.A(n_798),
.B(n_1007),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_796),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_SL g1925 ( 
.A(n_886),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_795),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_798),
.B(n_1007),
.Y(n_1927)
);

INVx3_ASAP7_75t_L g1928 ( 
.A(n_794),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_796),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_796),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_796),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_798),
.B(n_1007),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_798),
.B(n_1007),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_798),
.B(n_1007),
.Y(n_1934)
);

INVxp33_ASAP7_75t_L g1935 ( 
.A(n_1223),
.Y(n_1935)
);

NOR2xp33_ASAP7_75t_L g1936 ( 
.A(n_798),
.B(n_1007),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_798),
.B(n_1007),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_798),
.B(n_1007),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_798),
.B(n_1007),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1244),
.B(n_1246),
.Y(n_1940)
);

OR2x2_ASAP7_75t_L g1941 ( 
.A(n_1617),
.B(n_1721),
.Y(n_1941)
);

AOI221xp5_ASAP7_75t_L g1942 ( 
.A1(n_1262),
.A2(n_1553),
.B1(n_1566),
.B2(n_1550),
.C(n_1546),
.Y(n_1942)
);

NOR2x2_ASAP7_75t_L g1943 ( 
.A(n_1259),
.B(n_1612),
.Y(n_1943)
);

BUFx2_ASAP7_75t_L g1944 ( 
.A(n_1856),
.Y(n_1944)
);

INVxp67_ASAP7_75t_SL g1945 ( 
.A(n_1365),
.Y(n_1945)
);

NOR3x1_ASAP7_75t_L g1946 ( 
.A(n_1555),
.B(n_1561),
.C(n_1593),
.Y(n_1946)
);

AOI22xp33_ASAP7_75t_L g1947 ( 
.A1(n_1668),
.A2(n_1570),
.B1(n_1586),
.B2(n_1573),
.Y(n_1947)
);

INVx4_ASAP7_75t_L g1948 ( 
.A(n_1248),
.Y(n_1948)
);

NOR3xp33_ASAP7_75t_L g1949 ( 
.A(n_1591),
.B(n_1601),
.C(n_1596),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1272),
.B(n_1279),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1248),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1501),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1613),
.B(n_1618),
.Y(n_1953)
);

NOR2xp33_ASAP7_75t_L g1954 ( 
.A(n_1628),
.B(n_1643),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1645),
.B(n_1654),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1318),
.B(n_1296),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_SL g1957 ( 
.A(n_1399),
.B(n_1630),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1673),
.A2(n_1726),
.B1(n_1744),
.B2(n_1696),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1746),
.B(n_1753),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1782),
.B(n_1813),
.Y(n_1960)
);

OAI22xp33_ASAP7_75t_L g1961 ( 
.A1(n_1245),
.A2(n_1253),
.B1(n_1551),
.B2(n_1254),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1825),
.B(n_1837),
.Y(n_1962)
);

AO22x1_ASAP7_75t_L g1963 ( 
.A1(n_1845),
.A2(n_1849),
.B1(n_1904),
.B2(n_1897),
.Y(n_1963)
);

BUFx6f_ASAP7_75t_L g1964 ( 
.A(n_1258),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1488),
.B(n_1515),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1249),
.B(n_1243),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1505),
.Y(n_1967)
);

O2A1O1Ixp5_ASAP7_75t_L g1968 ( 
.A1(n_1257),
.A2(n_1274),
.B(n_1256),
.C(n_1648),
.Y(n_1968)
);

AOI22xp33_ASAP7_75t_L g1969 ( 
.A1(n_1910),
.A2(n_1923),
.B1(n_1932),
.B2(n_1911),
.Y(n_1969)
);

OAI22xp5_ASAP7_75t_L g1970 ( 
.A1(n_1934),
.A2(n_1936),
.B1(n_1559),
.B2(n_1564),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1263),
.B(n_1610),
.Y(n_1971)
);

A2O1A1Ixp33_ASAP7_75t_L g1972 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1568),
.C(n_1557),
.Y(n_1972)
);

INVx2_ASAP7_75t_L g1973 ( 
.A(n_1250),
.Y(n_1973)
);

NAND2xp33_ASAP7_75t_L g1974 ( 
.A(n_1294),
.B(n_1285),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1585),
.B(n_1588),
.Y(n_1975)
);

NOR2xp33_ASAP7_75t_L g1976 ( 
.A(n_1927),
.B(n_1933),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1937),
.B(n_1938),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1594),
.B(n_1595),
.Y(n_1978)
);

CKINVDCx5p33_ASAP7_75t_R g1979 ( 
.A(n_1684),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1598),
.B(n_1599),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1602),
.B(n_1604),
.Y(n_1981)
);

OR2x6_ASAP7_75t_L g1982 ( 
.A(n_1442),
.B(n_1876),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1939),
.B(n_1605),
.Y(n_1983)
);

OR2x2_ASAP7_75t_L g1984 ( 
.A(n_1289),
.B(n_1290),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1743),
.B(n_1755),
.Y(n_1985)
);

INVx3_ASAP7_75t_L g1986 ( 
.A(n_1747),
.Y(n_1986)
);

OR2x6_ASAP7_75t_L g1987 ( 
.A(n_1442),
.B(n_1876),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1258),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1624),
.B(n_1632),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1269),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1493),
.B(n_1459),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1646),
.B(n_1651),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1660),
.B(n_1663),
.Y(n_1993)
);

OR2x6_ASAP7_75t_L g1994 ( 
.A(n_1889),
.B(n_1259),
.Y(n_1994)
);

NOR2xp33_ASAP7_75t_L g1995 ( 
.A(n_1919),
.B(n_1922),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1281),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1295),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1665),
.B(n_1666),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1352),
.A2(n_1355),
.B(n_1354),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1667),
.B(n_1676),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1680),
.B(n_1687),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1298),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1255),
.A2(n_1698),
.B1(n_1702),
.B2(n_1694),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1878),
.B(n_1349),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1704),
.B(n_1710),
.Y(n_2005)
);

AOI22xp33_ASAP7_75t_L g2006 ( 
.A1(n_1725),
.A2(n_1842),
.B1(n_1715),
.B2(n_1717),
.Y(n_2006)
);

NAND2x1_ASAP7_75t_L g2007 ( 
.A(n_1495),
.B(n_1441),
.Y(n_2007)
);

INVxp67_ASAP7_75t_L g2008 ( 
.A(n_1336),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1305),
.Y(n_2009)
);

OAI22xp5_ASAP7_75t_L g2010 ( 
.A1(n_1713),
.A2(n_1718),
.B1(n_1728),
.B2(n_1722),
.Y(n_2010)
);

INVxp67_ASAP7_75t_SL g2011 ( 
.A(n_1615),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1554),
.B(n_1569),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1737),
.B(n_1745),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1749),
.B(n_1750),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1751),
.B(n_1754),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1760),
.B(n_1761),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1327),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1763),
.A2(n_1772),
.B1(n_1778),
.B2(n_1770),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1579),
.B(n_1580),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1780),
.B(n_1787),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_SL g2021 ( 
.A1(n_1769),
.A2(n_1790),
.B1(n_1802),
.B2(n_1791),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_R g2022 ( 
.A(n_1807),
.B(n_1855),
.Y(n_2022)
);

NAND2x1_ASAP7_75t_L g2023 ( 
.A(n_1261),
.B(n_1264),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1810),
.B(n_1829),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1831),
.B(n_1832),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1330),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1242),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1341),
.Y(n_2028)
);

A2O1A1Ixp33_ASAP7_75t_L g2029 ( 
.A1(n_1836),
.A2(n_1843),
.B(n_1844),
.C(n_1838),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1345),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1852),
.A2(n_1868),
.B1(n_1870),
.B2(n_1863),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1347),
.B(n_1299),
.Y(n_2032)
);

INVx3_ASAP7_75t_L g2033 ( 
.A(n_1242),
.Y(n_2033)
);

NOR2xp67_ASAP7_75t_L g2034 ( 
.A(n_1483),
.B(n_1597),
.Y(n_2034)
);

NAND2x1_ASAP7_75t_L g2035 ( 
.A(n_1266),
.B(n_1267),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1871),
.B(n_1873),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1348),
.Y(n_2037)
);

O2A1O1Ixp33_ASAP7_75t_L g2038 ( 
.A1(n_1881),
.A2(n_1890),
.B(n_1891),
.C(n_1887),
.Y(n_2038)
);

AND2x6_ASAP7_75t_L g2039 ( 
.A(n_1309),
.B(n_1487),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1892),
.B(n_1893),
.Y(n_2040)
);

O2A1O1Ixp5_ASAP7_75t_L g2041 ( 
.A1(n_1251),
.A2(n_1544),
.B(n_1578),
.C(n_1545),
.Y(n_2041)
);

AOI22xp33_ASAP7_75t_L g2042 ( 
.A1(n_1895),
.A2(n_1899),
.B1(n_1900),
.B2(n_1896),
.Y(n_2042)
);

AOI22xp33_ASAP7_75t_L g2043 ( 
.A1(n_1905),
.A2(n_1912),
.B1(n_1907),
.B2(n_1581),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1319),
.B(n_1619),
.Y(n_2044)
);

OR2x2_ASAP7_75t_L g2045 ( 
.A(n_1291),
.B(n_1287),
.Y(n_2045)
);

NOR2x1p5_ASAP7_75t_L g2046 ( 
.A(n_1445),
.B(n_1385),
.Y(n_2046)
);

OAI21xp5_ASAP7_75t_L g2047 ( 
.A1(n_1901),
.A2(n_1600),
.B(n_1587),
.Y(n_2047)
);

BUFx6f_ASAP7_75t_L g2048 ( 
.A(n_1258),
.Y(n_2048)
);

HB1xp67_ASAP7_75t_L g2049 ( 
.A(n_1656),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1380),
.Y(n_2050)
);

INVx2_ASAP7_75t_L g2051 ( 
.A(n_1382),
.Y(n_2051)
);

INVxp67_ASAP7_75t_L g2052 ( 
.A(n_1304),
.Y(n_2052)
);

AOI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_1527),
.A2(n_1278),
.B(n_1276),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_SL g2054 ( 
.A(n_1633),
.B(n_1712),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1590),
.B(n_1607),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1386),
.Y(n_2056)
);

CKINVDCx20_ASAP7_75t_R g2057 ( 
.A(n_1364),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1636),
.B(n_1639),
.Y(n_2058)
);

AND2x4_ASAP7_75t_L g2059 ( 
.A(n_1493),
.B(n_1430),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_1359),
.B(n_1368),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_1483),
.B(n_1506),
.Y(n_2061)
);

OAI22xp33_ASAP7_75t_L g2062 ( 
.A1(n_1358),
.A2(n_1360),
.B1(n_1367),
.B2(n_1362),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1411),
.Y(n_2063)
);

INVx5_ASAP7_75t_L g2064 ( 
.A(n_1612),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1767),
.B(n_1781),
.Y(n_2065)
);

NOR2xp67_ASAP7_75t_L g2066 ( 
.A(n_1483),
.B(n_1344),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1640),
.B(n_1641),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1672),
.B(n_1675),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1679),
.B(n_1693),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1565),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1723),
.B(n_1768),
.Y(n_2071)
);

AOI22x1_ASAP7_75t_L g2072 ( 
.A1(n_1417),
.A2(n_1440),
.B1(n_1449),
.B2(n_1427),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1616),
.Y(n_2073)
);

INVxp67_ASAP7_75t_L g2074 ( 
.A(n_1685),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1783),
.B(n_1788),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_SL g2076 ( 
.A(n_1826),
.B(n_1827),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1798),
.B(n_1823),
.Y(n_2077)
);

AO22x1_ASAP7_75t_L g2078 ( 
.A1(n_1730),
.A2(n_1739),
.B1(n_1357),
.B2(n_1297),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1894),
.B(n_1402),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1857),
.B(n_1915),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1622),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1302),
.A2(n_1308),
.B(n_1303),
.Y(n_2082)
);

OR2x6_ASAP7_75t_L g2083 ( 
.A(n_1889),
.B(n_1340),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_1450),
.B(n_1325),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_1623),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_1606),
.A2(n_1608),
.B1(n_1621),
.B2(n_1609),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1322),
.B(n_1311),
.Y(n_2087)
);

OR2x6_ASAP7_75t_L g2088 ( 
.A(n_1350),
.B(n_1534),
.Y(n_2088)
);

NOR3xp33_ASAP7_75t_L g2089 ( 
.A(n_1661),
.B(n_1293),
.C(n_1390),
.Y(n_2089)
);

NOR2x1_ASAP7_75t_R g2090 ( 
.A(n_1460),
.B(n_1543),
.Y(n_2090)
);

NOR2xp33_ASAP7_75t_SL g2091 ( 
.A(n_1653),
.B(n_1392),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1317),
.B(n_1314),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1629),
.B(n_1631),
.Y(n_2093)
);

NOR2xp67_ASAP7_75t_L g2094 ( 
.A(n_1403),
.B(n_1420),
.Y(n_2094)
);

BUFx12f_ASAP7_75t_L g2095 ( 
.A(n_1742),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1356),
.B(n_1372),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1642),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_1662),
.B(n_1674),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1652),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1683),
.B(n_1691),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1699),
.B(n_1706),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_L g2102 ( 
.A(n_1384),
.B(n_1727),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1729),
.B(n_1733),
.Y(n_2103)
);

INVx2_ASAP7_75t_L g2104 ( 
.A(n_1671),
.Y(n_2104)
);

OAI21xp33_ASAP7_75t_L g2105 ( 
.A1(n_1916),
.A2(n_1935),
.B(n_1394),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1735),
.B(n_1736),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_1748),
.B(n_1779),
.Y(n_2107)
);

NOR2xp67_ASAP7_75t_L g2108 ( 
.A(n_1525),
.B(n_1533),
.Y(n_2108)
);

NOR2x2_ASAP7_75t_L g2109 ( 
.A(n_1510),
.B(n_1511),
.Y(n_2109)
);

AND2x4_ASAP7_75t_L g2110 ( 
.A(n_1414),
.B(n_1418),
.Y(n_2110)
);

BUFx2_ASAP7_75t_L g2111 ( 
.A(n_1265),
.Y(n_2111)
);

AOI221xp5_ASAP7_75t_L g2112 ( 
.A1(n_1784),
.A2(n_1815),
.B1(n_1839),
.B2(n_1835),
.C(n_1834),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1853),
.B(n_1854),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1858),
.B(n_1865),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_SL g2115 ( 
.A(n_1307),
.B(n_1252),
.Y(n_2115)
);

OAI22x1_ASAP7_75t_SL g2116 ( 
.A1(n_1537),
.A2(n_1542),
.B1(n_1562),
.B2(n_1300),
.Y(n_2116)
);

BUFx6f_ASAP7_75t_L g2117 ( 
.A(n_1474),
.Y(n_2117)
);

AOI22xp33_ASAP7_75t_L g2118 ( 
.A1(n_1867),
.A2(n_1880),
.B1(n_1906),
.B2(n_1879),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1909),
.B(n_1913),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_SL g2120 ( 
.A(n_1343),
.B(n_1560),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1828),
.B(n_1331),
.Y(n_2121)
);

AOI22xp33_ASAP7_75t_L g2122 ( 
.A1(n_1366),
.A2(n_1422),
.B1(n_1439),
.B2(n_1688),
.Y(n_2122)
);

AND2x4_ASAP7_75t_L g2123 ( 
.A(n_1346),
.B(n_1363),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1455),
.B(n_1471),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_1369),
.B(n_1370),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1692),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1535),
.B(n_1321),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_SL g2128 ( 
.A(n_1331),
.B(n_1332),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_L g2129 ( 
.A(n_1371),
.B(n_1377),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1709),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1711),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1714),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_1378),
.B(n_1379),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_1381),
.B(n_1387),
.Y(n_2134)
);

OR2x2_ASAP7_75t_L g2135 ( 
.A(n_1757),
.B(n_1334),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_1388),
.B(n_1389),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_1724),
.Y(n_2137)
);

OAI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_1438),
.A2(n_1528),
.B(n_1415),
.Y(n_2138)
);

NOR2x2_ASAP7_75t_L g2139 ( 
.A(n_1268),
.B(n_1270),
.Y(n_2139)
);

NOR2xp33_ASAP7_75t_L g2140 ( 
.A(n_1342),
.B(n_1286),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_1265),
.Y(n_2141)
);

HB1xp67_ASAP7_75t_L g2142 ( 
.A(n_1429),
.Y(n_2142)
);

NAND2x1p5_ASAP7_75t_L g2143 ( 
.A(n_1361),
.B(n_1423),
.Y(n_2143)
);

AOI22xp5_ASAP7_75t_L g2144 ( 
.A1(n_1410),
.A2(n_1288),
.B1(n_1478),
.B2(n_1490),
.Y(n_2144)
);

NOR2xp33_ASAP7_75t_L g2145 ( 
.A(n_1567),
.B(n_1626),
.Y(n_2145)
);

AOI22xp33_ASAP7_75t_L g2146 ( 
.A1(n_1731),
.A2(n_1734),
.B1(n_1738),
.B2(n_1732),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1391),
.B(n_1398),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1758),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1400),
.B(n_1405),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1759),
.Y(n_2150)
);

INVx2_ASAP7_75t_SL g2151 ( 
.A(n_1644),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_1407),
.B(n_1408),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1762),
.B(n_1771),
.Y(n_2153)
);

AOI221xp5_ASAP7_75t_L g2154 ( 
.A1(n_1773),
.A2(n_1777),
.B1(n_1792),
.B2(n_1776),
.C(n_1775),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_1395),
.B(n_1658),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1756),
.B(n_1820),
.Y(n_2156)
);

AND2x2_ASAP7_75t_L g2157 ( 
.A(n_1451),
.B(n_1271),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_1872),
.B(n_1448),
.Y(n_2158)
);

BUFx3_ASAP7_75t_L g2159 ( 
.A(n_1644),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1799),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_L g2161 ( 
.A(n_1803),
.B(n_1804),
.Y(n_2161)
);

NOR2xp67_ASAP7_75t_SL g2162 ( 
.A(n_1634),
.B(n_1657),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1806),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1808),
.Y(n_2164)
);

INVxp67_ASAP7_75t_SL g2165 ( 
.A(n_1437),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1809),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1818),
.B(n_1830),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_1847),
.B(n_1848),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1375),
.B(n_1397),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1851),
.B(n_1859),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1861),
.B(n_1877),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_1883),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_1331),
.B(n_1332),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1884),
.B(n_1885),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_SL g2175 ( 
.A(n_1331),
.B(n_1332),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1898),
.B(n_1917),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1920),
.B(n_1926),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_1376),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1273),
.B(n_1275),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1479),
.Y(n_2180)
);

INVxp67_ASAP7_75t_L g2181 ( 
.A(n_1524),
.Y(n_2181)
);

AND2x6_ASAP7_75t_SL g2182 ( 
.A(n_1541),
.B(n_1540),
.Y(n_2182)
);

CKINVDCx5p33_ASAP7_75t_R g2183 ( 
.A(n_1549),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1284),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1292),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1332),
.B(n_1353),
.Y(n_2186)
);

OAI22xp5_ASAP7_75t_SL g2187 ( 
.A1(n_1882),
.A2(n_1531),
.B1(n_1526),
.B2(n_1530),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_1306),
.Y(n_2188)
);

AO22x1_ASAP7_75t_L g2189 ( 
.A1(n_1650),
.A2(n_1720),
.B1(n_1436),
.B2(n_1458),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1312),
.B(n_1313),
.Y(n_2190)
);

OAI21xp5_ASAP7_75t_L g2191 ( 
.A1(n_1473),
.A2(n_1421),
.B(n_1419),
.Y(n_2191)
);

AND2x2_ASAP7_75t_SL g2192 ( 
.A(n_1339),
.B(n_1416),
.Y(n_2192)
);

OR2x6_ASAP7_75t_L g2193 ( 
.A(n_1529),
.B(n_1650),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_SL g2194 ( 
.A(n_1353),
.B(n_1323),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_R g2195 ( 
.A(n_1494),
.B(n_1466),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1315),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_1404),
.B(n_1316),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_SL g2198 ( 
.A(n_1353),
.B(n_1328),
.Y(n_2198)
);

NOR2x2_ASAP7_75t_L g2199 ( 
.A(n_1324),
.B(n_1326),
.Y(n_2199)
);

AOI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_1572),
.A2(n_1833),
.B1(n_1841),
.B2(n_1766),
.Y(n_2200)
);

BUFx6f_ASAP7_75t_L g2201 ( 
.A(n_1474),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1329),
.Y(n_2202)
);

AOI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_1869),
.A2(n_1874),
.B1(n_1463),
.B2(n_1373),
.Y(n_2203)
);

AOI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_1485),
.A2(n_1523),
.B1(n_1930),
.B2(n_1929),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1335),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1338),
.B(n_1351),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_1556),
.A2(n_1574),
.B1(n_1924),
.B2(n_1918),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1563),
.B(n_1575),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_1584),
.A2(n_1931),
.B1(n_1814),
.B2(n_1812),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1589),
.Y(n_2210)
);

BUFx4f_ASAP7_75t_L g2211 ( 
.A(n_1720),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_1603),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1480),
.Y(n_2213)
);

INVx5_ASAP7_75t_L g2214 ( 
.A(n_1474),
.Y(n_2214)
);

BUFx3_ASAP7_75t_L g2215 ( 
.A(n_1774),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_1611),
.B(n_1614),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_SL g2217 ( 
.A(n_1577),
.B(n_1655),
.Y(n_2217)
);

OAI22xp5_ASAP7_75t_SL g2218 ( 
.A1(n_1489),
.A2(n_1508),
.B1(n_1491),
.B2(n_1514),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_SL g2219 ( 
.A(n_1353),
.B(n_1333),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_1620),
.B(n_1635),
.Y(n_2220)
);

NOR3xp33_ASAP7_75t_L g2221 ( 
.A(n_1456),
.B(n_1462),
.C(n_1538),
.Y(n_2221)
);

OR2x6_ASAP7_75t_L g2222 ( 
.A(n_1862),
.B(n_1866),
.Y(n_2222)
);

NAND2xp5_ASAP7_75t_L g2223 ( 
.A(n_1637),
.B(n_1638),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_1512),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1481),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1484),
.Y(n_2226)
);

NAND3xp33_ASAP7_75t_SL g2227 ( 
.A(n_1536),
.B(n_1486),
.C(n_1539),
.Y(n_2227)
);

CKINVDCx5p33_ASAP7_75t_R g2228 ( 
.A(n_1719),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_1512),
.Y(n_2229)
);

O2A1O1Ixp5_ASAP7_75t_L g2230 ( 
.A1(n_1532),
.A2(n_1482),
.B(n_1476),
.C(n_1496),
.Y(n_2230)
);

INVx5_ASAP7_75t_L g2231 ( 
.A(n_1512),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_1649),
.B(n_1659),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_1669),
.A2(n_1817),
.B1(n_1819),
.B2(n_1822),
.Y(n_2233)
);

NOR2xp33_ASAP7_75t_L g2234 ( 
.A(n_1670),
.B(n_1677),
.Y(n_2234)
);

NAND2xp5_ASAP7_75t_SL g2235 ( 
.A(n_1558),
.B(n_1647),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1681),
.B(n_1689),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1695),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_SL g2238 ( 
.A(n_1558),
.B(n_1647),
.Y(n_2238)
);

NAND3xp33_ASAP7_75t_L g2239 ( 
.A(n_1453),
.B(n_1454),
.C(n_1472),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_1705),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1260),
.B(n_1301),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1707),
.Y(n_2242)
);

NOR2x1p5_ASAP7_75t_L g2243 ( 
.A(n_1886),
.B(n_1282),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1716),
.B(n_1752),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_1764),
.B(n_1765),
.Y(n_2245)
);

OAI22xp5_ASAP7_75t_SL g2246 ( 
.A1(n_1446),
.A2(n_1516),
.B1(n_1517),
.B2(n_1860),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1789),
.B(n_1793),
.Y(n_2247)
);

NOR2xp33_ASAP7_75t_L g2248 ( 
.A(n_1795),
.B(n_1805),
.Y(n_2248)
);

BUFx12f_ASAP7_75t_L g2249 ( 
.A(n_1548),
.Y(n_2249)
);

AOI22xp33_ASAP7_75t_L g2250 ( 
.A1(n_1824),
.A2(n_1864),
.B1(n_1846),
.B2(n_1875),
.Y(n_2250)
);

AND2x2_ASAP7_75t_L g2251 ( 
.A(n_1908),
.B(n_1914),
.Y(n_2251)
);

NAND2x1p5_ASAP7_75t_L g2252 ( 
.A(n_1425),
.B(n_1558),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_SL g2253 ( 
.A(n_1260),
.B(n_1301),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_L g2254 ( 
.A1(n_1433),
.A2(n_1452),
.B1(n_1468),
.B2(n_1467),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_1434),
.B(n_1443),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1447),
.B(n_1457),
.Y(n_2256)
);

NOR2xp33_ASAP7_75t_L g2257 ( 
.A(n_1465),
.B(n_1470),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1374),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1426),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_1431),
.Y(n_2260)
);

AND2x2_ASAP7_75t_L g2261 ( 
.A(n_1383),
.B(n_1396),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_1401),
.B(n_1406),
.Y(n_2262)
);

NAND3xp33_ASAP7_75t_SL g2263 ( 
.A(n_1444),
.B(n_1475),
.C(n_1464),
.Y(n_2263)
);

NAND2x1_ASAP7_75t_L g2264 ( 
.A(n_1409),
.B(n_1413),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_SL g2265 ( 
.A(n_1260),
.B(n_1301),
.Y(n_2265)
);

OAI22xp33_ASAP7_75t_L g2266 ( 
.A1(n_1492),
.A2(n_1469),
.B1(n_1497),
.B2(n_1424),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_L g2267 ( 
.A(n_1432),
.B(n_1521),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_1393),
.B(n_1412),
.Y(n_2268)
);

OAI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_1498),
.A2(n_1502),
.B1(n_1507),
.B2(n_1519),
.Y(n_2269)
);

NAND2x1p5_ASAP7_75t_L g2270 ( 
.A(n_1647),
.B(n_1708),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1521),
.B(n_1500),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_1521),
.B(n_1435),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_1260),
.B(n_1301),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_L g2274 ( 
.A(n_1521),
.B(n_1518),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1552),
.B(n_1785),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_1428),
.B(n_1509),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1582),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_1625),
.A2(n_1697),
.B1(n_1627),
.B2(n_1903),
.Y(n_2278)
);

AOI22xp5_ASAP7_75t_L g2279 ( 
.A1(n_1703),
.A2(n_1794),
.B1(n_1797),
.B2(n_1461),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_1921),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_SL g2281 ( 
.A(n_1520),
.B(n_1925),
.C(n_1513),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_1708),
.B(n_1741),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1708),
.B(n_1741),
.Y(n_2283)
);

BUFx3_ASAP7_75t_L g2284 ( 
.A(n_1499),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_1552),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_1921),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1552),
.Y(n_2287)
);

BUFx3_ASAP7_75t_L g2288 ( 
.A(n_1548),
.Y(n_2288)
);

AND3x1_ASAP7_75t_L g2289 ( 
.A(n_1277),
.B(n_1310),
.C(n_1902),
.Y(n_2289)
);

AND2x6_ASAP7_75t_SL g2290 ( 
.A(n_1522),
.B(n_1320),
.Y(n_2290)
);

NOR2xp33_ASAP7_75t_L g2291 ( 
.A(n_1850),
.B(n_1888),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1552),
.Y(n_2292)
);

NOR2xp33_ASAP7_75t_R g2293 ( 
.A(n_1477),
.B(n_1928),
.Y(n_2293)
);

NOR2xp33_ASAP7_75t_L g2294 ( 
.A(n_1850),
.B(n_1888),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1741),
.B(n_1840),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_1800),
.B(n_1840),
.Y(n_2296)
);

AOI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_1504),
.A2(n_1786),
.B1(n_1796),
.B2(n_1503),
.Y(n_2297)
);

INVx5_ASAP7_75t_L g2298 ( 
.A(n_1800),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1664),
.Y(n_2299)
);

INVx3_ASAP7_75t_L g2300 ( 
.A(n_1664),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1664),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1800),
.B(n_1840),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_1811),
.A2(n_1821),
.B1(n_1816),
.B2(n_1571),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_1811),
.B(n_1821),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_1664),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_1811),
.B(n_1821),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1816),
.B(n_1785),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_1816),
.B(n_1785),
.Y(n_2308)
);

NOR2xp33_ASAP7_75t_L g2309 ( 
.A(n_1337),
.B(n_1547),
.Y(n_2309)
);

AOI22xp33_ASAP7_75t_L g2310 ( 
.A1(n_1785),
.A2(n_1801),
.B1(n_1583),
.B2(n_1592),
.Y(n_2310)
);

NAND2xp5_ASAP7_75t_SL g2311 ( 
.A(n_1576),
.B(n_1678),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1682),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_1700),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1686),
.Y(n_2314)
);

INVx2_ASAP7_75t_SL g2315 ( 
.A(n_1690),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_1701),
.B(n_1740),
.Y(n_2316)
);

OAI221xp5_ASAP7_75t_L g2317 ( 
.A1(n_1553),
.A2(n_1075),
.B1(n_1014),
.B2(n_1004),
.C(n_1244),
.Y(n_2317)
);

NOR3xp33_ASAP7_75t_L g2318 ( 
.A(n_1668),
.B(n_1014),
.C(n_1004),
.Y(n_2318)
);

AND3x1_ASAP7_75t_L g2319 ( 
.A(n_1478),
.B(n_888),
.C(n_1244),
.Y(n_2319)
);

INVx1_ASAP7_75t_L g2320 ( 
.A(n_1247),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1247),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2322)
);

NOR2xp33_ASAP7_75t_L g2323 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1501),
.Y(n_2324)
);

NAND2xp5_ASAP7_75t_L g2325 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2325)
);

AND2x2_ASAP7_75t_L g2326 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1247),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2330)
);

NAND3xp33_ASAP7_75t_L g2331 ( 
.A(n_1244),
.B(n_1014),
.C(n_1004),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1247),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1247),
.Y(n_2333)
);

AND2x2_ASAP7_75t_L g2334 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2336)
);

INVx2_ASAP7_75t_SL g2337 ( 
.A(n_1248),
.Y(n_2337)
);

AND2x6_ASAP7_75t_SL g2338 ( 
.A(n_1541),
.B(n_1525),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_1501),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2340)
);

INVx1_ASAP7_75t_L g2341 ( 
.A(n_1247),
.Y(n_2341)
);

OR2x6_ASAP7_75t_L g2342 ( 
.A(n_1442),
.B(n_1094),
.Y(n_2342)
);

INVx2_ASAP7_75t_SL g2343 ( 
.A(n_1248),
.Y(n_2343)
);

OR2x6_ASAP7_75t_L g2344 ( 
.A(n_1442),
.B(n_1094),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1501),
.Y(n_2347)
);

BUFx5_ASAP7_75t_L g2348 ( 
.A(n_1532),
.Y(n_2348)
);

AND2x2_ASAP7_75t_L g2349 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2350)
);

BUFx5_ASAP7_75t_L g2351 ( 
.A(n_1532),
.Y(n_2351)
);

AOI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_SL g2353 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_L g2354 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1247),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2356)
);

NOR2x1p5_ASAP7_75t_L g2357 ( 
.A(n_1399),
.B(n_401),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_1501),
.Y(n_2359)
);

NAND2xp33_ASAP7_75t_L g2360 ( 
.A(n_1630),
.B(n_1648),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2361)
);

A2O1A1Ixp33_ASAP7_75t_L g2362 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1546),
.C(n_1246),
.Y(n_2362)
);

NOR2xp33_ASAP7_75t_L g2363 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2364)
);

OR2x6_ASAP7_75t_L g2365 ( 
.A(n_1442),
.B(n_1094),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1247),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_R g2370 ( 
.A(n_1684),
.B(n_572),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2371)
);

AO22x1_ASAP7_75t_L g2372 ( 
.A1(n_1244),
.A2(n_1262),
.B1(n_1546),
.B2(n_1246),
.Y(n_2372)
);

OAI22xp5_ASAP7_75t_L g2373 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2373)
);

NOR2xp33_ASAP7_75t_L g2374 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_SL g2375 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2375)
);

AOI22xp5_ASAP7_75t_L g2376 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2376)
);

NAND2x1p5_ASAP7_75t_L g2377 ( 
.A(n_1747),
.B(n_1483),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_1501),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2382)
);

AOI22xp5_ASAP7_75t_L g2383 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_1247),
.Y(n_2385)
);

AO22x1_ASAP7_75t_L g2386 ( 
.A1(n_1244),
.A2(n_1262),
.B1(n_1546),
.B2(n_1246),
.Y(n_2386)
);

OAI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_1668),
.A2(n_1245),
.B1(n_1254),
.B2(n_1253),
.Y(n_2387)
);

AOI22xp5_ASAP7_75t_L g2388 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_1247),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_1501),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1501),
.Y(n_2391)
);

OAI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2393)
);

INVx8_ASAP7_75t_L g2394 ( 
.A(n_1876),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_L g2395 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_L g2396 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2396)
);

AOI21xp5_ASAP7_75t_L g2397 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_1247),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_1247),
.Y(n_2400)
);

BUFx3_ASAP7_75t_L g2401 ( 
.A(n_1876),
.Y(n_2401)
);

NAND2xp5_ASAP7_75t_L g2402 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_SL g2403 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2403)
);

AND2x6_ASAP7_75t_SL g2404 ( 
.A(n_1541),
.B(n_1525),
.Y(n_2404)
);

OAI221xp5_ASAP7_75t_L g2405 ( 
.A1(n_1553),
.A2(n_1075),
.B1(n_1014),
.B2(n_1004),
.C(n_1244),
.Y(n_2405)
);

OR2x2_ASAP7_75t_L g2406 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2407)
);

INVx2_ASAP7_75t_SL g2408 ( 
.A(n_1248),
.Y(n_2408)
);

AOI22xp33_ASAP7_75t_L g2409 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2409)
);

OAI21xp5_ASAP7_75t_L g2410 ( 
.A1(n_1630),
.A2(n_1014),
.B(n_1004),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_SL g2411 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_1501),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2413)
);

AOI22xp33_ASAP7_75t_L g2414 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2415)
);

AND2x6_ASAP7_75t_L g2416 ( 
.A(n_1299),
.B(n_1309),
.Y(n_2416)
);

OAI22xp5_ASAP7_75t_L g2417 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2417)
);

AND2x2_ASAP7_75t_L g2418 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2418)
);

NAND2xp5_ASAP7_75t_L g2419 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2420)
);

NOR3xp33_ASAP7_75t_L g2421 ( 
.A(n_1668),
.B(n_1014),
.C(n_1004),
.Y(n_2421)
);

NAND2xp5_ASAP7_75t_SL g2422 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_1247),
.Y(n_2423)
);

INVx1_ASAP7_75t_L g2424 ( 
.A(n_1247),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_1501),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_1247),
.Y(n_2426)
);

BUFx8_ASAP7_75t_L g2427 ( 
.A(n_1549),
.Y(n_2427)
);

OAI22xp5_ASAP7_75t_L g2428 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2430)
);

A2O1A1Ixp33_ASAP7_75t_L g2431 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1546),
.C(n_1246),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2433)
);

AOI22xp33_ASAP7_75t_L g2434 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_L g2435 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2435)
);

INVx3_ASAP7_75t_L g2436 ( 
.A(n_1747),
.Y(n_2436)
);

NOR2xp33_ASAP7_75t_L g2437 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2438)
);

NAND2xp33_ASAP7_75t_L g2439 ( 
.A(n_1630),
.B(n_1648),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2440)
);

AND2x2_ASAP7_75t_L g2441 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2442)
);

BUFx3_ASAP7_75t_L g2443 ( 
.A(n_1876),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2444)
);

A2O1A1Ixp33_ASAP7_75t_L g2445 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1546),
.C(n_1246),
.Y(n_2445)
);

HB1xp67_ASAP7_75t_L g2446 ( 
.A(n_1615),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2447)
);

INVx1_ASAP7_75t_L g2448 ( 
.A(n_1247),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_1501),
.Y(n_2449)
);

AOI22xp33_ASAP7_75t_L g2450 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2453)
);

OR2x2_ASAP7_75t_L g2454 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_1501),
.Y(n_2455)
);

O2A1O1Ixp5_ASAP7_75t_L g2456 ( 
.A1(n_1257),
.A2(n_1274),
.B(n_1256),
.C(n_1668),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_1258),
.Y(n_2457)
);

AOI22xp33_ASAP7_75t_L g2458 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2459)
);

CKINVDCx5p33_ASAP7_75t_R g2460 ( 
.A(n_1684),
.Y(n_2460)
);

OR2x6_ASAP7_75t_L g2461 ( 
.A(n_1442),
.B(n_1094),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_L g2462 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_1247),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2464)
);

BUFx3_ASAP7_75t_L g2465 ( 
.A(n_1876),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_1501),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_SL g2468 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_1247),
.Y(n_2469)
);

INVxp67_ASAP7_75t_L g2470 ( 
.A(n_1336),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_1247),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2473)
);

NAND2xp5_ASAP7_75t_L g2474 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_1248),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_1247),
.Y(n_2480)
);

INVx2_ASAP7_75t_SL g2481 ( 
.A(n_1248),
.Y(n_2481)
);

AOI21xp5_ASAP7_75t_L g2482 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2484)
);

AND2x2_ASAP7_75t_SL g2485 ( 
.A(n_1296),
.B(n_1244),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_SL g2486 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_1501),
.Y(n_2487)
);

BUFx3_ASAP7_75t_L g2488 ( 
.A(n_1876),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_SL g2489 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2489)
);

AOI22xp33_ASAP7_75t_L g2490 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_1247),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2493)
);

NAND2xp33_ASAP7_75t_L g2494 ( 
.A(n_1630),
.B(n_1648),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_1501),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2498)
);

AND2x6_ASAP7_75t_SL g2499 ( 
.A(n_1541),
.B(n_1525),
.Y(n_2499)
);

NOR2xp33_ASAP7_75t_L g2500 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_1247),
.Y(n_2501)
);

HB1xp67_ASAP7_75t_L g2502 ( 
.A(n_1615),
.Y(n_2502)
);

INVx2_ASAP7_75t_SL g2503 ( 
.A(n_1248),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_1501),
.Y(n_2504)
);

INVx2_ASAP7_75t_SL g2505 ( 
.A(n_1248),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2506)
);

AOI22xp5_ASAP7_75t_L g2507 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2507)
);

INVx5_ASAP7_75t_L g2508 ( 
.A(n_1259),
.Y(n_2508)
);

NAND2xp5_ASAP7_75t_L g2509 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2512)
);

NOR2xp33_ASAP7_75t_L g2513 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2513)
);

OAI22xp5_ASAP7_75t_L g2514 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_L g2515 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2516)
);

AOI22xp33_ASAP7_75t_L g2517 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2517)
);

NOR2xp33_ASAP7_75t_L g2518 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2519)
);

INVx2_ASAP7_75t_SL g2520 ( 
.A(n_1248),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_1247),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_1501),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_SL g2523 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_1247),
.Y(n_2524)
);

AOI22xp33_ASAP7_75t_L g2525 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_1501),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_1247),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_SL g2528 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2528)
);

NAND3xp33_ASAP7_75t_L g2529 ( 
.A(n_1244),
.B(n_1014),
.C(n_1004),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2531)
);

NOR2xp33_ASAP7_75t_L g2532 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_1247),
.Y(n_2533)
);

AND2x2_ASAP7_75t_L g2534 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_SL g2535 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_SL g2537 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_SL g2538 ( 
.A(n_1653),
.B(n_556),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2539)
);

AOI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2540)
);

AOI22xp33_ASAP7_75t_L g2541 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_1501),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_1247),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2544)
);

AND2x2_ASAP7_75t_L g2545 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2545)
);

OR2x2_ASAP7_75t_L g2546 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_SL g2547 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2547)
);

AOI21xp5_ASAP7_75t_L g2548 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_1684),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_1247),
.Y(n_2552)
);

INVx8_ASAP7_75t_L g2553 ( 
.A(n_1876),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_SL g2554 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_SL g2555 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2555)
);

OAI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_1247),
.Y(n_2557)
);

INVx2_ASAP7_75t_SL g2558 ( 
.A(n_1248),
.Y(n_2558)
);

AO22x1_ASAP7_75t_L g2559 ( 
.A1(n_1244),
.A2(n_1262),
.B1(n_1546),
.B2(n_1246),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_L g2560 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2560)
);

CKINVDCx20_ASAP7_75t_R g2561 ( 
.A(n_1364),
.Y(n_2561)
);

OAI22xp5_ASAP7_75t_L g2562 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2563)
);

NOR2xp33_ASAP7_75t_L g2564 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2564)
);

NOR2x1_ASAP7_75t_L g2565 ( 
.A(n_1288),
.B(n_405),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2566)
);

AND2x2_ASAP7_75t_L g2567 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_1247),
.Y(n_2569)
);

NOR2x1p5_ASAP7_75t_L g2570 ( 
.A(n_1399),
.B(n_401),
.Y(n_2570)
);

AOI22xp33_ASAP7_75t_L g2571 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_1247),
.Y(n_2572)
);

BUFx2_ASAP7_75t_L g2573 ( 
.A(n_1856),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2574)
);

NAND2xp5_ASAP7_75t_L g2575 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2576)
);

NAND2x1p5_ASAP7_75t_L g2577 ( 
.A(n_1747),
.B(n_1483),
.Y(n_2577)
);

AOI22xp33_ASAP7_75t_SL g2578 ( 
.A1(n_1553),
.A2(n_601),
.B1(n_1246),
.B2(n_1244),
.Y(n_2578)
);

INVx2_ASAP7_75t_SL g2579 ( 
.A(n_1248),
.Y(n_2579)
);

NOR2xp33_ASAP7_75t_L g2580 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2580)
);

NOR2xp33_ASAP7_75t_L g2581 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2581)
);

AOI22xp33_ASAP7_75t_L g2582 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2582)
);

OR2x2_ASAP7_75t_L g2583 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2583)
);

AOI21xp5_ASAP7_75t_L g2584 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_SL g2585 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_1501),
.Y(n_2587)
);

AOI22xp5_ASAP7_75t_L g2588 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2590)
);

AOI21xp5_ASAP7_75t_L g2591 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2592)
);

AND2x4_ASAP7_75t_L g2593 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2593)
);

AND2x2_ASAP7_75t_SL g2594 ( 
.A(n_1296),
.B(n_1244),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2595)
);

INVx2_ASAP7_75t_SL g2596 ( 
.A(n_1248),
.Y(n_2596)
);

AOI21xp5_ASAP7_75t_L g2597 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2597)
);

O2A1O1Ixp5_ASAP7_75t_L g2598 ( 
.A1(n_1257),
.A2(n_1274),
.B(n_1256),
.C(n_1668),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_1501),
.Y(n_2600)
);

HB1xp67_ASAP7_75t_L g2601 ( 
.A(n_1615),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_1501),
.Y(n_2602)
);

INVx2_ASAP7_75t_SL g2603 ( 
.A(n_1248),
.Y(n_2603)
);

AOI22xp33_ASAP7_75t_L g2604 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_1247),
.Y(n_2605)
);

NOR2xp33_ASAP7_75t_L g2606 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2606)
);

NOR2xp67_ASAP7_75t_L g2607 ( 
.A(n_1684),
.B(n_830),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_1876),
.Y(n_2610)
);

OR2x2_ASAP7_75t_L g2611 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2612)
);

AOI22xp33_ASAP7_75t_L g2613 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_1769),
.B(n_402),
.Y(n_2615)
);

BUFx6f_ASAP7_75t_L g2616 ( 
.A(n_1258),
.Y(n_2616)
);

O2A1O1Ixp5_ASAP7_75t_L g2617 ( 
.A1(n_1257),
.A2(n_1274),
.B(n_1256),
.C(n_1668),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_SL g2618 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2618)
);

O2A1O1Ixp33_ASAP7_75t_L g2619 ( 
.A1(n_1630),
.A2(n_1648),
.B(n_1668),
.C(n_1246),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2620)
);

AOI21xp5_ASAP7_75t_L g2621 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2622)
);

AOI222xp33_ASAP7_75t_L g2623 ( 
.A1(n_1244),
.A2(n_1550),
.B1(n_1262),
.B2(n_1553),
.C1(n_1546),
.C2(n_1246),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_1247),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2625)
);

INVx4_ASAP7_75t_L g2626 ( 
.A(n_1248),
.Y(n_2626)
);

INVx2_ASAP7_75t_SL g2627 ( 
.A(n_1248),
.Y(n_2627)
);

A2O1A1Ixp33_ASAP7_75t_L g2628 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1546),
.C(n_1246),
.Y(n_2628)
);

INVxp33_ASAP7_75t_SL g2629 ( 
.A(n_1882),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_L g2631 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2631)
);

NAND2xp33_ASAP7_75t_L g2632 ( 
.A(n_1630),
.B(n_1648),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_L g2634 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_L g2637 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_SL g2638 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2638)
);

AND2x4_ASAP7_75t_L g2639 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2639)
);

INVx4_ASAP7_75t_L g2640 ( 
.A(n_1248),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2641)
);

AOI22xp33_ASAP7_75t_L g2642 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2642)
);

INVxp67_ASAP7_75t_SL g2643 ( 
.A(n_1365),
.Y(n_2643)
);

A2O1A1Ixp33_ASAP7_75t_L g2644 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1546),
.C(n_1246),
.Y(n_2644)
);

INVx2_ASAP7_75t_SL g2645 ( 
.A(n_1248),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_SL g2646 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2646)
);

AOI22xp5_ASAP7_75t_L g2647 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2647)
);

CKINVDCx5p33_ASAP7_75t_R g2648 ( 
.A(n_1684),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2649)
);

BUFx6f_ASAP7_75t_SL g2650 ( 
.A(n_1493),
.Y(n_2650)
);

NOR3xp33_ASAP7_75t_L g2651 ( 
.A(n_1668),
.B(n_1014),
.C(n_1004),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_R g2652 ( 
.A(n_1684),
.B(n_572),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_1501),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_1501),
.Y(n_2654)
);

AOI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2655)
);

OAI22xp5_ASAP7_75t_L g2656 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_SL g2657 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2657)
);

AOI22xp5_ASAP7_75t_L g2658 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2658)
);

INVx3_ASAP7_75t_L g2659 ( 
.A(n_1747),
.Y(n_2659)
);

BUFx8_ASAP7_75t_L g2660 ( 
.A(n_1549),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_L g2661 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2661)
);

NOR2xp33_ASAP7_75t_L g2662 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2663)
);

INVxp67_ASAP7_75t_SL g2664 ( 
.A(n_1365),
.Y(n_2664)
);

AND2x4_ASAP7_75t_L g2665 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2668)
);

NAND2x1_ASAP7_75t_L g2669 ( 
.A(n_1501),
.B(n_818),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2670)
);

INVx3_ASAP7_75t_L g2671 ( 
.A(n_1747),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_1248),
.Y(n_2672)
);

AOI21xp5_ASAP7_75t_L g2673 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2673)
);

AOI22xp33_ASAP7_75t_L g2674 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_SL g2675 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_1501),
.Y(n_2676)
);

AOI22xp33_ASAP7_75t_L g2677 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2677)
);

OR2x2_ASAP7_75t_L g2678 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2678)
);

AOI22xp33_ASAP7_75t_L g2679 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2679)
);

AOI22xp5_ASAP7_75t_L g2680 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_1247),
.Y(n_2681)
);

O2A1O1Ixp33_ASAP7_75t_L g2682 ( 
.A1(n_1630),
.A2(n_1648),
.B(n_1668),
.C(n_1246),
.Y(n_2682)
);

NAND2x1_ASAP7_75t_L g2683 ( 
.A(n_1501),
.B(n_818),
.Y(n_2683)
);

AOI22xp33_ASAP7_75t_L g2684 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2684)
);

AOI221xp5_ASAP7_75t_SL g2685 ( 
.A1(n_1668),
.A2(n_1648),
.B1(n_1630),
.B2(n_1246),
.C(n_1546),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_1247),
.Y(n_2686)
);

NAND2xp5_ASAP7_75t_SL g2687 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_1247),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2690)
);

AND2x2_ASAP7_75t_L g2691 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2691)
);

INVx2_ASAP7_75t_SL g2692 ( 
.A(n_1248),
.Y(n_2692)
);

AOI22xp33_ASAP7_75t_L g2693 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2695)
);

INVx2_ASAP7_75t_L g2696 ( 
.A(n_1501),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2697)
);

NOR2xp33_ASAP7_75t_SL g2698 ( 
.A(n_1653),
.B(n_556),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2699)
);

BUFx3_ASAP7_75t_L g2700 ( 
.A(n_1876),
.Y(n_2700)
);

AOI22xp5_ASAP7_75t_L g2701 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2702)
);

BUFx6f_ASAP7_75t_L g2703 ( 
.A(n_1258),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2704)
);

AND3x1_ASAP7_75t_L g2705 ( 
.A(n_1478),
.B(n_888),
.C(n_1244),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_1247),
.Y(n_2706)
);

A2O1A1Ixp33_ASAP7_75t_L g2707 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1546),
.C(n_1246),
.Y(n_2707)
);

NAND2xp5_ASAP7_75t_L g2708 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2708)
);

CKINVDCx5p33_ASAP7_75t_R g2709 ( 
.A(n_1684),
.Y(n_2709)
);

INVx2_ASAP7_75t_SL g2710 ( 
.A(n_1248),
.Y(n_2710)
);

AND2x6_ASAP7_75t_SL g2711 ( 
.A(n_1541),
.B(n_1525),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_1247),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_SL g2714 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2714)
);

HB1xp67_ASAP7_75t_L g2715 ( 
.A(n_1615),
.Y(n_2715)
);

O2A1O1Ixp5_ASAP7_75t_L g2716 ( 
.A1(n_1257),
.A2(n_1274),
.B(n_1256),
.C(n_1668),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_1501),
.Y(n_2717)
);

NAND2xp5_ASAP7_75t_SL g2718 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2720)
);

NAND2x1_ASAP7_75t_L g2721 ( 
.A(n_1501),
.B(n_818),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_1247),
.Y(n_2723)
);

NAND2xp5_ASAP7_75t_L g2724 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_1247),
.Y(n_2725)
);

NOR2xp33_ASAP7_75t_L g2726 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2726)
);

INVx8_ASAP7_75t_L g2727 ( 
.A(n_1876),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2728)
);

AND2x2_ASAP7_75t_L g2729 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2729)
);

INVx3_ASAP7_75t_L g2730 ( 
.A(n_1747),
.Y(n_2730)
);

AOI21xp5_ASAP7_75t_L g2731 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2733)
);

OR2x2_ASAP7_75t_L g2734 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_SL g2735 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2735)
);

AOI221xp5_ASAP7_75t_L g2736 ( 
.A1(n_1244),
.A2(n_1546),
.B1(n_1550),
.B2(n_1262),
.C(n_1246),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2737)
);

O2A1O1Ixp5_ASAP7_75t_L g2738 ( 
.A1(n_1257),
.A2(n_1274),
.B(n_1256),
.C(n_1668),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_SL g2739 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2740)
);

INVxp67_ASAP7_75t_SL g2741 ( 
.A(n_1365),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2742)
);

AND2x6_ASAP7_75t_SL g2743 ( 
.A(n_1541),
.B(n_1525),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_SL g2744 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2744)
);

AOI22xp33_ASAP7_75t_L g2745 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_L g2746 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_R g2749 ( 
.A(n_1684),
.B(n_572),
.Y(n_2749)
);

O2A1O1Ixp33_ASAP7_75t_L g2750 ( 
.A1(n_1630),
.A2(n_1648),
.B(n_1668),
.C(n_1246),
.Y(n_2750)
);

AOI22xp5_ASAP7_75t_L g2751 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_1247),
.Y(n_2752)
);

INVx2_ASAP7_75t_SL g2753 ( 
.A(n_1248),
.Y(n_2753)
);

OAI22xp33_ASAP7_75t_L g2754 ( 
.A1(n_1668),
.A2(n_1245),
.B1(n_1254),
.B2(n_1253),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2756)
);

INVx2_ASAP7_75t_SL g2757 ( 
.A(n_1248),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_1247),
.Y(n_2761)
);

INVx4_ASAP7_75t_L g2762 ( 
.A(n_1248),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_SL g2765 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2766)
);

AOI22xp5_ASAP7_75t_L g2767 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2768)
);

BUFx4f_ASAP7_75t_L g2769 ( 
.A(n_1442),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_1684),
.Y(n_2770)
);

OR2x2_ASAP7_75t_L g2771 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2772)
);

CKINVDCx5p33_ASAP7_75t_R g2773 ( 
.A(n_1684),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_SL g2774 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2776)
);

AND2x4_ASAP7_75t_L g2777 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2777)
);

NOR2xp67_ASAP7_75t_SL g2778 ( 
.A(n_1483),
.B(n_402),
.Y(n_2778)
);

NAND2xp5_ASAP7_75t_L g2779 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2779)
);

NAND2x1_ASAP7_75t_L g2780 ( 
.A(n_1501),
.B(n_818),
.Y(n_2780)
);

NOR2xp33_ASAP7_75t_L g2781 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2782)
);

BUFx3_ASAP7_75t_L g2783 ( 
.A(n_1876),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2784)
);

NAND2xp5_ASAP7_75t_L g2785 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_1247),
.Y(n_2787)
);

AOI21xp5_ASAP7_75t_L g2788 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2789)
);

INVx2_ASAP7_75t_L g2790 ( 
.A(n_1501),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_1501),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_1501),
.Y(n_2792)
);

OR2x2_ASAP7_75t_L g2793 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_L g2795 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_1247),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2797)
);

NAND2x1p5_ASAP7_75t_L g2798 ( 
.A(n_1747),
.B(n_1483),
.Y(n_2798)
);

AOI22xp5_ASAP7_75t_L g2799 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1247),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_1501),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_1247),
.Y(n_2802)
);

BUFx3_ASAP7_75t_L g2803 ( 
.A(n_1876),
.Y(n_2803)
);

AND2x4_ASAP7_75t_L g2804 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_SL g2806 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_1501),
.Y(n_2807)
);

AOI22xp5_ASAP7_75t_L g2808 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2808)
);

NAND2xp5_ASAP7_75t_L g2809 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_1247),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2812)
);

INVx3_ASAP7_75t_L g2813 ( 
.A(n_1747),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_1247),
.Y(n_2814)
);

AOI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_L g2820 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2820)
);

AOI22xp5_ASAP7_75t_L g2821 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_1501),
.Y(n_2823)
);

NOR2xp33_ASAP7_75t_L g2824 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_1247),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_1247),
.Y(n_2826)
);

OR2x2_ASAP7_75t_L g2827 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2828)
);

AOI22xp5_ASAP7_75t_L g2829 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_1247),
.Y(n_2830)
);

INVx2_ASAP7_75t_L g2831 ( 
.A(n_1501),
.Y(n_2831)
);

NAND2xp5_ASAP7_75t_L g2832 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_1247),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_1247),
.Y(n_2835)
);

OAI21xp33_ASAP7_75t_L g2836 ( 
.A1(n_1244),
.A2(n_1262),
.B(n_1246),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_1247),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_1247),
.Y(n_2838)
);

AOI22xp5_ASAP7_75t_L g2839 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_L g2840 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2840)
);

AOI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_SL g2842 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2842)
);

OR2x2_ASAP7_75t_L g2843 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2843)
);

OAI21xp5_ASAP7_75t_L g2844 ( 
.A1(n_1630),
.A2(n_1014),
.B(n_1004),
.Y(n_2844)
);

NAND2xp5_ASAP7_75t_L g2845 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2845)
);

INVx3_ASAP7_75t_L g2846 ( 
.A(n_1747),
.Y(n_2846)
);

AOI22xp5_ASAP7_75t_L g2847 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2848)
);

BUFx5_ASAP7_75t_L g2849 ( 
.A(n_1532),
.Y(n_2849)
);

AO22x1_ASAP7_75t_L g2850 ( 
.A1(n_1244),
.A2(n_1262),
.B1(n_1546),
.B2(n_1246),
.Y(n_2850)
);

INVxp67_ASAP7_75t_L g2851 ( 
.A(n_1336),
.Y(n_2851)
);

INVx8_ASAP7_75t_L g2852 ( 
.A(n_1876),
.Y(n_2852)
);

A2O1A1Ixp33_ASAP7_75t_SL g2853 ( 
.A1(n_1244),
.A2(n_1007),
.B(n_1010),
.C(n_798),
.Y(n_2853)
);

INVx2_ASAP7_75t_SL g2854 ( 
.A(n_1248),
.Y(n_2854)
);

BUFx6f_ASAP7_75t_L g2855 ( 
.A(n_1258),
.Y(n_2855)
);

INVx2_ASAP7_75t_L g2856 ( 
.A(n_1501),
.Y(n_2856)
);

INVx1_ASAP7_75t_SL g2857 ( 
.A(n_1304),
.Y(n_2857)
);

INVx2_ASAP7_75t_SL g2858 ( 
.A(n_1248),
.Y(n_2858)
);

OR2x2_ASAP7_75t_L g2859 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2859)
);

AOI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2860)
);

NOR2xp33_ASAP7_75t_R g2861 ( 
.A(n_1684),
.B(n_572),
.Y(n_2861)
);

NAND2xp33_ASAP7_75t_L g2862 ( 
.A(n_1630),
.B(n_1648),
.Y(n_2862)
);

BUFx3_ASAP7_75t_L g2863 ( 
.A(n_1876),
.Y(n_2863)
);

OR2x2_ASAP7_75t_L g2864 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_1247),
.Y(n_2865)
);

INVx3_ASAP7_75t_L g2866 ( 
.A(n_1747),
.Y(n_2866)
);

AOI22xp5_ASAP7_75t_L g2867 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2867)
);

BUFx2_ASAP7_75t_L g2868 ( 
.A(n_1856),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_1247),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2870)
);

HB1xp67_ASAP7_75t_L g2871 ( 
.A(n_1615),
.Y(n_2871)
);

CKINVDCx20_ASAP7_75t_R g2872 ( 
.A(n_1364),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_1247),
.Y(n_2873)
);

AOI22xp5_ASAP7_75t_L g2874 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2875)
);

NOR2xp33_ASAP7_75t_L g2876 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_SL g2877 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2877)
);

NAND2x1p5_ASAP7_75t_L g2878 ( 
.A(n_1747),
.B(n_1483),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_SL g2880 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2880)
);

OAI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_1630),
.A2(n_1014),
.B(n_1004),
.Y(n_2881)
);

BUFx2_ASAP7_75t_L g2882 ( 
.A(n_1856),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_1247),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_1501),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_1247),
.Y(n_2886)
);

AOI22xp5_ASAP7_75t_L g2887 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_1247),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_L g2890 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2890)
);

NAND2x1_ASAP7_75t_L g2891 ( 
.A(n_1501),
.B(n_818),
.Y(n_2891)
);

INVx2_ASAP7_75t_SL g2892 ( 
.A(n_1248),
.Y(n_2892)
);

NOR2xp33_ASAP7_75t_L g2893 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_1501),
.Y(n_2895)
);

NOR2xp33_ASAP7_75t_L g2896 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2896)
);

AOI22xp33_ASAP7_75t_L g2897 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2898)
);

NAND2xp33_ASAP7_75t_L g2899 ( 
.A(n_1630),
.B(n_1648),
.Y(n_2899)
);

AOI21xp5_ASAP7_75t_L g2900 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2900)
);

OAI22xp5_ASAP7_75t_L g2901 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2901)
);

AOI22xp5_ASAP7_75t_L g2902 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2902)
);

AND2x6_ASAP7_75t_L g2903 ( 
.A(n_1299),
.B(n_1309),
.Y(n_2903)
);

AOI22xp33_ASAP7_75t_L g2904 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2904)
);

NAND2xp5_ASAP7_75t_L g2905 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2905)
);

BUFx3_ASAP7_75t_L g2906 ( 
.A(n_1876),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_1501),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2908)
);

NAND3xp33_ASAP7_75t_SL g2909 ( 
.A(n_1630),
.B(n_1648),
.C(n_1246),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_L g2910 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2910)
);

NAND2xp5_ASAP7_75t_L g2911 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2911)
);

INVx2_ASAP7_75t_SL g2912 ( 
.A(n_1248),
.Y(n_2912)
);

NAND2xp5_ASAP7_75t_L g2913 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2913)
);

CKINVDCx5p33_ASAP7_75t_R g2914 ( 
.A(n_1684),
.Y(n_2914)
);

INVx2_ASAP7_75t_L g2915 ( 
.A(n_1501),
.Y(n_2915)
);

NOR2xp33_ASAP7_75t_L g2916 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_L g2917 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_1247),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_SL g2919 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2919)
);

BUFx6f_ASAP7_75t_L g2920 ( 
.A(n_1258),
.Y(n_2920)
);

AOI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_1247),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_L g2924 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_1247),
.Y(n_2925)
);

INVx1_ASAP7_75t_L g2926 ( 
.A(n_1247),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2927)
);

BUFx2_ASAP7_75t_L g2928 ( 
.A(n_1856),
.Y(n_2928)
);

OR2x2_ASAP7_75t_L g2929 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2930)
);

INVx2_ASAP7_75t_L g2931 ( 
.A(n_1501),
.Y(n_2931)
);

OR2x2_ASAP7_75t_L g2932 ( 
.A(n_1617),
.B(n_1721),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_L g2933 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_L g2934 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_1247),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_1247),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2940)
);

NAND2xp5_ASAP7_75t_SL g2941 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_1247),
.Y(n_2943)
);

AOI22xp33_ASAP7_75t_SL g2944 ( 
.A1(n_1553),
.A2(n_601),
.B1(n_1246),
.B2(n_1244),
.Y(n_2944)
);

BUFx6f_ASAP7_75t_L g2945 ( 
.A(n_1258),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_SL g2946 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2946)
);

NAND3xp33_ASAP7_75t_L g2947 ( 
.A(n_1244),
.B(n_1014),
.C(n_1004),
.Y(n_2947)
);

OAI221xp5_ASAP7_75t_L g2948 ( 
.A1(n_1553),
.A2(n_1075),
.B1(n_1014),
.B2(n_1004),
.C(n_1244),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2949)
);

INVx2_ASAP7_75t_SL g2950 ( 
.A(n_1248),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_SL g2951 ( 
.A(n_1769),
.B(n_402),
.Y(n_2951)
);

AOI22xp33_ASAP7_75t_L g2952 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2953)
);

AOI22xp5_ASAP7_75t_L g2954 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_1769),
.B(n_402),
.Y(n_2955)
);

AOI21xp5_ASAP7_75t_L g2956 ( 
.A1(n_1274),
.A2(n_842),
.B(n_1352),
.Y(n_2956)
);

NOR2xp67_ASAP7_75t_L g2957 ( 
.A(n_1684),
.B(n_830),
.Y(n_2957)
);

AOI22xp33_ASAP7_75t_L g2958 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_1501),
.Y(n_2959)
);

NAND2xp5_ASAP7_75t_L g2960 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_1247),
.Y(n_2961)
);

NOR2xp33_ASAP7_75t_L g2962 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2962)
);

INVx2_ASAP7_75t_L g2963 ( 
.A(n_1501),
.Y(n_2963)
);

NOR2xp33_ASAP7_75t_L g2964 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2964)
);

OAI21xp5_ASAP7_75t_L g2965 ( 
.A1(n_1630),
.A2(n_1014),
.B(n_1004),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_1247),
.Y(n_2968)
);

BUFx3_ASAP7_75t_L g2969 ( 
.A(n_1876),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2970)
);

INVx2_ASAP7_75t_SL g2971 ( 
.A(n_1248),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2973)
);

NAND3xp33_ASAP7_75t_SL g2974 ( 
.A(n_1630),
.B(n_1648),
.C(n_1246),
.Y(n_2974)
);

AOI22xp33_ASAP7_75t_L g2975 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_L g2976 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_SL g2977 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2977)
);

NOR2xp33_ASAP7_75t_L g2978 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2978)
);

AND2x4_ASAP7_75t_L g2979 ( 
.A(n_1488),
.B(n_1515),
.Y(n_2979)
);

AOI22xp33_ASAP7_75t_L g2980 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2981)
);

NOR2xp33_ASAP7_75t_L g2982 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2983)
);

AOI22xp33_ASAP7_75t_L g2984 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2984)
);

AOI22xp33_ASAP7_75t_L g2985 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_1247),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_1247),
.Y(n_2987)
);

NAND2xp5_ASAP7_75t_L g2988 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2989)
);

AND2x2_ASAP7_75t_L g2990 ( 
.A(n_1249),
.B(n_1243),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_1501),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_L g2993 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_1244),
.B(n_1246),
.Y(n_2994)
);

AOI22xp5_ASAP7_75t_L g2995 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_SL g2997 ( 
.A(n_1318),
.B(n_1296),
.Y(n_2997)
);

INVx2_ASAP7_75t_L g2998 ( 
.A(n_1501),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_1501),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_SL g3000 ( 
.A(n_1318),
.B(n_1296),
.Y(n_3000)
);

AND2x2_ASAP7_75t_L g3001 ( 
.A(n_1249),
.B(n_1243),
.Y(n_3001)
);

AOI22xp5_ASAP7_75t_L g3002 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_1249),
.B(n_1243),
.Y(n_3003)
);

AND2x2_ASAP7_75t_L g3004 ( 
.A(n_1249),
.B(n_1243),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_1501),
.Y(n_3005)
);

AND2x2_ASAP7_75t_SL g3006 ( 
.A(n_1296),
.B(n_1244),
.Y(n_3006)
);

O2A1O1Ixp33_ASAP7_75t_L g3007 ( 
.A1(n_1630),
.A2(n_1648),
.B(n_1668),
.C(n_1246),
.Y(n_3007)
);

NAND2xp5_ASAP7_75t_L g3008 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_1318),
.B(n_1296),
.Y(n_3010)
);

NAND2xp33_ASAP7_75t_L g3011 ( 
.A(n_1630),
.B(n_1648),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_1501),
.Y(n_3012)
);

NAND2xp5_ASAP7_75t_L g3013 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_1501),
.Y(n_3014)
);

NOR3xp33_ASAP7_75t_L g3015 ( 
.A(n_1668),
.B(n_1014),
.C(n_1004),
.Y(n_3015)
);

NAND2xp5_ASAP7_75t_L g3016 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_1247),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_1488),
.B(n_1515),
.Y(n_3018)
);

INVx1_ASAP7_75t_L g3019 ( 
.A(n_1247),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_1247),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_SL g3021 ( 
.A(n_1318),
.B(n_1296),
.Y(n_3021)
);

NOR2xp33_ASAP7_75t_L g3022 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_1318),
.B(n_1296),
.Y(n_3023)
);

OAI22xp33_ASAP7_75t_L g3024 ( 
.A1(n_1668),
.A2(n_1245),
.B1(n_1254),
.B2(n_1253),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_1501),
.Y(n_3025)
);

NOR2xp33_ASAP7_75t_L g3026 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3026)
);

AOI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3028)
);

AND2x6_ASAP7_75t_SL g3029 ( 
.A(n_1541),
.B(n_1525),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_1247),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_1501),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3033)
);

INVx2_ASAP7_75t_L g3034 ( 
.A(n_1501),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_SL g3036 ( 
.A(n_1318),
.B(n_1296),
.Y(n_3036)
);

AND2x2_ASAP7_75t_L g3037 ( 
.A(n_1249),
.B(n_1243),
.Y(n_3037)
);

AOI22xp5_ASAP7_75t_L g3038 ( 
.A1(n_1244),
.A2(n_1246),
.B1(n_1546),
.B2(n_1262),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3039)
);

AOI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3041)
);

BUFx4f_ASAP7_75t_SL g3042 ( 
.A(n_1730),
.Y(n_3042)
);

AOI22xp33_ASAP7_75t_L g3043 ( 
.A1(n_1668),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3043)
);

NAND2xp5_ASAP7_75t_SL g3044 ( 
.A(n_1769),
.B(n_402),
.Y(n_3044)
);

INVx2_ASAP7_75t_SL g3045 ( 
.A(n_1248),
.Y(n_3045)
);

NAND2xp5_ASAP7_75t_L g3046 ( 
.A(n_1244),
.B(n_1246),
.Y(n_3046)
);

NAND2xp5_ASAP7_75t_SL g3047 ( 
.A(n_1318),
.B(n_1296),
.Y(n_3047)
);

AND3x1_ASAP7_75t_L g3048 ( 
.A(n_1478),
.B(n_888),
.C(n_1244),
.Y(n_3048)
);

INVx1_ASAP7_75t_L g3049 ( 
.A(n_1247),
.Y(n_3049)
);

NAND2xp33_ASAP7_75t_L g3050 ( 
.A(n_1949),
.B(n_2370),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2280),
.Y(n_3051)
);

AND2x4_ASAP7_75t_L g3052 ( 
.A(n_2047),
.B(n_2059),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2286),
.Y(n_3053)
);

OAI21xp33_ASAP7_75t_SL g3054 ( 
.A1(n_2112),
.A2(n_2118),
.B(n_2086),
.Y(n_3054)
);

BUFx6f_ASAP7_75t_L g3055 ( 
.A(n_2192),
.Y(n_3055)
);

NAND2xp5_ASAP7_75t_L g3056 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3057)
);

NOR2xp33_ASAP7_75t_L g3058 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_3024),
.B(n_1999),
.Y(n_3059)
);

AOI21xp5_ASAP7_75t_L g3060 ( 
.A1(n_2397),
.A2(n_2540),
.B(n_2482),
.Y(n_3060)
);

OAI321xp33_ASAP7_75t_L g3061 ( 
.A1(n_2373),
.A2(n_2514),
.A3(n_2417),
.B1(n_2556),
.B2(n_2428),
.C(n_2392),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3062)
);

OAI21xp5_ASAP7_75t_L g3063 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_3024),
.B(n_3006),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2348),
.Y(n_3065)
);

AOI21xp5_ASAP7_75t_L g3066 ( 
.A1(n_2548),
.A2(n_2591),
.B(n_2584),
.Y(n_3066)
);

INVx2_ASAP7_75t_L g3067 ( 
.A(n_2348),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3068)
);

OAI22xp5_ASAP7_75t_L g3069 ( 
.A1(n_1947),
.A2(n_2409),
.B1(n_2414),
.B2(n_2352),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_1961),
.B(n_2578),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3071)
);

NOR3xp33_ASAP7_75t_L g3072 ( 
.A(n_1942),
.B(n_2736),
.C(n_2656),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_SL g3073 ( 
.A(n_2944),
.B(n_2060),
.Y(n_3073)
);

HB1xp67_ASAP7_75t_L g3074 ( 
.A(n_2049),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2060),
.B(n_3006),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2348),
.Y(n_3076)
);

AOI21xp5_ASAP7_75t_L g3077 ( 
.A1(n_2597),
.A2(n_2673),
.B(n_2621),
.Y(n_3077)
);

BUFx8_ASAP7_75t_L g3078 ( 
.A(n_2650),
.Y(n_3078)
);

AOI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_1954),
.A2(n_1962),
.B1(n_2336),
.B2(n_2323),
.Y(n_3079)
);

AND2x2_ASAP7_75t_L g3080 ( 
.A(n_2685),
.B(n_2006),
.Y(n_3080)
);

NAND2xp33_ASAP7_75t_L g3081 ( 
.A(n_2370),
.B(n_2652),
.Y(n_3081)
);

BUFx6f_ASAP7_75t_L g3082 ( 
.A(n_2192),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_L g3083 ( 
.A(n_2114),
.B(n_1972),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_1962),
.B(n_2323),
.Y(n_3084)
);

INVx1_ASAP7_75t_SL g3085 ( 
.A(n_2139),
.Y(n_3085)
);

NAND2xp5_ASAP7_75t_SL g3086 ( 
.A(n_2376),
.B(n_2383),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2114),
.B(n_2086),
.Y(n_3087)
);

NOR2xp33_ASAP7_75t_L g3088 ( 
.A(n_2336),
.B(n_2354),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2006),
.B(n_1946),
.Y(n_3089)
);

A2O1A1Ixp33_ASAP7_75t_L g3090 ( 
.A1(n_2619),
.A2(n_2682),
.B(n_3007),
.C(n_2750),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2348),
.Y(n_3091)
);

AND2x2_ASAP7_75t_L g3092 ( 
.A(n_1957),
.B(n_2410),
.Y(n_3092)
);

AOI21xp5_ASAP7_75t_L g3093 ( 
.A1(n_2731),
.A2(n_2900),
.B(n_2788),
.Y(n_3093)
);

OAI21xp5_ASAP7_75t_L g3094 ( 
.A1(n_2617),
.A2(n_2738),
.B(n_2716),
.Y(n_3094)
);

O2A1O1Ixp33_ASAP7_75t_L g3095 ( 
.A1(n_2362),
.A2(n_2445),
.B(n_2628),
.C(n_2431),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2118),
.B(n_1976),
.Y(n_3096)
);

INVx4_ASAP7_75t_L g3097 ( 
.A(n_2214),
.Y(n_3097)
);

NOR2xp33_ASAP7_75t_L g3098 ( 
.A(n_2354),
.B(n_2363),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2348),
.Y(n_3099)
);

CKINVDCx5p33_ASAP7_75t_R g3100 ( 
.A(n_2652),
.Y(n_3100)
);

INVxp67_ASAP7_75t_L g3101 ( 
.A(n_2049),
.Y(n_3101)
);

BUFx3_ASAP7_75t_L g3102 ( 
.A(n_2394),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2348),
.Y(n_3103)
);

AOI22xp5_ASAP7_75t_L g3104 ( 
.A1(n_2363),
.A2(n_2374),
.B1(n_2380),
.B2(n_2371),
.Y(n_3104)
);

A2O1A1Ixp33_ASAP7_75t_L g3105 ( 
.A1(n_2038),
.A2(n_2707),
.B(n_2644),
.C(n_1968),
.Y(n_3105)
);

NOR2x1_ASAP7_75t_R g3106 ( 
.A(n_1979),
.B(n_2460),
.Y(n_3106)
);

A2O1A1Ixp33_ASAP7_75t_L g3107 ( 
.A1(n_2318),
.A2(n_2651),
.B(n_3015),
.C(n_2421),
.Y(n_3107)
);

NAND2xp5_ASAP7_75t_L g3108 ( 
.A(n_1976),
.B(n_1977),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_1977),
.B(n_1983),
.Y(n_3109)
);

NOR3xp33_ASAP7_75t_L g3110 ( 
.A(n_2562),
.B(n_2901),
.C(n_2405),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_1983),
.B(n_1993),
.Y(n_3111)
);

OAI22xp5_ASAP7_75t_L g3112 ( 
.A1(n_1947),
.A2(n_2409),
.B1(n_2414),
.B2(n_2352),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_1993),
.B(n_1995),
.Y(n_3113)
);

AND2x4_ASAP7_75t_L g3114 ( 
.A(n_2059),
.B(n_2287),
.Y(n_3114)
);

O2A1O1Ixp33_ASAP7_75t_L g3115 ( 
.A1(n_2029),
.A2(n_1970),
.B(n_1985),
.C(n_2317),
.Y(n_3115)
);

CKINVDCx5p33_ASAP7_75t_R g3116 ( 
.A(n_2749),
.Y(n_3116)
);

OAI21xp5_ASAP7_75t_L g3117 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_1995),
.B(n_2016),
.Y(n_3118)
);

AO21x1_ASAP7_75t_L g3119 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_3119)
);

AOI21x1_ASAP7_75t_L g3120 ( 
.A1(n_2079),
.A2(n_2044),
.B(n_1957),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2016),
.B(n_2018),
.Y(n_3121)
);

NOR2xp33_ASAP7_75t_L g3122 ( 
.A(n_2371),
.B(n_2374),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2351),
.Y(n_3123)
);

AOI21xp5_ASAP7_75t_L g3124 ( 
.A1(n_2921),
.A2(n_2956),
.B(n_2439),
.Y(n_3124)
);

AOI22xp33_ASAP7_75t_L g3125 ( 
.A1(n_2623),
.A2(n_2909),
.B1(n_2974),
.B2(n_1985),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2018),
.B(n_2031),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2031),
.B(n_2042),
.Y(n_3127)
);

NAND2xp5_ASAP7_75t_L g3128 ( 
.A(n_2042),
.B(n_2043),
.Y(n_3128)
);

OAI21xp5_ASAP7_75t_L g3129 ( 
.A1(n_2360),
.A2(n_2632),
.B(n_2494),
.Y(n_3129)
);

AOI21xp5_ASAP7_75t_L g3130 ( 
.A1(n_2862),
.A2(n_3011),
.B(n_2899),
.Y(n_3130)
);

INVxp67_ASAP7_75t_L g3131 ( 
.A(n_2446),
.Y(n_3131)
);

BUFx2_ASAP7_75t_L g3132 ( 
.A(n_2142),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2351),
.Y(n_3133)
);

INVx1_ASAP7_75t_L g3134 ( 
.A(n_2351),
.Y(n_3134)
);

AOI21xp5_ASAP7_75t_L g3135 ( 
.A1(n_1974),
.A2(n_2062),
.B(n_2098),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2043),
.B(n_2101),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_2388),
.B(n_2507),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2106),
.B(n_2107),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2113),
.B(n_2119),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_L g3140 ( 
.A(n_2010),
.B(n_2004),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_SL g3141 ( 
.A(n_2588),
.B(n_2647),
.Y(n_3141)
);

OR2x2_ASAP7_75t_L g3142 ( 
.A(n_2079),
.B(n_2044),
.Y(n_3142)
);

NOR2xp33_ASAP7_75t_L g3143 ( 
.A(n_2380),
.B(n_2395),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2351),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2004),
.B(n_2434),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_SL g3146 ( 
.A(n_2658),
.B(n_2680),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2395),
.B(n_2396),
.Y(n_3147)
);

AOI22xp5_ASAP7_75t_L g3148 ( 
.A1(n_2396),
.A2(n_2437),
.B1(n_2452),
.B2(n_2407),
.Y(n_3148)
);

INVx4_ASAP7_75t_L g3149 ( 
.A(n_2214),
.Y(n_3149)
);

AOI22x1_ASAP7_75t_L g3150 ( 
.A1(n_2844),
.A2(n_2881),
.B1(n_2965),
.B2(n_2053),
.Y(n_3150)
);

AOI21xp5_ASAP7_75t_L g3151 ( 
.A1(n_2062),
.A2(n_2353),
.B(n_1956),
.Y(n_3151)
);

AOI21xp5_ASAP7_75t_L g3152 ( 
.A1(n_1956),
.A2(n_2353),
.B(n_2329),
.Y(n_3152)
);

NAND2xp5_ASAP7_75t_L g3153 ( 
.A(n_2434),
.B(n_2442),
.Y(n_3153)
);

CKINVDCx6p67_ASAP7_75t_R g3154 ( 
.A(n_2214),
.Y(n_3154)
);

AOI22xp33_ASAP7_75t_L g3155 ( 
.A1(n_3039),
.A2(n_2437),
.B1(n_2452),
.B2(n_2407),
.Y(n_3155)
);

AOI21xp5_ASAP7_75t_L g3156 ( 
.A1(n_2329),
.A2(n_2382),
.B(n_2375),
.Y(n_3156)
);

AOI21xp5_ASAP7_75t_L g3157 ( 
.A1(n_2375),
.A2(n_2403),
.B(n_2382),
.Y(n_3157)
);

AOI21xp5_ASAP7_75t_L g3158 ( 
.A1(n_2403),
.A2(n_2422),
.B(n_2411),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2442),
.B(n_2450),
.Y(n_3159)
);

O2A1O1Ixp33_ASAP7_75t_L g3160 ( 
.A1(n_2948),
.A2(n_2853),
.B(n_2054),
.C(n_2075),
.Y(n_3160)
);

O2A1O1Ixp33_ASAP7_75t_L g3161 ( 
.A1(n_2853),
.A2(n_2054),
.B(n_2075),
.C(n_2065),
.Y(n_3161)
);

AOI21xp5_ASAP7_75t_L g3162 ( 
.A1(n_2411),
.A2(n_2440),
.B(n_2422),
.Y(n_3162)
);

AOI21xp5_ASAP7_75t_L g3163 ( 
.A1(n_2444),
.A2(n_2489),
.B(n_2477),
.Y(n_3163)
);

NAND2xp5_ASAP7_75t_L g3164 ( 
.A(n_2450),
.B(n_2458),
.Y(n_3164)
);

NOR2xp33_ASAP7_75t_L g3165 ( 
.A(n_2500),
.B(n_2512),
.Y(n_3165)
);

AOI21xp5_ASAP7_75t_L g3166 ( 
.A1(n_2444),
.A2(n_2486),
.B(n_2468),
.Y(n_3166)
);

AOI21xp5_ASAP7_75t_L g3167 ( 
.A1(n_2468),
.A2(n_2486),
.B(n_2477),
.Y(n_3167)
);

AOI21xp5_ASAP7_75t_L g3168 ( 
.A1(n_2489),
.A2(n_2496),
.B(n_2493),
.Y(n_3168)
);

AOI21xp5_ASAP7_75t_L g3169 ( 
.A1(n_2493),
.A2(n_2523),
.B(n_2496),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_2458),
.B(n_2490),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2701),
.B(n_2751),
.Y(n_3171)
);

NAND2xp5_ASAP7_75t_L g3172 ( 
.A(n_2490),
.B(n_2517),
.Y(n_3172)
);

NAND2xp5_ASAP7_75t_L g3173 ( 
.A(n_2517),
.B(n_2525),
.Y(n_3173)
);

OAI22xp5_ASAP7_75t_L g3174 ( 
.A1(n_2525),
.A2(n_2571),
.B1(n_2582),
.B2(n_2541),
.Y(n_3174)
);

NAND2xp5_ASAP7_75t_L g3175 ( 
.A(n_2541),
.B(n_2571),
.Y(n_3175)
);

AOI21xp5_ASAP7_75t_L g3176 ( 
.A1(n_2440),
.A2(n_2528),
.B(n_2523),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2582),
.B(n_2595),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_2528),
.A2(n_2537),
.B(n_2530),
.Y(n_3178)
);

AOI22xp5_ASAP7_75t_L g3179 ( 
.A1(n_2500),
.A2(n_2513),
.B1(n_2518),
.B2(n_2512),
.Y(n_3179)
);

AOI21xp5_ASAP7_75t_L g3180 ( 
.A1(n_2535),
.A2(n_2547),
.B(n_2537),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_2513),
.B(n_2518),
.Y(n_3181)
);

INVxp67_ASAP7_75t_L g3182 ( 
.A(n_2446),
.Y(n_3182)
);

A2O1A1Ixp33_ASAP7_75t_L g3183 ( 
.A1(n_2532),
.A2(n_2551),
.B(n_2564),
.C(n_2549),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2595),
.B(n_2604),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2849),
.Y(n_3185)
);

HB1xp67_ASAP7_75t_L g3186 ( 
.A(n_2502),
.Y(n_3186)
);

A2O1A1Ixp33_ASAP7_75t_L g3187 ( 
.A1(n_2532),
.A2(n_2551),
.B(n_2564),
.C(n_2549),
.Y(n_3187)
);

AOI21xp5_ASAP7_75t_L g3188 ( 
.A1(n_2530),
.A2(n_2554),
.B(n_2547),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2604),
.B(n_2613),
.Y(n_3189)
);

O2A1O1Ixp5_ASAP7_75t_L g3190 ( 
.A1(n_1971),
.A2(n_2372),
.B(n_2386),
.C(n_1963),
.Y(n_3190)
);

NAND2xp5_ASAP7_75t_L g3191 ( 
.A(n_2613),
.B(n_2642),
.Y(n_3191)
);

BUFx4f_ASAP7_75t_L g3192 ( 
.A(n_2416),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_2033),
.Y(n_3193)
);

A2O1A1Ixp33_ASAP7_75t_L g3194 ( 
.A1(n_2580),
.A2(n_2606),
.B(n_2634),
.C(n_2581),
.Y(n_3194)
);

NAND2x1p5_ASAP7_75t_L g3195 ( 
.A(n_2007),
.B(n_2194),
.Y(n_3195)
);

A2O1A1Ixp33_ASAP7_75t_L g3196 ( 
.A1(n_2580),
.A2(n_2606),
.B(n_2634),
.C(n_2581),
.Y(n_3196)
);

O2A1O1Ixp5_ASAP7_75t_L g3197 ( 
.A1(n_1971),
.A2(n_2850),
.B(n_2559),
.C(n_2065),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_2642),
.B(n_2655),
.Y(n_3198)
);

INVx11_ASAP7_75t_L g3199 ( 
.A(n_2249),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_2102),
.B(n_2032),
.Y(n_3200)
);

NOR2xp33_ASAP7_75t_L g3201 ( 
.A(n_2661),
.B(n_2662),
.Y(n_3201)
);

OAI22xp5_ASAP7_75t_L g3202 ( 
.A1(n_2655),
.A2(n_2677),
.B1(n_2679),
.B2(n_2674),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2102),
.B(n_2032),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2674),
.B(n_2677),
.Y(n_3204)
);

INVx2_ASAP7_75t_SL g3205 ( 
.A(n_2214),
.Y(n_3205)
);

NOR2xp33_ASAP7_75t_L g3206 ( 
.A(n_2661),
.B(n_2662),
.Y(n_3206)
);

AO21x1_ASAP7_75t_L g3207 ( 
.A1(n_2535),
.A2(n_2555),
.B(n_2554),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2679),
.B(n_2684),
.Y(n_3208)
);

NOR3xp33_ASAP7_75t_L g3209 ( 
.A(n_2331),
.B(n_2947),
.C(n_2529),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_2555),
.A2(n_2585),
.B(n_2568),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2849),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_SL g3212 ( 
.A(n_2767),
.B(n_2776),
.Y(n_3212)
);

AOI21xp5_ASAP7_75t_L g3213 ( 
.A1(n_2568),
.A2(n_2586),
.B(n_2585),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2849),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2849),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_2586),
.A2(n_2618),
.B(n_2614),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2230),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_L g3218 ( 
.A(n_2684),
.B(n_2693),
.Y(n_3218)
);

NOR2xp33_ASAP7_75t_L g3219 ( 
.A(n_2699),
.B(n_2726),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_2614),
.A2(n_2622),
.B(n_2618),
.Y(n_3220)
);

BUFx8_ASAP7_75t_L g3221 ( 
.A(n_2650),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2693),
.B(n_2745),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2745),
.B(n_2784),
.Y(n_3223)
);

OAI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_2784),
.A2(n_2897),
.B1(n_2904),
.B2(n_2860),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2039),
.Y(n_3225)
);

OAI22xp5_ASAP7_75t_L g3226 ( 
.A1(n_2860),
.A2(n_2904),
.B1(n_2952),
.B2(n_2897),
.Y(n_3226)
);

AOI21x1_ASAP7_75t_L g3227 ( 
.A1(n_2622),
.A2(n_2638),
.B(n_2636),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_2636),
.A2(n_2657),
.B(n_2646),
.Y(n_3228)
);

AOI21xp5_ASAP7_75t_L g3229 ( 
.A1(n_2646),
.A2(n_2668),
.B(n_2657),
.Y(n_3229)
);

NAND3xp33_ASAP7_75t_L g3230 ( 
.A(n_2952),
.B(n_2975),
.C(n_2958),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2072),
.Y(n_3231)
);

OAI21xp5_ASAP7_75t_L g3232 ( 
.A1(n_2638),
.A2(n_2675),
.B(n_2668),
.Y(n_3232)
);

AOI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_2675),
.A2(n_2718),
.B(n_2690),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_2799),
.B(n_2808),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2039),
.Y(n_3235)
);

AOI21xp5_ASAP7_75t_L g3236 ( 
.A1(n_2690),
.A2(n_2718),
.B(n_2714),
.Y(n_3236)
);

OAI21xp33_ASAP7_75t_L g3237 ( 
.A1(n_2958),
.A2(n_2980),
.B(n_2975),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2980),
.B(n_2984),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_2714),
.A2(n_2744),
.B(n_2739),
.Y(n_3239)
);

NAND2xp5_ASAP7_75t_L g3240 ( 
.A(n_2984),
.B(n_2985),
.Y(n_3240)
);

NOR2xp33_ASAP7_75t_L g3241 ( 
.A(n_2699),
.B(n_2726),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_2735),
.A2(n_2744),
.B(n_2739),
.Y(n_3242)
);

NOR2xp67_ASAP7_75t_L g3243 ( 
.A(n_2227),
.B(n_2125),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_2687),
.A2(n_2765),
.B(n_2735),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_2985),
.B(n_3040),
.Y(n_3245)
);

OAI21xp5_ASAP7_75t_L g3246 ( 
.A1(n_2687),
.A2(n_2766),
.B(n_2765),
.Y(n_3246)
);

BUFx4f_ASAP7_75t_L g3247 ( 
.A(n_2416),
.Y(n_3247)
);

INVxp67_ASAP7_75t_L g3248 ( 
.A(n_2502),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_L g3249 ( 
.A(n_2781),
.B(n_2789),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3040),
.B(n_3043),
.Y(n_3250)
);

INVxp67_ASAP7_75t_L g3251 ( 
.A(n_2601),
.Y(n_3251)
);

AOI21xp5_ASAP7_75t_L g3252 ( 
.A1(n_2766),
.A2(n_2774),
.B(n_2772),
.Y(n_3252)
);

OAI21xp5_ASAP7_75t_L g3253 ( 
.A1(n_2772),
.A2(n_2775),
.B(n_2774),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3043),
.B(n_2416),
.Y(n_3254)
);

AOI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_2775),
.A2(n_2817),
.B(n_2806),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_2416),
.B(n_2903),
.Y(n_3256)
);

NOR3xp33_ASAP7_75t_L g3257 ( 
.A(n_2076),
.B(n_2789),
.C(n_2781),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2039),
.Y(n_3258)
);

AOI21xp33_ASAP7_75t_L g3259 ( 
.A1(n_2824),
.A2(n_2876),
.B(n_2870),
.Y(n_3259)
);

AOI22xp5_ASAP7_75t_L g3260 ( 
.A1(n_2824),
.A2(n_2876),
.B1(n_2893),
.B2(n_2870),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_2815),
.B(n_2821),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_2829),
.B(n_2839),
.Y(n_3262)
);

A2O1A1Ixp33_ASAP7_75t_L g3263 ( 
.A1(n_2893),
.A2(n_2908),
.B(n_2916),
.C(n_2896),
.Y(n_3263)
);

AOI22xp33_ASAP7_75t_L g3264 ( 
.A1(n_3039),
.A2(n_2908),
.B1(n_2916),
.B2(n_2896),
.Y(n_3264)
);

NAND2xp5_ASAP7_75t_L g3265 ( 
.A(n_2416),
.B(n_2903),
.Y(n_3265)
);

AOI21x1_ASAP7_75t_L g3266 ( 
.A1(n_2806),
.A2(n_2842),
.B(n_2817),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2039),
.Y(n_3267)
);

AOI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_2842),
.A2(n_2919),
.B(n_2880),
.Y(n_3268)
);

INVxp67_ASAP7_75t_L g3269 ( 
.A(n_2601),
.Y(n_3269)
);

CKINVDCx11_ASAP7_75t_R g3270 ( 
.A(n_2057),
.Y(n_3270)
);

OAI21xp5_ASAP7_75t_L g3271 ( 
.A1(n_2877),
.A2(n_2919),
.B(n_2880),
.Y(n_3271)
);

OAI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_2877),
.A2(n_2946),
.B(n_2941),
.Y(n_3272)
);

O2A1O1Ixp33_ASAP7_75t_L g3273 ( 
.A1(n_2076),
.A2(n_2962),
.B(n_2964),
.C(n_2924),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_2941),
.A2(n_2970),
.B(n_2946),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_2903),
.B(n_1950),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_2903),
.B(n_1984),
.Y(n_3276)
);

AOI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_2924),
.A2(n_2964),
.B1(n_2967),
.B2(n_2962),
.Y(n_3277)
);

AOI21xp5_ASAP7_75t_L g3278 ( 
.A1(n_2970),
.A2(n_2997),
.B(n_2977),
.Y(n_3278)
);

AOI21xp5_ASAP7_75t_L g3279 ( 
.A1(n_2977),
.A2(n_3000),
.B(n_2997),
.Y(n_3279)
);

AOI21xp5_ASAP7_75t_L g3280 ( 
.A1(n_3000),
.A2(n_3021),
.B(n_3010),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_SL g3281 ( 
.A(n_2841),
.B(n_2847),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_2903),
.B(n_2003),
.Y(n_3282)
);

NOR2xp33_ASAP7_75t_L g3283 ( 
.A(n_2967),
.B(n_2973),
.Y(n_3283)
);

BUFx4f_ASAP7_75t_L g3284 ( 
.A(n_2039),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_3010),
.B(n_3021),
.Y(n_3285)
);

AOI21xp33_ASAP7_75t_L g3286 ( 
.A1(n_2973),
.A2(n_2982),
.B(n_2978),
.Y(n_3286)
);

OR2x2_ASAP7_75t_L g3287 ( 
.A(n_3023),
.B(n_3036),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_SL g3288 ( 
.A(n_2867),
.B(n_2874),
.Y(n_3288)
);

NOR2xp33_ASAP7_75t_L g3289 ( 
.A(n_2978),
.B(n_2982),
.Y(n_3289)
);

NOR2xp67_ASAP7_75t_L g3290 ( 
.A(n_2129),
.B(n_2133),
.Y(n_3290)
);

INVx2_ASAP7_75t_SL g3291 ( 
.A(n_2231),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_L g3292 ( 
.A(n_3023),
.B(n_3036),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_SL g3293 ( 
.A(n_2887),
.B(n_2902),
.Y(n_3293)
);

OAI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3047),
.A2(n_2138),
.B(n_2082),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_2143),
.B(n_2092),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2087),
.Y(n_3296)
);

AOI21xp5_ASAP7_75t_L g3297 ( 
.A1(n_3047),
.A2(n_2136),
.B(n_2134),
.Y(n_3297)
);

NOR2xp33_ASAP7_75t_L g3298 ( 
.A(n_3022),
.B(n_3026),
.Y(n_3298)
);

HB1xp67_ASAP7_75t_L g3299 ( 
.A(n_2715),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_1975),
.B(n_1978),
.Y(n_3300)
);

BUFx2_ASAP7_75t_L g3301 ( 
.A(n_2142),
.Y(n_3301)
);

OAI21xp33_ASAP7_75t_L g3302 ( 
.A1(n_1958),
.A2(n_1969),
.B(n_3022),
.Y(n_3302)
);

AOI21xp5_ASAP7_75t_L g3303 ( 
.A1(n_2147),
.A2(n_2152),
.B(n_2149),
.Y(n_3303)
);

OAI22xp5_ASAP7_75t_L g3304 ( 
.A1(n_2954),
.A2(n_2996),
.B1(n_3002),
.B2(n_2995),
.Y(n_3304)
);

AOI21xp5_ASAP7_75t_L g3305 ( 
.A1(n_2124),
.A2(n_2087),
.B(n_2084),
.Y(n_3305)
);

NAND2x1p5_ASAP7_75t_L g3306 ( 
.A(n_2194),
.B(n_2198),
.Y(n_3306)
);

AOI21xp5_ASAP7_75t_L g3307 ( 
.A1(n_2096),
.A2(n_2266),
.B(n_2173),
.Y(n_3307)
);

AOI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_2266),
.A2(n_2173),
.B(n_2128),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_SL g3309 ( 
.A(n_3027),
.B(n_3038),
.Y(n_3309)
);

NAND2x1p5_ASAP7_75t_L g3310 ( 
.A(n_2198),
.B(n_2219),
.Y(n_3310)
);

AOI21x1_ASAP7_75t_L g3311 ( 
.A1(n_2219),
.A2(n_2120),
.B(n_2241),
.Y(n_3311)
);

OAI22xp5_ASAP7_75t_L g3312 ( 
.A1(n_1958),
.A2(n_1969),
.B1(n_3026),
.B2(n_1940),
.Y(n_3312)
);

AOI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_2128),
.A2(n_2186),
.B(n_2175),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_2175),
.A2(n_2186),
.B(n_2269),
.Y(n_3314)
);

OAI21xp5_ASAP7_75t_L g3315 ( 
.A1(n_2122),
.A2(n_1981),
.B(n_1980),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_1996),
.Y(n_3316)
);

AOI21xp5_ASAP7_75t_L g3317 ( 
.A1(n_2269),
.A2(n_2253),
.B(n_2241),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_L g3318 ( 
.A(n_1953),
.B(n_1955),
.Y(n_3318)
);

BUFx2_ASAP7_75t_L g3319 ( 
.A(n_2199),
.Y(n_3319)
);

NOR2xp33_ASAP7_75t_L g3320 ( 
.A(n_1959),
.B(n_1960),
.Y(n_3320)
);

INVxp67_ASAP7_75t_L g3321 ( 
.A(n_2715),
.Y(n_3321)
);

OAI22xp5_ASAP7_75t_L g3322 ( 
.A1(n_2322),
.A2(n_3033),
.B1(n_3035),
.B2(n_3032),
.Y(n_3322)
);

AOI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_2325),
.A2(n_2327),
.B1(n_2335),
.B2(n_2330),
.Y(n_3323)
);

AOI21xp5_ASAP7_75t_L g3324 ( 
.A1(n_2253),
.A2(n_2273),
.B(n_2265),
.Y(n_3324)
);

BUFx3_ASAP7_75t_L g3325 ( 
.A(n_2394),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_1989),
.B(n_1992),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_2265),
.A2(n_2275),
.B(n_2273),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_2275),
.A2(n_2122),
.B(n_2263),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_1998),
.B(n_2000),
.Y(n_3329)
);

OAI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_2001),
.A2(n_2013),
.B(n_2005),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_SL g3331 ( 
.A(n_2045),
.B(n_2115),
.Y(n_3331)
);

AOI21xp5_ASAP7_75t_L g3332 ( 
.A1(n_2121),
.A2(n_2191),
.B(n_2120),
.Y(n_3332)
);

INVx4_ASAP7_75t_L g3333 ( 
.A(n_2231),
.Y(n_3333)
);

AND2x2_ASAP7_75t_L g3334 ( 
.A(n_2143),
.B(n_1966),
.Y(n_3334)
);

AOI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_2121),
.A2(n_2213),
.B(n_2180),
.Y(n_3335)
);

AOI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_2669),
.A2(n_2721),
.B(n_2683),
.Y(n_3336)
);

NOR2x1p5_ASAP7_75t_L g3337 ( 
.A(n_2281),
.B(n_2165),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_SL g3338 ( 
.A(n_2319),
.B(n_2705),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_2014),
.B(n_2015),
.Y(n_3339)
);

OAI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_2020),
.A2(n_2025),
.B(n_2024),
.Y(n_3340)
);

AOI22xp5_ASAP7_75t_L g3341 ( 
.A1(n_2340),
.A2(n_2346),
.B1(n_2350),
.B2(n_2345),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2036),
.B(n_2040),
.Y(n_3342)
);

O2A1O1Ixp33_ASAP7_75t_L g3343 ( 
.A1(n_3028),
.A2(n_3046),
.B(n_3041),
.C(n_2356),
.Y(n_3343)
);

AND2x4_ASAP7_75t_L g3344 ( 
.A(n_2292),
.B(n_2299),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_L g3345 ( 
.A(n_2358),
.B(n_2361),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2017),
.Y(n_3346)
);

NOR2xp33_ASAP7_75t_SL g3347 ( 
.A(n_2778),
.B(n_2091),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_L g3348 ( 
.A(n_2364),
.B(n_2366),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2368),
.B(n_2381),
.Y(n_3349)
);

CKINVDCx20_ASAP7_75t_R g3350 ( 
.A(n_2561),
.Y(n_3350)
);

HB1xp67_ASAP7_75t_L g3351 ( 
.A(n_2871),
.Y(n_3351)
);

NOR2xp33_ASAP7_75t_L g3352 ( 
.A(n_2384),
.B(n_2393),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_2399),
.B(n_2402),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_2326),
.B(n_2334),
.Y(n_3354)
);

O2A1O1Ixp33_ASAP7_75t_L g3355 ( 
.A1(n_2415),
.A2(n_2419),
.B(n_2429),
.C(n_2420),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_2430),
.B(n_2432),
.Y(n_3356)
);

NAND2xp5_ASAP7_75t_L g3357 ( 
.A(n_2433),
.B(n_2435),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_SL g3358 ( 
.A(n_3048),
.B(n_2094),
.Y(n_3358)
);

AND2x4_ASAP7_75t_L g3359 ( 
.A(n_2301),
.B(n_2285),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_2438),
.B(n_2447),
.Y(n_3360)
);

AOI21xp5_ASAP7_75t_L g3361 ( 
.A1(n_2780),
.A2(n_2891),
.B(n_2267),
.Y(n_3361)
);

NOR2xp33_ASAP7_75t_L g3362 ( 
.A(n_2451),
.B(n_2453),
.Y(n_3362)
);

INVx1_ASAP7_75t_SL g3363 ( 
.A(n_2857),
.Y(n_3363)
);

NAND2xp5_ASAP7_75t_L g3364 ( 
.A(n_2459),
.B(n_2462),
.Y(n_3364)
);

INVx2_ASAP7_75t_SL g3365 ( 
.A(n_2231),
.Y(n_3365)
);

O2A1O1Ixp33_ASAP7_75t_L g3366 ( 
.A1(n_2464),
.A2(n_2466),
.B(n_2473),
.C(n_2471),
.Y(n_3366)
);

AND2x2_ASAP7_75t_L g3367 ( 
.A(n_2349),
.B(n_2367),
.Y(n_3367)
);

NOR2xp33_ASAP7_75t_L g3368 ( 
.A(n_2474),
.B(n_2475),
.Y(n_3368)
);

OAI21xp5_ASAP7_75t_L g3369 ( 
.A1(n_2476),
.A2(n_2483),
.B(n_2478),
.Y(n_3369)
);

INVx1_ASAP7_75t_L g3370 ( 
.A(n_2056),
.Y(n_3370)
);

INVxp67_ASAP7_75t_SL g3371 ( 
.A(n_2871),
.Y(n_3371)
);

AND2x2_ASAP7_75t_L g3372 ( 
.A(n_2378),
.B(n_2418),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_2484),
.A2(n_2495),
.B(n_2492),
.Y(n_3373)
);

AO21x1_ASAP7_75t_L g3374 ( 
.A1(n_2089),
.A2(n_2277),
.B(n_2498),
.Y(n_3374)
);

NAND2xp5_ASAP7_75t_L g3375 ( 
.A(n_2506),
.B(n_2509),
.Y(n_3375)
);

O2A1O1Ixp33_ASAP7_75t_L g3376 ( 
.A1(n_2510),
.A2(n_2511),
.B(n_2516),
.C(n_2515),
.Y(n_3376)
);

OAI21xp33_ASAP7_75t_L g3377 ( 
.A1(n_2519),
.A2(n_2536),
.B(n_2531),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_2441),
.B(n_2534),
.Y(n_3378)
);

BUFx2_ASAP7_75t_L g3379 ( 
.A(n_2011),
.Y(n_3379)
);

AOI22xp5_ASAP7_75t_L g3380 ( 
.A1(n_2539),
.A2(n_2544),
.B1(n_2563),
.B2(n_2560),
.Y(n_3380)
);

OAI22xp5_ASAP7_75t_L g3381 ( 
.A1(n_2566),
.A2(n_2575),
.B1(n_2576),
.B2(n_2574),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_SL g3382 ( 
.A(n_2144),
.B(n_2589),
.Y(n_3382)
);

AND2x2_ASAP7_75t_L g3383 ( 
.A(n_2545),
.B(n_2567),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_SL g3384 ( 
.A(n_2590),
.B(n_2592),
.Y(n_3384)
);

NOR2xp67_ASAP7_75t_L g3385 ( 
.A(n_2207),
.B(n_2209),
.Y(n_3385)
);

BUFx6f_ASAP7_75t_L g3386 ( 
.A(n_2300),
.Y(n_3386)
);

NOR3xp33_ASAP7_75t_L g3387 ( 
.A(n_2599),
.B(n_2609),
.C(n_2608),
.Y(n_3387)
);

BUFx4f_ASAP7_75t_L g3388 ( 
.A(n_2377),
.Y(n_3388)
);

AOI33xp33_ASAP7_75t_L g3389 ( 
.A1(n_2691),
.A2(n_2704),
.A3(n_2729),
.B1(n_2747),
.B2(n_2733),
.B3(n_2720),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_2612),
.A2(n_2625),
.B(n_2620),
.Y(n_3390)
);

AOI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_2630),
.A2(n_2633),
.B1(n_2635),
.B2(n_2631),
.Y(n_3391)
);

OAI21xp5_ASAP7_75t_L g3392 ( 
.A1(n_2637),
.A2(n_2649),
.B(n_2641),
.Y(n_3392)
);

O2A1O1Ixp33_ASAP7_75t_SL g3393 ( 
.A1(n_2670),
.A2(n_2785),
.B(n_2795),
.C(n_2746),
.Y(n_3393)
);

AOI21xp33_ASAP7_75t_L g3394 ( 
.A1(n_2663),
.A2(n_2667),
.B(n_2666),
.Y(n_3394)
);

AOI21xp5_ASAP7_75t_L g3395 ( 
.A1(n_2689),
.A2(n_2695),
.B(n_2694),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_2697),
.B(n_3016),
.Y(n_3396)
);

AO21x1_ASAP7_75t_L g3397 ( 
.A1(n_2702),
.A2(n_2713),
.B(n_2708),
.Y(n_3397)
);

INVx11_ASAP7_75t_L g3398 ( 
.A(n_2427),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_2719),
.A2(n_2724),
.B(n_2722),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_L g3400 ( 
.A(n_2728),
.B(n_2732),
.Y(n_3400)
);

AOI21xp5_ASAP7_75t_L g3401 ( 
.A1(n_2737),
.A2(n_2742),
.B(n_2740),
.Y(n_3401)
);

AOI21xp5_ASAP7_75t_L g3402 ( 
.A1(n_2748),
.A2(n_2756),
.B(n_2755),
.Y(n_3402)
);

AOI21xp5_ASAP7_75t_L g3403 ( 
.A1(n_2759),
.A2(n_2763),
.B(n_2760),
.Y(n_3403)
);

O2A1O1Ixp33_ASAP7_75t_L g3404 ( 
.A1(n_2768),
.A2(n_2779),
.B(n_2786),
.C(n_2782),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_2758),
.B(n_2818),
.Y(n_3405)
);

AOI21x1_ASAP7_75t_L g3406 ( 
.A1(n_2023),
.A2(n_2035),
.B(n_2264),
.Y(n_3406)
);

AOI21xp5_ASAP7_75t_L g3407 ( 
.A1(n_2794),
.A2(n_2805),
.B(n_2797),
.Y(n_3407)
);

AOI21xp5_ASAP7_75t_L g3408 ( 
.A1(n_2809),
.A2(n_2812),
.B(n_2810),
.Y(n_3408)
);

OR2x2_ASAP7_75t_L g3409 ( 
.A(n_1941),
.B(n_2406),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_2816),
.B(n_2819),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_2820),
.B(n_2822),
.Y(n_3411)
);

O2A1O1Ixp5_ASAP7_75t_L g3412 ( 
.A1(n_2189),
.A2(n_2828),
.B(n_2834),
.C(n_2832),
.Y(n_3412)
);

AOI21xp5_ASAP7_75t_L g3413 ( 
.A1(n_2840),
.A2(n_2848),
.B(n_2845),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2875),
.B(n_2879),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2073),
.Y(n_3415)
);

AOI21xp5_ASAP7_75t_L g3416 ( 
.A1(n_2885),
.A2(n_2890),
.B(n_2888),
.Y(n_3416)
);

OAI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_2894),
.A2(n_2905),
.B(n_2898),
.Y(n_3417)
);

AOI21xp5_ASAP7_75t_L g3418 ( 
.A1(n_2910),
.A2(n_2913),
.B(n_2911),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_2917),
.B(n_2922),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_SL g3420 ( 
.A(n_2927),
.B(n_2930),
.Y(n_3420)
);

AOI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_2933),
.A2(n_2936),
.B(n_2934),
.Y(n_3421)
);

NOR2xp67_ASAP7_75t_L g3422 ( 
.A(n_2233),
.B(n_1986),
.Y(n_3422)
);

OAI21x1_ASAP7_75t_L g3423 ( 
.A1(n_2300),
.A2(n_2305),
.B(n_1986),
.Y(n_3423)
);

NAND2xp5_ASAP7_75t_SL g3424 ( 
.A(n_2937),
.B(n_2938),
.Y(n_3424)
);

AOI21xp5_ASAP7_75t_L g3425 ( 
.A1(n_2940),
.A2(n_2953),
.B(n_2942),
.Y(n_3425)
);

A2O1A1Ixp33_ASAP7_75t_L g3426 ( 
.A1(n_2960),
.A2(n_2966),
.B(n_2976),
.C(n_2972),
.Y(n_3426)
);

OAI21xp33_ASAP7_75t_L g3427 ( 
.A1(n_2981),
.A2(n_2988),
.B(n_2983),
.Y(n_3427)
);

NOR2xp33_ASAP7_75t_L g3428 ( 
.A(n_2989),
.B(n_2991),
.Y(n_3428)
);

AOI21xp33_ASAP7_75t_L g3429 ( 
.A1(n_2993),
.A2(n_3008),
.B(n_2994),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3009),
.A2(n_3013),
.B(n_2278),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_2454),
.B(n_2546),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_L g3432 ( 
.A(n_2008),
.B(n_2470),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_2583),
.B(n_2611),
.Y(n_3433)
);

CKINVDCx5p33_ASAP7_75t_R g3434 ( 
.A(n_2749),
.Y(n_3434)
);

BUFx4f_ASAP7_75t_L g3435 ( 
.A(n_2377),
.Y(n_3435)
);

AOI21xp5_ASAP7_75t_L g3436 ( 
.A1(n_2259),
.A2(n_2260),
.B(n_2239),
.Y(n_3436)
);

INVx3_ASAP7_75t_L g3437 ( 
.A(n_2436),
.Y(n_3437)
);

NOR2xp33_ASAP7_75t_L g3438 ( 
.A(n_2851),
.B(n_2949),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_2081),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_2678),
.B(n_2734),
.Y(n_3440)
);

NAND2xp5_ASAP7_75t_L g3441 ( 
.A(n_2771),
.B(n_2793),
.Y(n_3441)
);

NOR2xp33_ASAP7_75t_L g3442 ( 
.A(n_2990),
.B(n_3001),
.Y(n_3442)
);

NOR2xp33_ASAP7_75t_L g3443 ( 
.A(n_3003),
.B(n_3004),
.Y(n_3443)
);

CKINVDCx5p33_ASAP7_75t_R g3444 ( 
.A(n_2861),
.Y(n_3444)
);

HB1xp67_ASAP7_75t_L g3445 ( 
.A(n_2155),
.Y(n_3445)
);

AOI21xp5_ASAP7_75t_L g3446 ( 
.A1(n_2153),
.A2(n_2167),
.B(n_2161),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_2827),
.B(n_2843),
.Y(n_3447)
);

AND2x2_ASAP7_75t_L g3448 ( 
.A(n_3037),
.B(n_2012),
.Y(n_3448)
);

NOR2xp33_ASAP7_75t_L g3449 ( 
.A(n_2127),
.B(n_2859),
.Y(n_3449)
);

A2O1A1Ixp33_ASAP7_75t_L g3450 ( 
.A1(n_2034),
.A2(n_2570),
.B(n_2357),
.C(n_2232),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_2127),
.B(n_2864),
.Y(n_3451)
);

INVxp67_ASAP7_75t_L g3452 ( 
.A(n_2158),
.Y(n_3452)
);

AOI21xp5_ASAP7_75t_L g3453 ( 
.A1(n_2168),
.A2(n_2171),
.B(n_2170),
.Y(n_3453)
);

A2O1A1Ixp33_ASAP7_75t_L g3454 ( 
.A1(n_2232),
.A2(n_2234),
.B(n_2248),
.C(n_2279),
.Y(n_3454)
);

NAND2xp5_ASAP7_75t_L g3455 ( 
.A(n_2929),
.B(n_2932),
.Y(n_3455)
);

AOI21x1_ASAP7_75t_L g3456 ( 
.A1(n_2272),
.A2(n_2274),
.B(n_2307),
.Y(n_3456)
);

NAND3xp33_ASAP7_75t_L g3457 ( 
.A(n_2105),
.B(n_2204),
.C(n_2221),
.Y(n_3457)
);

NAND2xp5_ASAP7_75t_L g3458 ( 
.A(n_2132),
.B(n_2148),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_SL g3459 ( 
.A(n_2108),
.B(n_2123),
.Y(n_3459)
);

AOI21xp5_ASAP7_75t_L g3460 ( 
.A1(n_2174),
.A2(n_2177),
.B(n_2176),
.Y(n_3460)
);

OAI21xp33_ASAP7_75t_L g3461 ( 
.A1(n_2055),
.A2(n_2067),
.B(n_2058),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_SL g3462 ( 
.A(n_2123),
.B(n_2157),
.Y(n_3462)
);

BUFx3_ASAP7_75t_L g3463 ( 
.A(n_2394),
.Y(n_3463)
);

CKINVDCx20_ASAP7_75t_R g3464 ( 
.A(n_2872),
.Y(n_3464)
);

O2A1O1Ixp5_ASAP7_75t_L g3465 ( 
.A1(n_2615),
.A2(n_2955),
.B(n_3044),
.C(n_2951),
.Y(n_3465)
);

AOI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_2019),
.A2(n_2088),
.B1(n_2069),
.B2(n_2071),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_2150),
.Y(n_3467)
);

OAI21xp5_ASAP7_75t_L g3468 ( 
.A1(n_2250),
.A2(n_2254),
.B(n_1967),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_1952),
.B(n_2324),
.Y(n_3469)
);

AOI21xp5_ASAP7_75t_L g3470 ( 
.A1(n_2271),
.A2(n_2154),
.B(n_2146),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_2068),
.B(n_2077),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_2160),
.B(n_2164),
.Y(n_3472)
);

AOI21xp5_ASAP7_75t_L g3473 ( 
.A1(n_2146),
.A2(n_2659),
.B(n_2436),
.Y(n_3473)
);

INVx4_ASAP7_75t_L g3474 ( 
.A(n_2231),
.Y(n_3474)
);

AOI21xp5_ASAP7_75t_L g3475 ( 
.A1(n_2659),
.A2(n_2730),
.B(n_2671),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_2320),
.B(n_2321),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_2328),
.B(n_2332),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_2333),
.B(n_2341),
.Y(n_3478)
);

OAI22x1_ASAP7_75t_L g3479 ( 
.A1(n_2203),
.A2(n_1945),
.B1(n_2664),
.B2(n_2643),
.Y(n_3479)
);

NAND2xp5_ASAP7_75t_L g3480 ( 
.A(n_2355),
.B(n_2369),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_2813),
.A2(n_2866),
.B(n_2846),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_L g3482 ( 
.A(n_2385),
.B(n_2389),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_2398),
.B(n_2400),
.Y(n_3483)
);

OAI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2250),
.A2(n_2254),
.B(n_2339),
.Y(n_3484)
);

INVx2_ASAP7_75t_SL g3485 ( 
.A(n_2298),
.Y(n_3485)
);

O2A1O1Ixp33_ASAP7_75t_L g3486 ( 
.A1(n_2088),
.A2(n_2080),
.B(n_2181),
.C(n_2052),
.Y(n_3486)
);

AND2x4_ASAP7_75t_L g3487 ( 
.A(n_2866),
.B(n_2064),
.Y(n_3487)
);

AO21x1_ASAP7_75t_L g3488 ( 
.A1(n_2225),
.A2(n_2226),
.B(n_2423),
.Y(n_3488)
);

NOR2xp33_ASAP7_75t_SL g3489 ( 
.A(n_2538),
.B(n_2698),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_2424),
.B(n_2426),
.Y(n_3490)
);

NOR2x1_ASAP7_75t_L g3491 ( 
.A(n_2088),
.B(n_2565),
.Y(n_3491)
);

A2O1A1Ixp33_ASAP7_75t_L g3492 ( 
.A1(n_2234),
.A2(n_2248),
.B(n_2257),
.C(n_2255),
.Y(n_3492)
);

INVx3_ASAP7_75t_SL g3493 ( 
.A(n_2550),
.Y(n_3493)
);

NAND2x1_ASAP7_75t_L g3494 ( 
.A(n_2347),
.B(n_2359),
.Y(n_3494)
);

OAI21xp5_ASAP7_75t_L g3495 ( 
.A1(n_2379),
.A2(n_2391),
.B(n_2390),
.Y(n_3495)
);

AOI21xp5_ASAP7_75t_L g3496 ( 
.A1(n_2308),
.A2(n_2257),
.B(n_2255),
.Y(n_3496)
);

OAI21xp33_ASAP7_75t_L g3497 ( 
.A1(n_2195),
.A2(n_2158),
.B(n_2156),
.Y(n_3497)
);

OAI22xp5_ASAP7_75t_L g3498 ( 
.A1(n_2448),
.A2(n_2469),
.B1(n_2472),
.B2(n_2463),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_2412),
.A2(n_2449),
.B(n_2425),
.Y(n_3499)
);

AOI22xp33_ASAP7_75t_L g3500 ( 
.A1(n_2187),
.A2(n_1991),
.B1(n_2573),
.B2(n_1944),
.Y(n_3500)
);

A2O1A1Ixp33_ASAP7_75t_L g3501 ( 
.A1(n_2268),
.A2(n_1973),
.B(n_1997),
.C(n_1990),
.Y(n_3501)
);

AOI21xp5_ASAP7_75t_L g3502 ( 
.A1(n_2455),
.A2(n_2487),
.B(n_2467),
.Y(n_3502)
);

BUFx12f_ASAP7_75t_L g3503 ( 
.A(n_2427),
.Y(n_3503)
);

AOI22xp5_ASAP7_75t_L g3504 ( 
.A1(n_1991),
.A2(n_2218),
.B1(n_2140),
.B2(n_2156),
.Y(n_3504)
);

AND2x6_ASAP7_75t_L g3505 ( 
.A(n_2480),
.B(n_2491),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_2861),
.B(n_2064),
.Y(n_3506)
);

OAI21x1_ASAP7_75t_L g3507 ( 
.A1(n_2497),
.A2(n_2522),
.B(n_2504),
.Y(n_3507)
);

BUFx8_ASAP7_75t_SL g3508 ( 
.A(n_2769),
.Y(n_3508)
);

NAND2xp5_ASAP7_75t_SL g3509 ( 
.A(n_2064),
.B(n_2508),
.Y(n_3509)
);

NOR2xp33_ASAP7_75t_L g3510 ( 
.A(n_2629),
.B(n_2135),
.Y(n_3510)
);

OAI21xp5_ASAP7_75t_L g3511 ( 
.A1(n_2526),
.A2(n_2587),
.B(n_2542),
.Y(n_3511)
);

OAI21xp5_ASAP7_75t_L g3512 ( 
.A1(n_2600),
.A2(n_2653),
.B(n_2602),
.Y(n_3512)
);

AOI21xp5_ASAP7_75t_L g3513 ( 
.A1(n_2654),
.A2(n_2696),
.B(n_2676),
.Y(n_3513)
);

NAND2xp5_ASAP7_75t_L g3514 ( 
.A(n_2501),
.B(n_2521),
.Y(n_3514)
);

O2A1O1Ixp33_ASAP7_75t_L g3515 ( 
.A1(n_2074),
.A2(n_2311),
.B(n_2178),
.C(n_2741),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_L g3516 ( 
.A(n_2524),
.B(n_2527),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_L g3517 ( 
.A1(n_2533),
.A2(n_2552),
.B1(n_2557),
.B2(n_2543),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_2717),
.A2(n_2791),
.B(n_2790),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_2569),
.B(n_2572),
.Y(n_3519)
);

AOI22xp33_ASAP7_75t_L g3520 ( 
.A1(n_2868),
.A2(n_2882),
.B1(n_2928),
.B2(n_2140),
.Y(n_3520)
);

AOI22xp5_ASAP7_75t_L g3521 ( 
.A1(n_2145),
.A2(n_2197),
.B1(n_2246),
.B2(n_2116),
.Y(n_3521)
);

BUFx3_ASAP7_75t_L g3522 ( 
.A(n_2553),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_2145),
.B(n_2169),
.Y(n_3523)
);

AOI21x1_ASAP7_75t_L g3524 ( 
.A1(n_2605),
.A2(n_3049),
.B(n_2681),
.Y(n_3524)
);

AOI21xp5_ASAP7_75t_L g3525 ( 
.A1(n_2792),
.A2(n_2807),
.B(n_2801),
.Y(n_3525)
);

AND2x2_ASAP7_75t_L g3526 ( 
.A(n_2823),
.B(n_2831),
.Y(n_3526)
);

NAND2xp5_ASAP7_75t_SL g3527 ( 
.A(n_2064),
.B(n_2508),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_2169),
.B(n_2648),
.Y(n_3528)
);

INVx2_ASAP7_75t_SL g3529 ( 
.A(n_2298),
.Y(n_3529)
);

HB1xp67_ASAP7_75t_L g3530 ( 
.A(n_2178),
.Y(n_3530)
);

AOI21xp5_ASAP7_75t_L g3531 ( 
.A1(n_2856),
.A2(n_2895),
.B(n_2884),
.Y(n_3531)
);

AO21x1_ASAP7_75t_L g3532 ( 
.A1(n_2624),
.A2(n_2688),
.B(n_2686),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_SL g3533 ( 
.A(n_2508),
.B(n_1965),
.Y(n_3533)
);

AOI21xp5_ASAP7_75t_L g3534 ( 
.A1(n_2907),
.A2(n_2931),
.B(n_2915),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_2706),
.Y(n_3535)
);

O2A1O1Ixp5_ASAP7_75t_L g3536 ( 
.A1(n_2311),
.A2(n_2078),
.B(n_2238),
.C(n_2235),
.Y(n_3536)
);

O2A1O1Ixp33_ASAP7_75t_L g3537 ( 
.A1(n_2268),
.A2(n_2276),
.B(n_2197),
.C(n_2312),
.Y(n_3537)
);

INVx2_ASAP7_75t_SL g3538 ( 
.A(n_2298),
.Y(n_3538)
);

OAI21xp5_ASAP7_75t_L g3539 ( 
.A1(n_2959),
.A2(n_2992),
.B(n_2963),
.Y(n_3539)
);

OR2x6_ASAP7_75t_L g3540 ( 
.A(n_2577),
.B(n_2798),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_2712),
.B(n_2723),
.Y(n_3541)
);

AOI21xp5_ASAP7_75t_L g3542 ( 
.A1(n_2998),
.A2(n_3005),
.B(n_2999),
.Y(n_3542)
);

OAI21x1_ASAP7_75t_L g3543 ( 
.A1(n_3012),
.A2(n_3025),
.B(n_3014),
.Y(n_3543)
);

OAI22xp5_ASAP7_75t_L g3544 ( 
.A1(n_2725),
.A2(n_2761),
.B1(n_2787),
.B2(n_2752),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_2796),
.Y(n_3545)
);

AOI21xp5_ASAP7_75t_L g3546 ( 
.A1(n_3031),
.A2(n_3034),
.B(n_2009),
.Y(n_3546)
);

INVx4_ASAP7_75t_L g3547 ( 
.A(n_2298),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_2800),
.B(n_2802),
.Y(n_3548)
);

AOI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_2002),
.A2(n_2028),
.B(n_2026),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_2811),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_SL g3551 ( 
.A(n_2508),
.B(n_1965),
.Y(n_3551)
);

BUFx6f_ASAP7_75t_L g3552 ( 
.A(n_2577),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_2030),
.B(n_2037),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_L g3554 ( 
.A(n_2814),
.B(n_2825),
.Y(n_3554)
);

NOR3xp33_ASAP7_75t_L g3555 ( 
.A(n_2090),
.B(n_2626),
.C(n_1948),
.Y(n_3555)
);

CKINVDCx8_ASAP7_75t_R g3556 ( 
.A(n_2290),
.Y(n_3556)
);

CKINVDCx5p33_ASAP7_75t_R g3557 ( 
.A(n_2022),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_SL g3558 ( 
.A(n_2413),
.B(n_2593),
.Y(n_3558)
);

O2A1O1Ixp33_ASAP7_75t_L g3559 ( 
.A1(n_2314),
.A2(n_2303),
.B(n_2051),
.C(n_2063),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_L g3560 ( 
.A(n_2826),
.B(n_2830),
.Y(n_3560)
);

AOI22xp33_ASAP7_75t_L g3561 ( 
.A1(n_2193),
.A2(n_2593),
.B1(n_2639),
.B2(n_2413),
.Y(n_3561)
);

AOI21xp5_ASAP7_75t_L g3562 ( 
.A1(n_2050),
.A2(n_2085),
.B(n_2070),
.Y(n_3562)
);

OAI22xp5_ASAP7_75t_L g3563 ( 
.A1(n_2833),
.A2(n_2837),
.B1(n_2838),
.B2(n_2835),
.Y(n_3563)
);

AOI21xp5_ASAP7_75t_L g3564 ( 
.A1(n_2097),
.A2(n_2104),
.B(n_2099),
.Y(n_3564)
);

NOR2xp33_ASAP7_75t_L g3565 ( 
.A(n_2709),
.B(n_2770),
.Y(n_3565)
);

AOI21xp5_ASAP7_75t_L g3566 ( 
.A1(n_2126),
.A2(n_2131),
.B(n_2130),
.Y(n_3566)
);

NOR2xp33_ASAP7_75t_SL g3567 ( 
.A(n_2769),
.B(n_2217),
.Y(n_3567)
);

A2O1A1Ixp33_ASAP7_75t_L g3568 ( 
.A1(n_2137),
.A2(n_2172),
.B(n_2166),
.C(n_2163),
.Y(n_3568)
);

BUFx6f_ASAP7_75t_L g3569 ( 
.A(n_2798),
.Y(n_3569)
);

NOR2xp33_ASAP7_75t_L g3570 ( 
.A(n_2773),
.B(n_2914),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_2865),
.B(n_2869),
.Y(n_3571)
);

NOR2xp33_ASAP7_75t_L g3572 ( 
.A(n_2338),
.B(n_2404),
.Y(n_3572)
);

AOI21xp5_ASAP7_75t_L g3573 ( 
.A1(n_2190),
.A2(n_2208),
.B(n_2206),
.Y(n_3573)
);

OAI21xp33_ASAP7_75t_L g3574 ( 
.A1(n_2195),
.A2(n_2883),
.B(n_2873),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_2499),
.B(n_2711),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_2886),
.Y(n_3576)
);

AOI21xp5_ASAP7_75t_L g3577 ( 
.A1(n_2216),
.A2(n_2223),
.B(n_2220),
.Y(n_3577)
);

HB1xp67_ASAP7_75t_L g3578 ( 
.A(n_2302),
.Y(n_3578)
);

NOR2xp33_ASAP7_75t_R g3579 ( 
.A(n_2313),
.B(n_2553),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_2889),
.B(n_2918),
.Y(n_3580)
);

AOI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_2236),
.A2(n_2247),
.B(n_2244),
.Y(n_3581)
);

AND2x2_ASAP7_75t_L g3582 ( 
.A(n_2923),
.B(n_2925),
.Y(n_3582)
);

BUFx2_ASAP7_75t_L g3583 ( 
.A(n_2109),
.Y(n_3583)
);

HB1xp67_ASAP7_75t_L g3584 ( 
.A(n_2304),
.Y(n_3584)
);

CKINVDCx10_ASAP7_75t_R g3585 ( 
.A(n_1982),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_2926),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_2935),
.B(n_2939),
.Y(n_3587)
);

AOI21xp5_ASAP7_75t_L g3588 ( 
.A1(n_2256),
.A2(n_2961),
.B(n_2943),
.Y(n_3588)
);

OAI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_2240),
.A2(n_2986),
.B(n_2968),
.Y(n_3589)
);

O2A1O1Ixp33_ASAP7_75t_L g3590 ( 
.A1(n_2987),
.A2(n_3030),
.B(n_3020),
.C(n_3019),
.Y(n_3590)
);

OAI321xp33_ASAP7_75t_L g3591 ( 
.A1(n_2310),
.A2(n_3017),
.A3(n_2878),
.B1(n_2200),
.B2(n_2251),
.C(n_2179),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_2878),
.A2(n_2245),
.B(n_2261),
.Y(n_3592)
);

O2A1O1Ixp33_ASAP7_75t_SL g3593 ( 
.A1(n_2184),
.A2(n_2188),
.B(n_2185),
.C(n_2242),
.Y(n_3593)
);

AOI21xp5_ASAP7_75t_L g3594 ( 
.A1(n_2262),
.A2(n_2258),
.B(n_2210),
.Y(n_3594)
);

AOI21xp5_ASAP7_75t_L g3595 ( 
.A1(n_2196),
.A2(n_2205),
.B(n_2237),
.Y(n_3595)
);

NAND2xp5_ASAP7_75t_L g3596 ( 
.A(n_2202),
.B(n_2212),
.Y(n_3596)
);

BUFx2_ASAP7_75t_SL g3597 ( 
.A(n_2066),
.Y(n_3597)
);

NAND2xp5_ASAP7_75t_L g3598 ( 
.A(n_2639),
.B(n_2665),
.Y(n_3598)
);

INVx2_ASAP7_75t_L g3599 ( 
.A(n_1964),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_SL g3600 ( 
.A(n_2665),
.B(n_2764),
.Y(n_3600)
);

INVx3_ASAP7_75t_L g3601 ( 
.A(n_2764),
.Y(n_3601)
);

A2O1A1Ixp33_ASAP7_75t_L g3602 ( 
.A1(n_2777),
.A2(n_3018),
.B(n_2804),
.C(n_2979),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_1964),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_1964),
.Y(n_3604)
);

AOI21xp5_ASAP7_75t_L g3605 ( 
.A1(n_2110),
.A2(n_2211),
.B(n_2777),
.Y(n_3605)
);

INVx3_ASAP7_75t_L g3606 ( 
.A(n_2804),
.Y(n_3606)
);

INVx3_ASAP7_75t_L g3607 ( 
.A(n_2979),
.Y(n_3607)
);

AOI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_2110),
.A2(n_2211),
.B(n_3018),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_2743),
.B(n_3029),
.Y(n_3609)
);

NOR2xp67_ASAP7_75t_L g3610 ( 
.A(n_2061),
.B(n_2607),
.Y(n_3610)
);

AOI21xp5_ASAP7_75t_L g3611 ( 
.A1(n_2061),
.A2(n_2252),
.B(n_1994),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_1964),
.Y(n_3612)
);

OAI22xp5_ASAP7_75t_L g3613 ( 
.A1(n_2193),
.A2(n_1994),
.B1(n_2046),
.B2(n_2289),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_SL g3614 ( 
.A(n_2022),
.B(n_2957),
.Y(n_3614)
);

INVx1_ASAP7_75t_SL g3615 ( 
.A(n_2282),
.Y(n_3615)
);

AOI21xp5_ASAP7_75t_L g3616 ( 
.A1(n_2252),
.A2(n_1994),
.B(n_2295),
.Y(n_3616)
);

AOI21xp5_ASAP7_75t_L g3617 ( 
.A1(n_2283),
.A2(n_2193),
.B(n_2296),
.Y(n_3617)
);

AOI21xp5_ASAP7_75t_L g3618 ( 
.A1(n_2296),
.A2(n_2306),
.B(n_2083),
.Y(n_3618)
);

INVx3_ASAP7_75t_L g3619 ( 
.A(n_1988),
.Y(n_3619)
);

BUFx6f_ASAP7_75t_L g3620 ( 
.A(n_1988),
.Y(n_3620)
);

AND2x4_ASAP7_75t_L g3621 ( 
.A(n_2083),
.B(n_1982),
.Y(n_3621)
);

BUFx8_ASAP7_75t_L g3622 ( 
.A(n_2111),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_1988),
.Y(n_3623)
);

BUFx2_ASAP7_75t_L g3624 ( 
.A(n_2048),
.Y(n_3624)
);

HB1xp67_ASAP7_75t_L g3625 ( 
.A(n_2288),
.Y(n_3625)
);

AOI21xp5_ASAP7_75t_L g3626 ( 
.A1(n_2306),
.A2(n_2083),
.B(n_2270),
.Y(n_3626)
);

AOI21x1_ASAP7_75t_L g3627 ( 
.A1(n_2316),
.A2(n_2162),
.B(n_2222),
.Y(n_3627)
);

AND2x2_ASAP7_75t_L g3628 ( 
.A(n_2048),
.B(n_2117),
.Y(n_3628)
);

BUFx12f_ASAP7_75t_L g3629 ( 
.A(n_2660),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_2048),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_2270),
.A2(n_2945),
.B(n_2920),
.Y(n_3631)
);

O2A1O1Ixp33_ASAP7_75t_L g3632 ( 
.A1(n_1951),
.A2(n_2503),
.B(n_2971),
.C(n_2950),
.Y(n_3632)
);

AOI21xp5_ASAP7_75t_L g3633 ( 
.A1(n_2048),
.A2(n_2703),
.B(n_2616),
.Y(n_3633)
);

AOI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_2117),
.A2(n_2945),
.B(n_2920),
.Y(n_3634)
);

AND2x2_ASAP7_75t_L g3635 ( 
.A(n_2117),
.B(n_2201),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_2117),
.B(n_2201),
.Y(n_3636)
);

BUFx8_ASAP7_75t_SL g3637 ( 
.A(n_2183),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_2201),
.B(n_2224),
.Y(n_3638)
);

OAI22xp5_ASAP7_75t_L g3639 ( 
.A1(n_2297),
.A2(n_1987),
.B1(n_1982),
.B2(n_2222),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_L g3640 ( 
.A(n_2201),
.B(n_2224),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_2224),
.Y(n_3641)
);

NAND2x1p5_ASAP7_75t_L g3642 ( 
.A(n_1948),
.B(n_2626),
.Y(n_3642)
);

AOI21xp5_ASAP7_75t_L g3643 ( 
.A1(n_2224),
.A2(n_2616),
.B(n_2945),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_2229),
.B(n_2457),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_2229),
.B(n_2457),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_2229),
.A2(n_2945),
.B(n_2920),
.Y(n_3646)
);

INVx2_ASAP7_75t_SL g3647 ( 
.A(n_2229),
.Y(n_3647)
);

AOI21xp5_ASAP7_75t_L g3648 ( 
.A1(n_2457),
.A2(n_2920),
.B(n_2855),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_L g3649 ( 
.A(n_2457),
.B(n_2616),
.Y(n_3649)
);

O2A1O1Ixp33_ASAP7_75t_SL g3650 ( 
.A1(n_2315),
.A2(n_2558),
.B(n_2912),
.C(n_2892),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_2616),
.Y(n_3651)
);

NAND2xp5_ASAP7_75t_L g3652 ( 
.A(n_2703),
.B(n_2855),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_2703),
.B(n_2855),
.Y(n_3653)
);

O2A1O1Ixp33_ASAP7_75t_SL g3654 ( 
.A1(n_2151),
.A2(n_2520),
.B(n_2858),
.C(n_2854),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_2293),
.B(n_2855),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_2703),
.B(n_2640),
.Y(n_3656)
);

A2O1A1Ixp33_ASAP7_75t_L g3657 ( 
.A1(n_2309),
.A2(n_2627),
.B(n_2481),
.C(n_2757),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_SL g3658 ( 
.A(n_2293),
.B(n_2640),
.Y(n_3658)
);

OAI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_1987),
.A2(n_2222),
.B1(n_2365),
.B2(n_2344),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_2309),
.Y(n_3660)
);

NOR2xp33_ASAP7_75t_SL g3661 ( 
.A(n_1987),
.B(n_3042),
.Y(n_3661)
);

INVx2_ASAP7_75t_L g3662 ( 
.A(n_1943),
.Y(n_3662)
);

AOI22xp5_ASAP7_75t_L g3663 ( 
.A1(n_2095),
.A2(n_2461),
.B1(n_2365),
.B2(n_2344),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_2672),
.B(n_2762),
.Y(n_3664)
);

OAI22xp5_ASAP7_75t_L g3665 ( 
.A1(n_2342),
.A2(n_2461),
.B1(n_2365),
.B2(n_2344),
.Y(n_3665)
);

BUFx6f_ASAP7_75t_L g3666 ( 
.A(n_2553),
.Y(n_3666)
);

OAI22xp5_ASAP7_75t_L g3667 ( 
.A1(n_2342),
.A2(n_2461),
.B1(n_3045),
.B2(n_2603),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_2672),
.B(n_2762),
.Y(n_3668)
);

HB1xp67_ASAP7_75t_L g3669 ( 
.A(n_2284),
.Y(n_3669)
);

NAND2x1p5_ASAP7_75t_L g3670 ( 
.A(n_2243),
.B(n_2783),
.Y(n_3670)
);

NOR3xp33_ASAP7_75t_L g3671 ( 
.A(n_2337),
.B(n_2579),
.C(n_2753),
.Y(n_3671)
);

BUFx2_ASAP7_75t_L g3672 ( 
.A(n_2141),
.Y(n_3672)
);

NOR2xp33_ASAP7_75t_SL g3673 ( 
.A(n_3042),
.B(n_2342),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_2343),
.B(n_2596),
.Y(n_3674)
);

NAND2xp5_ASAP7_75t_L g3675 ( 
.A(n_2408),
.B(n_2479),
.Y(n_3675)
);

NOR2xp33_ASAP7_75t_L g3676 ( 
.A(n_2505),
.B(n_2645),
.Y(n_3676)
);

OAI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_2692),
.A2(n_2710),
.B1(n_2294),
.B2(n_2291),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_2159),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_SL g3679 ( 
.A(n_2291),
.B(n_2294),
.Y(n_3679)
);

AOI21x1_ASAP7_75t_L g3680 ( 
.A1(n_2182),
.A2(n_2852),
.B(n_2727),
.Y(n_3680)
);

AOI21xp5_ASAP7_75t_L g3681 ( 
.A1(n_2727),
.A2(n_2852),
.B(n_2906),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_2727),
.A2(n_2852),
.B(n_2863),
.Y(n_3682)
);

CKINVDCx10_ASAP7_75t_R g3683 ( 
.A(n_2660),
.Y(n_3683)
);

BUFx2_ASAP7_75t_SL g3684 ( 
.A(n_2401),
.Y(n_3684)
);

INVx1_ASAP7_75t_L g3685 ( 
.A(n_2443),
.Y(n_3685)
);

AND2x4_ASAP7_75t_L g3686 ( 
.A(n_2465),
.B(n_2488),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_2215),
.Y(n_3687)
);

O2A1O1Ixp33_ASAP7_75t_L g3688 ( 
.A1(n_2610),
.A2(n_2700),
.B(n_2803),
.C(n_2969),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_L g3689 ( 
.A(n_2228),
.B(n_2387),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3690)
);

INVx4_ASAP7_75t_L g3691 ( 
.A(n_2214),
.Y(n_3691)
);

NOR2xp33_ASAP7_75t_L g3692 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3692)
);

NAND2xp5_ASAP7_75t_L g3693 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3694)
);

NAND2xp5_ASAP7_75t_SL g3695 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3696)
);

OAI21xp5_ASAP7_75t_L g3697 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3697)
);

HB1xp67_ASAP7_75t_L g3698 ( 
.A(n_2049),
.Y(n_3698)
);

OAI21xp5_ASAP7_75t_L g3699 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3699)
);

INVx1_ASAP7_75t_L g3700 ( 
.A(n_2280),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3701)
);

OAI21xp5_ASAP7_75t_L g3702 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_L g3703 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_2280),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_2280),
.Y(n_3705)
);

AOI21xp33_ASAP7_75t_L g3706 ( 
.A1(n_2114),
.A2(n_2682),
.B(n_2619),
.Y(n_3706)
);

AOI21xp5_ASAP7_75t_L g3707 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3708)
);

CKINVDCx5p33_ASAP7_75t_R g3709 ( 
.A(n_2370),
.Y(n_3709)
);

AOI21xp5_ASAP7_75t_L g3710 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_SL g3712 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3712)
);

INVx2_ASAP7_75t_SL g3713 ( 
.A(n_2214),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_L g3714 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3714)
);

AOI21xp5_ASAP7_75t_L g3715 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3715)
);

OAI21xp5_ASAP7_75t_L g3716 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3716)
);

A2O1A1Ixp33_ASAP7_75t_L g3717 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3718)
);

BUFx6f_ASAP7_75t_L g3719 ( 
.A(n_2192),
.Y(n_3719)
);

AOI21x1_ASAP7_75t_L g3720 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_3720)
);

AOI21xp5_ASAP7_75t_L g3721 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3721)
);

INVxp67_ASAP7_75t_L g3722 ( 
.A(n_2049),
.Y(n_3722)
);

AO21x1_ASAP7_75t_L g3723 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_2100),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_L g3724 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3724)
);

AOI21xp5_ASAP7_75t_L g3725 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3725)
);

AOI21xp5_ASAP7_75t_L g3726 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3726)
);

OAI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3728)
);

NOR2xp33_ASAP7_75t_L g3729 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3730)
);

NOR2xp33_ASAP7_75t_L g3731 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3732)
);

NOR2xp33_ASAP7_75t_SL g3733 ( 
.A(n_2778),
.B(n_1653),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3734)
);

AOI21xp5_ASAP7_75t_L g3735 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3735)
);

NOR2xp33_ASAP7_75t_L g3736 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3738)
);

HB1xp67_ASAP7_75t_L g3739 ( 
.A(n_2049),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_2280),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_SL g3744 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3744)
);

AOI21xp5_ASAP7_75t_L g3745 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3748)
);

O2A1O1Ixp33_ASAP7_75t_SL g3749 ( 
.A1(n_2628),
.A2(n_1648),
.B(n_1630),
.C(n_2362),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_3750)
);

AO21x1_ASAP7_75t_L g3751 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_2100),
.Y(n_3751)
);

AOI22xp5_ASAP7_75t_L g3752 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3752)
);

HB1xp67_ASAP7_75t_L g3753 ( 
.A(n_2049),
.Y(n_3753)
);

AOI21xp5_ASAP7_75t_L g3754 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3754)
);

NOR2xp33_ASAP7_75t_L g3755 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3755)
);

NAND2xp5_ASAP7_75t_L g3756 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3757)
);

AOI21xp5_ASAP7_75t_L g3758 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3758)
);

O2A1O1Ixp5_ASAP7_75t_L g3759 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_3759)
);

INVx2_ASAP7_75t_L g3760 ( 
.A(n_2280),
.Y(n_3760)
);

AOI22xp5_ASAP7_75t_L g3761 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_L g3762 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3762)
);

INVxp67_ASAP7_75t_L g3763 ( 
.A(n_2049),
.Y(n_3763)
);

BUFx6f_ASAP7_75t_L g3764 ( 
.A(n_2192),
.Y(n_3764)
);

NAND2xp5_ASAP7_75t_L g3765 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3765)
);

NAND2x1_ASAP7_75t_L g3766 ( 
.A(n_2039),
.B(n_2086),
.Y(n_3766)
);

AOI22xp5_ASAP7_75t_L g3767 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3767)
);

AOI21x1_ASAP7_75t_L g3768 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3769)
);

O2A1O1Ixp33_ASAP7_75t_L g3770 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_3770)
);

AOI21xp5_ASAP7_75t_L g3771 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3771)
);

HB1xp67_ASAP7_75t_L g3772 ( 
.A(n_2049),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_L g3774 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3774)
);

AOI21xp5_ASAP7_75t_L g3775 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_2280),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_L g3781 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3781)
);

A2O1A1Ixp33_ASAP7_75t_L g3782 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_3782)
);

O2A1O1Ixp5_ASAP7_75t_L g3783 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_3783)
);

NAND2xp5_ASAP7_75t_L g3784 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3784)
);

OAI21xp5_ASAP7_75t_L g3785 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3786)
);

AOI21xp5_ASAP7_75t_L g3787 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_L g3788 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3788)
);

O2A1O1Ixp33_ASAP7_75t_L g3789 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_3789)
);

AOI21xp5_ASAP7_75t_L g3790 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3790)
);

A2O1A1Ixp33_ASAP7_75t_L g3791 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3794)
);

NAND2xp5_ASAP7_75t_L g3795 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3796)
);

AOI21x1_ASAP7_75t_L g3797 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_3797)
);

AOI21xp5_ASAP7_75t_L g3798 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3798)
);

NAND2xp5_ASAP7_75t_SL g3799 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3800)
);

OAI21x1_ASAP7_75t_L g3801 ( 
.A1(n_2138),
.A2(n_1968),
.B(n_846),
.Y(n_3801)
);

AND2x4_ASAP7_75t_L g3802 ( 
.A(n_2047),
.B(n_2059),
.Y(n_3802)
);

CKINVDCx5p33_ASAP7_75t_R g3803 ( 
.A(n_2370),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3804)
);

AOI22xp5_ASAP7_75t_L g3805 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3805)
);

AOI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3806)
);

AND2x2_ASAP7_75t_L g3807 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3807)
);

OAI21xp33_ASAP7_75t_L g3808 ( 
.A1(n_2623),
.A2(n_1246),
.B(n_1244),
.Y(n_3808)
);

OR2x2_ASAP7_75t_L g3809 ( 
.A(n_1957),
.B(n_2079),
.Y(n_3809)
);

OAI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3810)
);

INVxp67_ASAP7_75t_L g3811 ( 
.A(n_2049),
.Y(n_3811)
);

NOR2xp33_ASAP7_75t_L g3812 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3812)
);

AOI211xp5_ASAP7_75t_L g3813 ( 
.A1(n_2373),
.A2(n_2417),
.B(n_2428),
.C(n_2392),
.Y(n_3813)
);

NOR2xp33_ASAP7_75t_L g3814 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3814)
);

AOI21xp5_ASAP7_75t_L g3815 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3816)
);

O2A1O1Ixp33_ASAP7_75t_L g3817 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_3817)
);

NAND2xp5_ASAP7_75t_L g3818 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3820)
);

OAI22xp5_ASAP7_75t_L g3821 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3821)
);

AOI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3823)
);

AOI21xp5_ASAP7_75t_L g3824 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3824)
);

AOI21xp5_ASAP7_75t_L g3825 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3825)
);

AOI22xp5_ASAP7_75t_L g3826 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3827)
);

NAND2xp5_ASAP7_75t_L g3828 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_SL g3829 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3829)
);

NAND2xp5_ASAP7_75t_L g3830 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3830)
);

AOI21xp5_ASAP7_75t_L g3831 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3831)
);

O2A1O1Ixp5_ASAP7_75t_L g3832 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_3832)
);

AOI21xp5_ASAP7_75t_L g3833 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3833)
);

AOI22xp5_ASAP7_75t_L g3834 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3834)
);

HB1xp67_ASAP7_75t_L g3835 ( 
.A(n_2049),
.Y(n_3835)
);

NOR2xp33_ASAP7_75t_L g3836 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_2280),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3838)
);

OAI22x1_ASAP7_75t_L g3839 ( 
.A1(n_2376),
.A2(n_2383),
.B1(n_2507),
.B2(n_2388),
.Y(n_3839)
);

AOI21xp5_ASAP7_75t_L g3840 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3841)
);

NOR2xp33_ASAP7_75t_L g3842 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3842)
);

NAND2xp5_ASAP7_75t_L g3843 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3843)
);

AND2x2_ASAP7_75t_L g3844 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3844)
);

NOR3xp33_ASAP7_75t_L g3845 ( 
.A(n_1942),
.B(n_1014),
.C(n_1004),
.Y(n_3845)
);

AOI21xp5_ASAP7_75t_L g3846 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3846)
);

BUFx2_ASAP7_75t_L g3847 ( 
.A(n_2142),
.Y(n_3847)
);

INVx4_ASAP7_75t_L g3848 ( 
.A(n_2214),
.Y(n_3848)
);

AOI21xp5_ASAP7_75t_L g3849 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3849)
);

BUFx4f_ASAP7_75t_L g3850 ( 
.A(n_2192),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3851)
);

AOI22xp33_ASAP7_75t_L g3852 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_3852)
);

AOI21xp5_ASAP7_75t_L g3853 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3853)
);

NOR3xp33_ASAP7_75t_L g3854 ( 
.A(n_1942),
.B(n_1014),
.C(n_1004),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3855)
);

BUFx3_ASAP7_75t_L g3856 ( 
.A(n_2394),
.Y(n_3856)
);

AOI21xp5_ASAP7_75t_L g3857 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_2280),
.Y(n_3858)
);

AOI21xp5_ASAP7_75t_L g3859 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3859)
);

HB1xp67_ASAP7_75t_L g3860 ( 
.A(n_2049),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3862)
);

NOR2xp33_ASAP7_75t_L g3863 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3863)
);

INVxp67_ASAP7_75t_L g3864 ( 
.A(n_2049),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_L g3865 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3865)
);

AOI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3866)
);

AOI21xp5_ASAP7_75t_L g3867 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3867)
);

NAND2xp5_ASAP7_75t_L g3868 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3868)
);

INVx3_ASAP7_75t_L g3869 ( 
.A(n_2027),
.Y(n_3869)
);

OAI22xp5_ASAP7_75t_L g3870 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3870)
);

AOI21xp5_ASAP7_75t_L g3871 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3871)
);

AND2x2_ASAP7_75t_L g3872 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3872)
);

AOI21xp5_ASAP7_75t_L g3873 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3873)
);

O2A1O1Ixp5_ASAP7_75t_L g3874 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_3874)
);

BUFx6f_ASAP7_75t_L g3875 ( 
.A(n_2192),
.Y(n_3875)
);

NOR2xp33_ASAP7_75t_L g3876 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3876)
);

NOR2xp33_ASAP7_75t_L g3877 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3877)
);

AOI21xp5_ASAP7_75t_L g3878 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3878)
);

AND2x6_ASAP7_75t_L g3879 ( 
.A(n_1946),
.B(n_2278),
.Y(n_3879)
);

OAI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_SL g3881 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3882)
);

INVx11_ASAP7_75t_L g3883 ( 
.A(n_2249),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3884)
);

AOI21xp5_ASAP7_75t_L g3885 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_2280),
.Y(n_3886)
);

NAND2xp5_ASAP7_75t_L g3887 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3887)
);

AOI21xp5_ASAP7_75t_L g3888 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3888)
);

NAND2xp33_ASAP7_75t_L g3889 ( 
.A(n_1949),
.B(n_1630),
.Y(n_3889)
);

AOI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3890)
);

AND2x4_ASAP7_75t_L g3891 ( 
.A(n_2047),
.B(n_2059),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3893)
);

AOI21xp5_ASAP7_75t_L g3894 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3894)
);

BUFx6f_ASAP7_75t_L g3895 ( 
.A(n_2192),
.Y(n_3895)
);

OAI321xp33_ASAP7_75t_L g3896 ( 
.A1(n_2373),
.A2(n_1668),
.A3(n_2428),
.B1(n_2514),
.B2(n_2417),
.C(n_2392),
.Y(n_3896)
);

AOI22xp33_ASAP7_75t_SL g3897 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_2392),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3898)
);

AOI21xp5_ASAP7_75t_L g3899 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3899)
);

OAI21xp5_ASAP7_75t_L g3900 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3900)
);

AOI22xp5_ASAP7_75t_L g3901 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3901)
);

AOI21xp5_ASAP7_75t_L g3902 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3902)
);

NOR2xp33_ASAP7_75t_L g3903 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3903)
);

AOI21xp5_ASAP7_75t_L g3904 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3904)
);

AOI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3905)
);

INVx3_ASAP7_75t_L g3906 ( 
.A(n_2027),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3907)
);

HB1xp67_ASAP7_75t_L g3908 ( 
.A(n_2049),
.Y(n_3908)
);

AO21x1_ASAP7_75t_L g3909 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_2100),
.Y(n_3909)
);

AOI21xp5_ASAP7_75t_L g3910 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3910)
);

INVxp67_ASAP7_75t_L g3911 ( 
.A(n_2049),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3912)
);

AOI21xp5_ASAP7_75t_L g3913 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3913)
);

INVx2_ASAP7_75t_L g3914 ( 
.A(n_2280),
.Y(n_3914)
);

OAI21xp5_ASAP7_75t_L g3915 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3915)
);

NOR2xp33_ASAP7_75t_SL g3916 ( 
.A(n_2778),
.B(n_1653),
.Y(n_3916)
);

OAI22xp5_ASAP7_75t_L g3917 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3917)
);

INVx1_ASAP7_75t_SL g3918 ( 
.A(n_2139),
.Y(n_3918)
);

OAI21xp5_ASAP7_75t_L g3919 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_L g3920 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_L g3922 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3922)
);

AOI21xp5_ASAP7_75t_L g3923 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_L g3925 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3925)
);

INVx2_ASAP7_75t_SL g3926 ( 
.A(n_2214),
.Y(n_3926)
);

AOI22xp33_ASAP7_75t_L g3927 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3929)
);

AOI22xp5_ASAP7_75t_L g3930 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3930)
);

AOI21xp5_ASAP7_75t_L g3931 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3931)
);

OAI21xp5_ASAP7_75t_L g3932 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3932)
);

A2O1A1Ixp33_ASAP7_75t_L g3933 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_3933)
);

AND2x2_ASAP7_75t_L g3934 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3934)
);

NOR2xp33_ASAP7_75t_L g3935 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3935)
);

AOI21xp5_ASAP7_75t_L g3936 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3936)
);

AOI21x1_ASAP7_75t_L g3937 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_3937)
);

OAI21xp5_ASAP7_75t_L g3938 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3938)
);

NOR2xp33_ASAP7_75t_L g3939 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3939)
);

NOR2xp33_ASAP7_75t_L g3940 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3940)
);

INVx4_ASAP7_75t_L g3941 ( 
.A(n_2214),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3942)
);

AOI21xp5_ASAP7_75t_L g3943 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3943)
);

NOR2xp33_ASAP7_75t_L g3944 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3945)
);

AOI21xp5_ASAP7_75t_L g3946 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3946)
);

O2A1O1Ixp33_ASAP7_75t_L g3947 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_3947)
);

CKINVDCx10_ASAP7_75t_R g3948 ( 
.A(n_2650),
.Y(n_3948)
);

OAI22xp5_ASAP7_75t_L g3949 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_L g3950 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3950)
);

AOI21xp5_ASAP7_75t_L g3951 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_2192),
.Y(n_3952)
);

AND2x4_ASAP7_75t_L g3953 ( 
.A(n_2047),
.B(n_2059),
.Y(n_3953)
);

AOI22xp5_ASAP7_75t_L g3954 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3954)
);

AND2x4_ASAP7_75t_L g3955 ( 
.A(n_2047),
.B(n_2059),
.Y(n_3955)
);

OAI22xp5_ASAP7_75t_L g3956 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3956)
);

O2A1O1Ixp33_ASAP7_75t_L g3957 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3958)
);

OAI21xp5_ASAP7_75t_L g3959 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3959)
);

AND2x2_ASAP7_75t_SL g3960 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3960)
);

HB1xp67_ASAP7_75t_L g3961 ( 
.A(n_2049),
.Y(n_3961)
);

AOI21xp5_ASAP7_75t_L g3962 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3962)
);

OAI21xp5_ASAP7_75t_L g3963 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3963)
);

INVx3_ASAP7_75t_L g3964 ( 
.A(n_2027),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_L g3966 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3966)
);

AOI22xp5_ASAP7_75t_L g3967 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_L g3968 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3968)
);

AND2x4_ASAP7_75t_L g3969 ( 
.A(n_2047),
.B(n_2059),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3970)
);

NOR2xp33_ASAP7_75t_L g3971 ( 
.A(n_2836),
.B(n_1954),
.Y(n_3971)
);

AOI21xp5_ASAP7_75t_L g3972 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3972)
);

A2O1A1Ixp33_ASAP7_75t_L g3973 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3974)
);

AOI21xp5_ASAP7_75t_L g3975 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3975)
);

AOI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3976)
);

AND2x4_ASAP7_75t_L g3977 ( 
.A(n_2047),
.B(n_2059),
.Y(n_3977)
);

AOI21xp5_ASAP7_75t_L g3978 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3978)
);

AND2x2_ASAP7_75t_SL g3979 ( 
.A(n_2485),
.B(n_2594),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3980)
);

O2A1O1Ixp33_ASAP7_75t_L g3981 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_L g3982 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3984)
);

OAI21xp5_ASAP7_75t_L g3985 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_3985)
);

AOI21xp33_ASAP7_75t_L g3986 ( 
.A1(n_2114),
.A2(n_2682),
.B(n_2619),
.Y(n_3986)
);

AOI21xp5_ASAP7_75t_L g3987 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3987)
);

AOI21xp5_ASAP7_75t_L g3988 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3988)
);

HB1xp67_ASAP7_75t_L g3989 ( 
.A(n_2049),
.Y(n_3989)
);

AOI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3990)
);

AOI21xp5_ASAP7_75t_L g3991 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3991)
);

AOI21xp5_ASAP7_75t_L g3992 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_1961),
.B(n_2021),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_2387),
.B(n_2754),
.Y(n_3996)
);

INVx4_ASAP7_75t_L g3997 ( 
.A(n_2214),
.Y(n_3997)
);

INVx3_ASAP7_75t_L g3998 ( 
.A(n_2027),
.Y(n_3998)
);

INVx4_ASAP7_75t_L g3999 ( 
.A(n_2214),
.Y(n_3999)
);

INVx3_ASAP7_75t_L g4000 ( 
.A(n_2027),
.Y(n_4000)
);

NOR3xp33_ASAP7_75t_L g4001 ( 
.A(n_1942),
.B(n_1014),
.C(n_1004),
.Y(n_4001)
);

AOI21xp5_ASAP7_75t_L g4002 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4002)
);

BUFx8_ASAP7_75t_L g4003 ( 
.A(n_2650),
.Y(n_4003)
);

AOI21xp5_ASAP7_75t_L g4004 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4004)
);

A2O1A1Ixp33_ASAP7_75t_L g4005 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_4005)
);

AOI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4006)
);

INVx1_ASAP7_75t_SL g4007 ( 
.A(n_2139),
.Y(n_4007)
);

INVx3_ASAP7_75t_L g4008 ( 
.A(n_2027),
.Y(n_4008)
);

OAI21xp5_ASAP7_75t_L g4009 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4009)
);

HB1xp67_ASAP7_75t_L g4010 ( 
.A(n_2049),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_L g4011 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4011)
);

NOR2xp67_ASAP7_75t_L g4012 ( 
.A(n_2227),
.B(n_1597),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_L g4014 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4014)
);

AOI21xp5_ASAP7_75t_L g4015 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4015)
);

NOR2xp33_ASAP7_75t_L g4016 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4016)
);

AOI21xp5_ASAP7_75t_L g4017 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4017)
);

O2A1O1Ixp5_ASAP7_75t_L g4018 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_4018)
);

INVx3_ASAP7_75t_L g4019 ( 
.A(n_2027),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_2280),
.Y(n_4020)
);

BUFx6f_ASAP7_75t_L g4021 ( 
.A(n_2192),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4022)
);

O2A1O1Ixp5_ASAP7_75t_L g4023 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_4023)
);

AOI22xp33_ASAP7_75t_L g4024 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_4024)
);

NAND3xp33_ASAP7_75t_L g4025 ( 
.A(n_2623),
.B(n_1014),
.C(n_1004),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4026)
);

AOI21xp5_ASAP7_75t_L g4027 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4028)
);

NOR2x1_ASAP7_75t_L g4029 ( 
.A(n_2062),
.B(n_2093),
.Y(n_4029)
);

AOI21xp5_ASAP7_75t_L g4030 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4030)
);

HB1xp67_ASAP7_75t_L g4031 ( 
.A(n_2049),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4032)
);

AOI21xp5_ASAP7_75t_L g4033 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4033)
);

INVx5_ASAP7_75t_L g4034 ( 
.A(n_2039),
.Y(n_4034)
);

AOI21xp5_ASAP7_75t_L g4035 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_2280),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_L g4039 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_SL g4040 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4040)
);

BUFx6f_ASAP7_75t_L g4041 ( 
.A(n_2192),
.Y(n_4041)
);

INVx1_ASAP7_75t_SL g4042 ( 
.A(n_2139),
.Y(n_4042)
);

AOI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4044)
);

INVx2_ASAP7_75t_SL g4045 ( 
.A(n_2214),
.Y(n_4045)
);

NAND3xp33_ASAP7_75t_SL g4046 ( 
.A(n_2623),
.B(n_2736),
.C(n_1942),
.Y(n_4046)
);

AOI21xp5_ASAP7_75t_L g4047 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4047)
);

NOR2xp33_ASAP7_75t_L g4048 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4048)
);

INVx2_ASAP7_75t_SL g4049 ( 
.A(n_2214),
.Y(n_4049)
);

NOR2xp33_ASAP7_75t_L g4050 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4050)
);

BUFx6f_ASAP7_75t_L g4051 ( 
.A(n_2192),
.Y(n_4051)
);

NAND2xp5_ASAP7_75t_L g4052 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_L g4053 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_L g4055 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4055)
);

AOI21x1_ASAP7_75t_L g4056 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_4056)
);

NOR2xp33_ASAP7_75t_L g4057 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4058)
);

O2A1O1Ixp33_ASAP7_75t_L g4059 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4059)
);

INVxp67_ASAP7_75t_L g4060 ( 
.A(n_2049),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4061)
);

OAI21xp5_ASAP7_75t_L g4062 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4062)
);

OAI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4064)
);

INVxp67_ASAP7_75t_L g4065 ( 
.A(n_2049),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4066)
);

INVx3_ASAP7_75t_L g4067 ( 
.A(n_2027),
.Y(n_4067)
);

NOR2xp67_ASAP7_75t_L g4068 ( 
.A(n_2227),
.B(n_1597),
.Y(n_4068)
);

AND2x2_ASAP7_75t_L g4069 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4069)
);

AOI21xp5_ASAP7_75t_L g4070 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4070)
);

BUFx6f_ASAP7_75t_L g4071 ( 
.A(n_2192),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4073)
);

BUFx4f_ASAP7_75t_L g4074 ( 
.A(n_2192),
.Y(n_4074)
);

OAI22xp5_ASAP7_75t_L g4075 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4075)
);

AOI21xp5_ASAP7_75t_L g4076 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4076)
);

INVxp67_ASAP7_75t_L g4077 ( 
.A(n_2049),
.Y(n_4077)
);

NOR2xp33_ASAP7_75t_R g4078 ( 
.A(n_2313),
.B(n_830),
.Y(n_4078)
);

HB1xp67_ASAP7_75t_L g4079 ( 
.A(n_2049),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4080)
);

AOI21xp5_ASAP7_75t_L g4081 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4081)
);

AOI21xp5_ASAP7_75t_L g4082 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4082)
);

AOI21xp5_ASAP7_75t_L g4083 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4083)
);

OAI22xp5_ASAP7_75t_L g4084 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4084)
);

AND2x2_ASAP7_75t_L g4085 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4085)
);

BUFx6f_ASAP7_75t_L g4086 ( 
.A(n_2192),
.Y(n_4086)
);

OAI22xp5_ASAP7_75t_L g4087 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_L g4088 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4088)
);

AOI22xp5_ASAP7_75t_L g4089 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4089)
);

CKINVDCx6p67_ASAP7_75t_R g4090 ( 
.A(n_2214),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4091)
);

AOI21xp5_ASAP7_75t_L g4092 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4092)
);

NAND2xp5_ASAP7_75t_L g4093 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_L g4094 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4094)
);

NOR2xp33_ASAP7_75t_L g4095 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4095)
);

NAND2xp5_ASAP7_75t_L g4096 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4096)
);

OAI21xp5_ASAP7_75t_L g4097 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4098)
);

OAI22xp33_ASAP7_75t_SL g4099 ( 
.A1(n_1985),
.A2(n_1971),
.B1(n_1668),
.B2(n_1257),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_SL g4100 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_L g4101 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4101)
);

AOI21xp5_ASAP7_75t_L g4102 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_SL g4103 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4103)
);

AOI22xp5_ASAP7_75t_L g4104 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4104)
);

AOI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4106)
);

NOR2xp33_ASAP7_75t_L g4107 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4107)
);

NOR2xp33_ASAP7_75t_L g4108 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4108)
);

BUFx3_ASAP7_75t_L g4109 ( 
.A(n_2394),
.Y(n_4109)
);

HB1xp67_ASAP7_75t_L g4110 ( 
.A(n_2049),
.Y(n_4110)
);

INVx2_ASAP7_75t_L g4111 ( 
.A(n_2280),
.Y(n_4111)
);

AOI21xp5_ASAP7_75t_L g4112 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4112)
);

OAI22xp5_ASAP7_75t_L g4113 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4116)
);

A2O1A1Ixp33_ASAP7_75t_L g4117 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_4117)
);

OAI21xp5_ASAP7_75t_L g4118 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4118)
);

AOI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4119)
);

BUFx2_ASAP7_75t_L g4120 ( 
.A(n_2142),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_L g4121 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4121)
);

AOI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4124)
);

OAI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4125)
);

INVx2_ASAP7_75t_SL g4126 ( 
.A(n_2214),
.Y(n_4126)
);

AOI21xp5_ASAP7_75t_L g4127 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4127)
);

AOI222xp33_ASAP7_75t_L g4128 ( 
.A1(n_1942),
.A2(n_2736),
.B1(n_2428),
.B2(n_2392),
.C1(n_2514),
.C2(n_2417),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_L g4129 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_L g4130 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4130)
);

OAI21xp33_ASAP7_75t_L g4131 ( 
.A1(n_2623),
.A2(n_1246),
.B(n_1244),
.Y(n_4131)
);

INVx2_ASAP7_75t_L g4132 ( 
.A(n_2280),
.Y(n_4132)
);

OAI22x1_ASAP7_75t_L g4133 ( 
.A1(n_2376),
.A2(n_2383),
.B1(n_2507),
.B2(n_2388),
.Y(n_4133)
);

INVx2_ASAP7_75t_L g4134 ( 
.A(n_2280),
.Y(n_4134)
);

INVx2_ASAP7_75t_L g4135 ( 
.A(n_2280),
.Y(n_4135)
);

AND2x2_ASAP7_75t_L g4136 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4136)
);

AOI21xp5_ASAP7_75t_L g4137 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4137)
);

CKINVDCx5p33_ASAP7_75t_R g4138 ( 
.A(n_2370),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4139)
);

AOI21xp5_ASAP7_75t_L g4140 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4140)
);

AOI21xp5_ASAP7_75t_L g4141 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4141)
);

CKINVDCx5p33_ASAP7_75t_R g4142 ( 
.A(n_2370),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4143)
);

AND2x4_ASAP7_75t_L g4144 ( 
.A(n_2047),
.B(n_2059),
.Y(n_4144)
);

INVxp67_ASAP7_75t_L g4145 ( 
.A(n_2049),
.Y(n_4145)
);

OR2x2_ASAP7_75t_L g4146 ( 
.A(n_1957),
.B(n_2079),
.Y(n_4146)
);

INVx3_ASAP7_75t_L g4147 ( 
.A(n_2027),
.Y(n_4147)
);

NOR2xp33_ASAP7_75t_L g4148 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4148)
);

INVx2_ASAP7_75t_SL g4149 ( 
.A(n_2214),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4150)
);

AOI22xp33_ASAP7_75t_L g4151 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_SL g4152 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4152)
);

AOI21xp5_ASAP7_75t_L g4153 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4153)
);

BUFx6f_ASAP7_75t_L g4154 ( 
.A(n_2192),
.Y(n_4154)
);

AOI21xp5_ASAP7_75t_L g4155 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4155)
);

NAND2xp5_ASAP7_75t_L g4156 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4156)
);

O2A1O1Ixp33_ASAP7_75t_L g4157 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_L g4158 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4158)
);

INVx2_ASAP7_75t_L g4159 ( 
.A(n_2280),
.Y(n_4159)
);

INVxp67_ASAP7_75t_L g4160 ( 
.A(n_2049),
.Y(n_4160)
);

OAI21xp33_ASAP7_75t_L g4161 ( 
.A1(n_2623),
.A2(n_1246),
.B(n_1244),
.Y(n_4161)
);

AOI21xp5_ASAP7_75t_L g4162 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4163)
);

AOI211xp5_ASAP7_75t_L g4164 ( 
.A1(n_2373),
.A2(n_2417),
.B(n_2428),
.C(n_2392),
.Y(n_4164)
);

AOI21xp5_ASAP7_75t_L g4165 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4165)
);

NOR2xp33_ASAP7_75t_L g4166 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4166)
);

NAND2x1p5_ASAP7_75t_L g4167 ( 
.A(n_2093),
.B(n_2100),
.Y(n_4167)
);

OAI22xp5_ASAP7_75t_L g4168 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4168)
);

HB1xp67_ASAP7_75t_L g4169 ( 
.A(n_2049),
.Y(n_4169)
);

BUFx6f_ASAP7_75t_L g4170 ( 
.A(n_2192),
.Y(n_4170)
);

O2A1O1Ixp5_ASAP7_75t_L g4171 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_4171)
);

AOI21xp5_ASAP7_75t_L g4172 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_2280),
.Y(n_4174)
);

AOI22xp33_ASAP7_75t_L g4175 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4177)
);

AOI21xp5_ASAP7_75t_L g4178 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4178)
);

AOI22xp5_ASAP7_75t_L g4179 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4179)
);

AOI22xp5_ASAP7_75t_L g4180 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4180)
);

INVx4_ASAP7_75t_L g4181 ( 
.A(n_2214),
.Y(n_4181)
);

INVx1_ASAP7_75t_L g4182 ( 
.A(n_2280),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4183)
);

OAI22xp5_ASAP7_75t_L g4184 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_SL g4185 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4186)
);

NAND2xp5_ASAP7_75t_SL g4187 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4187)
);

BUFx3_ASAP7_75t_L g4188 ( 
.A(n_2394),
.Y(n_4188)
);

AOI21xp5_ASAP7_75t_L g4189 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4189)
);

AOI22xp33_ASAP7_75t_L g4190 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_4190)
);

A2O1A1Ixp33_ASAP7_75t_L g4191 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_4191)
);

OAI21xp5_ASAP7_75t_L g4192 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4192)
);

A2O1A1Ixp33_ASAP7_75t_L g4193 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4194)
);

AOI21xp5_ASAP7_75t_L g4195 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4195)
);

INVxp67_ASAP7_75t_L g4196 ( 
.A(n_2049),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_2280),
.Y(n_4197)
);

NAND2xp5_ASAP7_75t_L g4198 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4198)
);

AOI22xp5_ASAP7_75t_L g4199 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4201)
);

OAI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4203)
);

AOI21xp5_ASAP7_75t_L g4204 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4204)
);

AOI21xp33_ASAP7_75t_L g4205 ( 
.A1(n_2114),
.A2(n_2682),
.B(n_2619),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4206)
);

AOI22xp33_ASAP7_75t_SL g4207 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_2392),
.Y(n_4207)
);

A2O1A1Ixp33_ASAP7_75t_L g4208 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4209)
);

BUFx2_ASAP7_75t_L g4210 ( 
.A(n_2142),
.Y(n_4210)
);

O2A1O1Ixp33_ASAP7_75t_SL g4211 ( 
.A1(n_2628),
.A2(n_1648),
.B(n_1630),
.C(n_2362),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_SL g4212 ( 
.A(n_2778),
.B(n_1653),
.Y(n_4212)
);

OR2x2_ASAP7_75t_L g4213 ( 
.A(n_1957),
.B(n_2079),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_2280),
.Y(n_4214)
);

A2O1A1Ixp33_ASAP7_75t_L g4215 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_4215)
);

INVx2_ASAP7_75t_SL g4216 ( 
.A(n_2214),
.Y(n_4216)
);

AOI21xp33_ASAP7_75t_L g4217 ( 
.A1(n_2114),
.A2(n_2682),
.B(n_2619),
.Y(n_4217)
);

AOI22xp5_ASAP7_75t_L g4218 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4218)
);

AND2x4_ASAP7_75t_L g4219 ( 
.A(n_2047),
.B(n_2059),
.Y(n_4219)
);

AOI22xp33_ASAP7_75t_L g4220 ( 
.A1(n_2485),
.A2(n_3006),
.B1(n_2594),
.B2(n_1561),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_L g4221 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4221)
);

AND2x2_ASAP7_75t_L g4222 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4222)
);

AOI21xp5_ASAP7_75t_L g4223 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4223)
);

A2O1A1Ixp33_ASAP7_75t_L g4224 ( 
.A1(n_2619),
.A2(n_1246),
.B(n_1262),
.C(n_1244),
.Y(n_4224)
);

O2A1O1Ixp5_ASAP7_75t_L g4225 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_4225)
);

AND2x2_ASAP7_75t_L g4226 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4226)
);

NOR2xp33_ASAP7_75t_L g4227 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4227)
);

AOI21xp5_ASAP7_75t_L g4228 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4228)
);

NAND2xp5_ASAP7_75t_L g4229 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4229)
);

NAND2xp5_ASAP7_75t_L g4230 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4230)
);

OAI21xp5_ASAP7_75t_L g4231 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4231)
);

NOR2xp33_ASAP7_75t_L g4232 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4232)
);

AOI21xp5_ASAP7_75t_L g4233 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4233)
);

BUFx2_ASAP7_75t_L g4234 ( 
.A(n_2142),
.Y(n_4234)
);

INVx1_ASAP7_75t_L g4235 ( 
.A(n_2280),
.Y(n_4235)
);

AOI21xp5_ASAP7_75t_L g4236 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4236)
);

BUFx3_ASAP7_75t_L g4237 ( 
.A(n_2394),
.Y(n_4237)
);

AOI21xp5_ASAP7_75t_L g4238 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4238)
);

AOI21xp5_ASAP7_75t_L g4239 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4239)
);

INVx2_ASAP7_75t_SL g4240 ( 
.A(n_2214),
.Y(n_4240)
);

NOR2xp33_ASAP7_75t_L g4241 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4241)
);

AOI21xp5_ASAP7_75t_L g4242 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4242)
);

NOR2xp33_ASAP7_75t_L g4243 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4243)
);

AO21x1_ASAP7_75t_L g4244 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_2100),
.Y(n_4244)
);

INVx3_ASAP7_75t_L g4245 ( 
.A(n_2027),
.Y(n_4245)
);

O2A1O1Ixp33_ASAP7_75t_L g4246 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4246)
);

AO21x1_ASAP7_75t_L g4247 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_2100),
.Y(n_4247)
);

O2A1O1Ixp33_ASAP7_75t_L g4248 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4248)
);

NAND2xp5_ASAP7_75t_L g4249 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4249)
);

NOR2xp33_ASAP7_75t_L g4250 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4250)
);

O2A1O1Ixp33_ASAP7_75t_L g4251 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4251)
);

AOI21x1_ASAP7_75t_L g4252 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_4252)
);

AOI21xp5_ASAP7_75t_L g4253 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4253)
);

AOI21xp5_ASAP7_75t_L g4254 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4254)
);

OAI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4256)
);

BUFx8_ASAP7_75t_L g4257 ( 
.A(n_2650),
.Y(n_4257)
);

AOI21xp5_ASAP7_75t_L g4258 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4258)
);

AOI21x1_ASAP7_75t_L g4259 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_4259)
);

AOI22xp5_ASAP7_75t_L g4260 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4260)
);

AOI21xp5_ASAP7_75t_L g4261 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4261)
);

NOR2xp33_ASAP7_75t_L g4262 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4262)
);

NOR2x1_ASAP7_75t_R g4263 ( 
.A(n_1979),
.B(n_572),
.Y(n_4263)
);

NAND3xp33_ASAP7_75t_L g4264 ( 
.A(n_2623),
.B(n_1014),
.C(n_1004),
.Y(n_4264)
);

AOI21xp5_ASAP7_75t_L g4265 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4265)
);

AOI21xp5_ASAP7_75t_L g4266 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4266)
);

BUFx3_ASAP7_75t_L g4267 ( 
.A(n_2394),
.Y(n_4267)
);

CKINVDCx10_ASAP7_75t_R g4268 ( 
.A(n_2650),
.Y(n_4268)
);

AOI21x1_ASAP7_75t_L g4269 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_4269)
);

O2A1O1Ixp33_ASAP7_75t_L g4270 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4270)
);

O2A1O1Ixp5_ASAP7_75t_L g4271 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_1274),
.C(n_2100),
.Y(n_4271)
);

AOI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4272)
);

OAI21xp5_ASAP7_75t_L g4273 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4273)
);

AND2x4_ASAP7_75t_L g4274 ( 
.A(n_2047),
.B(n_2059),
.Y(n_4274)
);

AOI21x1_ASAP7_75t_L g4275 ( 
.A1(n_2093),
.A2(n_2103),
.B(n_2100),
.Y(n_4275)
);

BUFx2_ASAP7_75t_SL g4276 ( 
.A(n_2214),
.Y(n_4276)
);

NOR2xp33_ASAP7_75t_L g4277 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4277)
);

AOI22xp5_ASAP7_75t_L g4278 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4278)
);

INVx3_ASAP7_75t_L g4279 ( 
.A(n_2027),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_SL g4280 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4280)
);

AOI21xp5_ASAP7_75t_L g4281 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4281)
);

NAND2xp5_ASAP7_75t_L g4282 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4282)
);

HB1xp67_ASAP7_75t_L g4283 ( 
.A(n_2049),
.Y(n_4283)
);

BUFx2_ASAP7_75t_L g4284 ( 
.A(n_2142),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_L g4286 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4288)
);

AOI21xp5_ASAP7_75t_L g4289 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4289)
);

INVx4_ASAP7_75t_L g4290 ( 
.A(n_2214),
.Y(n_4290)
);

AOI21xp5_ASAP7_75t_L g4291 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_2485),
.B(n_2594),
.Y(n_4293)
);

AOI21xp5_ASAP7_75t_L g4294 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4294)
);

OAI21xp33_ASAP7_75t_L g4295 ( 
.A1(n_2623),
.A2(n_1246),
.B(n_1244),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4297)
);

AOI21xp5_ASAP7_75t_L g4298 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4298)
);

AO21x1_ASAP7_75t_L g4299 ( 
.A1(n_2093),
.A2(n_1257),
.B(n_2100),
.Y(n_4299)
);

AOI21xp5_ASAP7_75t_L g4300 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4300)
);

AOI21xp33_ASAP7_75t_L g4301 ( 
.A1(n_2114),
.A2(n_2682),
.B(n_2619),
.Y(n_4301)
);

INVx2_ASAP7_75t_SL g4302 ( 
.A(n_2214),
.Y(n_4302)
);

INVx1_ASAP7_75t_L g4303 ( 
.A(n_2280),
.Y(n_4303)
);

OR2x2_ASAP7_75t_SL g4304 ( 
.A(n_2909),
.B(n_2974),
.Y(n_4304)
);

AOI21xp5_ASAP7_75t_L g4305 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4306)
);

OR2x2_ASAP7_75t_L g4307 ( 
.A(n_1957),
.B(n_2079),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_L g4308 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4309)
);

NAND2xp5_ASAP7_75t_L g4310 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4310)
);

NAND2xp5_ASAP7_75t_L g4311 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4311)
);

OAI22xp5_ASAP7_75t_L g4312 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4312)
);

AOI21xp5_ASAP7_75t_L g4313 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4313)
);

NAND2xp33_ASAP7_75t_SL g4314 ( 
.A(n_2370),
.B(n_2652),
.Y(n_4314)
);

AOI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4315)
);

NOR2xp33_ASAP7_75t_L g4316 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4316)
);

OAI22xp5_ASAP7_75t_L g4317 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4317)
);

NOR2xp33_ASAP7_75t_L g4318 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4318)
);

NAND2xp5_ASAP7_75t_L g4319 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4319)
);

AOI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4320)
);

BUFx6f_ASAP7_75t_L g4321 ( 
.A(n_2192),
.Y(n_4321)
);

AOI21xp5_ASAP7_75t_L g4322 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4322)
);

OAI21xp5_ASAP7_75t_L g4323 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4323)
);

OR2x2_ASAP7_75t_L g4324 ( 
.A(n_1957),
.B(n_2079),
.Y(n_4324)
);

AOI21xp5_ASAP7_75t_L g4325 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4325)
);

NOR2xp33_ASAP7_75t_L g4326 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4326)
);

OAI21xp5_ASAP7_75t_L g4327 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4327)
);

INVx2_ASAP7_75t_SL g4328 ( 
.A(n_2214),
.Y(n_4328)
);

AOI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_SL g4330 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4330)
);

NOR2xp33_ASAP7_75t_L g4331 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4332)
);

OAI21xp5_ASAP7_75t_L g4333 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_SL g4334 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4334)
);

AND2x4_ASAP7_75t_L g4335 ( 
.A(n_2047),
.B(n_2059),
.Y(n_4335)
);

INVx3_ASAP7_75t_L g4336 ( 
.A(n_2027),
.Y(n_4336)
);

AOI22xp5_ASAP7_75t_L g4337 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4337)
);

OR2x2_ASAP7_75t_L g4338 ( 
.A(n_1957),
.B(n_2079),
.Y(n_4338)
);

AOI21xp5_ASAP7_75t_L g4339 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4339)
);

O2A1O1Ixp33_ASAP7_75t_L g4340 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4340)
);

AOI22xp5_ASAP7_75t_L g4341 ( 
.A1(n_1954),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4341)
);

AOI21xp5_ASAP7_75t_L g4342 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4342)
);

NOR2xp33_ASAP7_75t_L g4343 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4343)
);

AOI21xp5_ASAP7_75t_L g4344 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4345)
);

NOR2xp33_ASAP7_75t_L g4346 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4346)
);

AOI21xp5_ASAP7_75t_L g4347 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4347)
);

AOI21xp5_ASAP7_75t_L g4348 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4348)
);

OAI22xp5_ASAP7_75t_L g4349 ( 
.A1(n_1947),
.A2(n_1246),
.B1(n_1262),
.B2(n_1244),
.Y(n_4349)
);

INVx11_ASAP7_75t_L g4350 ( 
.A(n_2249),
.Y(n_4350)
);

BUFx6f_ASAP7_75t_L g4351 ( 
.A(n_2192),
.Y(n_4351)
);

BUFx6f_ASAP7_75t_L g4352 ( 
.A(n_2192),
.Y(n_4352)
);

OAI21xp5_ASAP7_75t_L g4353 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4353)
);

NOR2xp33_ASAP7_75t_L g4354 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4354)
);

NOR3xp33_ASAP7_75t_L g4355 ( 
.A(n_1942),
.B(n_1014),
.C(n_1004),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_2280),
.Y(n_4356)
);

NOR3xp33_ASAP7_75t_L g4357 ( 
.A(n_1942),
.B(n_1014),
.C(n_1004),
.Y(n_4357)
);

OAI21xp33_ASAP7_75t_L g4358 ( 
.A1(n_2623),
.A2(n_1246),
.B(n_1244),
.Y(n_4358)
);

BUFx12f_ASAP7_75t_L g4359 ( 
.A(n_2427),
.Y(n_4359)
);

INVxp33_ASAP7_75t_SL g4360 ( 
.A(n_2370),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4361)
);

INVx3_ASAP7_75t_L g4362 ( 
.A(n_2027),
.Y(n_4362)
);

AND2x4_ASAP7_75t_L g4363 ( 
.A(n_2047),
.B(n_2059),
.Y(n_4363)
);

OAI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_2041),
.A2(n_2598),
.B(n_2456),
.Y(n_4364)
);

O2A1O1Ixp33_ASAP7_75t_L g4365 ( 
.A1(n_2362),
.A2(n_1648),
.B(n_1630),
.C(n_1668),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_2280),
.Y(n_4366)
);

NAND2xp5_ASAP7_75t_L g4367 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_SL g4368 ( 
.A(n_1961),
.B(n_2021),
.Y(n_4368)
);

NOR2xp33_ASAP7_75t_L g4369 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4369)
);

NAND2xp5_ASAP7_75t_L g4370 ( 
.A(n_2387),
.B(n_2754),
.Y(n_4370)
);

NOR2xp33_ASAP7_75t_L g4371 ( 
.A(n_2836),
.B(n_1954),
.Y(n_4371)
);

AOI21xp5_ASAP7_75t_L g4372 ( 
.A1(n_1999),
.A2(n_2482),
.B(n_2397),
.Y(n_4372)
);

BUFx6f_ASAP7_75t_L g4373 ( 
.A(n_4034),
.Y(n_4373)
);

INVx2_ASAP7_75t_L g4374 ( 
.A(n_3053),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4366),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4366),
.Y(n_4376)
);

NOR2xp33_ASAP7_75t_L g4377 ( 
.A(n_4046),
.B(n_3808),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_3051),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_3053),
.Y(n_4379)
);

NOR2xp33_ASAP7_75t_L g4380 ( 
.A(n_3808),
.B(n_4131),
.Y(n_4380)
);

INVx1_ASAP7_75t_L g4381 ( 
.A(n_3051),
.Y(n_4381)
);

INVx2_ASAP7_75t_SL g4382 ( 
.A(n_4034),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_3700),
.Y(n_4383)
);

NAND2xp5_ASAP7_75t_L g4384 ( 
.A(n_3092),
.B(n_3303),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_3741),
.Y(n_4385)
);

HB1xp67_ASAP7_75t_L g4386 ( 
.A(n_3065),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_3741),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_SL g4388 ( 
.A(n_4128),
.B(n_3061),
.Y(n_4388)
);

HB1xp67_ASAP7_75t_L g4389 ( 
.A(n_3065),
.Y(n_4389)
);

BUFx3_ASAP7_75t_L g4390 ( 
.A(n_3284),
.Y(n_4390)
);

A2O1A1Ixp33_ASAP7_75t_L g4391 ( 
.A1(n_3130),
.A2(n_3129),
.B(n_3095),
.C(n_3054),
.Y(n_4391)
);

AND2x4_ASAP7_75t_L g4392 ( 
.A(n_4034),
.B(n_3067),
.Y(n_4392)
);

NAND2xp5_ASAP7_75t_L g4393 ( 
.A(n_3092),
.B(n_3303),
.Y(n_4393)
);

AO21x1_ASAP7_75t_L g4394 ( 
.A1(n_4099),
.A2(n_3112),
.B(n_3069),
.Y(n_4394)
);

BUFx3_ASAP7_75t_L g4395 ( 
.A(n_3284),
.Y(n_4395)
);

AOI22xp33_ASAP7_75t_L g4396 ( 
.A1(n_3072),
.A2(n_4131),
.B1(n_4295),
.B2(n_4161),
.Y(n_4396)
);

AOI22xp5_ASAP7_75t_L g4397 ( 
.A1(n_4161),
.A2(n_4358),
.B1(n_4295),
.B2(n_3727),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_3140),
.B(n_3121),
.Y(n_4398)
);

INVx2_ASAP7_75t_SL g4399 ( 
.A(n_4034),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_3741),
.B(n_3760),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_3140),
.B(n_3121),
.Y(n_4401)
);

NOR2xp33_ASAP7_75t_L g4402 ( 
.A(n_4358),
.B(n_3727),
.Y(n_4402)
);

INVx1_ASAP7_75t_L g4403 ( 
.A(n_3700),
.Y(n_4403)
);

NAND2xp5_ASAP7_75t_L g4404 ( 
.A(n_3809),
.B(n_4146),
.Y(n_4404)
);

AOI22xp5_ASAP7_75t_L g4405 ( 
.A1(n_3821),
.A2(n_3870),
.B1(n_3912),
.B2(n_3880),
.Y(n_4405)
);

INVx2_ASAP7_75t_L g4406 ( 
.A(n_3760),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_3704),
.Y(n_4407)
);

NAND2xp5_ASAP7_75t_L g4408 ( 
.A(n_3809),
.B(n_4146),
.Y(n_4408)
);

AOI22xp5_ASAP7_75t_L g4409 ( 
.A1(n_3821),
.A2(n_3870),
.B1(n_3912),
.B2(n_3880),
.Y(n_4409)
);

OR2x6_ASAP7_75t_L g4410 ( 
.A(n_3060),
.B(n_3066),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_3760),
.Y(n_4411)
);

INVx4_ASAP7_75t_L g4412 ( 
.A(n_3505),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_SL g4413 ( 
.A(n_4128),
.B(n_3061),
.Y(n_4413)
);

AND2x4_ASAP7_75t_L g4414 ( 
.A(n_3067),
.B(n_3091),
.Y(n_4414)
);

OAI21xp5_ASAP7_75t_L g4415 ( 
.A1(n_3717),
.A2(n_3791),
.B(n_3782),
.Y(n_4415)
);

HB1xp67_ASAP7_75t_L g4416 ( 
.A(n_3091),
.Y(n_4416)
);

INVx2_ASAP7_75t_L g4417 ( 
.A(n_3779),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_3779),
.B(n_3837),
.Y(n_4418)
);

AOI22x1_ASAP7_75t_L g4419 ( 
.A1(n_3130),
.A2(n_3129),
.B1(n_3124),
.B2(n_3151),
.Y(n_4419)
);

NOR2xp33_ASAP7_75t_L g4420 ( 
.A(n_3917),
.B(n_3949),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_3704),
.Y(n_4421)
);

NAND2xp5_ASAP7_75t_L g4422 ( 
.A(n_4213),
.B(n_4307),
.Y(n_4422)
);

AND2x4_ASAP7_75t_SL g4423 ( 
.A(n_3055),
.B(n_3082),
.Y(n_4423)
);

INVx2_ASAP7_75t_L g4424 ( 
.A(n_3779),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_3837),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_4213),
.B(n_4307),
.Y(n_4426)
);

AND2x2_ASAP7_75t_L g4427 ( 
.A(n_3837),
.B(n_3858),
.Y(n_4427)
);

OAI22xp5_ASAP7_75t_L g4428 ( 
.A1(n_3752),
.A2(n_3767),
.B1(n_3805),
.B2(n_3761),
.Y(n_4428)
);

INVx1_ASAP7_75t_L g4429 ( 
.A(n_3705),
.Y(n_4429)
);

INVx2_ASAP7_75t_L g4430 ( 
.A(n_3858),
.Y(n_4430)
);

AND3x1_ASAP7_75t_SL g4431 ( 
.A(n_3337),
.B(n_3660),
.C(n_3338),
.Y(n_4431)
);

AND2x4_ASAP7_75t_L g4432 ( 
.A(n_3099),
.B(n_3133),
.Y(n_4432)
);

INVx2_ASAP7_75t_SL g4433 ( 
.A(n_3099),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4356),
.Y(n_4434)
);

INVx1_ASAP7_75t_L g4435 ( 
.A(n_4356),
.Y(n_4435)
);

NOR2xp33_ASAP7_75t_L g4436 ( 
.A(n_3917),
.B(n_3949),
.Y(n_4436)
);

INVx8_ASAP7_75t_L g4437 ( 
.A(n_3505),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_SL g4438 ( 
.A(n_3125),
.B(n_3896),
.Y(n_4438)
);

BUFx12f_ASAP7_75t_L g4439 ( 
.A(n_3270),
.Y(n_4439)
);

BUFx3_ASAP7_75t_L g4440 ( 
.A(n_3284),
.Y(n_4440)
);

INVx2_ASAP7_75t_SL g4441 ( 
.A(n_3133),
.Y(n_4441)
);

BUFx6f_ASAP7_75t_L g4442 ( 
.A(n_3284),
.Y(n_4442)
);

CKINVDCx5p33_ASAP7_75t_R g4443 ( 
.A(n_3683),
.Y(n_4443)
);

BUFx4f_ASAP7_75t_L g4444 ( 
.A(n_3505),
.Y(n_4444)
);

INVx4_ASAP7_75t_L g4445 ( 
.A(n_3505),
.Y(n_4445)
);

AND3x1_ASAP7_75t_SL g4446 ( 
.A(n_3337),
.B(n_3660),
.C(n_3896),
.Y(n_4446)
);

INVx5_ASAP7_75t_L g4447 ( 
.A(n_3505),
.Y(n_4447)
);

AOI22xp33_ASAP7_75t_L g4448 ( 
.A1(n_3237),
.A2(n_3110),
.B1(n_3230),
.B2(n_3112),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_SL g4449 ( 
.A(n_3813),
.B(n_4164),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_SL g4450 ( 
.A(n_3813),
.B(n_4164),
.Y(n_4450)
);

NOR2xp33_ASAP7_75t_L g4451 ( 
.A(n_3956),
.B(n_4075),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4324),
.B(n_4338),
.Y(n_4452)
);

NAND2xp5_ASAP7_75t_L g4453 ( 
.A(n_4324),
.B(n_4338),
.Y(n_4453)
);

NAND2xp5_ASAP7_75t_L g4454 ( 
.A(n_3108),
.B(n_3109),
.Y(n_4454)
);

NOR4xp25_ASAP7_75t_SL g4455 ( 
.A(n_3068),
.B(n_3695),
.C(n_3712),
.D(n_3711),
.Y(n_4455)
);

O2A1O1Ixp33_ASAP7_75t_L g4456 ( 
.A1(n_3933),
.A2(n_3973),
.B(n_4117),
.C(n_4005),
.Y(n_4456)
);

BUFx6f_ASAP7_75t_SL g4457 ( 
.A(n_3621),
.Y(n_4457)
);

BUFx6f_ASAP7_75t_L g4458 ( 
.A(n_3766),
.Y(n_4458)
);

OR2x4_ASAP7_75t_L g4459 ( 
.A(n_3142),
.B(n_3055),
.Y(n_4459)
);

AO22x1_ASAP7_75t_L g4460 ( 
.A1(n_3069),
.A2(n_3202),
.B1(n_3224),
.B2(n_3174),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_3108),
.B(n_3109),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_3111),
.B(n_3113),
.Y(n_4462)
);

BUFx6f_ASAP7_75t_L g4463 ( 
.A(n_3766),
.Y(n_4463)
);

A2O1A1Ixp33_ASAP7_75t_L g4464 ( 
.A1(n_3054),
.A2(n_3237),
.B(n_3115),
.C(n_4191),
.Y(n_4464)
);

BUFx3_ASAP7_75t_L g4465 ( 
.A(n_3505),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_SL g4466 ( 
.A(n_3897),
.B(n_4207),
.Y(n_4466)
);

BUFx6f_ASAP7_75t_L g4467 ( 
.A(n_3247),
.Y(n_4467)
);

BUFx12f_ASAP7_75t_L g4468 ( 
.A(n_3557),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_L g4469 ( 
.A(n_3111),
.B(n_3113),
.Y(n_4469)
);

NOR2xp33_ASAP7_75t_L g4470 ( 
.A(n_3956),
.B(n_4075),
.Y(n_4470)
);

BUFx6f_ASAP7_75t_L g4471 ( 
.A(n_3192),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_3118),
.B(n_3136),
.Y(n_4472)
);

OR2x2_ASAP7_75t_L g4473 ( 
.A(n_4304),
.B(n_3287),
.Y(n_4473)
);

NAND2xp5_ASAP7_75t_L g4474 ( 
.A(n_3118),
.B(n_3136),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_3145),
.B(n_3096),
.Y(n_4475)
);

NOR2xp33_ASAP7_75t_L g4476 ( 
.A(n_4084),
.B(n_4087),
.Y(n_4476)
);

BUFx12f_ASAP7_75t_L g4477 ( 
.A(n_3100),
.Y(n_4477)
);

NOR2xp33_ASAP7_75t_L g4478 ( 
.A(n_4084),
.B(n_4087),
.Y(n_4478)
);

AOI22x1_ASAP7_75t_L g4479 ( 
.A1(n_3124),
.A2(n_3094),
.B1(n_4133),
.B2(n_3839),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_3886),
.B(n_3914),
.Y(n_4480)
);

BUFx4f_ASAP7_75t_SL g4481 ( 
.A(n_3503),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_3145),
.B(n_3096),
.Y(n_4482)
);

AOI21xp5_ASAP7_75t_L g4483 ( 
.A1(n_3690),
.A2(n_3707),
.B(n_3701),
.Y(n_4483)
);

BUFx6f_ASAP7_75t_L g4484 ( 
.A(n_3192),
.Y(n_4484)
);

INVx2_ASAP7_75t_SL g4485 ( 
.A(n_3185),
.Y(n_4485)
);

CKINVDCx6p67_ASAP7_75t_R g4486 ( 
.A(n_3585),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_3056),
.B(n_3057),
.Y(n_4487)
);

HB1xp67_ASAP7_75t_L g4488 ( 
.A(n_3215),
.Y(n_4488)
);

BUFx6f_ASAP7_75t_L g4489 ( 
.A(n_3192),
.Y(n_4489)
);

INVx4_ASAP7_75t_L g4490 ( 
.A(n_3505),
.Y(n_4490)
);

NAND2xp5_ASAP7_75t_SL g4491 ( 
.A(n_3315),
.B(n_3960),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_3056),
.B(n_3057),
.Y(n_4492)
);

BUFx3_ASAP7_75t_L g4493 ( 
.A(n_3052),
.Y(n_4493)
);

BUFx2_ASAP7_75t_L g4494 ( 
.A(n_3215),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_3693),
.B(n_3694),
.Y(n_4495)
);

AND2x4_ASAP7_75t_L g4496 ( 
.A(n_3225),
.B(n_3235),
.Y(n_4496)
);

INVx3_ASAP7_75t_SL g4497 ( 
.A(n_3540),
.Y(n_4497)
);

OAI21xp5_ASAP7_75t_L g4498 ( 
.A1(n_4193),
.A2(n_4215),
.B(n_4208),
.Y(n_4498)
);

BUFx2_ASAP7_75t_L g4499 ( 
.A(n_3076),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_3693),
.B(n_3694),
.Y(n_4500)
);

BUFx3_ASAP7_75t_L g4501 ( 
.A(n_3052),
.Y(n_4501)
);

NOR2xp33_ASAP7_75t_SL g4502 ( 
.A(n_3567),
.B(n_3733),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_SL g4503 ( 
.A(n_3315),
.B(n_3960),
.Y(n_4503)
);

OR2x6_ASAP7_75t_L g4504 ( 
.A(n_3060),
.B(n_3066),
.Y(n_4504)
);

INVx2_ASAP7_75t_SL g4505 ( 
.A(n_3103),
.Y(n_4505)
);

BUFx6f_ASAP7_75t_L g4506 ( 
.A(n_3192),
.Y(n_4506)
);

HB1xp67_ASAP7_75t_L g4507 ( 
.A(n_3214),
.Y(n_4507)
);

OR2x2_ASAP7_75t_L g4508 ( 
.A(n_4304),
.B(n_3287),
.Y(n_4508)
);

NAND2xp5_ASAP7_75t_SL g4509 ( 
.A(n_3960),
.B(n_3979),
.Y(n_4509)
);

AND2x4_ASAP7_75t_L g4510 ( 
.A(n_3225),
.B(n_3235),
.Y(n_4510)
);

NOR2xp33_ASAP7_75t_L g4511 ( 
.A(n_4113),
.B(n_4125),
.Y(n_4511)
);

AND2x6_ASAP7_75t_L g4512 ( 
.A(n_3055),
.B(n_3082),
.Y(n_4512)
);

CKINVDCx11_ASAP7_75t_R g4513 ( 
.A(n_3503),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_SL g4514 ( 
.A(n_3979),
.B(n_3304),
.Y(n_4514)
);

INVxp67_ASAP7_75t_L g4515 ( 
.A(n_3379),
.Y(n_4515)
);

OAI221xp5_ASAP7_75t_L g4516 ( 
.A1(n_3107),
.A2(n_4264),
.B1(n_4025),
.B2(n_3854),
.C(n_4001),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_3696),
.B(n_3703),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_SL g4518 ( 
.A(n_3979),
.B(n_3304),
.Y(n_4518)
);

INVx4_ASAP7_75t_L g4519 ( 
.A(n_3247),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_3696),
.B(n_3703),
.Y(n_4520)
);

NAND2xp5_ASAP7_75t_L g4521 ( 
.A(n_3714),
.B(n_3724),
.Y(n_4521)
);

AND2x4_ASAP7_75t_L g4522 ( 
.A(n_3258),
.B(n_3267),
.Y(n_4522)
);

NAND2xp5_ASAP7_75t_L g4523 ( 
.A(n_3714),
.B(n_3724),
.Y(n_4523)
);

NAND2xp5_ASAP7_75t_L g4524 ( 
.A(n_3728),
.B(n_3732),
.Y(n_4524)
);

NOR2xp33_ASAP7_75t_L g4525 ( 
.A(n_4113),
.B(n_4125),
.Y(n_4525)
);

A2O1A1Ixp33_ASAP7_75t_L g4526 ( 
.A1(n_4224),
.A2(n_3789),
.B(n_3817),
.C(n_3770),
.Y(n_4526)
);

BUFx6f_ASAP7_75t_L g4527 ( 
.A(n_3247),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4020),
.B(n_4038),
.Y(n_4528)
);

BUFx8_ASAP7_75t_L g4529 ( 
.A(n_3055),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_3728),
.B(n_3732),
.Y(n_4530)
);

A2O1A1Ixp33_ASAP7_75t_L g4531 ( 
.A1(n_3947),
.A2(n_3981),
.B(n_4246),
.C(n_3957),
.Y(n_4531)
);

NOR2xp67_ASAP7_75t_L g4532 ( 
.A(n_3142),
.B(n_3135),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_3734),
.B(n_3737),
.Y(n_4533)
);

NAND2xp5_ASAP7_75t_SL g4534 ( 
.A(n_3174),
.B(n_3202),
.Y(n_4534)
);

NOR2xp33_ASAP7_75t_L g4535 ( 
.A(n_4168),
.B(n_4184),
.Y(n_4535)
);

INVx2_ASAP7_75t_L g4536 ( 
.A(n_4020),
.Y(n_4536)
);

NAND2xp5_ASAP7_75t_L g4537 ( 
.A(n_3734),
.B(n_3737),
.Y(n_4537)
);

AO221x1_ASAP7_75t_L g4538 ( 
.A1(n_3224),
.A2(n_3226),
.B1(n_4184),
.B2(n_4194),
.C(n_4168),
.Y(n_4538)
);

NAND2xp5_ASAP7_75t_L g4539 ( 
.A(n_3740),
.B(n_3743),
.Y(n_4539)
);

AOI221xp5_ASAP7_75t_L g4540 ( 
.A1(n_3226),
.A2(n_4312),
.B1(n_4317),
.B2(n_4202),
.C(n_4194),
.Y(n_4540)
);

NAND3xp33_ASAP7_75t_SL g4541 ( 
.A(n_3257),
.B(n_3273),
.C(n_3767),
.Y(n_4541)
);

INVx5_ASAP7_75t_L g4542 ( 
.A(n_3055),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_SL g4543 ( 
.A(n_4099),
.B(n_4202),
.Y(n_4543)
);

INVx2_ASAP7_75t_L g4544 ( 
.A(n_4038),
.Y(n_4544)
);

OAI22xp5_ASAP7_75t_L g4545 ( 
.A1(n_3752),
.A2(n_3805),
.B1(n_3822),
.B2(n_3761),
.Y(n_4545)
);

BUFx6f_ASAP7_75t_L g4546 ( 
.A(n_3247),
.Y(n_4546)
);

NAND2xp5_ASAP7_75t_L g4547 ( 
.A(n_3740),
.B(n_3743),
.Y(n_4547)
);

BUFx6f_ASAP7_75t_L g4548 ( 
.A(n_3720),
.Y(n_4548)
);

AND2x4_ASAP7_75t_L g4549 ( 
.A(n_3258),
.B(n_3267),
.Y(n_4549)
);

NAND2xp5_ASAP7_75t_L g4550 ( 
.A(n_3747),
.B(n_3748),
.Y(n_4550)
);

AND2x4_ASAP7_75t_L g4551 ( 
.A(n_4363),
.B(n_3802),
.Y(n_4551)
);

BUFx6f_ASAP7_75t_L g4552 ( 
.A(n_3720),
.Y(n_4552)
);

NAND2xp5_ASAP7_75t_L g4553 ( 
.A(n_3747),
.B(n_3748),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_3756),
.B(n_3757),
.Y(n_4554)
);

AOI22xp5_ASAP7_75t_L g4555 ( 
.A1(n_4312),
.A2(n_4317),
.B1(n_4349),
.B2(n_3302),
.Y(n_4555)
);

NAND2xp5_ASAP7_75t_L g4556 ( 
.A(n_3756),
.B(n_3757),
.Y(n_4556)
);

INVx2_ASAP7_75t_L g4557 ( 
.A(n_4111),
.Y(n_4557)
);

AOI221x1_ASAP7_75t_L g4558 ( 
.A1(n_3230),
.A2(n_4205),
.B1(n_4217),
.B2(n_3986),
.C(n_3706),
.Y(n_4558)
);

OAI221xp5_ASAP7_75t_L g4559 ( 
.A1(n_4025),
.A2(n_4264),
.B1(n_4355),
.B2(n_4357),
.C(n_3845),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_3762),
.B(n_3765),
.Y(n_4560)
);

HB1xp67_ASAP7_75t_L g4561 ( 
.A(n_3134),
.Y(n_4561)
);

NAND2xp5_ASAP7_75t_L g4562 ( 
.A(n_3762),
.B(n_3765),
.Y(n_4562)
);

NOR2xp33_ASAP7_75t_L g4563 ( 
.A(n_4349),
.B(n_3302),
.Y(n_4563)
);

NAND2xp5_ASAP7_75t_L g4564 ( 
.A(n_3769),
.B(n_3774),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_3769),
.B(n_3774),
.Y(n_4565)
);

INVx2_ASAP7_75t_L g4566 ( 
.A(n_4111),
.Y(n_4566)
);

NAND2xp5_ASAP7_75t_L g4567 ( 
.A(n_3776),
.B(n_3777),
.Y(n_4567)
);

HB1xp67_ASAP7_75t_L g4568 ( 
.A(n_3134),
.Y(n_4568)
);

NAND2xp5_ASAP7_75t_L g4569 ( 
.A(n_3776),
.B(n_3777),
.Y(n_4569)
);

BUFx2_ASAP7_75t_L g4570 ( 
.A(n_3123),
.Y(n_4570)
);

HB1xp67_ASAP7_75t_L g4571 ( 
.A(n_3144),
.Y(n_4571)
);

OR2x2_ASAP7_75t_L g4572 ( 
.A(n_3059),
.B(n_3285),
.Y(n_4572)
);

NAND2xp5_ASAP7_75t_SL g4573 ( 
.A(n_3197),
.B(n_3290),
.Y(n_4573)
);

INVx2_ASAP7_75t_SL g4574 ( 
.A(n_3144),
.Y(n_4574)
);

INVx2_ASAP7_75t_L g4575 ( 
.A(n_4132),
.Y(n_4575)
);

INVxp67_ASAP7_75t_SL g4576 ( 
.A(n_3217),
.Y(n_4576)
);

INVx4_ASAP7_75t_L g4577 ( 
.A(n_3055),
.Y(n_4577)
);

AND2x4_ASAP7_75t_L g4578 ( 
.A(n_4363),
.B(n_3891),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_3780),
.B(n_3781),
.Y(n_4579)
);

NAND2xp5_ASAP7_75t_L g4580 ( 
.A(n_3780),
.B(n_3781),
.Y(n_4580)
);

INVx2_ASAP7_75t_L g4581 ( 
.A(n_4132),
.Y(n_4581)
);

OAI22xp5_ASAP7_75t_L g4582 ( 
.A1(n_3822),
.A2(n_3834),
.B1(n_3890),
.B2(n_3826),
.Y(n_4582)
);

BUFx4f_ASAP7_75t_L g4583 ( 
.A(n_3082),
.Y(n_4583)
);

AOI22xp33_ASAP7_75t_L g4584 ( 
.A1(n_3086),
.A2(n_3137),
.B1(n_3146),
.B2(n_3141),
.Y(n_4584)
);

HB1xp67_ASAP7_75t_L g4585 ( 
.A(n_3211),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_3784),
.B(n_3786),
.Y(n_4586)
);

OAI22xp5_ASAP7_75t_SL g4587 ( 
.A1(n_3155),
.A2(n_3264),
.B1(n_3165),
.B2(n_3181),
.Y(n_4587)
);

INVx5_ASAP7_75t_L g4588 ( 
.A(n_3082),
.Y(n_4588)
);

BUFx2_ASAP7_75t_L g4589 ( 
.A(n_3211),
.Y(n_4589)
);

INVx1_ASAP7_75t_SL g4590 ( 
.A(n_3379),
.Y(n_4590)
);

INVx5_ASAP7_75t_L g4591 ( 
.A(n_3082),
.Y(n_4591)
);

AND2x2_ASAP7_75t_L g4592 ( 
.A(n_4132),
.B(n_4134),
.Y(n_4592)
);

NAND2xp5_ASAP7_75t_L g4593 ( 
.A(n_3784),
.B(n_3786),
.Y(n_4593)
);

INVx1_ASAP7_75t_SL g4594 ( 
.A(n_3132),
.Y(n_4594)
);

INVx2_ASAP7_75t_L g4595 ( 
.A(n_4134),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_3788),
.B(n_3794),
.Y(n_4596)
);

BUFx2_ASAP7_75t_L g4597 ( 
.A(n_3214),
.Y(n_4597)
);

BUFx5_ASAP7_75t_L g4598 ( 
.A(n_3296),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_3788),
.B(n_3794),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_3795),
.B(n_3800),
.Y(n_4600)
);

BUFx6f_ASAP7_75t_L g4601 ( 
.A(n_3768),
.Y(n_4601)
);

AND2x4_ASAP7_75t_L g4602 ( 
.A(n_3891),
.B(n_3953),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_3795),
.B(n_3800),
.Y(n_4603)
);

CKINVDCx5p33_ASAP7_75t_R g4604 ( 
.A(n_3683),
.Y(n_4604)
);

AND2x4_ASAP7_75t_L g4605 ( 
.A(n_4363),
.B(n_3891),
.Y(n_4605)
);

BUFx4f_ASAP7_75t_L g4606 ( 
.A(n_3082),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_3804),
.B(n_3818),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_3804),
.B(n_3818),
.Y(n_4608)
);

BUFx6f_ASAP7_75t_L g4609 ( 
.A(n_3768),
.Y(n_4609)
);

HB1xp67_ASAP7_75t_L g4610 ( 
.A(n_3132),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_3819),
.B(n_3823),
.Y(n_4611)
);

OAI21xp5_ASAP7_75t_L g4612 ( 
.A1(n_3161),
.A2(n_3160),
.B(n_3759),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_3819),
.B(n_3823),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_4134),
.Y(n_4614)
);

NAND2x1_ASAP7_75t_L g4615 ( 
.A(n_3231),
.B(n_4029),
.Y(n_4615)
);

CKINVDCx14_ASAP7_75t_R g4616 ( 
.A(n_4078),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4135),
.Y(n_4617)
);

INVx5_ASAP7_75t_L g4618 ( 
.A(n_3719),
.Y(n_4618)
);

NAND2xp5_ASAP7_75t_L g4619 ( 
.A(n_3827),
.B(n_3828),
.Y(n_4619)
);

NOR2xp33_ASAP7_75t_L g4620 ( 
.A(n_3075),
.B(n_3382),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_3827),
.B(n_3828),
.Y(n_4621)
);

BUFx10_ASAP7_75t_L g4622 ( 
.A(n_3621),
.Y(n_4622)
);

CKINVDCx5p33_ASAP7_75t_R g4623 ( 
.A(n_3637),
.Y(n_4623)
);

BUFx6f_ASAP7_75t_L g4624 ( 
.A(n_3797),
.Y(n_4624)
);

NOR2xp33_ASAP7_75t_L g4625 ( 
.A(n_3171),
.B(n_3212),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_3830),
.B(n_3841),
.Y(n_4626)
);

NAND2xp5_ASAP7_75t_L g4627 ( 
.A(n_3830),
.B(n_3841),
.Y(n_4627)
);

AND2x2_ASAP7_75t_L g4628 ( 
.A(n_4159),
.B(n_4174),
.Y(n_4628)
);

BUFx6f_ASAP7_75t_L g4629 ( 
.A(n_3797),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_3843),
.B(n_3862),
.Y(n_4630)
);

BUFx2_ASAP7_75t_L g4631 ( 
.A(n_3306),
.Y(n_4631)
);

NOR2xp33_ASAP7_75t_L g4632 ( 
.A(n_3234),
.B(n_3261),
.Y(n_4632)
);

INVx3_ASAP7_75t_L g4633 ( 
.A(n_3306),
.Y(n_4633)
);

NOR2xp33_ASAP7_75t_R g4634 ( 
.A(n_4314),
.B(n_3733),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_3843),
.B(n_3862),
.Y(n_4635)
);

AOI22xp33_ASAP7_75t_L g4636 ( 
.A1(n_3262),
.A2(n_3281),
.B1(n_3293),
.B2(n_3288),
.Y(n_4636)
);

HB1xp67_ASAP7_75t_L g4637 ( 
.A(n_3301),
.Y(n_4637)
);

AOI22xp5_ASAP7_75t_L g4638 ( 
.A1(n_3309),
.A2(n_3889),
.B1(n_3834),
.B2(n_3826),
.Y(n_4638)
);

BUFx4f_ASAP7_75t_SL g4639 ( 
.A(n_3503),
.Y(n_4639)
);

INVx1_ASAP7_75t_SL g4640 ( 
.A(n_3301),
.Y(n_4640)
);

INVx2_ASAP7_75t_L g4641 ( 
.A(n_4159),
.Y(n_4641)
);

NAND2xp5_ASAP7_75t_L g4642 ( 
.A(n_3865),
.B(n_3868),
.Y(n_4642)
);

NAND2xp33_ASAP7_75t_SL g4643 ( 
.A(n_3839),
.B(n_4133),
.Y(n_4643)
);

INVxp67_ASAP7_75t_SL g4644 ( 
.A(n_3217),
.Y(n_4644)
);

AND2x2_ASAP7_75t_L g4645 ( 
.A(n_4159),
.B(n_4174),
.Y(n_4645)
);

NAND2xp5_ASAP7_75t_L g4646 ( 
.A(n_3865),
.B(n_3868),
.Y(n_4646)
);

INVx1_ASAP7_75t_SL g4647 ( 
.A(n_3847),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_3884),
.B(n_3887),
.Y(n_4648)
);

CKINVDCx5p33_ASAP7_75t_R g4649 ( 
.A(n_3948),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_3884),
.B(n_3887),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_3892),
.B(n_3898),
.Y(n_4651)
);

NAND2xp5_ASAP7_75t_L g4652 ( 
.A(n_3892),
.B(n_3898),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_3907),
.B(n_3920),
.Y(n_4653)
);

HB1xp67_ASAP7_75t_L g4654 ( 
.A(n_3847),
.Y(n_4654)
);

NAND2xp5_ASAP7_75t_L g4655 ( 
.A(n_3907),
.B(n_3920),
.Y(n_4655)
);

AND2x4_ASAP7_75t_L g4656 ( 
.A(n_3953),
.B(n_3955),
.Y(n_4656)
);

NAND2xp5_ASAP7_75t_SL g4657 ( 
.A(n_3290),
.B(n_3243),
.Y(n_4657)
);

HB1xp67_ASAP7_75t_SL g4658 ( 
.A(n_3078),
.Y(n_4658)
);

INVx2_ASAP7_75t_L g4659 ( 
.A(n_4174),
.Y(n_4659)
);

INVx3_ASAP7_75t_L g4660 ( 
.A(n_3306),
.Y(n_4660)
);

INVx3_ASAP7_75t_L g4661 ( 
.A(n_3310),
.Y(n_4661)
);

BUFx3_ASAP7_75t_L g4662 ( 
.A(n_3953),
.Y(n_4662)
);

INVx3_ASAP7_75t_L g4663 ( 
.A(n_3310),
.Y(n_4663)
);

INVxp67_ASAP7_75t_SL g4664 ( 
.A(n_3217),
.Y(n_4664)
);

NOR2xp33_ASAP7_75t_L g4665 ( 
.A(n_3073),
.B(n_3890),
.Y(n_4665)
);

A2O1A1Ixp33_ASAP7_75t_L g4666 ( 
.A1(n_4059),
.A2(n_4248),
.B(n_4251),
.C(n_4157),
.Y(n_4666)
);

BUFx2_ASAP7_75t_L g4667 ( 
.A(n_3310),
.Y(n_4667)
);

CKINVDCx14_ASAP7_75t_R g4668 ( 
.A(n_3350),
.Y(n_4668)
);

OR2x6_ASAP7_75t_L g4669 ( 
.A(n_3077),
.B(n_3093),
.Y(n_4669)
);

NOR2x1p5_ASAP7_75t_L g4670 ( 
.A(n_3083),
.B(n_3950),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_SL g4671 ( 
.A(n_3243),
.B(n_3190),
.Y(n_4671)
);

INVxp67_ASAP7_75t_L g4672 ( 
.A(n_3530),
.Y(n_4672)
);

NOR2xp33_ASAP7_75t_L g4673 ( 
.A(n_3901),
.B(n_3930),
.Y(n_4673)
);

INVx3_ASAP7_75t_L g4674 ( 
.A(n_3423),
.Y(n_4674)
);

AOI21xp5_ASAP7_75t_L g4675 ( 
.A1(n_3690),
.A2(n_3707),
.B(n_3701),
.Y(n_4675)
);

AOI221xp5_ASAP7_75t_L g4676 ( 
.A1(n_3312),
.A2(n_3286),
.B1(n_3259),
.B2(n_4211),
.C(n_3749),
.Y(n_4676)
);

NAND2xp5_ASAP7_75t_L g4677 ( 
.A(n_3921),
.B(n_3922),
.Y(n_4677)
);

INVx2_ASAP7_75t_SL g4678 ( 
.A(n_3955),
.Y(n_4678)
);

NAND2xp5_ASAP7_75t_L g4679 ( 
.A(n_3921),
.B(n_3922),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_L g4680 ( 
.A(n_3924),
.B(n_3925),
.Y(n_4680)
);

NAND2xp5_ASAP7_75t_L g4681 ( 
.A(n_3924),
.B(n_3925),
.Y(n_4681)
);

BUFx3_ASAP7_75t_L g4682 ( 
.A(n_3955),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_SL g4683 ( 
.A(n_3105),
.B(n_4270),
.Y(n_4683)
);

INVx3_ASAP7_75t_L g4684 ( 
.A(n_3423),
.Y(n_4684)
);

A2O1A1Ixp33_ASAP7_75t_L g4685 ( 
.A1(n_4365),
.A2(n_4340),
.B(n_4029),
.C(n_3090),
.Y(n_4685)
);

AND2x4_ASAP7_75t_L g4686 ( 
.A(n_4363),
.B(n_3969),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_3942),
.B(n_3945),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_L g4688 ( 
.A(n_3942),
.B(n_3945),
.Y(n_4688)
);

NAND2xp5_ASAP7_75t_SL g4689 ( 
.A(n_3297),
.B(n_3412),
.Y(n_4689)
);

INVxp67_ASAP7_75t_SL g4690 ( 
.A(n_3488),
.Y(n_4690)
);

AOI22xp33_ASAP7_75t_SL g4691 ( 
.A1(n_3208),
.A2(n_3312),
.B1(n_3692),
.B2(n_3058),
.Y(n_4691)
);

INVx3_ASAP7_75t_L g4692 ( 
.A(n_3311),
.Y(n_4692)
);

INVx2_ASAP7_75t_SL g4693 ( 
.A(n_3969),
.Y(n_4693)
);

BUFx6f_ASAP7_75t_L g4694 ( 
.A(n_3937),
.Y(n_4694)
);

CKINVDCx5p33_ASAP7_75t_R g4695 ( 
.A(n_3948),
.Y(n_4695)
);

NAND2x1p5_ASAP7_75t_L g4696 ( 
.A(n_3801),
.B(n_3231),
.Y(n_4696)
);

AOI22xp33_ASAP7_75t_L g4697 ( 
.A1(n_3729),
.A2(n_3731),
.B1(n_3755),
.B2(n_3736),
.Y(n_4697)
);

HB1xp67_ASAP7_75t_L g4698 ( 
.A(n_4120),
.Y(n_4698)
);

CKINVDCx5p33_ASAP7_75t_R g4699 ( 
.A(n_4268),
.Y(n_4699)
);

NAND3xp33_ASAP7_75t_L g4700 ( 
.A(n_3901),
.B(n_3954),
.C(n_3930),
.Y(n_4700)
);

AND3x1_ASAP7_75t_SL g4701 ( 
.A(n_3685),
.B(n_3744),
.C(n_3738),
.Y(n_4701)
);

CKINVDCx5p33_ASAP7_75t_R g4702 ( 
.A(n_4268),
.Y(n_4702)
);

AO22x1_ASAP7_75t_L g4703 ( 
.A1(n_3208),
.A2(n_3094),
.B1(n_3697),
.B2(n_3063),
.Y(n_4703)
);

INVx1_ASAP7_75t_SL g4704 ( 
.A(n_4120),
.Y(n_4704)
);

AO22x1_ASAP7_75t_L g4705 ( 
.A1(n_3063),
.A2(n_3699),
.B1(n_3702),
.B2(n_3697),
.Y(n_4705)
);

INVx4_ASAP7_75t_L g4706 ( 
.A(n_3719),
.Y(n_4706)
);

NOR2xp33_ASAP7_75t_L g4707 ( 
.A(n_3954),
.B(n_3967),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_3950),
.B(n_3958),
.Y(n_4708)
);

INVxp67_ASAP7_75t_SL g4709 ( 
.A(n_3488),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_3958),
.B(n_3965),
.Y(n_4710)
);

AND2x4_ASAP7_75t_L g4711 ( 
.A(n_3969),
.B(n_3977),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_L g4712 ( 
.A(n_3965),
.B(n_3966),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_3966),
.B(n_3970),
.Y(n_4713)
);

BUFx2_ASAP7_75t_L g4714 ( 
.A(n_4167),
.Y(n_4714)
);

NAND2xp5_ASAP7_75t_L g4715 ( 
.A(n_3970),
.B(n_3974),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_SL g4716 ( 
.A(n_3083),
.B(n_4012),
.Y(n_4716)
);

NOR2xp33_ASAP7_75t_R g4717 ( 
.A(n_3916),
.B(n_4212),
.Y(n_4717)
);

CKINVDCx14_ASAP7_75t_R g4718 ( 
.A(n_3464),
.Y(n_4718)
);

HB1xp67_ASAP7_75t_L g4719 ( 
.A(n_4210),
.Y(n_4719)
);

BUFx2_ASAP7_75t_L g4720 ( 
.A(n_4167),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_L g4721 ( 
.A(n_3974),
.B(n_3980),
.Y(n_4721)
);

BUFx3_ASAP7_75t_L g4722 ( 
.A(n_3969),
.Y(n_4722)
);

BUFx3_ASAP7_75t_L g4723 ( 
.A(n_3977),
.Y(n_4723)
);

AOI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_3708),
.A2(n_3715),
.B(n_3710),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_3980),
.B(n_3982),
.Y(n_4725)
);

CKINVDCx6p67_ASAP7_75t_R g4726 ( 
.A(n_3585),
.Y(n_4726)
);

AND3x1_ASAP7_75t_SL g4727 ( 
.A(n_3685),
.B(n_3829),
.C(n_3799),
.Y(n_4727)
);

HB1xp67_ASAP7_75t_L g4728 ( 
.A(n_4210),
.Y(n_4728)
);

INVx5_ASAP7_75t_L g4729 ( 
.A(n_3719),
.Y(n_4729)
);

NAND2xp5_ASAP7_75t_SL g4730 ( 
.A(n_4012),
.B(n_4068),
.Y(n_4730)
);

AND2x4_ASAP7_75t_L g4731 ( 
.A(n_3977),
.B(n_4144),
.Y(n_4731)
);

NAND2xp5_ASAP7_75t_L g4732 ( 
.A(n_3982),
.B(n_3983),
.Y(n_4732)
);

BUFx3_ASAP7_75t_L g4733 ( 
.A(n_3977),
.Y(n_4733)
);

AND2x6_ASAP7_75t_L g4734 ( 
.A(n_3719),
.B(n_3764),
.Y(n_4734)
);

HB1xp67_ASAP7_75t_L g4735 ( 
.A(n_4234),
.Y(n_4735)
);

NAND2xp5_ASAP7_75t_SL g4736 ( 
.A(n_4068),
.B(n_3706),
.Y(n_4736)
);

CKINVDCx20_ASAP7_75t_R g4737 ( 
.A(n_3508),
.Y(n_4737)
);

CKINVDCx20_ASAP7_75t_R g4738 ( 
.A(n_3078),
.Y(n_4738)
);

BUFx3_ASAP7_75t_L g4739 ( 
.A(n_4144),
.Y(n_4739)
);

NAND2xp5_ASAP7_75t_L g4740 ( 
.A(n_3983),
.B(n_3984),
.Y(n_4740)
);

BUFx4f_ASAP7_75t_L g4741 ( 
.A(n_3719),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_3984),
.B(n_3995),
.Y(n_4742)
);

INVx3_ASAP7_75t_L g4743 ( 
.A(n_3311),
.Y(n_4743)
);

NAND2xp5_ASAP7_75t_L g4744 ( 
.A(n_3995),
.B(n_3996),
.Y(n_4744)
);

AOI21xp5_ASAP7_75t_L g4745 ( 
.A1(n_3708),
.A2(n_3715),
.B(n_3710),
.Y(n_4745)
);

AND2x4_ASAP7_75t_L g4746 ( 
.A(n_4144),
.B(n_4219),
.Y(n_4746)
);

INVx3_ASAP7_75t_L g4747 ( 
.A(n_4056),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_3996),
.B(n_4011),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_4011),
.B(n_4014),
.Y(n_4749)
);

AOI22xp5_ASAP7_75t_L g4750 ( 
.A1(n_3967),
.A2(n_4089),
.B1(n_4104),
.B2(n_4006),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_4014),
.B(n_4026),
.Y(n_4751)
);

O2A1O1Ixp33_ASAP7_75t_L g4752 ( 
.A1(n_4368),
.A2(n_3855),
.B(n_3881),
.C(n_3851),
.Y(n_4752)
);

AOI22xp33_ASAP7_75t_L g4753 ( 
.A1(n_3773),
.A2(n_3814),
.B1(n_3836),
.B2(n_3812),
.Y(n_4753)
);

AOI22xp5_ASAP7_75t_L g4754 ( 
.A1(n_4006),
.A2(n_4104),
.B1(n_4179),
.B2(n_4089),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4026),
.B(n_4032),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4182),
.Y(n_4756)
);

OR2x6_ASAP7_75t_L g4757 ( 
.A(n_3077),
.B(n_3093),
.Y(n_4757)
);

AOI21xp5_ASAP7_75t_L g4758 ( 
.A1(n_3721),
.A2(n_3726),
.B(n_3725),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4182),
.Y(n_4759)
);

A2O1A1Ixp33_ASAP7_75t_L g4760 ( 
.A1(n_4364),
.A2(n_3702),
.B(n_3716),
.C(n_3699),
.Y(n_4760)
);

AND3x2_ASAP7_75t_SL g4761 ( 
.A(n_3231),
.B(n_3662),
.C(n_3070),
.Y(n_4761)
);

OR2x6_ASAP7_75t_L g4762 ( 
.A(n_3721),
.B(n_3725),
.Y(n_4762)
);

BUFx2_ASAP7_75t_L g4763 ( 
.A(n_4234),
.Y(n_4763)
);

NOR2xp33_ASAP7_75t_L g4764 ( 
.A(n_4179),
.B(n_4180),
.Y(n_4764)
);

INVxp67_ASAP7_75t_L g4765 ( 
.A(n_4284),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_L g4766 ( 
.A(n_4032),
.B(n_4036),
.Y(n_4766)
);

INVx5_ASAP7_75t_L g4767 ( 
.A(n_3719),
.Y(n_4767)
);

AND3x1_ASAP7_75t_SL g4768 ( 
.A(n_3993),
.B(n_4022),
.C(n_3994),
.Y(n_4768)
);

INVx6_ASAP7_75t_L g4769 ( 
.A(n_3764),
.Y(n_4769)
);

INVx2_ASAP7_75t_SL g4770 ( 
.A(n_4219),
.Y(n_4770)
);

NAND2xp5_ASAP7_75t_SL g4771 ( 
.A(n_3986),
.B(n_4205),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4036),
.B(n_4039),
.Y(n_4772)
);

INVx1_ASAP7_75t_SL g4773 ( 
.A(n_4284),
.Y(n_4773)
);

BUFx2_ASAP7_75t_L g4774 ( 
.A(n_4219),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4039),
.B(n_4052),
.Y(n_4775)
);

OAI221xp5_ASAP7_75t_L g4776 ( 
.A1(n_4180),
.A2(n_4260),
.B1(n_4278),
.B2(n_4218),
.C(n_4199),
.Y(n_4776)
);

INVx1_ASAP7_75t_SL g4777 ( 
.A(n_3615),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4197),
.Y(n_4778)
);

INVx1_ASAP7_75t_L g4779 ( 
.A(n_4197),
.Y(n_4779)
);

INVx1_ASAP7_75t_L g4780 ( 
.A(n_4214),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_4214),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_L g4782 ( 
.A(n_4052),
.B(n_4053),
.Y(n_4782)
);

NOR2xp33_ASAP7_75t_L g4783 ( 
.A(n_4199),
.B(n_4218),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4053),
.B(n_4055),
.Y(n_4784)
);

NOR2x1p5_ASAP7_75t_L g4785 ( 
.A(n_4061),
.B(n_4101),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_SL g4786 ( 
.A(n_4217),
.B(n_4301),
.Y(n_4786)
);

OR2x6_ASAP7_75t_L g4787 ( 
.A(n_3726),
.B(n_3730),
.Y(n_4787)
);

NOR2xp33_ASAP7_75t_R g4788 ( 
.A(n_3916),
.B(n_4212),
.Y(n_4788)
);

INVx1_ASAP7_75t_L g4789 ( 
.A(n_4235),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4235),
.Y(n_4790)
);

XOR2xp5_ASAP7_75t_L g4791 ( 
.A(n_3079),
.B(n_3104),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4303),
.Y(n_4792)
);

AND2x2_ASAP7_75t_L g4793 ( 
.A(n_3200),
.B(n_3203),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4303),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4055),
.B(n_4058),
.Y(n_4795)
);

AOI22xp33_ASAP7_75t_L g4796 ( 
.A1(n_3842),
.A2(n_3876),
.B1(n_3877),
.B2(n_3863),
.Y(n_4796)
);

AOI22xp5_ASAP7_75t_L g4797 ( 
.A1(n_4260),
.A2(n_4337),
.B1(n_4341),
.B2(n_4278),
.Y(n_4797)
);

NAND2xp5_ASAP7_75t_L g4798 ( 
.A(n_4058),
.B(n_4061),
.Y(n_4798)
);

BUFx3_ASAP7_75t_L g4799 ( 
.A(n_4274),
.Y(n_4799)
);

INVx2_ASAP7_75t_L g4800 ( 
.A(n_3524),
.Y(n_4800)
);

INVx2_ASAP7_75t_L g4801 ( 
.A(n_3524),
.Y(n_4801)
);

INVx2_ASAP7_75t_L g4802 ( 
.A(n_3296),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_SL g4803 ( 
.A(n_4301),
.B(n_3750),
.Y(n_4803)
);

NOR2xp67_ASAP7_75t_L g4804 ( 
.A(n_3328),
.B(n_3305),
.Y(n_4804)
);

AOI22xp5_ASAP7_75t_L g4805 ( 
.A1(n_4337),
.A2(n_4341),
.B1(n_3935),
.B2(n_3939),
.Y(n_4805)
);

NAND2xp5_ASAP7_75t_L g4806 ( 
.A(n_4064),
.B(n_4066),
.Y(n_4806)
);

INVx1_ASAP7_75t_L g4807 ( 
.A(n_3532),
.Y(n_4807)
);

AO21x2_ASAP7_75t_L g4808 ( 
.A1(n_4372),
.A2(n_3735),
.B(n_3730),
.Y(n_4808)
);

NAND2xp5_ASAP7_75t_L g4809 ( 
.A(n_4064),
.B(n_4066),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_3532),
.Y(n_4810)
);

INVx3_ASAP7_75t_L g4811 ( 
.A(n_4252),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4088),
.B(n_4093),
.Y(n_4812)
);

NAND2xp5_ASAP7_75t_SL g4813 ( 
.A(n_3852),
.B(n_3927),
.Y(n_4813)
);

AND2x4_ASAP7_75t_L g4814 ( 
.A(n_4274),
.B(n_4335),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_4088),
.B(n_4093),
.Y(n_4815)
);

AOI22xp5_ASAP7_75t_L g4816 ( 
.A1(n_3903),
.A2(n_3944),
.B1(n_3968),
.B2(n_3940),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_3200),
.B(n_3203),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_SL g4818 ( 
.A(n_4024),
.B(n_4151),
.Y(n_4818)
);

AND2x2_ASAP7_75t_L g4819 ( 
.A(n_3294),
.B(n_3232),
.Y(n_4819)
);

BUFx8_ASAP7_75t_L g4820 ( 
.A(n_3764),
.Y(n_4820)
);

AO22x1_ASAP7_75t_L g4821 ( 
.A1(n_3716),
.A2(n_3810),
.B1(n_3900),
.B2(n_3785),
.Y(n_4821)
);

OA22x2_ASAP7_75t_L g4822 ( 
.A1(n_4037),
.A2(n_4040),
.B1(n_4103),
.B2(n_4100),
.Y(n_4822)
);

INVx3_ASAP7_75t_L g4823 ( 
.A(n_4252),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_SL g4824 ( 
.A(n_4175),
.B(n_4190),
.Y(n_4824)
);

BUFx2_ASAP7_75t_L g4825 ( 
.A(n_4335),
.Y(n_4825)
);

INVx3_ASAP7_75t_L g4826 ( 
.A(n_4259),
.Y(n_4826)
);

AND3x1_ASAP7_75t_L g4827 ( 
.A(n_3567),
.B(n_3661),
.C(n_3673),
.Y(n_4827)
);

OAI21xp33_ASAP7_75t_L g4828 ( 
.A1(n_3971),
.A2(n_4048),
.B(n_4016),
.Y(n_4828)
);

AND2x4_ASAP7_75t_L g4829 ( 
.A(n_3114),
.B(n_3117),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_3294),
.B(n_3232),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4094),
.B(n_4096),
.Y(n_4831)
);

INVx3_ASAP7_75t_L g4832 ( 
.A(n_4259),
.Y(n_4832)
);

AND2x4_ASAP7_75t_SL g4833 ( 
.A(n_3764),
.B(n_3875),
.Y(n_4833)
);

INVx2_ASAP7_75t_SL g4834 ( 
.A(n_3195),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_4094),
.B(n_4096),
.Y(n_4835)
);

NOR2x1_ASAP7_75t_L g4836 ( 
.A(n_3059),
.B(n_3785),
.Y(n_4836)
);

INVx4_ASAP7_75t_L g4837 ( 
.A(n_3764),
.Y(n_4837)
);

INVx2_ASAP7_75t_SL g4838 ( 
.A(n_3195),
.Y(n_4838)
);

INVx1_ASAP7_75t_SL g4839 ( 
.A(n_3615),
.Y(n_4839)
);

OAI22xp5_ASAP7_75t_L g4840 ( 
.A1(n_3079),
.A2(n_3148),
.B1(n_3179),
.B2(n_3104),
.Y(n_4840)
);

AOI22xp33_ASAP7_75t_L g4841 ( 
.A1(n_4057),
.A2(n_4095),
.B1(n_4108),
.B2(n_4107),
.Y(n_4841)
);

AND2x4_ASAP7_75t_L g4842 ( 
.A(n_3114),
.B(n_3117),
.Y(n_4842)
);

BUFx3_ASAP7_75t_L g4843 ( 
.A(n_3764),
.Y(n_4843)
);

AOI22xp5_ASAP7_75t_L g4844 ( 
.A1(n_4050),
.A2(n_4148),
.B1(n_4166),
.B2(n_4158),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_4098),
.B(n_4101),
.Y(n_4845)
);

AO22x1_ASAP7_75t_L g4846 ( 
.A1(n_3810),
.A2(n_3900),
.B1(n_3919),
.B2(n_3915),
.Y(n_4846)
);

INVx1_ASAP7_75t_SL g4847 ( 
.A(n_3409),
.Y(n_4847)
);

BUFx8_ASAP7_75t_L g4848 ( 
.A(n_3875),
.Y(n_4848)
);

INVx5_ASAP7_75t_L g4849 ( 
.A(n_3875),
.Y(n_4849)
);

HB1xp67_ASAP7_75t_L g4850 ( 
.A(n_4269),
.Y(n_4850)
);

NAND2xp5_ASAP7_75t_L g4851 ( 
.A(n_4098),
.B(n_4106),
.Y(n_4851)
);

INVx5_ASAP7_75t_L g4852 ( 
.A(n_3875),
.Y(n_4852)
);

HB1xp67_ASAP7_75t_L g4853 ( 
.A(n_4269),
.Y(n_4853)
);

INVx3_ASAP7_75t_L g4854 ( 
.A(n_4275),
.Y(n_4854)
);

AND2x4_ASAP7_75t_L g4855 ( 
.A(n_3114),
.B(n_4275),
.Y(n_4855)
);

AOI22xp33_ASAP7_75t_L g4856 ( 
.A1(n_4201),
.A2(n_4221),
.B1(n_4227),
.B2(n_4209),
.Y(n_4856)
);

CKINVDCx5p33_ASAP7_75t_R g4857 ( 
.A(n_3398),
.Y(n_4857)
);

BUFx6f_ASAP7_75t_L g4858 ( 
.A(n_3875),
.Y(n_4858)
);

OR2x6_ASAP7_75t_L g4859 ( 
.A(n_3735),
.B(n_3742),
.Y(n_4859)
);

BUFx4f_ASAP7_75t_L g4860 ( 
.A(n_3875),
.Y(n_4860)
);

CKINVDCx8_ASAP7_75t_R g4861 ( 
.A(n_4276),
.Y(n_4861)
);

NAND2xp5_ASAP7_75t_L g4862 ( 
.A(n_4106),
.B(n_4115),
.Y(n_4862)
);

OR2x2_ASAP7_75t_L g4863 ( 
.A(n_3285),
.B(n_3292),
.Y(n_4863)
);

AND2x2_ASAP7_75t_L g4864 ( 
.A(n_3246),
.B(n_3253),
.Y(n_4864)
);

NOR2xp67_ASAP7_75t_L g4865 ( 
.A(n_3328),
.B(n_3305),
.Y(n_4865)
);

INVx5_ASAP7_75t_L g4866 ( 
.A(n_3895),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4115),
.B(n_4116),
.Y(n_4867)
);

AND2x4_ASAP7_75t_L g4868 ( 
.A(n_3114),
.B(n_3313),
.Y(n_4868)
);

INVx3_ASAP7_75t_L g4869 ( 
.A(n_3895),
.Y(n_4869)
);

OAI22xp5_ASAP7_75t_L g4870 ( 
.A1(n_3148),
.A2(n_3260),
.B1(n_3277),
.B2(n_3179),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4116),
.B(n_4121),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_SL g4872 ( 
.A(n_4220),
.B(n_3430),
.Y(n_4872)
);

NOR2xp67_ASAP7_75t_L g4873 ( 
.A(n_3120),
.B(n_3335),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4121),
.B(n_4129),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4129),
.B(n_4130),
.Y(n_4875)
);

NAND2xp5_ASAP7_75t_L g4876 ( 
.A(n_4130),
.B(n_4139),
.Y(n_4876)
);

AOI22xp5_ASAP7_75t_L g4877 ( 
.A1(n_4232),
.A2(n_4243),
.B1(n_4250),
.B2(n_4241),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_L g4878 ( 
.A(n_4139),
.B(n_4143),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4143),
.B(n_4156),
.Y(n_4879)
);

INVx3_ASAP7_75t_L g4880 ( 
.A(n_3895),
.Y(n_4880)
);

NAND2xp5_ASAP7_75t_L g4881 ( 
.A(n_4156),
.B(n_4163),
.Y(n_4881)
);

BUFx2_ASAP7_75t_L g4882 ( 
.A(n_3915),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4163),
.B(n_4173),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_L g4884 ( 
.A(n_4173),
.B(n_4176),
.Y(n_4884)
);

AOI211xp5_ASAP7_75t_L g4885 ( 
.A1(n_4124),
.A2(n_4185),
.B(n_4187),
.C(n_4152),
.Y(n_4885)
);

NAND2x1p5_ASAP7_75t_L g4886 ( 
.A(n_3801),
.B(n_3718),
.Y(n_4886)
);

HB1xp67_ASAP7_75t_L g4887 ( 
.A(n_3120),
.Y(n_4887)
);

AOI22xp5_ASAP7_75t_L g4888 ( 
.A1(n_4262),
.A2(n_4316),
.B1(n_4318),
.B2(n_4277),
.Y(n_4888)
);

NAND2xp5_ASAP7_75t_L g4889 ( 
.A(n_4176),
.B(n_4198),
.Y(n_4889)
);

NOR2xp33_ASAP7_75t_L g4890 ( 
.A(n_4280),
.B(n_4330),
.Y(n_4890)
);

A2O1A1Ixp33_ASAP7_75t_L g4891 ( 
.A1(n_4353),
.A2(n_4364),
.B(n_3932),
.C(n_3938),
.Y(n_4891)
);

BUFx6f_ASAP7_75t_L g4892 ( 
.A(n_3895),
.Y(n_4892)
);

AOI22xp5_ASAP7_75t_L g4893 ( 
.A1(n_4326),
.A2(n_4343),
.B1(n_4346),
.B2(n_4331),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4198),
.B(n_4200),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_3246),
.B(n_3253),
.Y(n_4895)
);

BUFx6f_ASAP7_75t_L g4896 ( 
.A(n_3895),
.Y(n_4896)
);

BUFx2_ASAP7_75t_L g4897 ( 
.A(n_3919),
.Y(n_4897)
);

AOI22xp5_ASAP7_75t_L g4898 ( 
.A1(n_4354),
.A2(n_4369),
.B1(n_4371),
.B2(n_4334),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4200),
.B(n_4206),
.Y(n_4899)
);

NAND2xp5_ASAP7_75t_SL g4900 ( 
.A(n_3486),
.B(n_3374),
.Y(n_4900)
);

BUFx3_ASAP7_75t_L g4901 ( 
.A(n_3895),
.Y(n_4901)
);

INVx3_ASAP7_75t_L g4902 ( 
.A(n_4351),
.Y(n_4902)
);

INVx2_ASAP7_75t_SL g4903 ( 
.A(n_3552),
.Y(n_4903)
);

HB1xp67_ASAP7_75t_L g4904 ( 
.A(n_3456),
.Y(n_4904)
);

BUFx4f_ASAP7_75t_SL g4905 ( 
.A(n_3629),
.Y(n_4905)
);

CKINVDCx5p33_ASAP7_75t_R g4906 ( 
.A(n_3398),
.Y(n_4906)
);

NAND2xp5_ASAP7_75t_SL g4907 ( 
.A(n_3374),
.B(n_3062),
.Y(n_4907)
);

BUFx6f_ASAP7_75t_L g4908 ( 
.A(n_3952),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4206),
.B(n_4229),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4229),
.B(n_4230),
.Y(n_4910)
);

BUFx3_ASAP7_75t_L g4911 ( 
.A(n_3952),
.Y(n_4911)
);

AOI22xp33_ASAP7_75t_L g4912 ( 
.A1(n_3153),
.A2(n_3164),
.B1(n_3170),
.B2(n_3159),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_SL g4913 ( 
.A(n_3062),
.B(n_3792),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_SL g4914 ( 
.A(n_3792),
.B(n_3807),
.Y(n_4914)
);

BUFx6f_ASAP7_75t_L g4915 ( 
.A(n_3952),
.Y(n_4915)
);

NOR2xp33_ASAP7_75t_L g4916 ( 
.A(n_3259),
.B(n_3286),
.Y(n_4916)
);

OR2x6_ASAP7_75t_L g4917 ( 
.A(n_3742),
.B(n_3745),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_3316),
.Y(n_4918)
);

BUFx6f_ASAP7_75t_L g4919 ( 
.A(n_3952),
.Y(n_4919)
);

BUFx8_ASAP7_75t_SL g4920 ( 
.A(n_3629),
.Y(n_4920)
);

XOR2xp5_ASAP7_75t_L g4921 ( 
.A(n_3260),
.B(n_3277),
.Y(n_4921)
);

NOR2xp33_ASAP7_75t_SL g4922 ( 
.A(n_3347),
.B(n_3183),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_3316),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4230),
.B(n_4249),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4249),
.B(n_4282),
.Y(n_4925)
);

AO221x1_ASAP7_75t_L g4926 ( 
.A1(n_3479),
.A2(n_4041),
.B1(n_4051),
.B2(n_4021),
.C(n_3952),
.Y(n_4926)
);

BUFx4f_ASAP7_75t_SL g4927 ( 
.A(n_3629),
.Y(n_4927)
);

AOI221xp5_ASAP7_75t_L g4928 ( 
.A1(n_3187),
.A2(n_3263),
.B1(n_3196),
.B2(n_3194),
.C(n_3322),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_3271),
.B(n_3272),
.Y(n_4929)
);

NAND2xp5_ASAP7_75t_L g4930 ( 
.A(n_4282),
.B(n_4285),
.Y(n_4930)
);

NAND2xp5_ASAP7_75t_L g4931 ( 
.A(n_4285),
.B(n_4286),
.Y(n_4931)
);

BUFx2_ASAP7_75t_L g4932 ( 
.A(n_3932),
.Y(n_4932)
);

INVx2_ASAP7_75t_L g4933 ( 
.A(n_3227),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4286),
.B(n_4287),
.Y(n_4934)
);

BUFx4f_ASAP7_75t_SL g4935 ( 
.A(n_4359),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4287),
.B(n_4296),
.Y(n_4936)
);

BUFx4f_ASAP7_75t_L g4937 ( 
.A(n_4021),
.Y(n_4937)
);

CKINVDCx5p33_ASAP7_75t_R g4938 ( 
.A(n_4359),
.Y(n_4938)
);

O2A1O1Ixp33_ASAP7_75t_L g4939 ( 
.A1(n_3393),
.A2(n_3358),
.B(n_3159),
.C(n_3164),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4296),
.B(n_4297),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_3227),
.Y(n_4941)
);

INVx2_ASAP7_75t_L g4942 ( 
.A(n_3266),
.Y(n_4942)
);

INVx1_ASAP7_75t_L g4943 ( 
.A(n_3346),
.Y(n_4943)
);

CKINVDCx5p33_ASAP7_75t_R g4944 ( 
.A(n_4359),
.Y(n_4944)
);

INVx2_ASAP7_75t_SL g4945 ( 
.A(n_3552),
.Y(n_4945)
);

CKINVDCx5p33_ASAP7_75t_R g4946 ( 
.A(n_3579),
.Y(n_4946)
);

OR2x6_ASAP7_75t_L g4947 ( 
.A(n_3745),
.B(n_3746),
.Y(n_4947)
);

BUFx2_ASAP7_75t_L g4948 ( 
.A(n_3938),
.Y(n_4948)
);

AOI22xp5_ASAP7_75t_L g4949 ( 
.A1(n_3084),
.A2(n_3098),
.B1(n_3122),
.B2(n_3088),
.Y(n_4949)
);

INVxp67_ASAP7_75t_SL g4950 ( 
.A(n_3723),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_SL g4951 ( 
.A(n_3807),
.B(n_3844),
.Y(n_4951)
);

INVx5_ASAP7_75t_L g4952 ( 
.A(n_4041),
.Y(n_4952)
);

CKINVDCx5p33_ASAP7_75t_R g4953 ( 
.A(n_3116),
.Y(n_4953)
);

BUFx2_ASAP7_75t_L g4954 ( 
.A(n_3959),
.Y(n_4954)
);

INVx2_ASAP7_75t_L g4955 ( 
.A(n_3266),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_3346),
.Y(n_4956)
);

CKINVDCx20_ASAP7_75t_R g4957 ( 
.A(n_3078),
.Y(n_4957)
);

HB1xp67_ASAP7_75t_L g4958 ( 
.A(n_3456),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4297),
.B(n_4306),
.Y(n_4959)
);

AND2x2_ASAP7_75t_L g4960 ( 
.A(n_3271),
.B(n_3272),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4306),
.B(n_4308),
.Y(n_4961)
);

BUFx2_ASAP7_75t_L g4962 ( 
.A(n_3959),
.Y(n_4962)
);

INVxp67_ASAP7_75t_L g4963 ( 
.A(n_3074),
.Y(n_4963)
);

BUFx2_ASAP7_75t_L g4964 ( 
.A(n_3963),
.Y(n_4964)
);

BUFx2_ASAP7_75t_L g4965 ( 
.A(n_3963),
.Y(n_4965)
);

AND2x4_ASAP7_75t_L g4966 ( 
.A(n_3313),
.B(n_3324),
.Y(n_4966)
);

AND2x2_ASAP7_75t_SL g4967 ( 
.A(n_3850),
.B(n_4074),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4308),
.B(n_4309),
.Y(n_4968)
);

INVx2_ASAP7_75t_L g4969 ( 
.A(n_3150),
.Y(n_4969)
);

INVx2_ASAP7_75t_L g4970 ( 
.A(n_3150),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_SL g4971 ( 
.A(n_3844),
.B(n_3861),
.Y(n_4971)
);

INVxp33_ASAP7_75t_L g4972 ( 
.A(n_3449),
.Y(n_4972)
);

NOR2xp33_ASAP7_75t_L g4973 ( 
.A(n_3377),
.B(n_3427),
.Y(n_4973)
);

AND3x1_ASAP7_75t_SL g4974 ( 
.A(n_3143),
.B(n_3201),
.C(n_3147),
.Y(n_4974)
);

NOR2xp67_ASAP7_75t_L g4975 ( 
.A(n_3335),
.B(n_3436),
.Y(n_4975)
);

AND2x2_ASAP7_75t_L g4976 ( 
.A(n_3295),
.B(n_3292),
.Y(n_4976)
);

AND2x4_ASAP7_75t_L g4977 ( 
.A(n_3324),
.B(n_3327),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4309),
.B(n_4310),
.Y(n_4978)
);

BUFx2_ASAP7_75t_L g4979 ( 
.A(n_3985),
.Y(n_4979)
);

NOR2xp33_ASAP7_75t_L g4980 ( 
.A(n_3377),
.B(n_3427),
.Y(n_4980)
);

INVxp67_ASAP7_75t_L g4981 ( 
.A(n_3186),
.Y(n_4981)
);

HB1xp67_ASAP7_75t_L g4982 ( 
.A(n_3299),
.Y(n_4982)
);

INVx4_ASAP7_75t_L g4983 ( 
.A(n_4041),
.Y(n_4983)
);

HB1xp67_ASAP7_75t_L g4984 ( 
.A(n_3351),
.Y(n_4984)
);

INVx2_ASAP7_75t_L g4985 ( 
.A(n_3370),
.Y(n_4985)
);

INVx4_ASAP7_75t_L g4986 ( 
.A(n_4051),
.Y(n_4986)
);

AOI21xp5_ASAP7_75t_L g4987 ( 
.A1(n_3746),
.A2(n_3758),
.B(n_3754),
.Y(n_4987)
);

BUFx4f_ASAP7_75t_SL g4988 ( 
.A(n_3493),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4310),
.B(n_4311),
.Y(n_4989)
);

INVx2_ASAP7_75t_L g4990 ( 
.A(n_3415),
.Y(n_4990)
);

NAND2xp5_ASAP7_75t_L g4991 ( 
.A(n_4311),
.B(n_4319),
.Y(n_4991)
);

INVx2_ASAP7_75t_L g4992 ( 
.A(n_3439),
.Y(n_4992)
);

BUFx4f_ASAP7_75t_SL g4993 ( 
.A(n_3493),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_4319),
.B(n_4332),
.Y(n_4994)
);

INVxp67_ASAP7_75t_SL g4995 ( 
.A(n_3723),
.Y(n_4995)
);

BUFx12f_ASAP7_75t_L g4996 ( 
.A(n_3434),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_3467),
.Y(n_4997)
);

AOI22x1_ASAP7_75t_L g4998 ( 
.A1(n_3985),
.A2(n_4062),
.B1(n_4063),
.B2(n_4009),
.Y(n_4998)
);

CKINVDCx20_ASAP7_75t_R g4999 ( 
.A(n_3078),
.Y(n_4999)
);

NOR2xp33_ASAP7_75t_L g5000 ( 
.A(n_3206),
.B(n_3219),
.Y(n_5000)
);

NAND2xp5_ASAP7_75t_L g5001 ( 
.A(n_4332),
.B(n_4345),
.Y(n_5001)
);

INVx2_ASAP7_75t_L g5002 ( 
.A(n_3535),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_3535),
.Y(n_5003)
);

AND3x2_ASAP7_75t_SL g5004 ( 
.A(n_3662),
.B(n_3909),
.C(n_3751),
.Y(n_5004)
);

AOI22xp5_ASAP7_75t_L g5005 ( 
.A1(n_3241),
.A2(n_3249),
.B1(n_3289),
.B2(n_3283),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_3545),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4345),
.B(n_4361),
.Y(n_5007)
);

AOI21x1_ASAP7_75t_L g5008 ( 
.A1(n_4372),
.A2(n_3758),
.B(n_3754),
.Y(n_5008)
);

AOI22xp5_ASAP7_75t_L g5009 ( 
.A1(n_3298),
.A2(n_3198),
.B1(n_3153),
.B2(n_3172),
.Y(n_5009)
);

NOR2xp33_ASAP7_75t_L g5010 ( 
.A(n_3331),
.B(n_3497),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_L g5011 ( 
.A(n_4361),
.B(n_4367),
.Y(n_5011)
);

NAND2xp5_ASAP7_75t_SL g5012 ( 
.A(n_3861),
.B(n_3872),
.Y(n_5012)
);

INVx1_ASAP7_75t_L g5013 ( 
.A(n_3550),
.Y(n_5013)
);

NOR2x1p5_ASAP7_75t_L g5014 ( 
.A(n_4367),
.B(n_4370),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4370),
.B(n_3138),
.Y(n_5015)
);

INVx2_ASAP7_75t_L g5016 ( 
.A(n_3550),
.Y(n_5016)
);

INVx2_ASAP7_75t_L g5017 ( 
.A(n_3576),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_3576),
.Y(n_5018)
);

CKINVDCx5p33_ASAP7_75t_R g5019 ( 
.A(n_3444),
.Y(n_5019)
);

AND3x1_ASAP7_75t_SL g5020 ( 
.A(n_3586),
.B(n_3209),
.C(n_3050),
.Y(n_5020)
);

INVx2_ASAP7_75t_L g5021 ( 
.A(n_3586),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_L g5022 ( 
.A(n_3138),
.B(n_3139),
.Y(n_5022)
);

NOR2xp33_ASAP7_75t_L g5023 ( 
.A(n_3497),
.B(n_3128),
.Y(n_5023)
);

INVx1_ASAP7_75t_L g5024 ( 
.A(n_3207),
.Y(n_5024)
);

NAND2xp5_ASAP7_75t_L g5025 ( 
.A(n_3139),
.B(n_3087),
.Y(n_5025)
);

INVx1_ASAP7_75t_L g5026 ( 
.A(n_3207),
.Y(n_5026)
);

BUFx2_ASAP7_75t_L g5027 ( 
.A(n_4009),
.Y(n_5027)
);

INVx5_ASAP7_75t_L g5028 ( 
.A(n_4071),
.Y(n_5028)
);

A2O1A1Ixp33_ASAP7_75t_L g5029 ( 
.A1(n_4333),
.A2(n_4353),
.B(n_4063),
.C(n_4097),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_3087),
.B(n_3126),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_3119),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_3119),
.Y(n_5032)
);

NAND2xp5_ASAP7_75t_L g5033 ( 
.A(n_3127),
.B(n_3064),
.Y(n_5033)
);

OR2x6_ASAP7_75t_L g5034 ( 
.A(n_4028),
.B(n_4030),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_3751),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_L g5036 ( 
.A(n_3064),
.B(n_3128),
.Y(n_5036)
);

CKINVDCx5p33_ASAP7_75t_R g5037 ( 
.A(n_3709),
.Y(n_5037)
);

INVx2_ASAP7_75t_L g5038 ( 
.A(n_3507),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_3152),
.B(n_3156),
.Y(n_5039)
);

A2O1A1Ixp33_ASAP7_75t_L g5040 ( 
.A1(n_4062),
.A2(n_4118),
.B(n_4192),
.C(n_4097),
.Y(n_5040)
);

HB1xp67_ASAP7_75t_L g5041 ( 
.A(n_3698),
.Y(n_5041)
);

INVx2_ASAP7_75t_L g5042 ( 
.A(n_3507),
.Y(n_5042)
);

NOR2xp33_ASAP7_75t_L g5043 ( 
.A(n_3322),
.B(n_3381),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_SL g5044 ( 
.A(n_3872),
.B(n_3882),
.Y(n_5044)
);

AOI22xp33_ASAP7_75t_L g5045 ( 
.A1(n_3170),
.A2(n_3172),
.B1(n_3175),
.B2(n_3173),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_3157),
.B(n_3158),
.Y(n_5046)
);

HB1xp67_ASAP7_75t_L g5047 ( 
.A(n_3739),
.Y(n_5047)
);

OR2x2_ASAP7_75t_L g5048 ( 
.A(n_3162),
.B(n_3163),
.Y(n_5048)
);

NAND2xp5_ASAP7_75t_SL g5049 ( 
.A(n_3882),
.B(n_3934),
.Y(n_5049)
);

BUFx12f_ASAP7_75t_L g5050 ( 
.A(n_3803),
.Y(n_5050)
);

INVx2_ASAP7_75t_L g5051 ( 
.A(n_3543),
.Y(n_5051)
);

AND2x4_ASAP7_75t_L g5052 ( 
.A(n_3327),
.B(n_3256),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_SL g5053 ( 
.A(n_3934),
.B(n_4044),
.Y(n_5053)
);

NOR3xp33_ASAP7_75t_L g5054 ( 
.A(n_3457),
.B(n_3832),
.C(n_3783),
.Y(n_5054)
);

BUFx8_ASAP7_75t_L g5055 ( 
.A(n_4071),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_SL g5056 ( 
.A(n_4044),
.B(n_4054),
.Y(n_5056)
);

INVx4_ASAP7_75t_L g5057 ( 
.A(n_4086),
.Y(n_5057)
);

NAND2xp5_ASAP7_75t_SL g5058 ( 
.A(n_4054),
.B(n_4069),
.Y(n_5058)
);

INVx1_ASAP7_75t_L g5059 ( 
.A(n_3909),
.Y(n_5059)
);

OAI22xp5_ASAP7_75t_L g5060 ( 
.A1(n_3323),
.A2(n_3341),
.B1(n_3391),
.B2(n_3380),
.Y(n_5060)
);

INVx1_ASAP7_75t_L g5061 ( 
.A(n_4244),
.Y(n_5061)
);

AOI22xp33_ASAP7_75t_L g5062 ( 
.A1(n_3173),
.A2(n_3175),
.B1(n_3184),
.B2(n_3177),
.Y(n_5062)
);

AOI22xp5_ASAP7_75t_L g5063 ( 
.A1(n_3222),
.A2(n_3223),
.B1(n_3177),
.B2(n_3189),
.Y(n_5063)
);

CKINVDCx6p67_ASAP7_75t_R g5064 ( 
.A(n_3493),
.Y(n_5064)
);

AND2x4_ASAP7_75t_L g5065 ( 
.A(n_3256),
.B(n_3265),
.Y(n_5065)
);

AND2x4_ASAP7_75t_L g5066 ( 
.A(n_3265),
.B(n_4118),
.Y(n_5066)
);

INVx2_ASAP7_75t_L g5067 ( 
.A(n_3874),
.Y(n_5067)
);

NAND2xp5_ASAP7_75t_L g5068 ( 
.A(n_3166),
.B(n_3167),
.Y(n_5068)
);

INVx1_ASAP7_75t_L g5069 ( 
.A(n_4244),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_3168),
.B(n_3169),
.Y(n_5070)
);

CKINVDCx5p33_ASAP7_75t_R g5071 ( 
.A(n_4138),
.Y(n_5071)
);

AND2x4_ASAP7_75t_L g5072 ( 
.A(n_4192),
.B(n_4231),
.Y(n_5072)
);

HB1xp67_ASAP7_75t_L g5073 ( 
.A(n_3753),
.Y(n_5073)
);

AND2x4_ASAP7_75t_L g5074 ( 
.A(n_4231),
.B(n_4255),
.Y(n_5074)
);

CKINVDCx6p67_ASAP7_75t_R g5075 ( 
.A(n_3154),
.Y(n_5075)
);

AND2x4_ASAP7_75t_L g5076 ( 
.A(n_4255),
.B(n_4273),
.Y(n_5076)
);

INVx1_ASAP7_75t_L g5077 ( 
.A(n_4247),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_SL g5078 ( 
.A(n_4069),
.B(n_4072),
.Y(n_5078)
);

AO22x1_ASAP7_75t_L g5079 ( 
.A1(n_4273),
.A2(n_4323),
.B1(n_4333),
.B2(n_4327),
.Y(n_5079)
);

AND2x4_ASAP7_75t_L g5080 ( 
.A(n_4323),
.B(n_4327),
.Y(n_5080)
);

BUFx12f_ASAP7_75t_L g5081 ( 
.A(n_4142),
.Y(n_5081)
);

BUFx4f_ASAP7_75t_L g5082 ( 
.A(n_4086),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_3176),
.B(n_3178),
.Y(n_5083)
);

AND2x2_ASAP7_75t_L g5084 ( 
.A(n_3295),
.B(n_3080),
.Y(n_5084)
);

INVx2_ASAP7_75t_L g5085 ( 
.A(n_4018),
.Y(n_5085)
);

NAND2xp33_ASAP7_75t_L g5086 ( 
.A(n_3184),
.B(n_3189),
.Y(n_5086)
);

NAND2xp5_ASAP7_75t_L g5087 ( 
.A(n_3180),
.B(n_3188),
.Y(n_5087)
);

INVx2_ASAP7_75t_L g5088 ( 
.A(n_4023),
.Y(n_5088)
);

INVx1_ASAP7_75t_SL g5089 ( 
.A(n_3409),
.Y(n_5089)
);

CKINVDCx20_ASAP7_75t_R g5090 ( 
.A(n_3221),
.Y(n_5090)
);

INVx1_ASAP7_75t_L g5091 ( 
.A(n_4247),
.Y(n_5091)
);

AO22x1_ASAP7_75t_L g5092 ( 
.A1(n_3879),
.A2(n_4073),
.B1(n_4085),
.B2(n_4072),
.Y(n_5092)
);

INVx1_ASAP7_75t_L g5093 ( 
.A(n_4299),
.Y(n_5093)
);

AND2x2_ASAP7_75t_L g5094 ( 
.A(n_3080),
.B(n_3210),
.Y(n_5094)
);

INVx2_ASAP7_75t_L g5095 ( 
.A(n_4171),
.Y(n_5095)
);

INVxp33_ASAP7_75t_SL g5096 ( 
.A(n_4263),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_SL g5097 ( 
.A(n_4073),
.B(n_4085),
.Y(n_5097)
);

AOI22xp33_ASAP7_75t_L g5098 ( 
.A1(n_3191),
.A2(n_3198),
.B1(n_3218),
.B2(n_3204),
.Y(n_5098)
);

AND2x2_ASAP7_75t_L g5099 ( 
.A(n_3213),
.B(n_3216),
.Y(n_5099)
);

AOI22xp33_ASAP7_75t_L g5100 ( 
.A1(n_3191),
.A2(n_3204),
.B1(n_3222),
.B2(n_3218),
.Y(n_5100)
);

BUFx12f_ASAP7_75t_L g5101 ( 
.A(n_3221),
.Y(n_5101)
);

CKINVDCx20_ASAP7_75t_R g5102 ( 
.A(n_3221),
.Y(n_5102)
);

AND2x2_ASAP7_75t_L g5103 ( 
.A(n_3220),
.B(n_3228),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_3229),
.B(n_3233),
.Y(n_5104)
);

AND3x1_ASAP7_75t_SL g5105 ( 
.A(n_3572),
.B(n_3609),
.C(n_3575),
.Y(n_5105)
);

HB1xp67_ASAP7_75t_L g5106 ( 
.A(n_3772),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_4299),
.Y(n_5107)
);

INVx2_ASAP7_75t_L g5108 ( 
.A(n_4225),
.Y(n_5108)
);

BUFx2_ASAP7_75t_L g5109 ( 
.A(n_3371),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_3236),
.B(n_3239),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_3589),
.Y(n_5111)
);

AND2x4_ASAP7_75t_L g5112 ( 
.A(n_3308),
.B(n_3314),
.Y(n_5112)
);

INVx2_ASAP7_75t_SL g5113 ( 
.A(n_3552),
.Y(n_5113)
);

BUFx8_ASAP7_75t_SL g5114 ( 
.A(n_3583),
.Y(n_5114)
);

AOI22xp5_ASAP7_75t_L g5115 ( 
.A1(n_3223),
.A2(n_3245),
.B1(n_3238),
.B2(n_3240),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_3589),
.Y(n_5116)
);

NAND2xp5_ASAP7_75t_SL g5117 ( 
.A(n_4136),
.B(n_4150),
.Y(n_5117)
);

HB1xp67_ASAP7_75t_L g5118 ( 
.A(n_3835),
.Y(n_5118)
);

INVxp67_ASAP7_75t_SL g5119 ( 
.A(n_4028),
.Y(n_5119)
);

HB1xp67_ASAP7_75t_L g5120 ( 
.A(n_3860),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_SL g5121 ( 
.A(n_4136),
.B(n_4150),
.Y(n_5121)
);

NOR3xp33_ASAP7_75t_L g5122 ( 
.A(n_3457),
.B(n_4271),
.C(n_3465),
.Y(n_5122)
);

AND2x4_ASAP7_75t_L g5123 ( 
.A(n_3308),
.B(n_3314),
.Y(n_5123)
);

AND2x4_ASAP7_75t_L g5124 ( 
.A(n_3317),
.B(n_3359),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_3242),
.B(n_3244),
.Y(n_5125)
);

NAND2x1_ASAP7_75t_L g5126 ( 
.A(n_3771),
.B(n_3775),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_L g5127 ( 
.A(n_3252),
.B(n_3255),
.Y(n_5127)
);

CKINVDCx5p33_ASAP7_75t_R g5128 ( 
.A(n_4360),
.Y(n_5128)
);

INVx1_ASAP7_75t_L g5129 ( 
.A(n_3317),
.Y(n_5129)
);

AOI22xp33_ASAP7_75t_L g5130 ( 
.A1(n_3238),
.A2(n_3240),
.B1(n_3250),
.B2(n_3245),
.Y(n_5130)
);

INVx1_ASAP7_75t_L g5131 ( 
.A(n_3498),
.Y(n_5131)
);

INVx1_ASAP7_75t_L g5132 ( 
.A(n_3498),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_3517),
.Y(n_5133)
);

NAND2x1p5_ASAP7_75t_L g5134 ( 
.A(n_3778),
.B(n_3787),
.Y(n_5134)
);

INVx1_ASAP7_75t_L g5135 ( 
.A(n_3517),
.Y(n_5135)
);

INVx4_ASAP7_75t_L g5136 ( 
.A(n_4154),
.Y(n_5136)
);

HB1xp67_ASAP7_75t_L g5137 ( 
.A(n_3908),
.Y(n_5137)
);

INVx2_ASAP7_75t_SL g5138 ( 
.A(n_3552),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_3268),
.B(n_3274),
.Y(n_5139)
);

INVx1_ASAP7_75t_L g5140 ( 
.A(n_3544),
.Y(n_5140)
);

AND2x2_ASAP7_75t_L g5141 ( 
.A(n_3278),
.B(n_3279),
.Y(n_5141)
);

AND2x6_ASAP7_75t_L g5142 ( 
.A(n_4154),
.B(n_4170),
.Y(n_5142)
);

AND2x2_ASAP7_75t_L g5143 ( 
.A(n_3280),
.B(n_4177),
.Y(n_5143)
);

NAND2xp5_ASAP7_75t_L g5144 ( 
.A(n_3397),
.B(n_3250),
.Y(n_5144)
);

NAND2xp5_ASAP7_75t_L g5145 ( 
.A(n_3397),
.B(n_4177),
.Y(n_5145)
);

A2O1A1Ixp33_ASAP7_75t_L g5146 ( 
.A1(n_3373),
.A2(n_3395),
.B(n_3399),
.C(n_3390),
.Y(n_5146)
);

AND2x4_ASAP7_75t_L g5147 ( 
.A(n_3359),
.B(n_3344),
.Y(n_5147)
);

AND2x2_ASAP7_75t_L g5148 ( 
.A(n_4222),
.B(n_4226),
.Y(n_5148)
);

NAND2xp5_ASAP7_75t_L g5149 ( 
.A(n_4222),
.B(n_4226),
.Y(n_5149)
);

NAND2xp5_ASAP7_75t_L g5150 ( 
.A(n_4256),
.B(n_4288),
.Y(n_5150)
);

NAND2x1p5_ASAP7_75t_L g5151 ( 
.A(n_3790),
.B(n_3793),
.Y(n_5151)
);

HB1xp67_ASAP7_75t_L g5152 ( 
.A(n_3961),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_3563),
.Y(n_5153)
);

AOI221xp5_ASAP7_75t_L g5154 ( 
.A1(n_3381),
.A2(n_3429),
.B1(n_3394),
.B2(n_3366),
.C(n_3376),
.Y(n_5154)
);

HB1xp67_ASAP7_75t_L g5155 ( 
.A(n_3989),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_4256),
.B(n_4288),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_SL g5157 ( 
.A(n_4293),
.B(n_3071),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_4293),
.B(n_3330),
.Y(n_5158)
);

INVx4_ASAP7_75t_L g5159 ( 
.A(n_4154),
.Y(n_5159)
);

AND2x2_ASAP7_75t_L g5160 ( 
.A(n_4170),
.B(n_4321),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_3330),
.B(n_3340),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_3340),
.B(n_3401),
.Y(n_5162)
);

AND2x2_ASAP7_75t_L g5163 ( 
.A(n_4170),
.B(n_4321),
.Y(n_5163)
);

INVx1_ASAP7_75t_SL g5164 ( 
.A(n_4010),
.Y(n_5164)
);

CKINVDCx5p33_ASAP7_75t_R g5165 ( 
.A(n_3199),
.Y(n_5165)
);

A2O1A1Ixp33_ASAP7_75t_L g5166 ( 
.A1(n_3402),
.A2(n_3407),
.B(n_3408),
.C(n_3403),
.Y(n_5166)
);

INVx1_ASAP7_75t_L g5167 ( 
.A(n_3458),
.Y(n_5167)
);

BUFx4f_ASAP7_75t_L g5168 ( 
.A(n_4170),
.Y(n_5168)
);

NOR2xp33_ASAP7_75t_L g5169 ( 
.A(n_3394),
.B(n_3429),
.Y(n_5169)
);

INVx4_ASAP7_75t_L g5170 ( 
.A(n_4321),
.Y(n_5170)
);

INVx1_ASAP7_75t_L g5171 ( 
.A(n_3458),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_3472),
.Y(n_5172)
);

NAND2xp5_ASAP7_75t_L g5173 ( 
.A(n_3413),
.B(n_3416),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_L g5174 ( 
.A(n_3418),
.B(n_3421),
.Y(n_5174)
);

CKINVDCx5p33_ASAP7_75t_R g5175 ( 
.A(n_3199),
.Y(n_5175)
);

INVx2_ASAP7_75t_L g5176 ( 
.A(n_3582),
.Y(n_5176)
);

NAND2xp5_ASAP7_75t_L g5177 ( 
.A(n_3425),
.B(n_3300),
.Y(n_5177)
);

NAND2xp5_ASAP7_75t_L g5178 ( 
.A(n_3300),
.B(n_3326),
.Y(n_5178)
);

BUFx2_ASAP7_75t_L g5179 ( 
.A(n_4321),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_SL g5180 ( 
.A(n_3071),
.B(n_3574),
.Y(n_5180)
);

INVx1_ASAP7_75t_SL g5181 ( 
.A(n_4031),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_3326),
.B(n_3329),
.Y(n_5182)
);

INVx1_ASAP7_75t_L g5183 ( 
.A(n_3472),
.Y(n_5183)
);

INVx1_ASAP7_75t_L g5184 ( 
.A(n_3476),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_3476),
.Y(n_5185)
);

INVx2_ASAP7_75t_SL g5186 ( 
.A(n_3552),
.Y(n_5186)
);

INVx1_ASAP7_75t_L g5187 ( 
.A(n_3477),
.Y(n_5187)
);

HB1xp67_ASAP7_75t_L g5188 ( 
.A(n_4079),
.Y(n_5188)
);

INVx1_ASAP7_75t_L g5189 ( 
.A(n_3477),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_3478),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_SL g5191 ( 
.A(n_3574),
.B(n_3466),
.Y(n_5191)
);

AOI22xp33_ASAP7_75t_L g5192 ( 
.A1(n_3387),
.A2(n_3089),
.B1(n_3320),
.B2(n_3318),
.Y(n_5192)
);

INVxp67_ASAP7_75t_L g5193 ( 
.A(n_4110),
.Y(n_5193)
);

NOR2xp33_ASAP7_75t_L g5194 ( 
.A(n_3689),
.B(n_3323),
.Y(n_5194)
);

NAND2xp5_ASAP7_75t_SL g5195 ( 
.A(n_3466),
.B(n_3591),
.Y(n_5195)
);

BUFx8_ASAP7_75t_SL g5196 ( 
.A(n_3583),
.Y(n_5196)
);

NAND2xp5_ASAP7_75t_L g5197 ( 
.A(n_3329),
.B(n_3339),
.Y(n_5197)
);

NAND2xp5_ASAP7_75t_SL g5198 ( 
.A(n_3591),
.B(n_3282),
.Y(n_5198)
);

INVx1_ASAP7_75t_L g5199 ( 
.A(n_3478),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_3339),
.B(n_3342),
.Y(n_5200)
);

AOI22xp5_ASAP7_75t_L g5201 ( 
.A1(n_3352),
.A2(n_3353),
.B1(n_3368),
.B2(n_3362),
.Y(n_5201)
);

INVx1_ASAP7_75t_L g5202 ( 
.A(n_3480),
.Y(n_5202)
);

INVx2_ASAP7_75t_SL g5203 ( 
.A(n_3552),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_3482),
.Y(n_5204)
);

NAND2xp5_ASAP7_75t_L g5205 ( 
.A(n_3342),
.B(n_3341),
.Y(n_5205)
);

NOR2xp33_ASAP7_75t_L g5206 ( 
.A(n_3689),
.B(n_3380),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_3482),
.Y(n_5207)
);

BUFx4f_ASAP7_75t_L g5208 ( 
.A(n_4352),
.Y(n_5208)
);

HB1xp67_ASAP7_75t_L g5209 ( 
.A(n_4169),
.Y(n_5209)
);

INVx1_ASAP7_75t_L g5210 ( 
.A(n_3483),
.Y(n_5210)
);

NOR2x1_ASAP7_75t_L g5211 ( 
.A(n_3491),
.B(n_3307),
.Y(n_5211)
);

AND2x4_ASAP7_75t_L g5212 ( 
.A(n_3359),
.B(n_3601),
.Y(n_5212)
);

NOR2xp33_ASAP7_75t_R g5213 ( 
.A(n_3081),
.B(n_3347),
.Y(n_5213)
);

INVx3_ASAP7_75t_L g5214 ( 
.A(n_3193),
.Y(n_5214)
);

XOR2xp5_ASAP7_75t_L g5215 ( 
.A(n_3504),
.B(n_3391),
.Y(n_5215)
);

NAND2xp5_ASAP7_75t_L g5216 ( 
.A(n_3332),
.B(n_3345),
.Y(n_5216)
);

INVx8_ASAP7_75t_L g5217 ( 
.A(n_3540),
.Y(n_5217)
);

NAND2xp5_ASAP7_75t_L g5218 ( 
.A(n_3348),
.B(n_3349),
.Y(n_5218)
);

OR2x2_ASAP7_75t_L g5219 ( 
.A(n_3282),
.B(n_3275),
.Y(n_5219)
);

AOI22xp5_ASAP7_75t_L g5220 ( 
.A1(n_3410),
.A2(n_3428),
.B1(n_3089),
.B2(n_3879),
.Y(n_5220)
);

INVx3_ASAP7_75t_L g5221 ( 
.A(n_3193),
.Y(n_5221)
);

CKINVDCx5p33_ASAP7_75t_R g5222 ( 
.A(n_3883),
.Y(n_5222)
);

NAND2xp5_ASAP7_75t_L g5223 ( 
.A(n_3348),
.B(n_3349),
.Y(n_5223)
);

OR2x6_ASAP7_75t_L g5224 ( 
.A(n_4030),
.B(n_4033),
.Y(n_5224)
);

INVx1_ASAP7_75t_SL g5225 ( 
.A(n_4283),
.Y(n_5225)
);

BUFx6f_ASAP7_75t_L g5226 ( 
.A(n_3850),
.Y(n_5226)
);

AOI22xp33_ASAP7_75t_L g5227 ( 
.A1(n_3461),
.A2(n_3879),
.B1(n_3392),
.B2(n_3417),
.Y(n_5227)
);

BUFx2_ASAP7_75t_L g5228 ( 
.A(n_3479),
.Y(n_5228)
);

CKINVDCx16_ASAP7_75t_R g5229 ( 
.A(n_3489),
.Y(n_5229)
);

INVx4_ASAP7_75t_L g5230 ( 
.A(n_3850),
.Y(n_5230)
);

AND2x4_ASAP7_75t_L g5231 ( 
.A(n_3359),
.B(n_3601),
.Y(n_5231)
);

NAND2xp5_ASAP7_75t_L g5232 ( 
.A(n_3356),
.B(n_3357),
.Y(n_5232)
);

OAI21xp5_ASAP7_75t_L g5233 ( 
.A1(n_3307),
.A2(n_3454),
.B(n_3796),
.Y(n_5233)
);

HB1xp67_ASAP7_75t_L g5234 ( 
.A(n_3627),
.Y(n_5234)
);

BUFx2_ASAP7_75t_L g5235 ( 
.A(n_3275),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_3490),
.Y(n_5236)
);

BUFx4f_ASAP7_75t_L g5237 ( 
.A(n_3879),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_3356),
.B(n_3357),
.Y(n_5238)
);

CKINVDCx20_ASAP7_75t_R g5239 ( 
.A(n_3221),
.Y(n_5239)
);

NAND2x1p5_ASAP7_75t_L g5240 ( 
.A(n_3798),
.B(n_3806),
.Y(n_5240)
);

AND2x2_ASAP7_75t_L g5241 ( 
.A(n_3850),
.B(n_4074),
.Y(n_5241)
);

NAND2xp5_ASAP7_75t_L g5242 ( 
.A(n_3360),
.B(n_3364),
.Y(n_5242)
);

CKINVDCx14_ASAP7_75t_R g5243 ( 
.A(n_3565),
.Y(n_5243)
);

BUFx2_ASAP7_75t_L g5244 ( 
.A(n_3276),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_L g5245 ( 
.A(n_3360),
.B(n_3364),
.Y(n_5245)
);

BUFx4f_ASAP7_75t_SL g5246 ( 
.A(n_4003),
.Y(n_5246)
);

INVx1_ASAP7_75t_L g5247 ( 
.A(n_3490),
.Y(n_5247)
);

HB1xp67_ASAP7_75t_L g5248 ( 
.A(n_3627),
.Y(n_5248)
);

NAND2xp5_ASAP7_75t_L g5249 ( 
.A(n_3375),
.B(n_3396),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_3375),
.B(n_3396),
.Y(n_5250)
);

NAND2xp5_ASAP7_75t_L g5251 ( 
.A(n_3400),
.B(n_3411),
.Y(n_5251)
);

AND2x2_ASAP7_75t_L g5252 ( 
.A(n_4074),
.B(n_3276),
.Y(n_5252)
);

BUFx12f_ASAP7_75t_L g5253 ( 
.A(n_4003),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_3514),
.Y(n_5254)
);

BUFx4f_ASAP7_75t_SL g5255 ( 
.A(n_4003),
.Y(n_5255)
);

NAND2xp5_ASAP7_75t_L g5256 ( 
.A(n_3400),
.B(n_3411),
.Y(n_5256)
);

CKINVDCx5p33_ASAP7_75t_R g5257 ( 
.A(n_3883),
.Y(n_5257)
);

INVx1_ASAP7_75t_L g5258 ( 
.A(n_3514),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_L g5259 ( 
.A(n_3414),
.B(n_3419),
.Y(n_5259)
);

NAND2x1_ASAP7_75t_L g5260 ( 
.A(n_3815),
.B(n_3816),
.Y(n_5260)
);

NAND2xp5_ASAP7_75t_L g5261 ( 
.A(n_3414),
.B(n_3419),
.Y(n_5261)
);

BUFx2_ASAP7_75t_L g5262 ( 
.A(n_3254),
.Y(n_5262)
);

NAND2xp5_ASAP7_75t_SL g5263 ( 
.A(n_3343),
.B(n_3355),
.Y(n_5263)
);

INVx1_ASAP7_75t_L g5264 ( 
.A(n_3516),
.Y(n_5264)
);

NOR2xp33_ASAP7_75t_L g5265 ( 
.A(n_3426),
.B(n_3384),
.Y(n_5265)
);

HB1xp67_ASAP7_75t_L g5266 ( 
.A(n_3385),
.Y(n_5266)
);

BUFx6f_ASAP7_75t_L g5267 ( 
.A(n_4074),
.Y(n_5267)
);

NAND2xp33_ASAP7_75t_L g5268 ( 
.A(n_3879),
.B(n_3450),
.Y(n_5268)
);

NAND2xp5_ASAP7_75t_L g5269 ( 
.A(n_3369),
.B(n_3392),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_3516),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_3369),
.B(n_3417),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_3446),
.B(n_3453),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_SL g5273 ( 
.A(n_3404),
.B(n_3385),
.Y(n_5273)
);

INVx1_ASAP7_75t_L g5274 ( 
.A(n_3519),
.Y(n_5274)
);

HB1xp67_ASAP7_75t_L g5275 ( 
.A(n_3422),
.Y(n_5275)
);

BUFx2_ASAP7_75t_L g5276 ( 
.A(n_3879),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_3334),
.B(n_3553),
.Y(n_5277)
);

AND2x2_ASAP7_75t_L g5278 ( 
.A(n_3334),
.B(n_3553),
.Y(n_5278)
);

NOR2xp33_ASAP7_75t_L g5279 ( 
.A(n_3420),
.B(n_3424),
.Y(n_5279)
);

NOR2x1_ASAP7_75t_L g5280 ( 
.A(n_3491),
.B(n_3422),
.Y(n_5280)
);

CKINVDCx20_ASAP7_75t_R g5281 ( 
.A(n_4003),
.Y(n_5281)
);

NAND2xp5_ASAP7_75t_L g5282 ( 
.A(n_3460),
.B(n_3431),
.Y(n_5282)
);

INVx1_ASAP7_75t_L g5283 ( 
.A(n_3541),
.Y(n_5283)
);

NAND2xp5_ASAP7_75t_L g5284 ( 
.A(n_3431),
.B(n_3433),
.Y(n_5284)
);

CKINVDCx5p33_ASAP7_75t_R g5285 ( 
.A(n_4350),
.Y(n_5285)
);

HB1xp67_ASAP7_75t_L g5286 ( 
.A(n_3101),
.Y(n_5286)
);

NAND2xp5_ASAP7_75t_L g5287 ( 
.A(n_3433),
.B(n_3440),
.Y(n_5287)
);

BUFx3_ASAP7_75t_L g5288 ( 
.A(n_3621),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_3440),
.B(n_3441),
.Y(n_5289)
);

NAND2xp5_ASAP7_75t_L g5290 ( 
.A(n_3441),
.B(n_3447),
.Y(n_5290)
);

AOI22xp5_ASAP7_75t_L g5291 ( 
.A1(n_3879),
.A2(n_3461),
.B1(n_3451),
.B2(n_3523),
.Y(n_5291)
);

INVx5_ASAP7_75t_L g5292 ( 
.A(n_3540),
.Y(n_5292)
);

NAND2xp5_ASAP7_75t_L g5293 ( 
.A(n_3447),
.B(n_3455),
.Y(n_5293)
);

BUFx3_ASAP7_75t_L g5294 ( 
.A(n_3621),
.Y(n_5294)
);

AOI22xp5_ASAP7_75t_L g5295 ( 
.A1(n_3879),
.A2(n_3918),
.B1(n_4007),
.B2(n_3085),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_3455),
.B(n_3496),
.Y(n_5296)
);

BUFx3_ASAP7_75t_L g5297 ( 
.A(n_4257),
.Y(n_5297)
);

INVxp67_ASAP7_75t_SL g5298 ( 
.A(n_4033),
.Y(n_5298)
);

AOI22xp5_ASAP7_75t_L g5299 ( 
.A1(n_3085),
.A2(n_3918),
.B1(n_4042),
.B2(n_4007),
.Y(n_5299)
);

BUFx8_ASAP7_75t_L g5300 ( 
.A(n_3319),
.Y(n_5300)
);

CKINVDCx5p33_ASAP7_75t_R g5301 ( 
.A(n_4350),
.Y(n_5301)
);

NAND2xp5_ASAP7_75t_L g5302 ( 
.A(n_3470),
.B(n_3492),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_3548),
.B(n_3554),
.Y(n_5303)
);

CKINVDCx5p33_ASAP7_75t_R g5304 ( 
.A(n_3556),
.Y(n_5304)
);

BUFx2_ASAP7_75t_L g5305 ( 
.A(n_3468),
.Y(n_5305)
);

NAND2xp5_ASAP7_75t_L g5306 ( 
.A(n_3548),
.B(n_3554),
.Y(n_5306)
);

NAND2xp5_ASAP7_75t_L g5307 ( 
.A(n_3560),
.B(n_3571),
.Y(n_5307)
);

HB1xp67_ASAP7_75t_L g5308 ( 
.A(n_3131),
.Y(n_5308)
);

NAND2xp5_ASAP7_75t_L g5309 ( 
.A(n_3580),
.B(n_3587),
.Y(n_5309)
);

CKINVDCx11_ASAP7_75t_R g5310 ( 
.A(n_3556),
.Y(n_5310)
);

AND2x4_ASAP7_75t_SL g5311 ( 
.A(n_3540),
.B(n_3569),
.Y(n_5311)
);

INVxp67_ASAP7_75t_SL g5312 ( 
.A(n_4035),
.Y(n_5312)
);

INVx1_ASAP7_75t_L g5313 ( 
.A(n_3587),
.Y(n_5313)
);

NAND2xp5_ASAP7_75t_L g5314 ( 
.A(n_3617),
.B(n_3588),
.Y(n_5314)
);

NAND2xp5_ASAP7_75t_L g5315 ( 
.A(n_3617),
.B(n_4035),
.Y(n_5315)
);

OR2x6_ASAP7_75t_L g5316 ( 
.A(n_4043),
.B(n_4047),
.Y(n_5316)
);

AND2x4_ASAP7_75t_L g5317 ( 
.A(n_3601),
.B(n_3606),
.Y(n_5317)
);

INVx2_ASAP7_75t_SL g5318 ( 
.A(n_3569),
.Y(n_5318)
);

INVx1_ASAP7_75t_L g5319 ( 
.A(n_3590),
.Y(n_5319)
);

INVx5_ASAP7_75t_L g5320 ( 
.A(n_3540),
.Y(n_5320)
);

AND2x4_ASAP7_75t_L g5321 ( 
.A(n_3601),
.B(n_3606),
.Y(n_5321)
);

AND2x4_ASAP7_75t_L g5322 ( 
.A(n_3606),
.B(n_3607),
.Y(n_5322)
);

CKINVDCx5p33_ASAP7_75t_R g5323 ( 
.A(n_3570),
.Y(n_5323)
);

INVx1_ASAP7_75t_L g5324 ( 
.A(n_3568),
.Y(n_5324)
);

INVx1_ASAP7_75t_L g5325 ( 
.A(n_3549),
.Y(n_5325)
);

NAND2xp5_ASAP7_75t_L g5326 ( 
.A(n_4043),
.B(n_4047),
.Y(n_5326)
);

NAND2xp5_ASAP7_75t_L g5327 ( 
.A(n_4070),
.B(n_4076),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_4070),
.B(n_4076),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_4080),
.B(n_4081),
.Y(n_5329)
);

INVx1_ASAP7_75t_SL g5330 ( 
.A(n_3363),
.Y(n_5330)
);

INVx1_ASAP7_75t_L g5331 ( 
.A(n_4080),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_4081),
.B(n_4082),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_L g5333 ( 
.A(n_4082),
.B(n_4083),
.Y(n_5333)
);

INVx1_ASAP7_75t_L g5334 ( 
.A(n_4083),
.Y(n_5334)
);

INVx1_ASAP7_75t_L g5335 ( 
.A(n_4091),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_4091),
.B(n_4092),
.Y(n_5336)
);

HB1xp67_ASAP7_75t_L g5337 ( 
.A(n_3182),
.Y(n_5337)
);

NAND2xp5_ASAP7_75t_L g5338 ( 
.A(n_4092),
.B(n_4102),
.Y(n_5338)
);

INVx1_ASAP7_75t_L g5339 ( 
.A(n_3562),
.Y(n_5339)
);

NAND2xp5_ASAP7_75t_L g5340 ( 
.A(n_4102),
.B(n_4294),
.Y(n_5340)
);

NOR2xp33_ASAP7_75t_R g5341 ( 
.A(n_3489),
.B(n_3661),
.Y(n_5341)
);

BUFx4f_ASAP7_75t_L g5342 ( 
.A(n_3569),
.Y(n_5342)
);

NAND2xp5_ASAP7_75t_L g5343 ( 
.A(n_4294),
.B(n_4298),
.Y(n_5343)
);

OAI22xp5_ASAP7_75t_L g5344 ( 
.A1(n_3521),
.A2(n_4042),
.B1(n_3504),
.B2(n_3452),
.Y(n_5344)
);

NAND2xp5_ASAP7_75t_L g5345 ( 
.A(n_4298),
.B(n_4300),
.Y(n_5345)
);

OAI21x1_ASAP7_75t_L g5346 ( 
.A1(n_4300),
.A2(n_4313),
.B(n_4305),
.Y(n_5346)
);

NOR2xp33_ASAP7_75t_L g5347 ( 
.A(n_3462),
.B(n_3319),
.Y(n_5347)
);

NAND2xp5_ASAP7_75t_L g5348 ( 
.A(n_4305),
.B(n_4313),
.Y(n_5348)
);

BUFx4f_ASAP7_75t_SL g5349 ( 
.A(n_4257),
.Y(n_5349)
);

CKINVDCx5p33_ASAP7_75t_R g5350 ( 
.A(n_4257),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_3564),
.Y(n_5351)
);

AND3x2_ASAP7_75t_SL g5352 ( 
.A(n_3662),
.B(n_3612),
.C(n_3599),
.Y(n_5352)
);

OAI22xp5_ASAP7_75t_L g5353 ( 
.A1(n_3521),
.A2(n_3500),
.B1(n_3363),
.B2(n_3471),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_4315),
.B(n_4320),
.Y(n_5354)
);

NAND2xp5_ASAP7_75t_L g5355 ( 
.A(n_4315),
.B(n_4320),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_3566),
.Y(n_5356)
);

AOI22xp33_ASAP7_75t_L g5357 ( 
.A1(n_3354),
.A2(n_3372),
.B1(n_3378),
.B2(n_3367),
.Y(n_5357)
);

INVx1_ASAP7_75t_L g5358 ( 
.A(n_3495),
.Y(n_5358)
);

NOR2xp33_ASAP7_75t_L g5359 ( 
.A(n_3459),
.B(n_3442),
.Y(n_5359)
);

HB1xp67_ASAP7_75t_L g5360 ( 
.A(n_3248),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_3495),
.Y(n_5361)
);

INVx1_ASAP7_75t_L g5362 ( 
.A(n_3511),
.Y(n_5362)
);

NAND2xp5_ASAP7_75t_L g5363 ( 
.A(n_4322),
.B(n_4325),
.Y(n_5363)
);

NAND2xp5_ASAP7_75t_L g5364 ( 
.A(n_4322),
.B(n_4325),
.Y(n_5364)
);

BUFx8_ASAP7_75t_L g5365 ( 
.A(n_3569),
.Y(n_5365)
);

AND2x4_ASAP7_75t_L g5366 ( 
.A(n_3606),
.B(n_3607),
.Y(n_5366)
);

NAND2xp5_ASAP7_75t_L g5367 ( 
.A(n_4329),
.B(n_4339),
.Y(n_5367)
);

NAND2xp5_ASAP7_75t_L g5368 ( 
.A(n_4329),
.B(n_4339),
.Y(n_5368)
);

NAND2xp5_ASAP7_75t_L g5369 ( 
.A(n_4342),
.B(n_4344),
.Y(n_5369)
);

CKINVDCx6p67_ASAP7_75t_R g5370 ( 
.A(n_3154),
.Y(n_5370)
);

INVx1_ASAP7_75t_L g5371 ( 
.A(n_3511),
.Y(n_5371)
);

INVx1_ASAP7_75t_L g5372 ( 
.A(n_3512),
.Y(n_5372)
);

INVx1_ASAP7_75t_L g5373 ( 
.A(n_3512),
.Y(n_5373)
);

INVx2_ASAP7_75t_SL g5374 ( 
.A(n_3569),
.Y(n_5374)
);

INVx1_ASAP7_75t_L g5375 ( 
.A(n_3539),
.Y(n_5375)
);

AND2x4_ASAP7_75t_SL g5376 ( 
.A(n_3569),
.B(n_3487),
.Y(n_5376)
);

NAND2xp5_ASAP7_75t_L g5377 ( 
.A(n_4342),
.B(n_4344),
.Y(n_5377)
);

BUFx12f_ASAP7_75t_L g5378 ( 
.A(n_4257),
.Y(n_5378)
);

HB1xp67_ASAP7_75t_L g5379 ( 
.A(n_3251),
.Y(n_5379)
);

NAND2xp5_ASAP7_75t_L g5380 ( 
.A(n_4347),
.B(n_4348),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_3539),
.Y(n_5381)
);

BUFx2_ASAP7_75t_L g5382 ( 
.A(n_3468),
.Y(n_5382)
);

BUFx3_ASAP7_75t_L g5383 ( 
.A(n_3663),
.Y(n_5383)
);

NAND2xp33_ASAP7_75t_L g5384 ( 
.A(n_3666),
.B(n_3555),
.Y(n_5384)
);

INVx1_ASAP7_75t_L g5385 ( 
.A(n_4347),
.Y(n_5385)
);

OR2x6_ASAP7_75t_L g5386 ( 
.A(n_4348),
.B(n_3820),
.Y(n_5386)
);

BUFx2_ASAP7_75t_L g5387 ( 
.A(n_3484),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_3824),
.B(n_3825),
.Y(n_5388)
);

INVx1_ASAP7_75t_L g5389 ( 
.A(n_3831),
.Y(n_5389)
);

INVx1_ASAP7_75t_L g5390 ( 
.A(n_3833),
.Y(n_5390)
);

INVx5_ASAP7_75t_L g5391 ( 
.A(n_3386),
.Y(n_5391)
);

INVxp67_ASAP7_75t_SL g5392 ( 
.A(n_3838),
.Y(n_5392)
);

BUFx4f_ASAP7_75t_L g5393 ( 
.A(n_4090),
.Y(n_5393)
);

BUFx2_ASAP7_75t_L g5394 ( 
.A(n_3484),
.Y(n_5394)
);

A2O1A1Ixp33_ASAP7_75t_L g5395 ( 
.A1(n_3840),
.A2(n_3849),
.B(n_3853),
.C(n_3846),
.Y(n_5395)
);

NAND2xp5_ASAP7_75t_L g5396 ( 
.A(n_3857),
.B(n_3859),
.Y(n_5396)
);

INVx1_ASAP7_75t_L g5397 ( 
.A(n_3596),
.Y(n_5397)
);

NAND2xp5_ASAP7_75t_L g5398 ( 
.A(n_3866),
.B(n_3867),
.Y(n_5398)
);

NAND2xp5_ASAP7_75t_L g5399 ( 
.A(n_3871),
.B(n_3873),
.Y(n_5399)
);

INVxp67_ASAP7_75t_L g5400 ( 
.A(n_3445),
.Y(n_5400)
);

NAND2x1p5_ASAP7_75t_L g5401 ( 
.A(n_3878),
.B(n_3885),
.Y(n_5401)
);

NOR2xp33_ASAP7_75t_L g5402 ( 
.A(n_3443),
.B(n_3598),
.Y(n_5402)
);

AND2x4_ASAP7_75t_L g5403 ( 
.A(n_3607),
.B(n_3888),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_3596),
.Y(n_5404)
);

INVx1_ASAP7_75t_L g5405 ( 
.A(n_3593),
.Y(n_5405)
);

NAND2xp5_ASAP7_75t_SL g5406 ( 
.A(n_3592),
.B(n_3594),
.Y(n_5406)
);

NAND2xp5_ASAP7_75t_L g5407 ( 
.A(n_3893),
.B(n_3894),
.Y(n_5407)
);

AOI22xp5_ASAP7_75t_L g5408 ( 
.A1(n_3438),
.A2(n_3432),
.B1(n_3448),
.B2(n_3367),
.Y(n_5408)
);

BUFx3_ASAP7_75t_L g5409 ( 
.A(n_3663),
.Y(n_5409)
);

NAND2xp5_ASAP7_75t_L g5410 ( 
.A(n_3899),
.B(n_3902),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_3494),
.Y(n_5411)
);

AND2x4_ASAP7_75t_L g5412 ( 
.A(n_3607),
.B(n_3904),
.Y(n_5412)
);

INVx2_ASAP7_75t_SL g5413 ( 
.A(n_3388),
.Y(n_5413)
);

AOI211xp5_ASAP7_75t_L g5414 ( 
.A1(n_3639),
.A2(n_3537),
.B(n_3613),
.C(n_3665),
.Y(n_5414)
);

INVx1_ASAP7_75t_SL g5415 ( 
.A(n_3578),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_3494),
.Y(n_5416)
);

INVx6_ASAP7_75t_L g5417 ( 
.A(n_3487),
.Y(n_5417)
);

NAND2xp5_ASAP7_75t_L g5418 ( 
.A(n_3905),
.B(n_3910),
.Y(n_5418)
);

NAND2xp5_ASAP7_75t_L g5419 ( 
.A(n_3913),
.B(n_3923),
.Y(n_5419)
);

NOR2xp33_ASAP7_75t_L g5420 ( 
.A(n_3598),
.B(n_3584),
.Y(n_5420)
);

INVx1_ASAP7_75t_L g5421 ( 
.A(n_3928),
.Y(n_5421)
);

NOR2xp33_ASAP7_75t_SL g5422 ( 
.A(n_3673),
.B(n_4263),
.Y(n_5422)
);

NAND2xp5_ASAP7_75t_L g5423 ( 
.A(n_3929),
.B(n_3931),
.Y(n_5423)
);

HB1xp67_ASAP7_75t_L g5424 ( 
.A(n_3269),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_L g5425 ( 
.A(n_3936),
.B(n_3943),
.Y(n_5425)
);

OR2x2_ASAP7_75t_L g5426 ( 
.A(n_3946),
.B(n_3951),
.Y(n_5426)
);

NAND2xp5_ASAP7_75t_SL g5427 ( 
.A(n_3389),
.B(n_3515),
.Y(n_5427)
);

AOI221xp5_ASAP7_75t_L g5428 ( 
.A1(n_3321),
.A2(n_3911),
.B1(n_3722),
.B2(n_3763),
.C(n_3811),
.Y(n_5428)
);

NAND2xp5_ASAP7_75t_L g5429 ( 
.A(n_3962),
.B(n_3972),
.Y(n_5429)
);

NAND2xp5_ASAP7_75t_L g5430 ( 
.A(n_3975),
.B(n_3976),
.Y(n_5430)
);

INVx1_ASAP7_75t_L g5431 ( 
.A(n_3978),
.Y(n_5431)
);

OAI221xp5_ASAP7_75t_L g5432 ( 
.A1(n_3987),
.A2(n_4162),
.B1(n_4203),
.B2(n_4204),
.C(n_4155),
.Y(n_5432)
);

INVx1_ASAP7_75t_L g5433 ( 
.A(n_3988),
.Y(n_5433)
);

OR2x6_ASAP7_75t_L g5434 ( 
.A(n_3990),
.B(n_3991),
.Y(n_5434)
);

BUFx2_ASAP7_75t_L g5435 ( 
.A(n_3864),
.Y(n_5435)
);

INVx1_ASAP7_75t_L g5436 ( 
.A(n_3992),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_4002),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_4004),
.B(n_4013),
.Y(n_5438)
);

INVxp67_ASAP7_75t_L g5439 ( 
.A(n_3469),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_4015),
.Y(n_5440)
);

OAI22xp5_ASAP7_75t_SL g5441 ( 
.A1(n_3520),
.A2(n_3639),
.B1(n_3528),
.B2(n_3561),
.Y(n_5441)
);

HB1xp67_ASAP7_75t_L g5442 ( 
.A(n_4060),
.Y(n_5442)
);

NAND2xp5_ASAP7_75t_L g5443 ( 
.A(n_4017),
.B(n_4027),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_4105),
.B(n_4112),
.Y(n_5444)
);

HB1xp67_ASAP7_75t_L g5445 ( 
.A(n_4065),
.Y(n_5445)
);

AND2x2_ASAP7_75t_SL g5446 ( 
.A(n_3388),
.B(n_3435),
.Y(n_5446)
);

NAND2xp5_ASAP7_75t_L g5447 ( 
.A(n_4114),
.B(n_4119),
.Y(n_5447)
);

INVx1_ASAP7_75t_L g5448 ( 
.A(n_4122),
.Y(n_5448)
);

O2A1O1Ixp33_ASAP7_75t_L g5449 ( 
.A1(n_3501),
.A2(n_3657),
.B(n_3559),
.C(n_3677),
.Y(n_5449)
);

INVx1_ASAP7_75t_L g5450 ( 
.A(n_4123),
.Y(n_5450)
);

BUFx3_ASAP7_75t_L g5451 ( 
.A(n_3665),
.Y(n_5451)
);

CKINVDCx5p33_ASAP7_75t_R g5452 ( 
.A(n_3669),
.Y(n_5452)
);

INVx1_ASAP7_75t_SL g5453 ( 
.A(n_3624),
.Y(n_5453)
);

BUFx2_ASAP7_75t_L g5454 ( 
.A(n_4077),
.Y(n_5454)
);

NAND2xp5_ASAP7_75t_L g5455 ( 
.A(n_4127),
.B(n_4137),
.Y(n_5455)
);

NAND2xp5_ASAP7_75t_SL g5456 ( 
.A(n_3473),
.B(n_3618),
.Y(n_5456)
);

NAND2xp5_ASAP7_75t_SL g5457 ( 
.A(n_3618),
.B(n_3616),
.Y(n_5457)
);

BUFx4f_ASAP7_75t_L g5458 ( 
.A(n_4090),
.Y(n_5458)
);

CKINVDCx5p33_ASAP7_75t_R g5459 ( 
.A(n_3684),
.Y(n_5459)
);

NAND2xp5_ASAP7_75t_L g5460 ( 
.A(n_4140),
.B(n_4141),
.Y(n_5460)
);

BUFx3_ASAP7_75t_L g5461 ( 
.A(n_3622),
.Y(n_5461)
);

INVx1_ASAP7_75t_L g5462 ( 
.A(n_4153),
.Y(n_5462)
);

AOI22xp33_ASAP7_75t_L g5463 ( 
.A1(n_3354),
.A2(n_3378),
.B1(n_3383),
.B2(n_3372),
.Y(n_5463)
);

NOR2xp33_ASAP7_75t_L g5464 ( 
.A(n_3679),
.B(n_3448),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_4165),
.B(n_4172),
.Y(n_5465)
);

HB1xp67_ASAP7_75t_L g5466 ( 
.A(n_4145),
.Y(n_5466)
);

BUFx3_ASAP7_75t_L g5467 ( 
.A(n_3622),
.Y(n_5467)
);

NAND2xp5_ASAP7_75t_L g5468 ( 
.A(n_4178),
.B(n_4183),
.Y(n_5468)
);

INVx2_ASAP7_75t_SL g5469 ( 
.A(n_3388),
.Y(n_5469)
);

INVx2_ASAP7_75t_L g5470 ( 
.A(n_4374),
.Y(n_5470)
);

INVx5_ASAP7_75t_L g5471 ( 
.A(n_4447),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_4794),
.Y(n_5472)
);

O2A1O1Ixp33_ASAP7_75t_L g5473 ( 
.A1(n_4516),
.A2(n_3677),
.B(n_3602),
.C(n_3613),
.Y(n_5473)
);

CKINVDCx5p33_ASAP7_75t_R g5474 ( 
.A(n_4623),
.Y(n_5474)
);

O2A1O1Ixp33_ASAP7_75t_L g5475 ( 
.A1(n_4516),
.A2(n_3536),
.B(n_3667),
.C(n_3659),
.Y(n_5475)
);

O2A1O1Ixp33_ASAP7_75t_L g5476 ( 
.A1(n_4559),
.A2(n_3667),
.B(n_3659),
.C(n_3558),
.Y(n_5476)
);

INVx2_ASAP7_75t_L g5477 ( 
.A(n_4374),
.Y(n_5477)
);

AND2x4_ASAP7_75t_L g5478 ( 
.A(n_4868),
.B(n_4186),
.Y(n_5478)
);

AND2x4_ASAP7_75t_L g5479 ( 
.A(n_4868),
.B(n_4189),
.Y(n_5479)
);

INVx1_ASAP7_75t_L g5480 ( 
.A(n_4794),
.Y(n_5480)
);

AOI22xp33_ASAP7_75t_L g5481 ( 
.A1(n_4377),
.A2(n_3405),
.B1(n_3383),
.B2(n_3510),
.Y(n_5481)
);

INVx2_ASAP7_75t_L g5482 ( 
.A(n_4374),
.Y(n_5482)
);

INVx2_ASAP7_75t_L g5483 ( 
.A(n_4374),
.Y(n_5483)
);

AOI22xp33_ASAP7_75t_L g5484 ( 
.A1(n_4377),
.A2(n_3405),
.B1(n_3600),
.B2(n_3506),
.Y(n_5484)
);

OAI22xp5_ASAP7_75t_L g5485 ( 
.A1(n_4396),
.A2(n_5201),
.B1(n_4397),
.B2(n_4753),
.Y(n_5485)
);

AOI22xp33_ASAP7_75t_L g5486 ( 
.A1(n_4380),
.A2(n_4160),
.B1(n_4196),
.B2(n_4292),
.Y(n_5486)
);

INVx5_ASAP7_75t_L g5487 ( 
.A(n_4447),
.Y(n_5487)
);

NOR2xp33_ASAP7_75t_L g5488 ( 
.A(n_4559),
.B(n_3533),
.Y(n_5488)
);

INVx1_ASAP7_75t_L g5489 ( 
.A(n_4794),
.Y(n_5489)
);

OAI22xp5_ASAP7_75t_L g5490 ( 
.A1(n_4396),
.A2(n_3388),
.B1(n_3435),
.B2(n_3611),
.Y(n_5490)
);

NOR2x1_ASAP7_75t_L g5491 ( 
.A(n_5263),
.B(n_4195),
.Y(n_5491)
);

NAND2x1p5_ASAP7_75t_L g5492 ( 
.A(n_4447),
.B(n_4223),
.Y(n_5492)
);

AOI21xp5_ASAP7_75t_L g5493 ( 
.A1(n_4483),
.A2(n_4233),
.B(n_4228),
.Y(n_5493)
);

AOI21xp5_ASAP7_75t_L g5494 ( 
.A1(n_4675),
.A2(n_4238),
.B(n_4236),
.Y(n_5494)
);

NAND2xp5_ASAP7_75t_L g5495 ( 
.A(n_5216),
.B(n_4239),
.Y(n_5495)
);

INVx1_ASAP7_75t_SL g5496 ( 
.A(n_4777),
.Y(n_5496)
);

CKINVDCx16_ASAP7_75t_R g5497 ( 
.A(n_4658),
.Y(n_5497)
);

INVx1_ASAP7_75t_L g5498 ( 
.A(n_4792),
.Y(n_5498)
);

AOI22xp33_ASAP7_75t_L g5499 ( 
.A1(n_4380),
.A2(n_4388),
.B1(n_4413),
.B2(n_4402),
.Y(n_5499)
);

HB1xp67_ASAP7_75t_L g5500 ( 
.A(n_4887),
.Y(n_5500)
);

INVx4_ASAP7_75t_L g5501 ( 
.A(n_4447),
.Y(n_5501)
);

NAND2xp5_ASAP7_75t_SL g5502 ( 
.A(n_4928),
.B(n_4242),
.Y(n_5502)
);

AOI22xp33_ASAP7_75t_L g5503 ( 
.A1(n_4388),
.A2(n_4254),
.B1(n_4265),
.B2(n_4291),
.Y(n_5503)
);

INVx6_ASAP7_75t_L g5504 ( 
.A(n_4529),
.Y(n_5504)
);

BUFx12f_ASAP7_75t_L g5505 ( 
.A(n_4443),
.Y(n_5505)
);

AOI221x1_ASAP7_75t_L g5506 ( 
.A1(n_5054),
.A2(n_4258),
.B1(n_4289),
.B2(n_4281),
.C(n_4253),
.Y(n_5506)
);

CKINVDCx16_ASAP7_75t_R g5507 ( 
.A(n_4658),
.Y(n_5507)
);

NAND2xp5_ASAP7_75t_L g5508 ( 
.A(n_5216),
.B(n_4261),
.Y(n_5508)
);

BUFx2_ASAP7_75t_SL g5509 ( 
.A(n_4861),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_4792),
.Y(n_5510)
);

OAI22xp5_ASAP7_75t_L g5511 ( 
.A1(n_5201),
.A2(n_3435),
.B1(n_3611),
.B2(n_3680),
.Y(n_5511)
);

HB1xp67_ASAP7_75t_L g5512 ( 
.A(n_4887),
.Y(n_5512)
);

INVx2_ASAP7_75t_L g5513 ( 
.A(n_4379),
.Y(n_5513)
);

OAI21x1_ASAP7_75t_SL g5514 ( 
.A1(n_4415),
.A2(n_3361),
.B(n_3336),
.Y(n_5514)
);

NOR2xp33_ASAP7_75t_L g5515 ( 
.A(n_4828),
.B(n_3551),
.Y(n_5515)
);

AOI22xp33_ASAP7_75t_L g5516 ( 
.A1(n_4413),
.A2(n_4272),
.B1(n_4266),
.B2(n_3671),
.Y(n_5516)
);

INVx1_ASAP7_75t_L g5517 ( 
.A(n_4792),
.Y(n_5517)
);

OAI22xp5_ASAP7_75t_SL g5518 ( 
.A1(n_4697),
.A2(n_3670),
.B1(n_3687),
.B2(n_3672),
.Y(n_5518)
);

AOI22xp5_ASAP7_75t_L g5519 ( 
.A1(n_4625),
.A2(n_3610),
.B1(n_3608),
.B2(n_3605),
.Y(n_5519)
);

AND2x2_ASAP7_75t_L g5520 ( 
.A(n_5112),
.B(n_3599),
.Y(n_5520)
);

BUFx2_ASAP7_75t_SL g5521 ( 
.A(n_4861),
.Y(n_5521)
);

INVx1_ASAP7_75t_SL g5522 ( 
.A(n_4777),
.Y(n_5522)
);

INVx1_ASAP7_75t_SL g5523 ( 
.A(n_4839),
.Y(n_5523)
);

NAND2xp5_ASAP7_75t_L g5524 ( 
.A(n_4384),
.B(n_4393),
.Y(n_5524)
);

AOI22xp5_ASAP7_75t_L g5525 ( 
.A1(n_4625),
.A2(n_3610),
.B1(n_3605),
.B2(n_3608),
.Y(n_5525)
);

INVx2_ASAP7_75t_L g5526 ( 
.A(n_4379),
.Y(n_5526)
);

INVx2_ASAP7_75t_L g5527 ( 
.A(n_4379),
.Y(n_5527)
);

BUFx6f_ASAP7_75t_L g5528 ( 
.A(n_4444),
.Y(n_5528)
);

BUFx12f_ASAP7_75t_L g5529 ( 
.A(n_4443),
.Y(n_5529)
);

AOI21xp5_ASAP7_75t_L g5530 ( 
.A1(n_4724),
.A2(n_3435),
.B(n_3361),
.Y(n_5530)
);

INVx2_ASAP7_75t_SL g5531 ( 
.A(n_5292),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_4792),
.Y(n_5532)
);

O2A1O1Ixp5_ASAP7_75t_L g5533 ( 
.A1(n_5263),
.A2(n_3527),
.B(n_3509),
.C(n_3336),
.Y(n_5533)
);

BUFx6f_ASAP7_75t_L g5534 ( 
.A(n_4444),
.Y(n_5534)
);

NOR2xp33_ASAP7_75t_L g5535 ( 
.A(n_4828),
.B(n_3680),
.Y(n_5535)
);

BUFx6f_ASAP7_75t_L g5536 ( 
.A(n_4444),
.Y(n_5536)
);

INVx2_ASAP7_75t_L g5537 ( 
.A(n_4379),
.Y(n_5537)
);

CKINVDCx20_ASAP7_75t_R g5538 ( 
.A(n_5310),
.Y(n_5538)
);

AND2x2_ASAP7_75t_L g5539 ( 
.A(n_5112),
.B(n_3599),
.Y(n_5539)
);

INVx6_ASAP7_75t_L g5540 ( 
.A(n_4529),
.Y(n_5540)
);

CKINVDCx5p33_ASAP7_75t_R g5541 ( 
.A(n_4623),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_4385),
.Y(n_5542)
);

NAND2xp5_ASAP7_75t_SL g5543 ( 
.A(n_4928),
.B(n_3626),
.Y(n_5543)
);

O2A1O1Ixp33_ASAP7_75t_L g5544 ( 
.A1(n_4438),
.A2(n_3650),
.B(n_3658),
.C(n_3654),
.Y(n_5544)
);

AOI21xp33_ASAP7_75t_L g5545 ( 
.A1(n_4456),
.A2(n_3632),
.B(n_3678),
.Y(n_5545)
);

A2O1A1Ixp33_ASAP7_75t_SL g5546 ( 
.A1(n_4415),
.A2(n_3676),
.B(n_3678),
.C(n_3687),
.Y(n_5546)
);

CKINVDCx20_ASAP7_75t_R g5547 ( 
.A(n_5310),
.Y(n_5547)
);

BUFx6f_ASAP7_75t_L g5548 ( 
.A(n_4444),
.Y(n_5548)
);

AND2x2_ASAP7_75t_L g5549 ( 
.A(n_5112),
.B(n_3612),
.Y(n_5549)
);

OAI21xp33_ASAP7_75t_L g5550 ( 
.A1(n_4584),
.A2(n_3674),
.B(n_3675),
.Y(n_5550)
);

OR2x6_ASAP7_75t_L g5551 ( 
.A(n_4437),
.B(n_3626),
.Y(n_5551)
);

INVxp67_ASAP7_75t_L g5552 ( 
.A(n_4610),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4375),
.Y(n_5553)
);

INVx2_ASAP7_75t_L g5554 ( 
.A(n_4385),
.Y(n_5554)
);

OAI22x1_ASAP7_75t_L g5555 ( 
.A1(n_4479),
.A2(n_3655),
.B1(n_3678),
.B2(n_3672),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_4375),
.Y(n_5556)
);

BUFx6f_ASAP7_75t_L g5557 ( 
.A(n_4444),
.Y(n_5557)
);

AOI22xp33_ASAP7_75t_L g5558 ( 
.A1(n_4402),
.A2(n_3614),
.B1(n_3622),
.B2(n_3526),
.Y(n_5558)
);

BUFx6f_ASAP7_75t_L g5559 ( 
.A(n_4447),
.Y(n_5559)
);

INVx1_ASAP7_75t_L g5560 ( 
.A(n_4376),
.Y(n_5560)
);

INVx1_ASAP7_75t_L g5561 ( 
.A(n_4376),
.Y(n_5561)
);

INVx2_ASAP7_75t_L g5562 ( 
.A(n_4385),
.Y(n_5562)
);

INVx1_ASAP7_75t_L g5563 ( 
.A(n_4378),
.Y(n_5563)
);

INVx1_ASAP7_75t_L g5564 ( 
.A(n_4378),
.Y(n_5564)
);

O2A1O1Ixp33_ASAP7_75t_L g5565 ( 
.A1(n_4438),
.A2(n_3688),
.B(n_3675),
.C(n_3674),
.Y(n_5565)
);

AOI22xp33_ASAP7_75t_L g5566 ( 
.A1(n_4449),
.A2(n_3622),
.B1(n_3526),
.B2(n_3687),
.Y(n_5566)
);

NAND2xp33_ASAP7_75t_L g5567 ( 
.A(n_4464),
.B(n_3666),
.Y(n_5567)
);

BUFx6f_ASAP7_75t_L g5568 ( 
.A(n_4447),
.Y(n_5568)
);

INVx1_ASAP7_75t_L g5569 ( 
.A(n_4381),
.Y(n_5569)
);

BUFx6f_ASAP7_75t_L g5570 ( 
.A(n_4447),
.Y(n_5570)
);

BUFx2_ASAP7_75t_L g5571 ( 
.A(n_5124),
.Y(n_5571)
);

BUFx3_ASAP7_75t_L g5572 ( 
.A(n_5292),
.Y(n_5572)
);

INVx1_ASAP7_75t_L g5573 ( 
.A(n_4381),
.Y(n_5573)
);

INVx2_ASAP7_75t_L g5574 ( 
.A(n_4385),
.Y(n_5574)
);

O2A1O1Ixp33_ASAP7_75t_L g5575 ( 
.A1(n_4449),
.A2(n_3664),
.B(n_3668),
.C(n_3670),
.Y(n_5575)
);

INVxp67_ASAP7_75t_SL g5576 ( 
.A(n_5272),
.Y(n_5576)
);

NAND2x1p5_ASAP7_75t_L g5577 ( 
.A(n_4447),
.B(n_3487),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_4383),
.Y(n_5578)
);

CKINVDCx6p67_ASAP7_75t_R g5579 ( 
.A(n_5101),
.Y(n_5579)
);

BUFx2_ASAP7_75t_L g5580 ( 
.A(n_5124),
.Y(n_5580)
);

NAND2xp5_ASAP7_75t_L g5581 ( 
.A(n_4393),
.B(n_3546),
.Y(n_5581)
);

INVx2_ASAP7_75t_L g5582 ( 
.A(n_4387),
.Y(n_5582)
);

AND2x2_ASAP7_75t_L g5583 ( 
.A(n_5112),
.B(n_3612),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_5043),
.B(n_3573),
.Y(n_5584)
);

AOI21xp5_ASAP7_75t_L g5585 ( 
.A1(n_4745),
.A2(n_3481),
.B(n_3475),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_4383),
.Y(n_5586)
);

BUFx6f_ASAP7_75t_L g5587 ( 
.A(n_4373),
.Y(n_5587)
);

AO32x1_ASAP7_75t_L g5588 ( 
.A1(n_4807),
.A2(n_4810),
.A3(n_5032),
.B1(n_5031),
.B2(n_5035),
.Y(n_5588)
);

OAI22xp5_ASAP7_75t_L g5589 ( 
.A1(n_4397),
.A2(n_3670),
.B1(n_4276),
.B2(n_3102),
.Y(n_5589)
);

NOR2xp33_ASAP7_75t_L g5590 ( 
.A(n_4898),
.B(n_3603),
.Y(n_5590)
);

AOI221xp5_ASAP7_75t_L g5591 ( 
.A1(n_4540),
.A2(n_3581),
.B1(n_3577),
.B2(n_3518),
.C(n_3542),
.Y(n_5591)
);

INVx2_ASAP7_75t_SL g5592 ( 
.A(n_5292),
.Y(n_5592)
);

INVx2_ASAP7_75t_L g5593 ( 
.A(n_4387),
.Y(n_5593)
);

AO22x1_ASAP7_75t_L g5594 ( 
.A1(n_4612),
.A2(n_3487),
.B1(n_3102),
.B2(n_4267),
.Y(n_5594)
);

INVx2_ASAP7_75t_L g5595 ( 
.A(n_4406),
.Y(n_5595)
);

HB1xp67_ASAP7_75t_L g5596 ( 
.A(n_4386),
.Y(n_5596)
);

INVx1_ASAP7_75t_L g5597 ( 
.A(n_4403),
.Y(n_5597)
);

AOI21xp5_ASAP7_75t_L g5598 ( 
.A1(n_4745),
.A2(n_3437),
.B(n_3595),
.Y(n_5598)
);

NAND2xp5_ASAP7_75t_L g5599 ( 
.A(n_5043),
.B(n_3869),
.Y(n_5599)
);

NOR2xp33_ASAP7_75t_L g5600 ( 
.A(n_4898),
.B(n_3603),
.Y(n_5600)
);

NAND2xp5_ASAP7_75t_L g5601 ( 
.A(n_5169),
.B(n_3869),
.Y(n_5601)
);

CKINVDCx16_ASAP7_75t_R g5602 ( 
.A(n_4439),
.Y(n_5602)
);

AO221x2_ASAP7_75t_L g5603 ( 
.A1(n_5215),
.A2(n_3604),
.B1(n_3641),
.B2(n_3623),
.C(n_3630),
.Y(n_5603)
);

INVx3_ASAP7_75t_L g5604 ( 
.A(n_4674),
.Y(n_5604)
);

INVx4_ASAP7_75t_L g5605 ( 
.A(n_4519),
.Y(n_5605)
);

AOI21xp5_ASAP7_75t_L g5606 ( 
.A1(n_4758),
.A2(n_3437),
.B(n_3499),
.Y(n_5606)
);

NAND2xp5_ASAP7_75t_L g5607 ( 
.A(n_5169),
.B(n_3906),
.Y(n_5607)
);

AND2x2_ASAP7_75t_L g5608 ( 
.A(n_5112),
.B(n_3630),
.Y(n_5608)
);

AND2x2_ASAP7_75t_L g5609 ( 
.A(n_5123),
.B(n_3630),
.Y(n_5609)
);

INVx1_ASAP7_75t_L g5610 ( 
.A(n_4403),
.Y(n_5610)
);

INVx3_ASAP7_75t_L g5611 ( 
.A(n_4674),
.Y(n_5611)
);

OR2x2_ASAP7_75t_L g5612 ( 
.A(n_4807),
.B(n_3651),
.Y(n_5612)
);

INVx1_ASAP7_75t_L g5613 ( 
.A(n_4407),
.Y(n_5613)
);

HB1xp67_ASAP7_75t_L g5614 ( 
.A(n_4386),
.Y(n_5614)
);

AOI21xp5_ASAP7_75t_L g5615 ( 
.A1(n_4758),
.A2(n_3437),
.B(n_3502),
.Y(n_5615)
);

INVx1_ASAP7_75t_SL g5616 ( 
.A(n_4839),
.Y(n_5616)
);

AOI221xp5_ASAP7_75t_L g5617 ( 
.A1(n_4540),
.A2(n_3531),
.B1(n_3513),
.B2(n_3525),
.C(n_3534),
.Y(n_5617)
);

NAND2xp5_ASAP7_75t_L g5618 ( 
.A(n_4572),
.B(n_3906),
.Y(n_5618)
);

BUFx8_ASAP7_75t_L g5619 ( 
.A(n_5101),
.Y(n_5619)
);

NAND2xp5_ASAP7_75t_L g5620 ( 
.A(n_4572),
.B(n_3906),
.Y(n_5620)
);

AOI21xp5_ASAP7_75t_L g5621 ( 
.A1(n_4987),
.A2(n_3631),
.B(n_3633),
.Y(n_5621)
);

NAND2xp5_ASAP7_75t_L g5622 ( 
.A(n_4572),
.B(n_3964),
.Y(n_5622)
);

INVx4_ASAP7_75t_L g5623 ( 
.A(n_4519),
.Y(n_5623)
);

AOI22xp33_ASAP7_75t_L g5624 ( 
.A1(n_4450),
.A2(n_3597),
.B1(n_3684),
.B2(n_3625),
.Y(n_5624)
);

BUFx2_ASAP7_75t_L g5625 ( 
.A(n_4855),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_SL g5626 ( 
.A(n_4638),
.B(n_3664),
.Y(n_5626)
);

INVx4_ASAP7_75t_L g5627 ( 
.A(n_4519),
.Y(n_5627)
);

INVx1_ASAP7_75t_L g5628 ( 
.A(n_4407),
.Y(n_5628)
);

CKINVDCx20_ASAP7_75t_R g5629 ( 
.A(n_4513),
.Y(n_5629)
);

NAND2xp5_ASAP7_75t_L g5630 ( 
.A(n_5205),
.B(n_3964),
.Y(n_5630)
);

O2A1O1Ixp33_ASAP7_75t_L g5631 ( 
.A1(n_4450),
.A2(n_3668),
.B(n_3656),
.C(n_3681),
.Y(n_5631)
);

AND2x2_ASAP7_75t_L g5632 ( 
.A(n_5123),
.B(n_3651),
.Y(n_5632)
);

AOI222xp33_ASAP7_75t_L g5633 ( 
.A1(n_4587),
.A2(n_3106),
.B1(n_3686),
.B2(n_3102),
.C1(n_3856),
.C2(n_4109),
.Y(n_5633)
);

BUFx2_ASAP7_75t_L g5634 ( 
.A(n_4855),
.Y(n_5634)
);

AOI22xp33_ASAP7_75t_L g5635 ( 
.A1(n_4700),
.A2(n_3597),
.B1(n_3686),
.B2(n_3666),
.Y(n_5635)
);

NOR2xp33_ASAP7_75t_L g5636 ( 
.A(n_4844),
.B(n_3604),
.Y(n_5636)
);

NAND2xp5_ASAP7_75t_L g5637 ( 
.A(n_5205),
.B(n_3964),
.Y(n_5637)
);

INVx1_ASAP7_75t_L g5638 ( 
.A(n_4421),
.Y(n_5638)
);

INVx6_ASAP7_75t_L g5639 ( 
.A(n_4529),
.Y(n_5639)
);

HB1xp67_ASAP7_75t_L g5640 ( 
.A(n_4389),
.Y(n_5640)
);

NOR2xp33_ASAP7_75t_L g5641 ( 
.A(n_4844),
.B(n_3623),
.Y(n_5641)
);

INVx1_ASAP7_75t_L g5642 ( 
.A(n_4421),
.Y(n_5642)
);

AOI22xp33_ASAP7_75t_SL g5643 ( 
.A1(n_4538),
.A2(n_4428),
.B1(n_4582),
.B2(n_4545),
.Y(n_5643)
);

CKINVDCx6p67_ASAP7_75t_R g5644 ( 
.A(n_5101),
.Y(n_5644)
);

BUFx2_ASAP7_75t_L g5645 ( 
.A(n_4855),
.Y(n_5645)
);

BUFx12f_ASAP7_75t_L g5646 ( 
.A(n_4604),
.Y(n_5646)
);

AND2x2_ASAP7_75t_L g5647 ( 
.A(n_5123),
.B(n_3651),
.Y(n_5647)
);

CKINVDCx11_ASAP7_75t_R g5648 ( 
.A(n_4486),
.Y(n_5648)
);

INVx3_ASAP7_75t_L g5649 ( 
.A(n_4674),
.Y(n_5649)
);

O2A1O1Ixp33_ASAP7_75t_L g5650 ( 
.A1(n_4752),
.A2(n_3656),
.B(n_3681),
.C(n_3682),
.Y(n_5650)
);

OAI22xp5_ASAP7_75t_L g5651 ( 
.A1(n_4697),
.A2(n_4109),
.B1(n_3463),
.B2(n_3856),
.Y(n_5651)
);

INVx4_ASAP7_75t_L g5652 ( 
.A(n_4519),
.Y(n_5652)
);

OAI22xp5_ASAP7_75t_L g5653 ( 
.A1(n_4753),
.A2(n_4841),
.B1(n_4856),
.B2(n_4796),
.Y(n_5653)
);

NAND2xp5_ASAP7_75t_L g5654 ( 
.A(n_4398),
.B(n_3998),
.Y(n_5654)
);

OAI22xp5_ASAP7_75t_L g5655 ( 
.A1(n_4796),
.A2(n_4109),
.B1(n_3463),
.B2(n_3856),
.Y(n_5655)
);

NOR2xp33_ASAP7_75t_L g5656 ( 
.A(n_4816),
.B(n_3641),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_4429),
.Y(n_5657)
);

AND2x2_ASAP7_75t_L g5658 ( 
.A(n_5123),
.B(n_3998),
.Y(n_5658)
);

HB1xp67_ASAP7_75t_L g5659 ( 
.A(n_4389),
.Y(n_5659)
);

NAND2xp5_ASAP7_75t_L g5660 ( 
.A(n_4398),
.B(n_3998),
.Y(n_5660)
);

AOI21xp5_ASAP7_75t_L g5661 ( 
.A1(n_4987),
.A2(n_3631),
.B(n_3633),
.Y(n_5661)
);

INVx3_ASAP7_75t_SL g5662 ( 
.A(n_4967),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_4411),
.Y(n_5663)
);

OAI22xp5_ASAP7_75t_L g5664 ( 
.A1(n_4841),
.A2(n_3522),
.B1(n_3463),
.B2(n_4267),
.Y(n_5664)
);

OAI22xp5_ASAP7_75t_L g5665 ( 
.A1(n_4856),
.A2(n_5192),
.B1(n_4877),
.B2(n_4888),
.Y(n_5665)
);

BUFx3_ASAP7_75t_L g5666 ( 
.A(n_5292),
.Y(n_5666)
);

BUFx2_ASAP7_75t_L g5667 ( 
.A(n_4855),
.Y(n_5667)
);

INVx2_ASAP7_75t_L g5668 ( 
.A(n_4411),
.Y(n_5668)
);

INVx2_ASAP7_75t_SL g5669 ( 
.A(n_5292),
.Y(n_5669)
);

OAI21x1_ASAP7_75t_L g5670 ( 
.A1(n_5008),
.A2(n_3406),
.B(n_4336),
.Y(n_5670)
);

INVx2_ASAP7_75t_SL g5671 ( 
.A(n_5292),
.Y(n_5671)
);

OAI22xp5_ASAP7_75t_L g5672 ( 
.A1(n_5192),
.A2(n_3522),
.B1(n_4188),
.B2(n_4267),
.Y(n_5672)
);

BUFx3_ASAP7_75t_L g5673 ( 
.A(n_5320),
.Y(n_5673)
);

A2O1A1Ixp33_ASAP7_75t_L g5674 ( 
.A1(n_4456),
.A2(n_3682),
.B(n_3634),
.C(n_3648),
.Y(n_5674)
);

NAND2xp5_ASAP7_75t_SL g5675 ( 
.A(n_4638),
.B(n_4000),
.Y(n_5675)
);

INVx4_ASAP7_75t_L g5676 ( 
.A(n_4519),
.Y(n_5676)
);

AND2x2_ASAP7_75t_L g5677 ( 
.A(n_5123),
.B(n_4000),
.Y(n_5677)
);

OAI22xp5_ASAP7_75t_L g5678 ( 
.A1(n_4816),
.A2(n_3522),
.B1(n_3325),
.B2(n_4188),
.Y(n_5678)
);

INVx3_ASAP7_75t_L g5679 ( 
.A(n_4674),
.Y(n_5679)
);

NOR2xp67_ASAP7_75t_SL g5680 ( 
.A(n_5101),
.B(n_3097),
.Y(n_5680)
);

O2A1O1Ixp33_ASAP7_75t_L g5681 ( 
.A1(n_4752),
.A2(n_4464),
.B(n_4498),
.C(n_4526),
.Y(n_5681)
);

AOI21xp5_ASAP7_75t_L g5682 ( 
.A1(n_5272),
.A2(n_3634),
.B(n_3643),
.Y(n_5682)
);

INVx1_ASAP7_75t_L g5683 ( 
.A(n_4429),
.Y(n_5683)
);

CKINVDCx5p33_ASAP7_75t_R g5684 ( 
.A(n_4604),
.Y(n_5684)
);

INVx3_ASAP7_75t_L g5685 ( 
.A(n_4674),
.Y(n_5685)
);

AOI22xp5_ASAP7_75t_L g5686 ( 
.A1(n_4632),
.A2(n_3686),
.B1(n_3666),
.B2(n_4188),
.Y(n_5686)
);

O2A1O1Ixp33_ASAP7_75t_L g5687 ( 
.A1(n_4526),
.A2(n_3642),
.B(n_3653),
.C(n_3652),
.Y(n_5687)
);

BUFx2_ASAP7_75t_L g5688 ( 
.A(n_4855),
.Y(n_5688)
);

OAI22xp5_ASAP7_75t_L g5689 ( 
.A1(n_4877),
.A2(n_3325),
.B1(n_4237),
.B2(n_3149),
.Y(n_5689)
);

BUFx2_ASAP7_75t_L g5690 ( 
.A(n_4855),
.Y(n_5690)
);

INVx3_ASAP7_75t_L g5691 ( 
.A(n_4684),
.Y(n_5691)
);

CKINVDCx6p67_ASAP7_75t_R g5692 ( 
.A(n_5253),
.Y(n_5692)
);

OAI22xp5_ASAP7_75t_L g5693 ( 
.A1(n_4893),
.A2(n_3325),
.B1(n_4237),
.B2(n_3149),
.Y(n_5693)
);

AOI21xp5_ASAP7_75t_L g5694 ( 
.A1(n_5146),
.A2(n_3643),
.B(n_3646),
.Y(n_5694)
);

INVx4_ASAP7_75t_L g5695 ( 
.A(n_4467),
.Y(n_5695)
);

INVx1_ASAP7_75t_L g5696 ( 
.A(n_4434),
.Y(n_5696)
);

BUFx4f_ASAP7_75t_L g5697 ( 
.A(n_5446),
.Y(n_5697)
);

HB1xp67_ASAP7_75t_L g5698 ( 
.A(n_4416),
.Y(n_5698)
);

INVx1_ASAP7_75t_SL g5699 ( 
.A(n_4590),
.Y(n_5699)
);

INVx2_ASAP7_75t_L g5700 ( 
.A(n_4417),
.Y(n_5700)
);

INVx1_ASAP7_75t_L g5701 ( 
.A(n_4434),
.Y(n_5701)
);

NOR2xp33_ASAP7_75t_L g5702 ( 
.A(n_4888),
.B(n_3624),
.Y(n_5702)
);

INVx2_ASAP7_75t_L g5703 ( 
.A(n_4417),
.Y(n_5703)
);

A2O1A1Ixp33_ASAP7_75t_L g5704 ( 
.A1(n_4685),
.A2(n_3646),
.B(n_3648),
.C(n_4237),
.Y(n_5704)
);

INVx2_ASAP7_75t_SL g5705 ( 
.A(n_5320),
.Y(n_5705)
);

NAND2xp5_ASAP7_75t_L g5706 ( 
.A(n_4401),
.B(n_4362),
.Y(n_5706)
);

O2A1O1Ixp33_ASAP7_75t_L g5707 ( 
.A1(n_4541),
.A2(n_3642),
.B(n_3652),
.C(n_3649),
.Y(n_5707)
);

AOI21xp5_ASAP7_75t_L g5708 ( 
.A1(n_5146),
.A2(n_3097),
.B(n_4290),
.Y(n_5708)
);

NAND2xp5_ASAP7_75t_L g5709 ( 
.A(n_4401),
.B(n_4336),
.Y(n_5709)
);

AOI21xp5_ASAP7_75t_L g5710 ( 
.A1(n_5166),
.A2(n_3097),
.B(n_4290),
.Y(n_5710)
);

INVx1_ASAP7_75t_L g5711 ( 
.A(n_4435),
.Y(n_5711)
);

CKINVDCx20_ASAP7_75t_R g5712 ( 
.A(n_4513),
.Y(n_5712)
);

BUFx10_ASAP7_75t_L g5713 ( 
.A(n_4967),
.Y(n_5713)
);

OAI22xp5_ASAP7_75t_L g5714 ( 
.A1(n_4893),
.A2(n_3097),
.B1(n_4290),
.B2(n_3149),
.Y(n_5714)
);

INVx3_ASAP7_75t_L g5715 ( 
.A(n_4684),
.Y(n_5715)
);

NAND2xp5_ASAP7_75t_L g5716 ( 
.A(n_5177),
.B(n_4245),
.Y(n_5716)
);

AND2x6_ASAP7_75t_L g5717 ( 
.A(n_4465),
.B(n_4279),
.Y(n_5717)
);

NAND2xp5_ASAP7_75t_L g5718 ( 
.A(n_5177),
.B(n_4245),
.Y(n_5718)
);

OA21x2_ASAP7_75t_L g5719 ( 
.A1(n_5346),
.A2(n_3406),
.B(n_3649),
.Y(n_5719)
);

INVx1_ASAP7_75t_L g5720 ( 
.A(n_4435),
.Y(n_5720)
);

A2O1A1Ixp33_ASAP7_75t_L g5721 ( 
.A1(n_4685),
.A2(n_4391),
.B(n_4436),
.C(n_4420),
.Y(n_5721)
);

AOI22xp5_ASAP7_75t_L g5722 ( 
.A1(n_4632),
.A2(n_3686),
.B1(n_3666),
.B2(n_3642),
.Y(n_5722)
);

NOR2xp33_ASAP7_75t_L g5723 ( 
.A(n_4541),
.B(n_3640),
.Y(n_5723)
);

INVx2_ASAP7_75t_L g5724 ( 
.A(n_4424),
.Y(n_5724)
);

NOR2xp33_ASAP7_75t_L g5725 ( 
.A(n_4730),
.B(n_3640),
.Y(n_5725)
);

NOR2xp33_ASAP7_75t_L g5726 ( 
.A(n_4730),
.B(n_3638),
.Y(n_5726)
);

INVx3_ASAP7_75t_L g5727 ( 
.A(n_4684),
.Y(n_5727)
);

HB1xp67_ASAP7_75t_L g5728 ( 
.A(n_4416),
.Y(n_5728)
);

OAI21xp5_ASAP7_75t_L g5729 ( 
.A1(n_4531),
.A2(n_4328),
.B(n_4302),
.Y(n_5729)
);

A2O1A1Ixp33_ASAP7_75t_L g5730 ( 
.A1(n_4391),
.A2(n_4328),
.B(n_4302),
.C(n_3205),
.Y(n_5730)
);

AOI21xp5_ASAP7_75t_L g5731 ( 
.A1(n_5166),
.A2(n_4290),
.B(n_3149),
.Y(n_5731)
);

INVx3_ASAP7_75t_L g5732 ( 
.A(n_4684),
.Y(n_5732)
);

CKINVDCx11_ASAP7_75t_R g5733 ( 
.A(n_4486),
.Y(n_5733)
);

AND2x4_ASAP7_75t_SL g5734 ( 
.A(n_5230),
.B(n_3474),
.Y(n_5734)
);

NOR2xp33_ASAP7_75t_L g5735 ( 
.A(n_4716),
.B(n_3636),
.Y(n_5735)
);

INVx3_ASAP7_75t_L g5736 ( 
.A(n_4684),
.Y(n_5736)
);

NOR2xp33_ASAP7_75t_L g5737 ( 
.A(n_4716),
.B(n_3636),
.Y(n_5737)
);

AOI222xp33_ASAP7_75t_L g5738 ( 
.A1(n_4587),
.A2(n_3106),
.B1(n_3666),
.B2(n_3635),
.C1(n_3628),
.C2(n_4181),
.Y(n_5738)
);

BUFx3_ASAP7_75t_L g5739 ( 
.A(n_5320),
.Y(n_5739)
);

NOR2xp33_ASAP7_75t_L g5740 ( 
.A(n_4805),
.B(n_3645),
.Y(n_5740)
);

O2A1O1Ixp33_ASAP7_75t_L g5741 ( 
.A1(n_5273),
.A2(n_3653),
.B(n_3645),
.C(n_3644),
.Y(n_5741)
);

NOR2x1_ASAP7_75t_L g5742 ( 
.A(n_4612),
.B(n_5173),
.Y(n_5742)
);

AOI22xp5_ASAP7_75t_L g5743 ( 
.A1(n_4665),
.A2(n_3635),
.B1(n_3628),
.B2(n_3713),
.Y(n_5743)
);

INVx1_ASAP7_75t_SL g5744 ( 
.A(n_4590),
.Y(n_5744)
);

NAND2xp5_ASAP7_75t_SL g5745 ( 
.A(n_4405),
.B(n_4245),
.Y(n_5745)
);

NAND2x1p5_ASAP7_75t_L g5746 ( 
.A(n_5320),
.B(n_3848),
.Y(n_5746)
);

AOI21xp5_ASAP7_75t_L g5747 ( 
.A1(n_5395),
.A2(n_3848),
.B(n_4181),
.Y(n_5747)
);

NAND2xp5_ASAP7_75t_SL g5748 ( 
.A(n_4405),
.B(n_4245),
.Y(n_5748)
);

O2A1O1Ixp33_ASAP7_75t_L g5749 ( 
.A1(n_5273),
.A2(n_3644),
.B(n_3638),
.C(n_4240),
.Y(n_5749)
);

A2O1A1Ixp33_ASAP7_75t_L g5750 ( 
.A1(n_4420),
.A2(n_4436),
.B(n_4470),
.C(n_4451),
.Y(n_5750)
);

OAI21xp5_ASAP7_75t_L g5751 ( 
.A1(n_4531),
.A2(n_3205),
.B(n_3291),
.Y(n_5751)
);

INVx3_ASAP7_75t_L g5752 ( 
.A(n_4496),
.Y(n_5752)
);

NAND2xp5_ASAP7_75t_SL g5753 ( 
.A(n_4409),
.B(n_4008),
.Y(n_5753)
);

AOI21xp5_ASAP7_75t_L g5754 ( 
.A1(n_5395),
.A2(n_3547),
.B(n_3333),
.Y(n_5754)
);

NAND2xp5_ASAP7_75t_L g5755 ( 
.A(n_5144),
.B(n_4279),
.Y(n_5755)
);

A2O1A1Ixp33_ASAP7_75t_L g5756 ( 
.A1(n_4451),
.A2(n_3291),
.B(n_4240),
.C(n_3365),
.Y(n_5756)
);

INVx3_ASAP7_75t_L g5757 ( 
.A(n_4496),
.Y(n_5757)
);

O2A1O1Ixp33_ASAP7_75t_L g5758 ( 
.A1(n_4683),
.A2(n_4216),
.B(n_3365),
.C(n_4149),
.Y(n_5758)
);

NOR2x1_ASAP7_75t_L g5759 ( 
.A(n_5173),
.B(n_4019),
.Y(n_5759)
);

INVx2_ASAP7_75t_SL g5760 ( 
.A(n_5320),
.Y(n_5760)
);

NOR2xp33_ASAP7_75t_L g5761 ( 
.A(n_4805),
.B(n_3619),
.Y(n_5761)
);

INVx2_ASAP7_75t_L g5762 ( 
.A(n_4424),
.Y(n_5762)
);

INVx2_ASAP7_75t_L g5763 ( 
.A(n_4424),
.Y(n_5763)
);

INVx2_ASAP7_75t_L g5764 ( 
.A(n_4425),
.Y(n_5764)
);

AO32x2_ASAP7_75t_L g5765 ( 
.A1(n_5060),
.A2(n_4678),
.A3(n_4770),
.B1(n_4693),
.B2(n_4574),
.Y(n_5765)
);

BUFx2_ASAP7_75t_L g5766 ( 
.A(n_5052),
.Y(n_5766)
);

INVx1_ASAP7_75t_SL g5767 ( 
.A(n_4594),
.Y(n_5767)
);

HB1xp67_ASAP7_75t_L g5768 ( 
.A(n_4488),
.Y(n_5768)
);

NAND2xp5_ASAP7_75t_L g5769 ( 
.A(n_5296),
.B(n_4019),
.Y(n_5769)
);

INVx4_ASAP7_75t_L g5770 ( 
.A(n_4467),
.Y(n_5770)
);

AOI21xp5_ASAP7_75t_L g5771 ( 
.A1(n_4762),
.A2(n_3333),
.B(n_3474),
.Y(n_5771)
);

BUFx2_ASAP7_75t_L g5772 ( 
.A(n_5052),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_4425),
.Y(n_5773)
);

AOI22xp5_ASAP7_75t_L g5774 ( 
.A1(n_4665),
.A2(n_3926),
.B1(n_4149),
.B2(n_3485),
.Y(n_5774)
);

INVx5_ASAP7_75t_L g5775 ( 
.A(n_4437),
.Y(n_5775)
);

HB1xp67_ASAP7_75t_L g5776 ( 
.A(n_4488),
.Y(n_5776)
);

INVx2_ASAP7_75t_L g5777 ( 
.A(n_4430),
.Y(n_5777)
);

NAND2xp5_ASAP7_75t_L g5778 ( 
.A(n_5296),
.B(n_4147),
.Y(n_5778)
);

A2O1A1Ixp33_ASAP7_75t_L g5779 ( 
.A1(n_4470),
.A2(n_4216),
.B(n_4045),
.C(n_3485),
.Y(n_5779)
);

AOI21xp5_ASAP7_75t_L g5780 ( 
.A1(n_4762),
.A2(n_4859),
.B(n_4787),
.Y(n_5780)
);

NAND2xp5_ASAP7_75t_L g5781 ( 
.A(n_5282),
.B(n_4147),
.Y(n_5781)
);

CKINVDCx16_ASAP7_75t_R g5782 ( 
.A(n_4439),
.Y(n_5782)
);

O2A1O1Ixp5_ASAP7_75t_SL g5783 ( 
.A1(n_4689),
.A2(n_4067),
.B(n_4019),
.C(n_3619),
.Y(n_5783)
);

BUFx2_ASAP7_75t_L g5784 ( 
.A(n_5052),
.Y(n_5784)
);

NAND2xp5_ASAP7_75t_L g5785 ( 
.A(n_5282),
.B(n_4067),
.Y(n_5785)
);

O2A1O1Ixp33_ASAP7_75t_L g5786 ( 
.A1(n_4683),
.A2(n_3713),
.B(n_4126),
.C(n_3529),
.Y(n_5786)
);

NOR2xp33_ASAP7_75t_L g5787 ( 
.A(n_5194),
.B(n_3619),
.Y(n_5787)
);

AND2x2_ASAP7_75t_L g5788 ( 
.A(n_5262),
.B(n_5235),
.Y(n_5788)
);

BUFx12f_ASAP7_75t_L g5789 ( 
.A(n_4649),
.Y(n_5789)
);

BUFx2_ASAP7_75t_L g5790 ( 
.A(n_5403),
.Y(n_5790)
);

INVx3_ASAP7_75t_L g5791 ( 
.A(n_4496),
.Y(n_5791)
);

OAI22xp5_ASAP7_75t_L g5792 ( 
.A1(n_4409),
.A2(n_3333),
.B1(n_3474),
.B2(n_4181),
.Y(n_5792)
);

NAND2x1_ASAP7_75t_SL g5793 ( 
.A(n_5211),
.B(n_3619),
.Y(n_5793)
);

NAND2xp5_ASAP7_75t_L g5794 ( 
.A(n_4863),
.B(n_3620),
.Y(n_5794)
);

NOR2xp33_ASAP7_75t_L g5795 ( 
.A(n_5194),
.B(n_5206),
.Y(n_5795)
);

AOI21xp5_ASAP7_75t_L g5796 ( 
.A1(n_4762),
.A2(n_3333),
.B(n_3474),
.Y(n_5796)
);

NOR2xp33_ASAP7_75t_L g5797 ( 
.A(n_5206),
.B(n_3620),
.Y(n_5797)
);

O2A1O1Ixp33_ASAP7_75t_L g5798 ( 
.A1(n_5060),
.A2(n_3529),
.B(n_3538),
.C(n_4126),
.Y(n_5798)
);

O2A1O1Ixp5_ASAP7_75t_SL g5799 ( 
.A1(n_4689),
.A2(n_4771),
.B(n_4786),
.C(n_4900),
.Y(n_5799)
);

AND3x1_ASAP7_75t_SL g5800 ( 
.A(n_4776),
.B(n_4181),
.C(n_3547),
.Y(n_5800)
);

BUFx2_ASAP7_75t_L g5801 ( 
.A(n_5403),
.Y(n_5801)
);

AOI21xp5_ASAP7_75t_L g5802 ( 
.A1(n_4762),
.A2(n_3848),
.B(n_3547),
.Y(n_5802)
);

NAND2xp5_ASAP7_75t_SL g5803 ( 
.A(n_5154),
.B(n_3848),
.Y(n_5803)
);

AND2x2_ASAP7_75t_L g5804 ( 
.A(n_5262),
.B(n_3620),
.Y(n_5804)
);

A2O1A1Ixp33_ASAP7_75t_L g5805 ( 
.A1(n_4476),
.A2(n_3538),
.B(n_4049),
.C(n_4045),
.Y(n_5805)
);

NOR2xp33_ASAP7_75t_L g5806 ( 
.A(n_4620),
.B(n_3620),
.Y(n_5806)
);

INVxp33_ASAP7_75t_SL g5807 ( 
.A(n_4649),
.Y(n_5807)
);

BUFx2_ASAP7_75t_L g5808 ( 
.A(n_5403),
.Y(n_5808)
);

AOI22xp33_ASAP7_75t_L g5809 ( 
.A1(n_4700),
.A2(n_3547),
.B1(n_3999),
.B2(n_3997),
.Y(n_5809)
);

AOI22xp33_ASAP7_75t_L g5810 ( 
.A1(n_4776),
.A2(n_3999),
.B1(n_3997),
.B2(n_3691),
.Y(n_5810)
);

HB1xp67_ASAP7_75t_L g5811 ( 
.A(n_5109),
.Y(n_5811)
);

OAI21xp33_ASAP7_75t_L g5812 ( 
.A1(n_4584),
.A2(n_3926),
.B(n_4049),
.Y(n_5812)
);

OAI221xp5_ASAP7_75t_L g5813 ( 
.A1(n_4636),
.A2(n_3691),
.B1(n_3941),
.B2(n_3997),
.C(n_3999),
.Y(n_5813)
);

AOI21xp5_ASAP7_75t_L g5814 ( 
.A1(n_4762),
.A2(n_3691),
.B(n_3941),
.Y(n_5814)
);

NAND2xp5_ASAP7_75t_L g5815 ( 
.A(n_4863),
.B(n_3620),
.Y(n_5815)
);

NAND2xp5_ASAP7_75t_L g5816 ( 
.A(n_4863),
.B(n_3620),
.Y(n_5816)
);

INVx4_ASAP7_75t_L g5817 ( 
.A(n_4467),
.Y(n_5817)
);

NOR2xp33_ASAP7_75t_L g5818 ( 
.A(n_4620),
.B(n_3647),
.Y(n_5818)
);

INVxp67_ASAP7_75t_SL g5819 ( 
.A(n_4904),
.Y(n_5819)
);

AOI21xp5_ASAP7_75t_L g5820 ( 
.A1(n_4762),
.A2(n_3691),
.B(n_3941),
.Y(n_5820)
);

AO21x1_ASAP7_75t_L g5821 ( 
.A1(n_4543),
.A2(n_3941),
.B(n_3997),
.Y(n_5821)
);

A2O1A1Ixp33_ASAP7_75t_L g5822 ( 
.A1(n_4476),
.A2(n_3647),
.B(n_3999),
.C(n_4478),
.Y(n_5822)
);

NOR2x1_ASAP7_75t_SL g5823 ( 
.A(n_5320),
.B(n_4465),
.Y(n_5823)
);

AOI22xp33_ASAP7_75t_L g5824 ( 
.A1(n_4538),
.A2(n_4707),
.B1(n_4764),
.B2(n_4673),
.Y(n_5824)
);

BUFx12f_ASAP7_75t_L g5825 ( 
.A(n_4695),
.Y(n_5825)
);

AOI21xp5_ASAP7_75t_L g5826 ( 
.A1(n_4762),
.A2(n_4859),
.B(n_4787),
.Y(n_5826)
);

HB1xp67_ASAP7_75t_L g5827 ( 
.A(n_5109),
.Y(n_5827)
);

BUFx2_ASAP7_75t_L g5828 ( 
.A(n_5403),
.Y(n_5828)
);

OR2x2_ASAP7_75t_L g5829 ( 
.A(n_4810),
.B(n_5235),
.Y(n_5829)
);

NAND2x1_ASAP7_75t_L g5830 ( 
.A(n_4412),
.B(n_4445),
.Y(n_5830)
);

OR2x6_ASAP7_75t_L g5831 ( 
.A(n_4437),
.B(n_5217),
.Y(n_5831)
);

OR2x2_ASAP7_75t_L g5832 ( 
.A(n_4810),
.B(n_5244),
.Y(n_5832)
);

NAND2xp5_ASAP7_75t_L g5833 ( 
.A(n_5269),
.B(n_5271),
.Y(n_5833)
);

NOR2xp33_ASAP7_75t_L g5834 ( 
.A(n_4922),
.B(n_4736),
.Y(n_5834)
);

OAI22xp33_ASAP7_75t_L g5835 ( 
.A1(n_4922),
.A2(n_4822),
.B1(n_4750),
.B2(n_4797),
.Y(n_5835)
);

OAI22xp5_ASAP7_75t_L g5836 ( 
.A1(n_4555),
.A2(n_4636),
.B1(n_4949),
.B2(n_5005),
.Y(n_5836)
);

INVx2_ASAP7_75t_SL g5837 ( 
.A(n_5217),
.Y(n_5837)
);

AOI21xp5_ASAP7_75t_L g5838 ( 
.A1(n_4787),
.A2(n_4917),
.B(n_4859),
.Y(n_5838)
);

INVx1_ASAP7_75t_SL g5839 ( 
.A(n_4594),
.Y(n_5839)
);

AOI22xp5_ASAP7_75t_L g5840 ( 
.A1(n_4890),
.A2(n_4921),
.B1(n_4791),
.B2(n_4707),
.Y(n_5840)
);

NAND2xp5_ASAP7_75t_L g5841 ( 
.A(n_5269),
.B(n_5271),
.Y(n_5841)
);

INVx3_ASAP7_75t_L g5842 ( 
.A(n_4496),
.Y(n_5842)
);

NAND2xp5_ASAP7_75t_L g5843 ( 
.A(n_4475),
.B(n_4482),
.Y(n_5843)
);

OAI22xp5_ASAP7_75t_L g5844 ( 
.A1(n_4555),
.A2(n_4949),
.B1(n_5005),
.B2(n_4448),
.Y(n_5844)
);

BUFx12f_ASAP7_75t_L g5845 ( 
.A(n_4695),
.Y(n_5845)
);

INVx2_ASAP7_75t_SL g5846 ( 
.A(n_5217),
.Y(n_5846)
);

CKINVDCx11_ASAP7_75t_R g5847 ( 
.A(n_4486),
.Y(n_5847)
);

O2A1O1Ixp5_ASAP7_75t_SL g5848 ( 
.A1(n_4771),
.A2(n_4786),
.B(n_4900),
.C(n_4736),
.Y(n_5848)
);

BUFx12f_ASAP7_75t_L g5849 ( 
.A(n_4699),
.Y(n_5849)
);

AOI21xp5_ASAP7_75t_L g5850 ( 
.A1(n_4787),
.A2(n_4917),
.B(n_4859),
.Y(n_5850)
);

BUFx12f_ASAP7_75t_L g5851 ( 
.A(n_4699),
.Y(n_5851)
);

AOI21xp5_ASAP7_75t_L g5852 ( 
.A1(n_4787),
.A2(n_4917),
.B(n_4859),
.Y(n_5852)
);

BUFx2_ASAP7_75t_L g5853 ( 
.A(n_5403),
.Y(n_5853)
);

NOR2xp33_ASAP7_75t_L g5854 ( 
.A(n_4890),
.B(n_5265),
.Y(n_5854)
);

NAND2xp5_ASAP7_75t_L g5855 ( 
.A(n_4475),
.B(n_4482),
.Y(n_5855)
);

OAI21x1_ASAP7_75t_SL g5856 ( 
.A1(n_5230),
.A2(n_5449),
.B(n_4394),
.Y(n_5856)
);

BUFx2_ASAP7_75t_L g5857 ( 
.A(n_5403),
.Y(n_5857)
);

NAND2xp5_ASAP7_75t_L g5858 ( 
.A(n_5025),
.B(n_5161),
.Y(n_5858)
);

NOR2xp67_ASAP7_75t_SL g5859 ( 
.A(n_5253),
.B(n_5378),
.Y(n_5859)
);

BUFx4_ASAP7_75t_SL g5860 ( 
.A(n_4737),
.Y(n_5860)
);

O2A1O1Ixp5_ASAP7_75t_L g5861 ( 
.A1(n_4705),
.A2(n_4821),
.B(n_5079),
.C(n_4846),
.Y(n_5861)
);

NAND2xp5_ASAP7_75t_L g5862 ( 
.A(n_5025),
.B(n_5161),
.Y(n_5862)
);

OAI22xp5_ASAP7_75t_L g5863 ( 
.A1(n_4448),
.A2(n_4822),
.B1(n_4921),
.B2(n_4791),
.Y(n_5863)
);

BUFx8_ASAP7_75t_L g5864 ( 
.A(n_5253),
.Y(n_5864)
);

INVx3_ASAP7_75t_L g5865 ( 
.A(n_4510),
.Y(n_5865)
);

INVx4_ASAP7_75t_L g5866 ( 
.A(n_4467),
.Y(n_5866)
);

NOR2xp33_ASAP7_75t_L g5867 ( 
.A(n_5265),
.B(n_4791),
.Y(n_5867)
);

OAI22xp5_ASAP7_75t_L g5868 ( 
.A1(n_4822),
.A2(n_4921),
.B1(n_4750),
.B2(n_4797),
.Y(n_5868)
);

OR2x6_ASAP7_75t_L g5869 ( 
.A(n_5217),
.B(n_5434),
.Y(n_5869)
);

OAI221xp5_ASAP7_75t_L g5870 ( 
.A1(n_4666),
.A2(n_4754),
.B1(n_4885),
.B2(n_4428),
.C(n_4582),
.Y(n_5870)
);

OR2x4_ASAP7_75t_L g5871 ( 
.A(n_4478),
.B(n_4511),
.Y(n_5871)
);

BUFx2_ASAP7_75t_SL g5872 ( 
.A(n_4861),
.Y(n_5872)
);

AOI21xp5_ASAP7_75t_L g5873 ( 
.A1(n_4787),
.A2(n_4917),
.B(n_4859),
.Y(n_5873)
);

NAND2xp5_ASAP7_75t_SL g5874 ( 
.A(n_5154),
.B(n_4394),
.Y(n_5874)
);

CKINVDCx11_ASAP7_75t_R g5875 ( 
.A(n_4726),
.Y(n_5875)
);

O2A1O1Ixp33_ASAP7_75t_L g5876 ( 
.A1(n_4666),
.A2(n_4885),
.B(n_4803),
.C(n_4872),
.Y(n_5876)
);

INVx1_ASAP7_75t_SL g5877 ( 
.A(n_4640),
.Y(n_5877)
);

CKINVDCx5p33_ASAP7_75t_R g5878 ( 
.A(n_4439),
.Y(n_5878)
);

AND2x4_ASAP7_75t_L g5879 ( 
.A(n_4510),
.B(n_4522),
.Y(n_5879)
);

BUFx2_ASAP7_75t_L g5880 ( 
.A(n_5412),
.Y(n_5880)
);

BUFx12f_ASAP7_75t_L g5881 ( 
.A(n_4702),
.Y(n_5881)
);

AND2x4_ASAP7_75t_L g5882 ( 
.A(n_4510),
.B(n_4522),
.Y(n_5882)
);

HB1xp67_ASAP7_75t_L g5883 ( 
.A(n_5109),
.Y(n_5883)
);

BUFx4f_ASAP7_75t_L g5884 ( 
.A(n_5446),
.Y(n_5884)
);

A2O1A1Ixp33_ASAP7_75t_L g5885 ( 
.A1(n_4511),
.A2(n_4535),
.B(n_4525),
.C(n_4563),
.Y(n_5885)
);

INVx4_ASAP7_75t_L g5886 ( 
.A(n_4467),
.Y(n_5886)
);

BUFx2_ASAP7_75t_L g5887 ( 
.A(n_5412),
.Y(n_5887)
);

OR2x6_ASAP7_75t_SL g5888 ( 
.A(n_4840),
.B(n_4870),
.Y(n_5888)
);

AOI22xp5_ASAP7_75t_L g5889 ( 
.A1(n_4673),
.A2(n_4764),
.B1(n_4783),
.B2(n_4545),
.Y(n_5889)
);

NAND2xp5_ASAP7_75t_SL g5890 ( 
.A(n_4394),
.B(n_5054),
.Y(n_5890)
);

NAND2xp5_ASAP7_75t_L g5891 ( 
.A(n_5030),
.B(n_5094),
.Y(n_5891)
);

O2A1O1Ixp33_ASAP7_75t_L g5892 ( 
.A1(n_4803),
.A2(n_4872),
.B(n_4813),
.C(n_4824),
.Y(n_5892)
);

O2A1O1Ixp33_ASAP7_75t_SL g5893 ( 
.A1(n_4466),
.A2(n_4534),
.B(n_4671),
.C(n_4543),
.Y(n_5893)
);

CKINVDCx5p33_ASAP7_75t_R g5894 ( 
.A(n_4439),
.Y(n_5894)
);

AOI22xp33_ASAP7_75t_L g5895 ( 
.A1(n_4538),
.A2(n_4783),
.B1(n_4535),
.B2(n_4525),
.Y(n_5895)
);

NAND2xp5_ASAP7_75t_L g5896 ( 
.A(n_5030),
.B(n_5094),
.Y(n_5896)
);

INVx4_ASAP7_75t_L g5897 ( 
.A(n_4467),
.Y(n_5897)
);

A2O1A1Ixp33_ASAP7_75t_SL g5898 ( 
.A1(n_4455),
.A2(n_5122),
.B(n_4563),
.C(n_5233),
.Y(n_5898)
);

HAxp5_ASAP7_75t_L g5899 ( 
.A(n_4785),
.B(n_5014),
.CON(n_5899),
.SN(n_5899)
);

NAND2xp5_ASAP7_75t_L g5900 ( 
.A(n_5162),
.B(n_4916),
.Y(n_5900)
);

AOI22xp33_ASAP7_75t_L g5901 ( 
.A1(n_4840),
.A2(n_4870),
.B1(n_4534),
.B2(n_4822),
.Y(n_5901)
);

INVx3_ASAP7_75t_L g5902 ( 
.A(n_4510),
.Y(n_5902)
);

CKINVDCx5p33_ASAP7_75t_R g5903 ( 
.A(n_4702),
.Y(n_5903)
);

INVx3_ASAP7_75t_L g5904 ( 
.A(n_4522),
.Y(n_5904)
);

INVx2_ASAP7_75t_SL g5905 ( 
.A(n_5217),
.Y(n_5905)
);

NAND2xp5_ASAP7_75t_L g5906 ( 
.A(n_5162),
.B(n_4916),
.Y(n_5906)
);

INVx3_ASAP7_75t_L g5907 ( 
.A(n_4522),
.Y(n_5907)
);

NOR2xp33_ASAP7_75t_L g5908 ( 
.A(n_4973),
.B(n_4980),
.Y(n_5908)
);

INVxp67_ASAP7_75t_L g5909 ( 
.A(n_4610),
.Y(n_5909)
);

NAND2xp5_ASAP7_75t_SL g5910 ( 
.A(n_4676),
.B(n_4754),
.Y(n_5910)
);

A2O1A1Ixp33_ASAP7_75t_SL g5911 ( 
.A1(n_4455),
.A2(n_5122),
.B(n_5233),
.C(n_4980),
.Y(n_5911)
);

O2A1O1Ixp33_ASAP7_75t_L g5912 ( 
.A1(n_4813),
.A2(n_4824),
.B(n_4818),
.C(n_4760),
.Y(n_5912)
);

NOR2xp33_ASAP7_75t_L g5913 ( 
.A(n_4973),
.B(n_5220),
.Y(n_5913)
);

CKINVDCx20_ASAP7_75t_R g5914 ( 
.A(n_4920),
.Y(n_5914)
);

NAND2xp5_ASAP7_75t_SL g5915 ( 
.A(n_4676),
.B(n_5302),
.Y(n_5915)
);

BUFx2_ASAP7_75t_L g5916 ( 
.A(n_5412),
.Y(n_5916)
);

OR2x2_ASAP7_75t_L g5917 ( 
.A(n_5315),
.B(n_5129),
.Y(n_5917)
);

OAI21x1_ASAP7_75t_SL g5918 ( 
.A1(n_5230),
.A2(n_5449),
.B(n_4939),
.Y(n_5918)
);

INVx3_ASAP7_75t_L g5919 ( 
.A(n_4522),
.Y(n_5919)
);

INVx3_ASAP7_75t_L g5920 ( 
.A(n_4522),
.Y(n_5920)
);

AOI22xp5_ASAP7_75t_L g5921 ( 
.A1(n_4818),
.A2(n_5215),
.B1(n_4466),
.B2(n_4518),
.Y(n_5921)
);

OAI22xp5_ASAP7_75t_L g5922 ( 
.A1(n_5220),
.A2(n_5215),
.B1(n_5000),
.B2(n_4691),
.Y(n_5922)
);

INVx5_ASAP7_75t_L g5923 ( 
.A(n_4412),
.Y(n_5923)
);

HB1xp67_ASAP7_75t_L g5924 ( 
.A(n_4904),
.Y(n_5924)
);

OAI21xp33_ASAP7_75t_L g5925 ( 
.A1(n_4691),
.A2(n_5302),
.B(n_5227),
.Y(n_5925)
);

BUFx2_ASAP7_75t_L g5926 ( 
.A(n_5412),
.Y(n_5926)
);

OAI221xp5_ASAP7_75t_L g5927 ( 
.A1(n_4479),
.A2(n_4643),
.B1(n_5227),
.B2(n_4518),
.C(n_4514),
.Y(n_5927)
);

AOI22xp5_ASAP7_75t_L g5928 ( 
.A1(n_4514),
.A2(n_4643),
.B1(n_4768),
.B2(n_5291),
.Y(n_5928)
);

AOI22xp5_ASAP7_75t_L g5929 ( 
.A1(n_4768),
.A2(n_5291),
.B1(n_5010),
.B2(n_5268),
.Y(n_5929)
);

INVx5_ASAP7_75t_L g5930 ( 
.A(n_4412),
.Y(n_5930)
);

NOR2xp33_ASAP7_75t_SL g5931 ( 
.A(n_5446),
.B(n_4502),
.Y(n_5931)
);

AOI221xp5_ASAP7_75t_L g5932 ( 
.A1(n_4460),
.A2(n_5000),
.B1(n_5023),
.B2(n_4939),
.C(n_4703),
.Y(n_5932)
);

OAI222xp33_ASAP7_75t_L g5933 ( 
.A1(n_4503),
.A2(n_4491),
.B1(n_4509),
.B2(n_5195),
.C1(n_4479),
.C2(n_5009),
.Y(n_5933)
);

AOI21xp5_ASAP7_75t_L g5934 ( 
.A1(n_4787),
.A2(n_4917),
.B(n_4859),
.Y(n_5934)
);

AOI222xp33_ASAP7_75t_L g5935 ( 
.A1(n_4460),
.A2(n_5268),
.B1(n_5441),
.B2(n_5086),
.C1(n_5023),
.C2(n_4503),
.Y(n_5935)
);

A2O1A1Ixp33_ASAP7_75t_L g5936 ( 
.A1(n_5237),
.A2(n_4491),
.B(n_4891),
.C(n_4760),
.Y(n_5936)
);

BUFx12f_ASAP7_75t_L g5937 ( 
.A(n_4857),
.Y(n_5937)
);

NOR2xp33_ASAP7_75t_L g5938 ( 
.A(n_5266),
.B(n_5010),
.Y(n_5938)
);

AOI21xp5_ASAP7_75t_L g5939 ( 
.A1(n_4917),
.A2(n_5034),
.B(n_4947),
.Y(n_5939)
);

A2O1A1Ixp33_ASAP7_75t_L g5940 ( 
.A1(n_5237),
.A2(n_5029),
.B(n_5040),
.C(n_4891),
.Y(n_5940)
);

INVx3_ASAP7_75t_L g5941 ( 
.A(n_4549),
.Y(n_5941)
);

INVx4_ASAP7_75t_L g5942 ( 
.A(n_4467),
.Y(n_5942)
);

AOI22xp33_ASAP7_75t_SL g5943 ( 
.A1(n_4419),
.A2(n_5237),
.B1(n_5276),
.B2(n_5229),
.Y(n_5943)
);

OAI22xp5_ASAP7_75t_L g5944 ( 
.A1(n_5237),
.A2(n_5229),
.B1(n_5009),
.B2(n_5295),
.Y(n_5944)
);

INVx1_ASAP7_75t_SL g5945 ( 
.A(n_4640),
.Y(n_5945)
);

AND2x4_ASAP7_75t_L g5946 ( 
.A(n_4549),
.B(n_5412),
.Y(n_5946)
);

NOR2xp33_ASAP7_75t_L g5947 ( 
.A(n_5266),
.B(n_4671),
.Y(n_5947)
);

BUFx10_ASAP7_75t_L g5948 ( 
.A(n_4967),
.Y(n_5948)
);

BUFx2_ASAP7_75t_L g5949 ( 
.A(n_5412),
.Y(n_5949)
);

A2O1A1Ixp33_ASAP7_75t_L g5950 ( 
.A1(n_5237),
.A2(n_5040),
.B(n_5029),
.C(n_4509),
.Y(n_5950)
);

AOI21xp5_ASAP7_75t_L g5951 ( 
.A1(n_4917),
.A2(n_5034),
.B(n_4947),
.Y(n_5951)
);

CKINVDCx20_ASAP7_75t_R g5952 ( 
.A(n_4920),
.Y(n_5952)
);

AOI22xp33_ASAP7_75t_L g5953 ( 
.A1(n_5441),
.A2(n_5344),
.B1(n_4419),
.B2(n_5086),
.Y(n_5953)
);

OAI21xp5_ASAP7_75t_L g5954 ( 
.A1(n_4558),
.A2(n_5174),
.B(n_4998),
.Y(n_5954)
);

AND2x4_ASAP7_75t_SL g5955 ( 
.A(n_5230),
.B(n_5226),
.Y(n_5955)
);

O2A1O1Ixp33_ASAP7_75t_L g5956 ( 
.A1(n_5344),
.A2(n_5427),
.B(n_5353),
.C(n_4573),
.Y(n_5956)
);

AND3x1_ASAP7_75t_SL g5957 ( 
.A(n_4670),
.B(n_5014),
.C(n_4785),
.Y(n_5957)
);

BUFx2_ASAP7_75t_L g5958 ( 
.A(n_4714),
.Y(n_5958)
);

OR2x4_ASAP7_75t_L g5959 ( 
.A(n_4473),
.B(n_4508),
.Y(n_5959)
);

INVx8_ASAP7_75t_L g5960 ( 
.A(n_4512),
.Y(n_5960)
);

AOI22x1_ASAP7_75t_L g5961 ( 
.A1(n_4950),
.A2(n_4995),
.B1(n_4882),
.B2(n_4932),
.Y(n_5961)
);

NOR2xp33_ASAP7_75t_L g5962 ( 
.A(n_4573),
.B(n_5427),
.Y(n_5962)
);

BUFx6f_ASAP7_75t_L g5963 ( 
.A(n_4458),
.Y(n_5963)
);

NAND2xp5_ASAP7_75t_SL g5964 ( 
.A(n_4967),
.B(n_4657),
.Y(n_5964)
);

NOR2xp33_ASAP7_75t_L g5965 ( 
.A(n_4473),
.B(n_4508),
.Y(n_5965)
);

INVx4_ASAP7_75t_L g5966 ( 
.A(n_4467),
.Y(n_5966)
);

AOI22xp5_ASAP7_75t_L g5967 ( 
.A1(n_4460),
.A2(n_5353),
.B1(n_4502),
.B2(n_4974),
.Y(n_5967)
);

AOI21xp5_ASAP7_75t_L g5968 ( 
.A1(n_4947),
.A2(n_5224),
.B(n_5034),
.Y(n_5968)
);

NAND2x1p5_ASAP7_75t_L g5969 ( 
.A(n_4412),
.B(n_4445),
.Y(n_5969)
);

O2A1O1Ixp33_ASAP7_75t_L g5970 ( 
.A1(n_5195),
.A2(n_5191),
.B(n_5174),
.C(n_5279),
.Y(n_5970)
);

NOR2xp33_ASAP7_75t_L g5971 ( 
.A(n_4473),
.B(n_4508),
.Y(n_5971)
);

BUFx2_ASAP7_75t_L g5972 ( 
.A(n_4714),
.Y(n_5972)
);

O2A1O1Ixp33_ASAP7_75t_L g5973 ( 
.A1(n_5191),
.A2(n_5279),
.B(n_5198),
.C(n_4657),
.Y(n_5973)
);

AOI21xp5_ASAP7_75t_L g5974 ( 
.A1(n_4947),
.A2(n_5224),
.B(n_5034),
.Y(n_5974)
);

BUFx6f_ASAP7_75t_L g5975 ( 
.A(n_4458),
.Y(n_5975)
);

AOI21xp5_ASAP7_75t_L g5976 ( 
.A1(n_4947),
.A2(n_5224),
.B(n_5034),
.Y(n_5976)
);

CKINVDCx11_ASAP7_75t_R g5977 ( 
.A(n_4726),
.Y(n_5977)
);

OR2x2_ASAP7_75t_L g5978 ( 
.A(n_5315),
.B(n_5129),
.Y(n_5978)
);

BUFx6f_ASAP7_75t_L g5979 ( 
.A(n_4458),
.Y(n_5979)
);

BUFx6f_ASAP7_75t_L g5980 ( 
.A(n_4458),
.Y(n_5980)
);

HB1xp67_ASAP7_75t_L g5981 ( 
.A(n_4958),
.Y(n_5981)
);

HB1xp67_ASAP7_75t_L g5982 ( 
.A(n_4958),
.Y(n_5982)
);

HB1xp67_ASAP7_75t_L g5983 ( 
.A(n_4507),
.Y(n_5983)
);

HB1xp67_ASAP7_75t_L g5984 ( 
.A(n_4507),
.Y(n_5984)
);

BUFx6f_ASAP7_75t_L g5985 ( 
.A(n_4458),
.Y(n_5985)
);

O2A1O1Ixp33_ASAP7_75t_L g5986 ( 
.A1(n_5198),
.A2(n_4907),
.B(n_5223),
.C(n_5218),
.Y(n_5986)
);

BUFx6f_ASAP7_75t_L g5987 ( 
.A(n_4458),
.Y(n_5987)
);

OAI22xp33_ASAP7_75t_L g5988 ( 
.A1(n_5295),
.A2(n_4972),
.B1(n_4558),
.B2(n_5276),
.Y(n_5988)
);

INVx2_ASAP7_75t_SL g5989 ( 
.A(n_4493),
.Y(n_5989)
);

O2A1O1Ixp33_ASAP7_75t_L g5990 ( 
.A1(n_4907),
.A2(n_5218),
.B(n_5232),
.C(n_5223),
.Y(n_5990)
);

INVx2_ASAP7_75t_SL g5991 ( 
.A(n_4493),
.Y(n_5991)
);

BUFx2_ASAP7_75t_L g5992 ( 
.A(n_4714),
.Y(n_5992)
);

BUFx3_ASAP7_75t_L g5993 ( 
.A(n_5461),
.Y(n_5993)
);

INVx2_ASAP7_75t_SL g5994 ( 
.A(n_4493),
.Y(n_5994)
);

AOI22xp33_ASAP7_75t_L g5995 ( 
.A1(n_4419),
.A2(n_4670),
.B1(n_4972),
.B2(n_5305),
.Y(n_5995)
);

HB1xp67_ASAP7_75t_L g5996 ( 
.A(n_4561),
.Y(n_5996)
);

AOI22xp33_ASAP7_75t_L g5997 ( 
.A1(n_5305),
.A2(n_5387),
.B1(n_5394),
.B2(n_5382),
.Y(n_5997)
);

BUFx6f_ASAP7_75t_L g5998 ( 
.A(n_4458),
.Y(n_5998)
);

AOI21xp5_ASAP7_75t_L g5999 ( 
.A1(n_4947),
.A2(n_5224),
.B(n_5034),
.Y(n_5999)
);

NAND2xp5_ASAP7_75t_L g6000 ( 
.A(n_5283),
.B(n_4404),
.Y(n_6000)
);

AOI221xp5_ASAP7_75t_L g6001 ( 
.A1(n_4703),
.A2(n_4821),
.B1(n_5079),
.B2(n_4846),
.C(n_4705),
.Y(n_6001)
);

NAND2xp5_ASAP7_75t_SL g6002 ( 
.A(n_4532),
.B(n_5414),
.Y(n_6002)
);

AOI22xp33_ASAP7_75t_L g6003 ( 
.A1(n_5305),
.A2(n_5387),
.B1(n_5394),
.B2(n_5382),
.Y(n_6003)
);

NAND2x1p5_ASAP7_75t_L g6004 ( 
.A(n_4412),
.B(n_4445),
.Y(n_6004)
);

HB1xp67_ASAP7_75t_L g6005 ( 
.A(n_4561),
.Y(n_6005)
);

AOI22xp33_ASAP7_75t_L g6006 ( 
.A1(n_5382),
.A2(n_5394),
.B1(n_5387),
.B2(n_4998),
.Y(n_6006)
);

AOI21xp5_ASAP7_75t_L g6007 ( 
.A1(n_4947),
.A2(n_5224),
.B(n_5034),
.Y(n_6007)
);

BUFx6f_ASAP7_75t_L g6008 ( 
.A(n_4458),
.Y(n_6008)
);

HB1xp67_ASAP7_75t_L g6009 ( 
.A(n_4568),
.Y(n_6009)
);

O2A1O1Ixp33_ASAP7_75t_L g6010 ( 
.A1(n_5232),
.A2(n_5242),
.B(n_5245),
.C(n_5238),
.Y(n_6010)
);

AND2x4_ASAP7_75t_L g6011 ( 
.A(n_4551),
.B(n_4578),
.Y(n_6011)
);

BUFx6f_ASAP7_75t_L g6012 ( 
.A(n_4463),
.Y(n_6012)
);

AOI22xp33_ASAP7_75t_L g6013 ( 
.A1(n_4998),
.A2(n_5341),
.B1(n_5045),
.B2(n_5062),
.Y(n_6013)
);

BUFx6f_ASAP7_75t_L g6014 ( 
.A(n_4463),
.Y(n_6014)
);

NOR2xp33_ASAP7_75t_L g6015 ( 
.A(n_4472),
.B(n_4474),
.Y(n_6015)
);

HB1xp67_ASAP7_75t_L g6016 ( 
.A(n_4568),
.Y(n_6016)
);

INVx2_ASAP7_75t_SL g6017 ( 
.A(n_4493),
.Y(n_6017)
);

BUFx8_ASAP7_75t_SL g6018 ( 
.A(n_4737),
.Y(n_6018)
);

INVx3_ASAP7_75t_L g6019 ( 
.A(n_4633),
.Y(n_6019)
);

INVx1_ASAP7_75t_SL g6020 ( 
.A(n_4647),
.Y(n_6020)
);

NOR2xp33_ASAP7_75t_L g6021 ( 
.A(n_4472),
.B(n_4474),
.Y(n_6021)
);

A2O1A1Ixp33_ASAP7_75t_L g6022 ( 
.A1(n_5276),
.A2(n_4532),
.B(n_5414),
.C(n_5074),
.Y(n_6022)
);

NOR2xp33_ASAP7_75t_L g6023 ( 
.A(n_5180),
.B(n_5275),
.Y(n_6023)
);

AOI21xp5_ASAP7_75t_L g6024 ( 
.A1(n_5224),
.A2(n_5316),
.B(n_5326),
.Y(n_6024)
);

A2O1A1Ixp33_ASAP7_75t_L g6025 ( 
.A1(n_5072),
.A2(n_5076),
.B(n_5080),
.C(n_5074),
.Y(n_6025)
);

BUFx6f_ASAP7_75t_L g6026 ( 
.A(n_4463),
.Y(n_6026)
);

CKINVDCx5p33_ASAP7_75t_R g6027 ( 
.A(n_5323),
.Y(n_6027)
);

INVx4_ASAP7_75t_L g6028 ( 
.A(n_4471),
.Y(n_6028)
);

OAI21x1_ASAP7_75t_L g6029 ( 
.A1(n_5008),
.A2(n_5346),
.B(n_4886),
.Y(n_6029)
);

OR2x6_ASAP7_75t_L g6030 ( 
.A(n_5434),
.B(n_5224),
.Y(n_6030)
);

INVx1_ASAP7_75t_SL g6031 ( 
.A(n_4647),
.Y(n_6031)
);

NOR2xp33_ASAP7_75t_L g6032 ( 
.A(n_5180),
.B(n_5275),
.Y(n_6032)
);

NOR2xp33_ASAP7_75t_L g6033 ( 
.A(n_5036),
.B(n_5158),
.Y(n_6033)
);

O2A1O1Ixp5_ASAP7_75t_L g6034 ( 
.A1(n_4705),
.A2(n_4821),
.B(n_5079),
.C(n_4846),
.Y(n_6034)
);

INVx8_ASAP7_75t_L g6035 ( 
.A(n_4512),
.Y(n_6035)
);

OA21x2_ASAP7_75t_L g6036 ( 
.A1(n_5346),
.A2(n_5327),
.B(n_5326),
.Y(n_6036)
);

O2A1O1Ixp33_ASAP7_75t_L g6037 ( 
.A1(n_5238),
.A2(n_5245),
.B(n_5249),
.C(n_5242),
.Y(n_6037)
);

AOI21xp5_ASAP7_75t_L g6038 ( 
.A1(n_5316),
.A2(n_5328),
.B(n_5327),
.Y(n_6038)
);

OR2x2_ASAP7_75t_L g6039 ( 
.A(n_5129),
.B(n_5328),
.Y(n_6039)
);

INVx4_ASAP7_75t_L g6040 ( 
.A(n_4471),
.Y(n_6040)
);

AOI21xp5_ASAP7_75t_L g6041 ( 
.A1(n_5316),
.A2(n_5332),
.B(n_5329),
.Y(n_6041)
);

BUFx6f_ASAP7_75t_L g6042 ( 
.A(n_4463),
.Y(n_6042)
);

AOI22xp33_ASAP7_75t_SL g6043 ( 
.A1(n_4926),
.A2(n_5341),
.B1(n_4897),
.B2(n_4932),
.Y(n_6043)
);

A2O1A1Ixp33_ASAP7_75t_L g6044 ( 
.A1(n_5072),
.A2(n_5076),
.B(n_5080),
.C(n_5074),
.Y(n_6044)
);

INVx4_ASAP7_75t_L g6045 ( 
.A(n_4471),
.Y(n_6045)
);

INVx1_ASAP7_75t_SL g6046 ( 
.A(n_4704),
.Y(n_6046)
);

NAND2xp5_ASAP7_75t_L g6047 ( 
.A(n_4404),
.B(n_4408),
.Y(n_6047)
);

BUFx6f_ASAP7_75t_L g6048 ( 
.A(n_4463),
.Y(n_6048)
);

BUFx8_ASAP7_75t_SL g6049 ( 
.A(n_5253),
.Y(n_6049)
);

AOI22xp33_ASAP7_75t_L g6050 ( 
.A1(n_4912),
.A2(n_5062),
.B1(n_5098),
.B2(n_5045),
.Y(n_6050)
);

NAND2xp33_ASAP7_75t_L g6051 ( 
.A(n_5213),
.B(n_4634),
.Y(n_6051)
);

CKINVDCx5p33_ASAP7_75t_R g6052 ( 
.A(n_5323),
.Y(n_6052)
);

NAND2xp5_ASAP7_75t_L g6053 ( 
.A(n_4408),
.B(n_4422),
.Y(n_6053)
);

NAND2xp5_ASAP7_75t_L g6054 ( 
.A(n_4422),
.B(n_4426),
.Y(n_6054)
);

NOR2xp33_ASAP7_75t_L g6055 ( 
.A(n_5036),
.B(n_5158),
.Y(n_6055)
);

NOR2xp33_ASAP7_75t_L g6056 ( 
.A(n_5033),
.B(n_5015),
.Y(n_6056)
);

NAND2xp5_ASAP7_75t_L g6057 ( 
.A(n_4426),
.B(n_4452),
.Y(n_6057)
);

AO21x2_ASAP7_75t_L g6058 ( 
.A1(n_5329),
.A2(n_5333),
.B(n_5332),
.Y(n_6058)
);

O2A1O1Ixp33_ASAP7_75t_L g6059 ( 
.A1(n_5249),
.A2(n_5251),
.B(n_5256),
.C(n_5250),
.Y(n_6059)
);

NOR2xp33_ASAP7_75t_L g6060 ( 
.A(n_5033),
.B(n_5015),
.Y(n_6060)
);

NOR2xp33_ASAP7_75t_R g6061 ( 
.A(n_4616),
.B(n_4668),
.Y(n_6061)
);

NOR2xp67_ASAP7_75t_L g6062 ( 
.A(n_5234),
.B(n_5248),
.Y(n_6062)
);

INVx1_ASAP7_75t_SL g6063 ( 
.A(n_4704),
.Y(n_6063)
);

AOI22xp33_ASAP7_75t_L g6064 ( 
.A1(n_4912),
.A2(n_5100),
.B1(n_5130),
.B2(n_5098),
.Y(n_6064)
);

A2O1A1Ixp33_ASAP7_75t_L g6065 ( 
.A1(n_5072),
.A2(n_5076),
.B(n_5080),
.C(n_5074),
.Y(n_6065)
);

CKINVDCx5p33_ASAP7_75t_R g6066 ( 
.A(n_4616),
.Y(n_6066)
);

NAND2xp5_ASAP7_75t_L g6067 ( 
.A(n_4452),
.B(n_4453),
.Y(n_6067)
);

AND2x2_ASAP7_75t_SL g6068 ( 
.A(n_4965),
.B(n_5027),
.Y(n_6068)
);

AOI21xp5_ASAP7_75t_L g6069 ( 
.A1(n_5316),
.A2(n_5336),
.B(n_5333),
.Y(n_6069)
);

BUFx2_ASAP7_75t_L g6070 ( 
.A(n_4720),
.Y(n_6070)
);

NAND2xp5_ASAP7_75t_L g6071 ( 
.A(n_4453),
.B(n_5167),
.Y(n_6071)
);

INVx4_ASAP7_75t_L g6072 ( 
.A(n_4471),
.Y(n_6072)
);

NAND2xp5_ASAP7_75t_L g6073 ( 
.A(n_5167),
.B(n_5171),
.Y(n_6073)
);

NAND2xp5_ASAP7_75t_L g6074 ( 
.A(n_5171),
.B(n_5172),
.Y(n_6074)
);

A2O1A1Ixp33_ASAP7_75t_L g6075 ( 
.A1(n_5072),
.A2(n_5076),
.B(n_5080),
.C(n_5074),
.Y(n_6075)
);

INVx3_ASAP7_75t_L g6076 ( 
.A(n_4633),
.Y(n_6076)
);

INVx1_ASAP7_75t_SL g6077 ( 
.A(n_4773),
.Y(n_6077)
);

OR2x2_ASAP7_75t_L g6078 ( 
.A(n_5336),
.B(n_5338),
.Y(n_6078)
);

BUFx2_ASAP7_75t_L g6079 ( 
.A(n_4720),
.Y(n_6079)
);

NOR2xp33_ASAP7_75t_L g6080 ( 
.A(n_5383),
.B(n_5409),
.Y(n_6080)
);

OAI21xp5_ASAP7_75t_L g6081 ( 
.A1(n_4558),
.A2(n_4865),
.B(n_4804),
.Y(n_6081)
);

BUFx6f_ASAP7_75t_L g6082 ( 
.A(n_4463),
.Y(n_6082)
);

INVx5_ASAP7_75t_SL g6083 ( 
.A(n_5446),
.Y(n_6083)
);

AOI22xp5_ASAP7_75t_L g6084 ( 
.A1(n_4974),
.A2(n_5359),
.B1(n_4827),
.B2(n_5422),
.Y(n_6084)
);

NAND2x2_ASAP7_75t_L g6085 ( 
.A(n_5297),
.B(n_5383),
.Y(n_6085)
);

NAND2xp5_ASAP7_75t_L g6086 ( 
.A(n_5172),
.B(n_5183),
.Y(n_6086)
);

OAI22xp33_ASAP7_75t_SL g6087 ( 
.A1(n_4882),
.A2(n_4932),
.B1(n_4948),
.B2(n_4897),
.Y(n_6087)
);

BUFx6f_ASAP7_75t_L g6088 ( 
.A(n_4463),
.Y(n_6088)
);

AOI221xp5_ASAP7_75t_L g6089 ( 
.A1(n_4703),
.A2(n_4830),
.B1(n_4819),
.B2(n_4895),
.C(n_4864),
.Y(n_6089)
);

NAND2xp5_ASAP7_75t_L g6090 ( 
.A(n_5183),
.B(n_5184),
.Y(n_6090)
);

O2A1O1Ixp33_ASAP7_75t_L g6091 ( 
.A1(n_5250),
.A2(n_5256),
.B(n_5259),
.C(n_5251),
.Y(n_6091)
);

O2A1O1Ixp33_ASAP7_75t_SL g6092 ( 
.A1(n_5413),
.A2(n_5469),
.B(n_4738),
.C(n_4999),
.Y(n_6092)
);

BUFx6f_ASAP7_75t_L g6093 ( 
.A(n_4463),
.Y(n_6093)
);

O2A1O1Ixp33_ASAP7_75t_L g6094 ( 
.A1(n_5259),
.A2(n_5261),
.B(n_5456),
.C(n_5319),
.Y(n_6094)
);

AOI22xp5_ASAP7_75t_L g6095 ( 
.A1(n_5359),
.A2(n_4827),
.B1(n_5422),
.B2(n_5347),
.Y(n_6095)
);

INVx2_ASAP7_75t_SL g6096 ( 
.A(n_4501),
.Y(n_6096)
);

OAI22x1_ASAP7_75t_L g6097 ( 
.A1(n_4954),
.A2(n_4897),
.B1(n_4948),
.B2(n_4882),
.Y(n_6097)
);

NOR2xp33_ASAP7_75t_L g6098 ( 
.A(n_5383),
.B(n_5409),
.Y(n_6098)
);

BUFx2_ASAP7_75t_L g6099 ( 
.A(n_4631),
.Y(n_6099)
);

O2A1O1Ixp33_ASAP7_75t_L g6100 ( 
.A1(n_5261),
.A2(n_5456),
.B(n_5319),
.C(n_4979),
.Y(n_6100)
);

NAND2xp5_ASAP7_75t_L g6101 ( 
.A(n_5184),
.B(n_5185),
.Y(n_6101)
);

NAND2xp5_ASAP7_75t_L g6102 ( 
.A(n_5185),
.B(n_5187),
.Y(n_6102)
);

INVxp67_ASAP7_75t_L g6103 ( 
.A(n_4637),
.Y(n_6103)
);

INVx3_ASAP7_75t_L g6104 ( 
.A(n_4633),
.Y(n_6104)
);

NOR2x1_ASAP7_75t_L g6105 ( 
.A(n_5211),
.B(n_5280),
.Y(n_6105)
);

A2O1A1Ixp33_ASAP7_75t_L g6106 ( 
.A1(n_5072),
.A2(n_5076),
.B(n_5080),
.C(n_5074),
.Y(n_6106)
);

CKINVDCx6p67_ASAP7_75t_R g6107 ( 
.A(n_5378),
.Y(n_6107)
);

AND2x2_ASAP7_75t_SL g6108 ( 
.A(n_4964),
.B(n_4965),
.Y(n_6108)
);

NAND2xp5_ASAP7_75t_L g6109 ( 
.A(n_5187),
.B(n_5189),
.Y(n_6109)
);

NOR2x1_ASAP7_75t_L g6110 ( 
.A(n_5280),
.B(n_4836),
.Y(n_6110)
);

OAI22xp5_ASAP7_75t_L g6111 ( 
.A1(n_5100),
.A2(n_5130),
.B1(n_5115),
.B2(n_5063),
.Y(n_6111)
);

NAND2xp5_ASAP7_75t_L g6112 ( 
.A(n_5189),
.B(n_5190),
.Y(n_6112)
);

OAI211xp5_ASAP7_75t_SL g6113 ( 
.A1(n_5299),
.A2(n_5428),
.B(n_5400),
.C(n_5408),
.Y(n_6113)
);

NAND2xp5_ASAP7_75t_L g6114 ( 
.A(n_5190),
.B(n_5199),
.Y(n_6114)
);

AOI21xp5_ASAP7_75t_L g6115 ( 
.A1(n_5316),
.A2(n_5343),
.B(n_5340),
.Y(n_6115)
);

CKINVDCx11_ASAP7_75t_R g6116 ( 
.A(n_4726),
.Y(n_6116)
);

O2A1O1Ixp5_ASAP7_75t_L g6117 ( 
.A1(n_4950),
.A2(n_4995),
.B(n_5457),
.C(n_5076),
.Y(n_6117)
);

BUFx6f_ASAP7_75t_L g6118 ( 
.A(n_4966),
.Y(n_6118)
);

INVx4_ASAP7_75t_L g6119 ( 
.A(n_4471),
.Y(n_6119)
);

O2A1O1Ixp33_ASAP7_75t_L g6120 ( 
.A1(n_4948),
.A2(n_4962),
.B(n_4964),
.C(n_4954),
.Y(n_6120)
);

BUFx4f_ASAP7_75t_L g6121 ( 
.A(n_4471),
.Y(n_6121)
);

NOR2x1_ASAP7_75t_L g6122 ( 
.A(n_4836),
.B(n_4975),
.Y(n_6122)
);

INVx2_ASAP7_75t_SL g6123 ( 
.A(n_4501),
.Y(n_6123)
);

NOR2xp33_ASAP7_75t_L g6124 ( 
.A(n_5383),
.B(n_5409),
.Y(n_6124)
);

O2A1O1Ixp5_ASAP7_75t_L g6125 ( 
.A1(n_5457),
.A2(n_5072),
.B(n_5080),
.C(n_5092),
.Y(n_6125)
);

BUFx8_ASAP7_75t_SL g6126 ( 
.A(n_5378),
.Y(n_6126)
);

CKINVDCx8_ASAP7_75t_R g6127 ( 
.A(n_4542),
.Y(n_6127)
);

NAND2xp5_ASAP7_75t_L g6128 ( 
.A(n_5199),
.B(n_5202),
.Y(n_6128)
);

O2A1O1Ixp5_ASAP7_75t_L g6129 ( 
.A1(n_5092),
.A2(n_5085),
.B(n_5088),
.C(n_5067),
.Y(n_6129)
);

NAND3xp33_ASAP7_75t_L g6130 ( 
.A(n_4804),
.B(n_4865),
.C(n_4954),
.Y(n_6130)
);

AND2x4_ASAP7_75t_L g6131 ( 
.A(n_4578),
.B(n_4602),
.Y(n_6131)
);

CKINVDCx20_ASAP7_75t_R g6132 ( 
.A(n_4738),
.Y(n_6132)
);

INVx4_ASAP7_75t_L g6133 ( 
.A(n_4471),
.Y(n_6133)
);

INVx2_ASAP7_75t_L g6134 ( 
.A(n_4536),
.Y(n_6134)
);

OR2x6_ASAP7_75t_SL g6135 ( 
.A(n_5145),
.B(n_5219),
.Y(n_6135)
);

CKINVDCx6p67_ASAP7_75t_R g6136 ( 
.A(n_5378),
.Y(n_6136)
);

CKINVDCx16_ASAP7_75t_R g6137 ( 
.A(n_4717),
.Y(n_6137)
);

BUFx6f_ASAP7_75t_SL g6138 ( 
.A(n_5230),
.Y(n_6138)
);

NAND2xp5_ASAP7_75t_SL g6139 ( 
.A(n_5178),
.B(n_5182),
.Y(n_6139)
);

INVx4_ASAP7_75t_L g6140 ( 
.A(n_4471),
.Y(n_6140)
);

O2A1O1Ixp33_ASAP7_75t_L g6141 ( 
.A1(n_4964),
.A2(n_4965),
.B(n_4979),
.C(n_4962),
.Y(n_6141)
);

OAI21xp5_ASAP7_75t_L g6142 ( 
.A1(n_5406),
.A2(n_4979),
.B(n_4962),
.Y(n_6142)
);

INVx4_ASAP7_75t_L g6143 ( 
.A(n_4484),
.Y(n_6143)
);

OAI22xp5_ASAP7_75t_L g6144 ( 
.A1(n_5063),
.A2(n_5115),
.B1(n_4461),
.B2(n_4462),
.Y(n_6144)
);

NOR2xp33_ASAP7_75t_L g6145 ( 
.A(n_5409),
.B(n_5145),
.Y(n_6145)
);

NAND2xp5_ASAP7_75t_L g6146 ( 
.A(n_5202),
.B(n_5204),
.Y(n_6146)
);

CKINVDCx5p33_ASAP7_75t_R g6147 ( 
.A(n_4668),
.Y(n_6147)
);

NOR2xp33_ASAP7_75t_L g6148 ( 
.A(n_4487),
.B(n_4492),
.Y(n_6148)
);

NAND2xp5_ASAP7_75t_L g6149 ( 
.A(n_5204),
.B(n_5207),
.Y(n_6149)
);

O2A1O1Ixp33_ASAP7_75t_L g6150 ( 
.A1(n_5027),
.A2(n_5400),
.B(n_4461),
.C(n_4462),
.Y(n_6150)
);

NOR2xp33_ASAP7_75t_L g6151 ( 
.A(n_4487),
.B(n_4492),
.Y(n_6151)
);

AND2x4_ASAP7_75t_L g6152 ( 
.A(n_4602),
.B(n_4605),
.Y(n_6152)
);

AOI21xp5_ASAP7_75t_L g6153 ( 
.A1(n_5345),
.A2(n_5354),
.B(n_5348),
.Y(n_6153)
);

NOR2xp33_ASAP7_75t_L g6154 ( 
.A(n_4495),
.B(n_4500),
.Y(n_6154)
);

AOI22xp33_ASAP7_75t_L g6155 ( 
.A1(n_4717),
.A2(n_4788),
.B1(n_4830),
.B2(n_4819),
.Y(n_6155)
);

NAND2xp5_ASAP7_75t_L g6156 ( 
.A(n_5207),
.B(n_5210),
.Y(n_6156)
);

INVx2_ASAP7_75t_SL g6157 ( 
.A(n_4501),
.Y(n_6157)
);

NAND2xp5_ASAP7_75t_L g6158 ( 
.A(n_5210),
.B(n_5236),
.Y(n_6158)
);

AOI21xp5_ASAP7_75t_L g6159 ( 
.A1(n_5348),
.A2(n_5355),
.B(n_5354),
.Y(n_6159)
);

AOI21xp5_ASAP7_75t_L g6160 ( 
.A1(n_5355),
.A2(n_5364),
.B(n_5363),
.Y(n_6160)
);

NOR2xp33_ASAP7_75t_L g6161 ( 
.A(n_4495),
.B(n_4500),
.Y(n_6161)
);

BUFx2_ASAP7_75t_SL g6162 ( 
.A(n_5297),
.Y(n_6162)
);

BUFx4f_ASAP7_75t_L g6163 ( 
.A(n_4484),
.Y(n_6163)
);

OR2x6_ASAP7_75t_L g6164 ( 
.A(n_5434),
.B(n_5386),
.Y(n_6164)
);

HB1xp67_ASAP7_75t_L g6165 ( 
.A(n_4571),
.Y(n_6165)
);

NAND2xp5_ASAP7_75t_L g6166 ( 
.A(n_5236),
.B(n_5247),
.Y(n_6166)
);

AOI21xp5_ASAP7_75t_L g6167 ( 
.A1(n_5363),
.A2(n_5367),
.B(n_5364),
.Y(n_6167)
);

INVx4_ASAP7_75t_L g6168 ( 
.A(n_4484),
.Y(n_6168)
);

AND2x4_ASAP7_75t_L g6169 ( 
.A(n_4602),
.B(n_4605),
.Y(n_6169)
);

OR2x2_ASAP7_75t_L g6170 ( 
.A(n_5367),
.B(n_5368),
.Y(n_6170)
);

INVx2_ASAP7_75t_L g6171 ( 
.A(n_4544),
.Y(n_6171)
);

INVxp67_ASAP7_75t_SL g6172 ( 
.A(n_4576),
.Y(n_6172)
);

AOI22xp5_ASAP7_75t_L g6173 ( 
.A1(n_5347),
.A2(n_4727),
.B1(n_4701),
.B2(n_5299),
.Y(n_6173)
);

AND2x2_ASAP7_75t_L g6174 ( 
.A(n_4494),
.B(n_4976),
.Y(n_6174)
);

BUFx4f_ASAP7_75t_L g6175 ( 
.A(n_4484),
.Y(n_6175)
);

AOI21xp5_ASAP7_75t_L g6176 ( 
.A1(n_5368),
.A2(n_5377),
.B(n_5369),
.Y(n_6176)
);

BUFx6f_ASAP7_75t_L g6177 ( 
.A(n_4966),
.Y(n_6177)
);

NOR2xp33_ASAP7_75t_L g6178 ( 
.A(n_4517),
.B(n_4520),
.Y(n_6178)
);

NOR2xp33_ASAP7_75t_L g6179 ( 
.A(n_4517),
.B(n_4520),
.Y(n_6179)
);

AOI21xp5_ASAP7_75t_L g6180 ( 
.A1(n_5369),
.A2(n_5380),
.B(n_5377),
.Y(n_6180)
);

NAND2xp5_ASAP7_75t_L g6181 ( 
.A(n_5247),
.B(n_5254),
.Y(n_6181)
);

INVxp67_ASAP7_75t_L g6182 ( 
.A(n_4637),
.Y(n_6182)
);

AOI22xp33_ASAP7_75t_L g6183 ( 
.A1(n_4788),
.A2(n_4830),
.B1(n_4819),
.B2(n_4864),
.Y(n_6183)
);

O2A1O1Ixp33_ASAP7_75t_L g6184 ( 
.A1(n_5027),
.A2(n_4469),
.B(n_4454),
.C(n_5178),
.Y(n_6184)
);

INVx2_ASAP7_75t_SL g6185 ( 
.A(n_4501),
.Y(n_6185)
);

NAND2xp5_ASAP7_75t_L g6186 ( 
.A(n_5254),
.B(n_5258),
.Y(n_6186)
);

INVxp67_ASAP7_75t_L g6187 ( 
.A(n_4654),
.Y(n_6187)
);

CKINVDCx5p33_ASAP7_75t_R g6188 ( 
.A(n_4718),
.Y(n_6188)
);

CKINVDCx5p33_ASAP7_75t_R g6189 ( 
.A(n_4718),
.Y(n_6189)
);

AO32x2_ASAP7_75t_L g6190 ( 
.A1(n_4678),
.A2(n_4693),
.A3(n_4770),
.B1(n_4574),
.B2(n_4505),
.Y(n_6190)
);

BUFx2_ASAP7_75t_L g6191 ( 
.A(n_4667),
.Y(n_6191)
);

NAND2xp5_ASAP7_75t_SL g6192 ( 
.A(n_5182),
.B(n_5197),
.Y(n_6192)
);

HB1xp67_ASAP7_75t_L g6193 ( 
.A(n_4571),
.Y(n_6193)
);

CKINVDCx5p33_ASAP7_75t_R g6194 ( 
.A(n_5304),
.Y(n_6194)
);

O2A1O1Ixp33_ASAP7_75t_L g6195 ( 
.A1(n_4454),
.A2(n_4469),
.B(n_5200),
.C(n_5197),
.Y(n_6195)
);

INVx4_ASAP7_75t_L g6196 ( 
.A(n_4484),
.Y(n_6196)
);

INVx4_ASAP7_75t_L g6197 ( 
.A(n_4484),
.Y(n_6197)
);

AOI22xp33_ASAP7_75t_L g6198 ( 
.A1(n_4864),
.A2(n_4895),
.B1(n_4960),
.B2(n_4929),
.Y(n_6198)
);

BUFx6f_ASAP7_75t_L g6199 ( 
.A(n_4966),
.Y(n_6199)
);

OAI31xp33_ASAP7_75t_SL g6200 ( 
.A1(n_4895),
.A2(n_4929),
.A3(n_4960),
.B(n_4761),
.Y(n_6200)
);

AND2x4_ASAP7_75t_L g6201 ( 
.A(n_4605),
.B(n_4656),
.Y(n_6201)
);

OAI22xp5_ASAP7_75t_L g6202 ( 
.A1(n_5408),
.A2(n_4523),
.B1(n_4524),
.B2(n_4521),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_4494),
.B(n_4976),
.Y(n_6203)
);

OAI22xp5_ASAP7_75t_L g6204 ( 
.A1(n_4521),
.A2(n_4524),
.B1(n_4530),
.B2(n_4523),
.Y(n_6204)
);

INVx3_ASAP7_75t_SL g6205 ( 
.A(n_5075),
.Y(n_6205)
);

NAND2x1p5_ASAP7_75t_L g6206 ( 
.A(n_4490),
.B(n_4542),
.Y(n_6206)
);

AO21x1_ASAP7_75t_L g6207 ( 
.A1(n_4690),
.A2(n_4709),
.B(n_5035),
.Y(n_6207)
);

A2O1A1Ixp33_ASAP7_75t_L g6208 ( 
.A1(n_5067),
.A2(n_5085),
.B(n_5095),
.C(n_5088),
.Y(n_6208)
);

AOI21xp5_ASAP7_75t_L g6209 ( 
.A1(n_5380),
.A2(n_5298),
.B(n_5119),
.Y(n_6209)
);

NAND2xp5_ASAP7_75t_L g6210 ( 
.A(n_5258),
.B(n_5264),
.Y(n_6210)
);

OAI22x1_ASAP7_75t_L g6211 ( 
.A1(n_5228),
.A2(n_4690),
.B1(n_4709),
.B2(n_5059),
.Y(n_6211)
);

BUFx6f_ASAP7_75t_L g6212 ( 
.A(n_4966),
.Y(n_6212)
);

O2A1O1Ixp33_ASAP7_75t_L g6213 ( 
.A1(n_5200),
.A2(n_4530),
.B(n_4537),
.C(n_4533),
.Y(n_6213)
);

BUFx4f_ASAP7_75t_L g6214 ( 
.A(n_4484),
.Y(n_6214)
);

BUFx2_ASAP7_75t_L g6215 ( 
.A(n_4977),
.Y(n_6215)
);

AOI22xp5_ASAP7_75t_L g6216 ( 
.A1(n_4701),
.A2(n_4727),
.B1(n_4446),
.B2(n_5402),
.Y(n_6216)
);

AOI21xp5_ASAP7_75t_L g6217 ( 
.A1(n_5119),
.A2(n_5312),
.B(n_5298),
.Y(n_6217)
);

NAND2xp5_ASAP7_75t_L g6218 ( 
.A(n_5264),
.B(n_5270),
.Y(n_6218)
);

NAND2xp5_ASAP7_75t_L g6219 ( 
.A(n_5270),
.B(n_5274),
.Y(n_6219)
);

INVxp67_ASAP7_75t_SL g6220 ( 
.A(n_4576),
.Y(n_6220)
);

AOI21xp5_ASAP7_75t_L g6221 ( 
.A1(n_5312),
.A2(n_5392),
.B(n_5432),
.Y(n_6221)
);

AOI21xp5_ASAP7_75t_L g6222 ( 
.A1(n_5392),
.A2(n_5432),
.B(n_5386),
.Y(n_6222)
);

AND3x1_ASAP7_75t_L g6223 ( 
.A(n_5402),
.B(n_5428),
.C(n_5464),
.Y(n_6223)
);

OAI22xp5_ASAP7_75t_SL g6224 ( 
.A1(n_5243),
.A2(n_4999),
.B1(n_5090),
.B2(n_4957),
.Y(n_6224)
);

BUFx3_ASAP7_75t_L g6225 ( 
.A(n_5461),
.Y(n_6225)
);

BUFx6f_ASAP7_75t_L g6226 ( 
.A(n_4977),
.Y(n_6226)
);

A2O1A1Ixp33_ASAP7_75t_L g6227 ( 
.A1(n_5067),
.A2(n_5085),
.B(n_5095),
.C(n_5088),
.Y(n_6227)
);

BUFx2_ASAP7_75t_L g6228 ( 
.A(n_4977),
.Y(n_6228)
);

NAND2xp5_ASAP7_75t_SL g6229 ( 
.A(n_5067),
.B(n_5085),
.Y(n_6229)
);

OAI22xp5_ASAP7_75t_L g6230 ( 
.A1(n_4533),
.A2(n_4539),
.B1(n_4547),
.B2(n_4537),
.Y(n_6230)
);

BUFx3_ASAP7_75t_L g6231 ( 
.A(n_5461),
.Y(n_6231)
);

OAI21xp33_ASAP7_75t_L g6232 ( 
.A1(n_5039),
.A2(n_5068),
.B(n_5046),
.Y(n_6232)
);

AOI21xp5_ASAP7_75t_L g6233 ( 
.A1(n_5386),
.A2(n_4808),
.B(n_4504),
.Y(n_6233)
);

AOI21xp5_ASAP7_75t_L g6234 ( 
.A1(n_5386),
.A2(n_4808),
.B(n_4504),
.Y(n_6234)
);

OAI22xp5_ASAP7_75t_L g6235 ( 
.A1(n_4539),
.A2(n_4550),
.B1(n_4553),
.B2(n_4547),
.Y(n_6235)
);

INVx4_ASAP7_75t_L g6236 ( 
.A(n_4484),
.Y(n_6236)
);

AND2x2_ASAP7_75t_L g6237 ( 
.A(n_4976),
.B(n_4774),
.Y(n_6237)
);

A2O1A1Ixp33_ASAP7_75t_L g6238 ( 
.A1(n_5088),
.A2(n_5095),
.B(n_5108),
.C(n_4975),
.Y(n_6238)
);

INVxp67_ASAP7_75t_SL g6239 ( 
.A(n_4644),
.Y(n_6239)
);

INVx4_ASAP7_75t_L g6240 ( 
.A(n_4489),
.Y(n_6240)
);

INVx4_ASAP7_75t_L g6241 ( 
.A(n_4489),
.Y(n_6241)
);

AO21x2_ASAP7_75t_L g6242 ( 
.A1(n_5468),
.A2(n_5396),
.B(n_5388),
.Y(n_6242)
);

CKINVDCx8_ASAP7_75t_R g6243 ( 
.A(n_4542),
.Y(n_6243)
);

INVx4_ASAP7_75t_L g6244 ( 
.A(n_4489),
.Y(n_6244)
);

INVxp67_ASAP7_75t_L g6245 ( 
.A(n_4654),
.Y(n_6245)
);

BUFx6f_ASAP7_75t_L g6246 ( 
.A(n_4977),
.Y(n_6246)
);

OR2x2_ASAP7_75t_L g6247 ( 
.A(n_4933),
.B(n_4941),
.Y(n_6247)
);

BUFx12f_ASAP7_75t_L g6248 ( 
.A(n_4857),
.Y(n_6248)
);

INVx8_ASAP7_75t_L g6249 ( 
.A(n_4512),
.Y(n_6249)
);

AOI22xp33_ASAP7_75t_L g6250 ( 
.A1(n_4929),
.A2(n_4960),
.B1(n_5089),
.B2(n_4847),
.Y(n_6250)
);

A2O1A1Ixp33_ASAP7_75t_L g6251 ( 
.A1(n_5095),
.A2(n_5108),
.B(n_5314),
.C(n_5406),
.Y(n_6251)
);

BUFx4f_ASAP7_75t_L g6252 ( 
.A(n_4489),
.Y(n_6252)
);

BUFx2_ASAP7_75t_L g6253 ( 
.A(n_4977),
.Y(n_6253)
);

INVx4_ASAP7_75t_L g6254 ( 
.A(n_4489),
.Y(n_6254)
);

NOR2x1_ASAP7_75t_L g6255 ( 
.A(n_5031),
.B(n_5032),
.Y(n_6255)
);

HB1xp67_ASAP7_75t_L g6256 ( 
.A(n_4585),
.Y(n_6256)
);

A2O1A1Ixp33_ASAP7_75t_L g6257 ( 
.A1(n_5108),
.A2(n_5314),
.B(n_4761),
.C(n_4615),
.Y(n_6257)
);

O2A1O1Ixp33_ASAP7_75t_L g6258 ( 
.A1(n_4550),
.A2(n_4553),
.B(n_4556),
.C(n_4554),
.Y(n_6258)
);

BUFx12f_ASAP7_75t_L g6259 ( 
.A(n_4906),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_SL g6260 ( 
.A(n_5108),
.B(n_5022),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_4557),
.Y(n_6261)
);

CKINVDCx16_ASAP7_75t_R g6262 ( 
.A(n_4957),
.Y(n_6262)
);

AOI21xp5_ASAP7_75t_L g6263 ( 
.A1(n_5386),
.A2(n_4808),
.B(n_4504),
.Y(n_6263)
);

AOI21xp33_ASAP7_75t_L g6264 ( 
.A1(n_5039),
.A2(n_5068),
.B(n_5046),
.Y(n_6264)
);

BUFx6f_ASAP7_75t_L g6265 ( 
.A(n_4977),
.Y(n_6265)
);

INVx1_ASAP7_75t_SL g6266 ( 
.A(n_4773),
.Y(n_6266)
);

NOR2xp33_ASAP7_75t_L g6267 ( 
.A(n_4554),
.B(n_4556),
.Y(n_6267)
);

CKINVDCx20_ASAP7_75t_R g6268 ( 
.A(n_5090),
.Y(n_6268)
);

NAND2x1_ASAP7_75t_L g6269 ( 
.A(n_4490),
.B(n_4926),
.Y(n_6269)
);

NAND3xp33_ASAP7_75t_L g6270 ( 
.A(n_5070),
.B(n_5087),
.C(n_5083),
.Y(n_6270)
);

CKINVDCx20_ASAP7_75t_R g6271 ( 
.A(n_5102),
.Y(n_6271)
);

AOI21x1_ASAP7_75t_L g6272 ( 
.A1(n_5126),
.A2(n_5260),
.B(n_4873),
.Y(n_6272)
);

BUFx2_ASAP7_75t_L g6273 ( 
.A(n_4774),
.Y(n_6273)
);

AOI21xp5_ASAP7_75t_L g6274 ( 
.A1(n_5386),
.A2(n_4808),
.B(n_4504),
.Y(n_6274)
);

AOI21xp5_ASAP7_75t_L g6275 ( 
.A1(n_5386),
.A2(n_4808),
.B(n_4504),
.Y(n_6275)
);

NAND2xp5_ASAP7_75t_SL g6276 ( 
.A(n_5022),
.B(n_5070),
.Y(n_6276)
);

AND2x2_ASAP7_75t_L g6277 ( 
.A(n_4774),
.B(n_4825),
.Y(n_6277)
);

INVx4_ASAP7_75t_L g6278 ( 
.A(n_4489),
.Y(n_6278)
);

INVx2_ASAP7_75t_L g6279 ( 
.A(n_4557),
.Y(n_6279)
);

NAND2xp33_ASAP7_75t_L g6280 ( 
.A(n_5213),
.B(n_4634),
.Y(n_6280)
);

OAI22xp5_ASAP7_75t_L g6281 ( 
.A1(n_4560),
.A2(n_4564),
.B1(n_4565),
.B2(n_4562),
.Y(n_6281)
);

NOR2x1p5_ASAP7_75t_SL g6282 ( 
.A(n_5426),
.B(n_5331),
.Y(n_6282)
);

AOI22x1_ASAP7_75t_L g6283 ( 
.A1(n_5459),
.A2(n_5452),
.B1(n_5248),
.B2(n_5234),
.Y(n_6283)
);

OAI21xp5_ASAP7_75t_L g6284 ( 
.A1(n_5083),
.A2(n_5104),
.B(n_5087),
.Y(n_6284)
);

AOI21x1_ASAP7_75t_L g6285 ( 
.A1(n_5126),
.A2(n_5260),
.B(n_4873),
.Y(n_6285)
);

INVx2_ASAP7_75t_L g6286 ( 
.A(n_4566),
.Y(n_6286)
);

BUFx2_ASAP7_75t_L g6287 ( 
.A(n_4825),
.Y(n_6287)
);

A2O1A1Ixp33_ASAP7_75t_L g6288 ( 
.A1(n_4761),
.A2(n_4615),
.B(n_5110),
.C(n_5104),
.Y(n_6288)
);

A2O1A1Ixp33_ASAP7_75t_L g6289 ( 
.A1(n_4761),
.A2(n_4615),
.B(n_5125),
.C(n_5110),
.Y(n_6289)
);

BUFx6f_ASAP7_75t_L g6290 ( 
.A(n_4489),
.Y(n_6290)
);

AOI21xp5_ASAP7_75t_L g6291 ( 
.A1(n_4410),
.A2(n_4669),
.B(n_4504),
.Y(n_6291)
);

AO22x1_ASAP7_75t_L g6292 ( 
.A1(n_5300),
.A2(n_5459),
.B1(n_5297),
.B2(n_5241),
.Y(n_6292)
);

INVx2_ASAP7_75t_L g6293 ( 
.A(n_4566),
.Y(n_6293)
);

AND2x4_ASAP7_75t_L g6294 ( 
.A(n_4605),
.B(n_4656),
.Y(n_6294)
);

OAI22xp5_ASAP7_75t_L g6295 ( 
.A1(n_4560),
.A2(n_4564),
.B1(n_4565),
.B2(n_4562),
.Y(n_6295)
);

INVx2_ASAP7_75t_L g6296 ( 
.A(n_4566),
.Y(n_6296)
);

OR2x2_ASAP7_75t_L g6297 ( 
.A(n_4933),
.B(n_4941),
.Y(n_6297)
);

OAI21xp5_ASAP7_75t_L g6298 ( 
.A1(n_5125),
.A2(n_5139),
.B(n_5127),
.Y(n_6298)
);

NAND2xp5_ASAP7_75t_L g6299 ( 
.A(n_5313),
.B(n_4847),
.Y(n_6299)
);

INVx1_ASAP7_75t_SL g6300 ( 
.A(n_5330),
.Y(n_6300)
);

AND2x2_ASAP7_75t_L g6301 ( 
.A(n_4414),
.B(n_4432),
.Y(n_6301)
);

AOI21xp5_ASAP7_75t_L g6302 ( 
.A1(n_4410),
.A2(n_4669),
.B(n_4504),
.Y(n_6302)
);

CKINVDCx6p67_ASAP7_75t_R g6303 ( 
.A(n_5064),
.Y(n_6303)
);

O2A1O1Ixp33_ASAP7_75t_L g6304 ( 
.A1(n_4567),
.A2(n_4569),
.B(n_4580),
.C(n_4579),
.Y(n_6304)
);

AOI21xp5_ASAP7_75t_L g6305 ( 
.A1(n_4410),
.A2(n_4757),
.B(n_4669),
.Y(n_6305)
);

AO21x2_ASAP7_75t_L g6306 ( 
.A1(n_5468),
.A2(n_5396),
.B(n_5388),
.Y(n_6306)
);

BUFx2_ASAP7_75t_L g6307 ( 
.A(n_4660),
.Y(n_6307)
);

A2O1A1Ixp33_ASAP7_75t_L g6308 ( 
.A1(n_5127),
.A2(n_5139),
.B(n_5228),
.C(n_5099),
.Y(n_6308)
);

AOI22xp33_ASAP7_75t_L g6309 ( 
.A1(n_5089),
.A2(n_5464),
.B1(n_4569),
.B2(n_4580),
.Y(n_6309)
);

AOI22xp33_ASAP7_75t_SL g6310 ( 
.A1(n_4926),
.A2(n_5243),
.B1(n_5451),
.B2(n_5143),
.Y(n_6310)
);

BUFx6f_ASAP7_75t_L g6311 ( 
.A(n_4489),
.Y(n_6311)
);

OR2x6_ASAP7_75t_L g6312 ( 
.A(n_5434),
.B(n_4410),
.Y(n_6312)
);

INVx4_ASAP7_75t_L g6313 ( 
.A(n_4506),
.Y(n_6313)
);

NAND2xp5_ASAP7_75t_L g6314 ( 
.A(n_4802),
.B(n_5176),
.Y(n_6314)
);

INVx2_ASAP7_75t_L g6315 ( 
.A(n_4575),
.Y(n_6315)
);

CKINVDCx5p33_ASAP7_75t_R g6316 ( 
.A(n_5304),
.Y(n_6316)
);

INVx2_ASAP7_75t_L g6317 ( 
.A(n_4575),
.Y(n_6317)
);

AOI21xp5_ASAP7_75t_L g6318 ( 
.A1(n_4410),
.A2(n_4757),
.B(n_4669),
.Y(n_6318)
);

BUFx2_ASAP7_75t_L g6319 ( 
.A(n_4661),
.Y(n_6319)
);

BUFx6f_ASAP7_75t_L g6320 ( 
.A(n_4506),
.Y(n_6320)
);

A2O1A1Ixp33_ASAP7_75t_L g6321 ( 
.A1(n_5228),
.A2(n_5099),
.B(n_5141),
.C(n_5103),
.Y(n_6321)
);

NAND2xp5_ASAP7_75t_SL g6322 ( 
.A(n_4829),
.B(n_4842),
.Y(n_6322)
);

O2A1O1Ixp33_ASAP7_75t_L g6323 ( 
.A1(n_4567),
.A2(n_4579),
.B(n_4593),
.C(n_4586),
.Y(n_6323)
);

A2O1A1Ixp33_ASAP7_75t_L g6324 ( 
.A1(n_5099),
.A2(n_5103),
.B(n_5141),
.C(n_5048),
.Y(n_6324)
);

NOR2xp33_ASAP7_75t_L g6325 ( 
.A(n_4586),
.B(n_4593),
.Y(n_6325)
);

BUFx2_ASAP7_75t_L g6326 ( 
.A(n_4661),
.Y(n_6326)
);

INVx1_ASAP7_75t_SL g6327 ( 
.A(n_5330),
.Y(n_6327)
);

OAI22xp5_ASAP7_75t_L g6328 ( 
.A1(n_4596),
.A2(n_4600),
.B1(n_4603),
.B2(n_4599),
.Y(n_6328)
);

NAND2xp5_ASAP7_75t_L g6329 ( 
.A(n_4802),
.B(n_5176),
.Y(n_6329)
);

NAND2x1p5_ASAP7_75t_L g6330 ( 
.A(n_4490),
.B(n_4542),
.Y(n_6330)
);

AOI22xp33_ASAP7_75t_L g6331 ( 
.A1(n_4596),
.A2(n_4600),
.B1(n_4607),
.B2(n_4603),
.Y(n_6331)
);

INVx2_ASAP7_75t_L g6332 ( 
.A(n_4581),
.Y(n_6332)
);

BUFx2_ASAP7_75t_L g6333 ( 
.A(n_4661),
.Y(n_6333)
);

INVx3_ASAP7_75t_L g6334 ( 
.A(n_4661),
.Y(n_6334)
);

INVx3_ASAP7_75t_L g6335 ( 
.A(n_4661),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_4802),
.B(n_5176),
.Y(n_6336)
);

BUFx2_ASAP7_75t_L g6337 ( 
.A(n_4663),
.Y(n_6337)
);

BUFx6f_ASAP7_75t_L g6338 ( 
.A(n_4506),
.Y(n_6338)
);

OAI22xp5_ASAP7_75t_L g6339 ( 
.A1(n_4599),
.A2(n_4608),
.B1(n_4611),
.B2(n_4607),
.Y(n_6339)
);

INVx3_ASAP7_75t_SL g6340 ( 
.A(n_5075),
.Y(n_6340)
);

BUFx6f_ASAP7_75t_L g6341 ( 
.A(n_4506),
.Y(n_6341)
);

HB1xp67_ASAP7_75t_L g6342 ( 
.A(n_4585),
.Y(n_6342)
);

AND2x2_ASAP7_75t_L g6343 ( 
.A(n_4414),
.B(n_4432),
.Y(n_6343)
);

BUFx3_ASAP7_75t_L g6344 ( 
.A(n_5461),
.Y(n_6344)
);

INVx2_ASAP7_75t_L g6345 ( 
.A(n_4581),
.Y(n_6345)
);

NAND2xp5_ASAP7_75t_SL g6346 ( 
.A(n_4829),
.B(n_4842),
.Y(n_6346)
);

NAND2xp5_ASAP7_75t_SL g6347 ( 
.A(n_4829),
.B(n_4842),
.Y(n_6347)
);

BUFx2_ASAP7_75t_L g6348 ( 
.A(n_4663),
.Y(n_6348)
);

AND2x2_ASAP7_75t_L g6349 ( 
.A(n_4414),
.B(n_4432),
.Y(n_6349)
);

INVx8_ASAP7_75t_L g6350 ( 
.A(n_4512),
.Y(n_6350)
);

NOR2x1_ASAP7_75t_L g6351 ( 
.A(n_5059),
.B(n_5061),
.Y(n_6351)
);

NAND2xp5_ASAP7_75t_SL g6352 ( 
.A(n_4829),
.B(n_4842),
.Y(n_6352)
);

AOI21xp5_ASAP7_75t_L g6353 ( 
.A1(n_4410),
.A2(n_4757),
.B(n_4669),
.Y(n_6353)
);

AOI21xp5_ASAP7_75t_L g6354 ( 
.A1(n_4669),
.A2(n_4757),
.B(n_5434),
.Y(n_6354)
);

O2A1O1Ixp33_ASAP7_75t_L g6355 ( 
.A1(n_4608),
.A2(n_4613),
.B(n_4619),
.C(n_4611),
.Y(n_6355)
);

HB1xp67_ASAP7_75t_L g6356 ( 
.A(n_4850),
.Y(n_6356)
);

INVx2_ASAP7_75t_L g6357 ( 
.A(n_4581),
.Y(n_6357)
);

BUFx6f_ASAP7_75t_L g6358 ( 
.A(n_4506),
.Y(n_6358)
);

INVx3_ASAP7_75t_L g6359 ( 
.A(n_4663),
.Y(n_6359)
);

O2A1O1Ixp33_ASAP7_75t_L g6360 ( 
.A1(n_4613),
.A2(n_4621),
.B(n_4626),
.C(n_4619),
.Y(n_6360)
);

CKINVDCx8_ASAP7_75t_R g6361 ( 
.A(n_4542),
.Y(n_6361)
);

AOI21xp5_ASAP7_75t_L g6362 ( 
.A1(n_4757),
.A2(n_5434),
.B(n_5399),
.Y(n_6362)
);

INVx2_ASAP7_75t_L g6363 ( 
.A(n_4581),
.Y(n_6363)
);

BUFx6f_ASAP7_75t_SL g6364 ( 
.A(n_4506),
.Y(n_6364)
);

AO32x2_ASAP7_75t_L g6365 ( 
.A1(n_4678),
.A2(n_4693),
.A3(n_4770),
.B1(n_4574),
.B2(n_4505),
.Y(n_6365)
);

O2A1O1Ixp33_ASAP7_75t_L g6366 ( 
.A1(n_4621),
.A2(n_4627),
.B(n_4630),
.C(n_4626),
.Y(n_6366)
);

AOI21xp5_ASAP7_75t_L g6367 ( 
.A1(n_4757),
.A2(n_5434),
.B(n_5399),
.Y(n_6367)
);

BUFx12f_ASAP7_75t_L g6368 ( 
.A(n_4906),
.Y(n_6368)
);

AND2x2_ASAP7_75t_L g6369 ( 
.A(n_4414),
.B(n_4432),
.Y(n_6369)
);

BUFx6f_ASAP7_75t_L g6370 ( 
.A(n_4506),
.Y(n_6370)
);

NOR2xp33_ASAP7_75t_L g6371 ( 
.A(n_4627),
.B(n_4630),
.Y(n_6371)
);

O2A1O1Ixp33_ASAP7_75t_L g6372 ( 
.A1(n_4635),
.A2(n_4646),
.B(n_4648),
.C(n_4642),
.Y(n_6372)
);

AND2x4_ASAP7_75t_L g6373 ( 
.A(n_4605),
.B(n_4656),
.Y(n_6373)
);

A2O1A1Ixp33_ASAP7_75t_SL g6374 ( 
.A1(n_4969),
.A2(n_4970),
.B(n_5431),
.C(n_5421),
.Y(n_6374)
);

CKINVDCx5p33_ASAP7_75t_R g6375 ( 
.A(n_4953),
.Y(n_6375)
);

AO31x2_ASAP7_75t_L g6376 ( 
.A1(n_5024),
.A2(n_5026),
.A3(n_5069),
.B(n_5061),
.Y(n_6376)
);

CKINVDCx16_ASAP7_75t_R g6377 ( 
.A(n_5102),
.Y(n_6377)
);

BUFx2_ASAP7_75t_L g6378 ( 
.A(n_4663),
.Y(n_6378)
);

BUFx4f_ASAP7_75t_L g6379 ( 
.A(n_4506),
.Y(n_6379)
);

NAND2xp5_ASAP7_75t_L g6380 ( 
.A(n_5084),
.B(n_5303),
.Y(n_6380)
);

INVxp67_ASAP7_75t_L g6381 ( 
.A(n_4698),
.Y(n_6381)
);

BUFx2_ASAP7_75t_L g6382 ( 
.A(n_4663),
.Y(n_6382)
);

INVx1_ASAP7_75t_SL g6383 ( 
.A(n_4763),
.Y(n_6383)
);

AND2x4_ASAP7_75t_L g6384 ( 
.A(n_4605),
.B(n_4656),
.Y(n_6384)
);

HB1xp67_ASAP7_75t_L g6385 ( 
.A(n_4850),
.Y(n_6385)
);

AOI221xp5_ASAP7_75t_L g6386 ( 
.A1(n_4635),
.A2(n_4642),
.B1(n_4650),
.B2(n_4648),
.C(n_4646),
.Y(n_6386)
);

AOI21xp5_ASAP7_75t_L g6387 ( 
.A1(n_5398),
.A2(n_5410),
.B(n_5407),
.Y(n_6387)
);

AOI22xp33_ASAP7_75t_L g6388 ( 
.A1(n_4650),
.A2(n_4652),
.B1(n_4653),
.B2(n_4651),
.Y(n_6388)
);

NOR2xp33_ASAP7_75t_L g6389 ( 
.A(n_4651),
.B(n_4652),
.Y(n_6389)
);

AOI21xp5_ASAP7_75t_L g6390 ( 
.A1(n_5398),
.A2(n_5410),
.B(n_5407),
.Y(n_6390)
);

AOI21xp5_ASAP7_75t_L g6391 ( 
.A1(n_5418),
.A2(n_5423),
.B(n_5419),
.Y(n_6391)
);

INVx2_ASAP7_75t_L g6392 ( 
.A(n_4595),
.Y(n_6392)
);

BUFx6f_ASAP7_75t_L g6393 ( 
.A(n_4527),
.Y(n_6393)
);

BUFx2_ASAP7_75t_L g6394 ( 
.A(n_4598),
.Y(n_6394)
);

AOI22xp5_ASAP7_75t_L g6395 ( 
.A1(n_4446),
.A2(n_5020),
.B1(n_4653),
.B2(n_4677),
.Y(n_6395)
);

O2A1O1Ixp33_ASAP7_75t_L g6396 ( 
.A1(n_4655),
.A2(n_4677),
.B(n_4680),
.C(n_4679),
.Y(n_6396)
);

INVx2_ASAP7_75t_L g6397 ( 
.A(n_4595),
.Y(n_6397)
);

NOR2xp33_ASAP7_75t_SL g6398 ( 
.A(n_5393),
.B(n_5458),
.Y(n_6398)
);

INVx8_ASAP7_75t_L g6399 ( 
.A(n_4512),
.Y(n_6399)
);

INVx2_ASAP7_75t_L g6400 ( 
.A(n_4595),
.Y(n_6400)
);

BUFx6f_ASAP7_75t_L g6401 ( 
.A(n_4527),
.Y(n_6401)
);

AOI21xp5_ASAP7_75t_L g6402 ( 
.A1(n_5418),
.A2(n_5423),
.B(n_5419),
.Y(n_6402)
);

HB1xp67_ASAP7_75t_L g6403 ( 
.A(n_4853),
.Y(n_6403)
);

NAND2xp5_ASAP7_75t_SL g6404 ( 
.A(n_4829),
.B(n_4842),
.Y(n_6404)
);

INVx2_ASAP7_75t_L g6405 ( 
.A(n_4595),
.Y(n_6405)
);

INVx2_ASAP7_75t_L g6406 ( 
.A(n_4614),
.Y(n_6406)
);

OAI22xp5_ASAP7_75t_L g6407 ( 
.A1(n_4655),
.A2(n_4679),
.B1(n_4681),
.B2(n_4680),
.Y(n_6407)
);

A2O1A1Ixp33_ASAP7_75t_L g6408 ( 
.A1(n_5103),
.A2(n_5141),
.B(n_5048),
.C(n_5077),
.Y(n_6408)
);

NAND2xp5_ASAP7_75t_L g6409 ( 
.A(n_5084),
.B(n_5303),
.Y(n_6409)
);

AOI22xp33_ASAP7_75t_L g6410 ( 
.A1(n_4681),
.A2(n_4688),
.B1(n_4710),
.B2(n_4687),
.Y(n_6410)
);

NOR2xp67_ASAP7_75t_SL g6411 ( 
.A(n_5297),
.B(n_4477),
.Y(n_6411)
);

NOR2xp33_ASAP7_75t_L g6412 ( 
.A(n_4687),
.B(n_4688),
.Y(n_6412)
);

BUFx3_ASAP7_75t_L g6413 ( 
.A(n_5467),
.Y(n_6413)
);

O2A1O1Ixp33_ASAP7_75t_L g6414 ( 
.A1(n_4708),
.A2(n_4710),
.B(n_4713),
.C(n_4712),
.Y(n_6414)
);

BUFx8_ASAP7_75t_SL g6415 ( 
.A(n_5239),
.Y(n_6415)
);

BUFx3_ASAP7_75t_L g6416 ( 
.A(n_5467),
.Y(n_6416)
);

INVx5_ASAP7_75t_L g6417 ( 
.A(n_4548),
.Y(n_6417)
);

A2O1A1Ixp33_ASAP7_75t_SL g6418 ( 
.A1(n_4969),
.A2(n_4970),
.B(n_5431),
.C(n_5421),
.Y(n_6418)
);

AOI21xp5_ASAP7_75t_L g6419 ( 
.A1(n_5425),
.A2(n_5430),
.B(n_5429),
.Y(n_6419)
);

INVx2_ASAP7_75t_L g6420 ( 
.A(n_4614),
.Y(n_6420)
);

NAND2xp5_ASAP7_75t_SL g6421 ( 
.A(n_4829),
.B(n_4842),
.Y(n_6421)
);

INVx2_ASAP7_75t_L g6422 ( 
.A(n_4614),
.Y(n_6422)
);

OAI22xp5_ASAP7_75t_L g6423 ( 
.A1(n_4708),
.A2(n_4712),
.B1(n_4715),
.B2(n_4713),
.Y(n_6423)
);

O2A1O1Ixp33_ASAP7_75t_L g6424 ( 
.A1(n_4715),
.A2(n_4721),
.B(n_4732),
.C(n_4725),
.Y(n_6424)
);

AOI21xp5_ASAP7_75t_L g6425 ( 
.A1(n_5425),
.A2(n_5430),
.B(n_5429),
.Y(n_6425)
);

AOI21xp5_ASAP7_75t_L g6426 ( 
.A1(n_5438),
.A2(n_5444),
.B(n_5443),
.Y(n_6426)
);

NAND2xp5_ASAP7_75t_L g6427 ( 
.A(n_5084),
.B(n_5306),
.Y(n_6427)
);

INVx3_ASAP7_75t_L g6428 ( 
.A(n_4686),
.Y(n_6428)
);

INVx3_ASAP7_75t_L g6429 ( 
.A(n_4686),
.Y(n_6429)
);

INVx2_ASAP7_75t_L g6430 ( 
.A(n_4614),
.Y(n_6430)
);

NAND2xp5_ASAP7_75t_SL g6431 ( 
.A(n_5066),
.B(n_5226),
.Y(n_6431)
);

BUFx6f_ASAP7_75t_L g6432 ( 
.A(n_4527),
.Y(n_6432)
);

INVx8_ASAP7_75t_L g6433 ( 
.A(n_4512),
.Y(n_6433)
);

CKINVDCx5p33_ASAP7_75t_R g6434 ( 
.A(n_4953),
.Y(n_6434)
);

AND2x2_ASAP7_75t_L g6435 ( 
.A(n_4414),
.B(n_4432),
.Y(n_6435)
);

OAI22xp5_ASAP7_75t_L g6436 ( 
.A1(n_4721),
.A2(n_4725),
.B1(n_4740),
.B2(n_4732),
.Y(n_6436)
);

NAND2xp5_ASAP7_75t_SL g6437 ( 
.A(n_5066),
.B(n_5226),
.Y(n_6437)
);

INVx2_ASAP7_75t_L g6438 ( 
.A(n_4617),
.Y(n_6438)
);

INVx4_ASAP7_75t_L g6439 ( 
.A(n_4527),
.Y(n_6439)
);

NAND2xp5_ASAP7_75t_L g6440 ( 
.A(n_5306),
.B(n_5307),
.Y(n_6440)
);

NOR2xp33_ASAP7_75t_L g6441 ( 
.A(n_4740),
.B(n_4742),
.Y(n_6441)
);

NAND2xp5_ASAP7_75t_L g6442 ( 
.A(n_5307),
.B(n_5309),
.Y(n_6442)
);

NAND2xp5_ASAP7_75t_SL g6443 ( 
.A(n_5066),
.B(n_5226),
.Y(n_6443)
);

OAI22xp5_ASAP7_75t_L g6444 ( 
.A1(n_4742),
.A2(n_4744),
.B1(n_4749),
.B2(n_4748),
.Y(n_6444)
);

AOI21x1_ASAP7_75t_L g6445 ( 
.A1(n_5438),
.A2(n_5444),
.B(n_5443),
.Y(n_6445)
);

CKINVDCx8_ASAP7_75t_R g6446 ( 
.A(n_4542),
.Y(n_6446)
);

INVx2_ASAP7_75t_L g6447 ( 
.A(n_4617),
.Y(n_6447)
);

HB1xp67_ASAP7_75t_L g6448 ( 
.A(n_4853),
.Y(n_6448)
);

AO22x1_ASAP7_75t_L g6449 ( 
.A1(n_5300),
.A2(n_5241),
.B1(n_5467),
.B2(n_5096),
.Y(n_6449)
);

OR2x6_ASAP7_75t_L g6450 ( 
.A(n_4382),
.B(n_4399),
.Y(n_6450)
);

INVxp67_ASAP7_75t_SL g6451 ( 
.A(n_4644),
.Y(n_6451)
);

AOI21xp5_ASAP7_75t_L g6452 ( 
.A1(n_5447),
.A2(n_5460),
.B(n_5455),
.Y(n_6452)
);

INVx4_ASAP7_75t_L g6453 ( 
.A(n_4527),
.Y(n_6453)
);

INVx2_ASAP7_75t_L g6454 ( 
.A(n_4617),
.Y(n_6454)
);

BUFx6f_ASAP7_75t_L g6455 ( 
.A(n_4527),
.Y(n_6455)
);

NOR2xp33_ASAP7_75t_L g6456 ( 
.A(n_4744),
.B(n_4748),
.Y(n_6456)
);

NOR2xp33_ASAP7_75t_L g6457 ( 
.A(n_4749),
.B(n_4751),
.Y(n_6457)
);

OR2x6_ASAP7_75t_L g6458 ( 
.A(n_4382),
.B(n_4399),
.Y(n_6458)
);

AND2x4_ASAP7_75t_L g6459 ( 
.A(n_4686),
.B(n_4711),
.Y(n_6459)
);

OAI21x1_ASAP7_75t_L g6460 ( 
.A1(n_4886),
.A2(n_5151),
.B(n_5134),
.Y(n_6460)
);

BUFx8_ASAP7_75t_L g6461 ( 
.A(n_4457),
.Y(n_6461)
);

O2A1O1Ixp5_ASAP7_75t_SL g6462 ( 
.A1(n_5024),
.A2(n_5026),
.B(n_5077),
.C(n_5069),
.Y(n_6462)
);

NOR2xp33_ASAP7_75t_L g6463 ( 
.A(n_4751),
.B(n_4755),
.Y(n_6463)
);

INVx5_ASAP7_75t_L g6464 ( 
.A(n_4548),
.Y(n_6464)
);

NAND2xp5_ASAP7_75t_L g6465 ( 
.A(n_5309),
.B(n_5131),
.Y(n_6465)
);

HB1xp67_ASAP7_75t_L g6466 ( 
.A(n_4698),
.Y(n_6466)
);

INVx2_ASAP7_75t_L g6467 ( 
.A(n_4617),
.Y(n_6467)
);

INVx5_ASAP7_75t_L g6468 ( 
.A(n_4548),
.Y(n_6468)
);

NAND2xp5_ASAP7_75t_L g6469 ( 
.A(n_5131),
.B(n_5132),
.Y(n_6469)
);

NAND2xp5_ASAP7_75t_L g6470 ( 
.A(n_5131),
.B(n_5132),
.Y(n_6470)
);

INVxp67_ASAP7_75t_L g6471 ( 
.A(n_4719),
.Y(n_6471)
);

NAND2xp5_ASAP7_75t_L g6472 ( 
.A(n_5132),
.B(n_5133),
.Y(n_6472)
);

AOI22xp33_ASAP7_75t_L g6473 ( 
.A1(n_4755),
.A2(n_4775),
.B1(n_4782),
.B2(n_4766),
.Y(n_6473)
);

NAND2xp5_ASAP7_75t_L g6474 ( 
.A(n_5133),
.B(n_5135),
.Y(n_6474)
);

HB1xp67_ASAP7_75t_L g6475 ( 
.A(n_4719),
.Y(n_6475)
);

BUFx6f_ASAP7_75t_L g6476 ( 
.A(n_4527),
.Y(n_6476)
);

AND2x4_ASAP7_75t_L g6477 ( 
.A(n_4711),
.B(n_4731),
.Y(n_6477)
);

AOI21xp5_ASAP7_75t_L g6478 ( 
.A1(n_5447),
.A2(n_5460),
.B(n_5455),
.Y(n_6478)
);

AND2x2_ASAP7_75t_SL g6479 ( 
.A(n_5241),
.B(n_5226),
.Y(n_6479)
);

OAI22xp33_ASAP7_75t_L g6480 ( 
.A1(n_4766),
.A2(n_4775),
.B1(n_4782),
.B2(n_4772),
.Y(n_6480)
);

BUFx4f_ASAP7_75t_L g6481 ( 
.A(n_4546),
.Y(n_6481)
);

NAND2xp5_ASAP7_75t_L g6482 ( 
.A(n_5133),
.B(n_5135),
.Y(n_6482)
);

HB1xp67_ASAP7_75t_L g6483 ( 
.A(n_4728),
.Y(n_6483)
);

OAI22xp5_ASAP7_75t_L g6484 ( 
.A1(n_4772),
.A2(n_4784),
.B1(n_4798),
.B2(n_4795),
.Y(n_6484)
);

AOI22xp5_ASAP7_75t_L g6485 ( 
.A1(n_5020),
.A2(n_4784),
.B1(n_4798),
.B2(n_4795),
.Y(n_6485)
);

NOR2xp67_ASAP7_75t_SL g6486 ( 
.A(n_4477),
.B(n_4996),
.Y(n_6486)
);

NAND2xp5_ASAP7_75t_SL g6487 ( 
.A(n_5066),
.B(n_5226),
.Y(n_6487)
);

NAND2xp5_ASAP7_75t_SL g6488 ( 
.A(n_5066),
.B(n_5226),
.Y(n_6488)
);

OAI22xp5_ASAP7_75t_L g6489 ( 
.A1(n_4806),
.A2(n_4809),
.B1(n_4815),
.B2(n_4812),
.Y(n_6489)
);

BUFx2_ASAP7_75t_L g6490 ( 
.A(n_4598),
.Y(n_6490)
);

NAND2x1p5_ASAP7_75t_L g6491 ( 
.A(n_4542),
.B(n_4588),
.Y(n_6491)
);

AOI21xp5_ASAP7_75t_L g6492 ( 
.A1(n_5465),
.A2(n_5151),
.B(n_5134),
.Y(n_6492)
);

NOR2xp33_ASAP7_75t_L g6493 ( 
.A(n_4806),
.B(n_4809),
.Y(n_6493)
);

A2O1A1Ixp33_ASAP7_75t_L g6494 ( 
.A1(n_5048),
.A2(n_5093),
.B(n_5107),
.C(n_5091),
.Y(n_6494)
);

INVx1_ASAP7_75t_SL g6495 ( 
.A(n_4763),
.Y(n_6495)
);

OR2x6_ASAP7_75t_L g6496 ( 
.A(n_5134),
.B(n_5151),
.Y(n_6496)
);

NAND2xp5_ASAP7_75t_L g6497 ( 
.A(n_5135),
.B(n_5140),
.Y(n_6497)
);

AOI222xp33_ASAP7_75t_L g6498 ( 
.A1(n_4812),
.A2(n_4845),
.B1(n_4831),
.B2(n_4851),
.C1(n_4835),
.C2(n_4815),
.Y(n_6498)
);

INVx4_ASAP7_75t_L g6499 ( 
.A(n_4546),
.Y(n_6499)
);

AOI21xp5_ASAP7_75t_L g6500 ( 
.A1(n_5465),
.A2(n_5151),
.B(n_5134),
.Y(n_6500)
);

OAI22x1_ASAP7_75t_L g6501 ( 
.A1(n_5091),
.A2(n_5093),
.B1(n_5107),
.B2(n_5352),
.Y(n_6501)
);

BUFx2_ASAP7_75t_L g6502 ( 
.A(n_4598),
.Y(n_6502)
);

BUFx2_ASAP7_75t_L g6503 ( 
.A(n_4598),
.Y(n_6503)
);

INVx4_ASAP7_75t_L g6504 ( 
.A(n_4546),
.Y(n_6504)
);

OAI22xp5_ASAP7_75t_L g6505 ( 
.A1(n_4831),
.A2(n_4835),
.B1(n_4851),
.B2(n_4845),
.Y(n_6505)
);

BUFx3_ASAP7_75t_L g6506 ( 
.A(n_5467),
.Y(n_6506)
);

A2O1A1Ixp33_ASAP7_75t_L g6507 ( 
.A1(n_5324),
.A2(n_4606),
.B(n_4741),
.C(n_4583),
.Y(n_6507)
);

CKINVDCx20_ASAP7_75t_R g6508 ( 
.A(n_5239),
.Y(n_6508)
);

O2A1O1Ixp33_ASAP7_75t_L g6509 ( 
.A1(n_4862),
.A2(n_4867),
.B(n_4874),
.C(n_4871),
.Y(n_6509)
);

OAI22xp5_ASAP7_75t_L g6510 ( 
.A1(n_4862),
.A2(n_4867),
.B1(n_4874),
.B2(n_4871),
.Y(n_6510)
);

AO32x2_ASAP7_75t_L g6511 ( 
.A1(n_4505),
.A2(n_4485),
.A3(n_4441),
.B1(n_4433),
.B2(n_4834),
.Y(n_6511)
);

BUFx2_ASAP7_75t_L g6512 ( 
.A(n_4598),
.Y(n_6512)
);

INVx2_ASAP7_75t_L g6513 ( 
.A(n_4641),
.Y(n_6513)
);

O2A1O1Ixp33_ASAP7_75t_L g6514 ( 
.A1(n_4875),
.A2(n_4876),
.B(n_4879),
.C(n_4878),
.Y(n_6514)
);

INVxp67_ASAP7_75t_L g6515 ( 
.A(n_4728),
.Y(n_6515)
);

A2O1A1Ixp33_ASAP7_75t_L g6516 ( 
.A1(n_5324),
.A2(n_4606),
.B(n_4741),
.C(n_4583),
.Y(n_6516)
);

BUFx2_ASAP7_75t_L g6517 ( 
.A(n_4598),
.Y(n_6517)
);

AND3x2_ASAP7_75t_L g6518 ( 
.A(n_4969),
.B(n_4970),
.C(n_5286),
.Y(n_6518)
);

BUFx2_ASAP7_75t_L g6519 ( 
.A(n_4598),
.Y(n_6519)
);

A2O1A1Ixp33_ASAP7_75t_L g6520 ( 
.A1(n_4583),
.A2(n_4741),
.B(n_4860),
.C(n_4606),
.Y(n_6520)
);

INVx2_ASAP7_75t_L g6521 ( 
.A(n_4641),
.Y(n_6521)
);

OAI21x1_ASAP7_75t_L g6522 ( 
.A1(n_4886),
.A2(n_5151),
.B(n_5134),
.Y(n_6522)
);

A2O1A1Ixp33_ASAP7_75t_L g6523 ( 
.A1(n_4583),
.A2(n_4741),
.B(n_4860),
.C(n_4606),
.Y(n_6523)
);

INVx2_ASAP7_75t_L g6524 ( 
.A(n_4641),
.Y(n_6524)
);

NOR2xp33_ASAP7_75t_L g6525 ( 
.A(n_4875),
.B(n_4876),
.Y(n_6525)
);

NAND2xp5_ASAP7_75t_L g6526 ( 
.A(n_5153),
.B(n_4793),
.Y(n_6526)
);

INVx1_ASAP7_75t_L g6527 ( 
.A(n_4756),
.Y(n_6527)
);

NAND2xp5_ASAP7_75t_L g6528 ( 
.A(n_4793),
.B(n_4817),
.Y(n_6528)
);

CKINVDCx11_ASAP7_75t_R g6529 ( 
.A(n_5281),
.Y(n_6529)
);

INVx1_ASAP7_75t_SL g6530 ( 
.A(n_4763),
.Y(n_6530)
);

OAI221xp5_ASAP7_75t_L g6531 ( 
.A1(n_4878),
.A2(n_4881),
.B1(n_4884),
.B2(n_4883),
.C(n_4879),
.Y(n_6531)
);

HB1xp67_ASAP7_75t_L g6532 ( 
.A(n_4735),
.Y(n_6532)
);

NAND2xp5_ASAP7_75t_SL g6533 ( 
.A(n_5066),
.B(n_5267),
.Y(n_6533)
);

INVx1_ASAP7_75t_L g6534 ( 
.A(n_4756),
.Y(n_6534)
);

AOI21xp5_ASAP7_75t_L g6535 ( 
.A1(n_5240),
.A2(n_5401),
.B(n_5334),
.Y(n_6535)
);

AOI21xp5_ASAP7_75t_L g6536 ( 
.A1(n_5240),
.A2(n_5401),
.B(n_5334),
.Y(n_6536)
);

NAND2xp5_ASAP7_75t_L g6537 ( 
.A(n_4793),
.B(n_4817),
.Y(n_6537)
);

BUFx12f_ASAP7_75t_L g6538 ( 
.A(n_4938),
.Y(n_6538)
);

OR2x6_ASAP7_75t_L g6539 ( 
.A(n_5240),
.B(n_5401),
.Y(n_6539)
);

NOR2xp33_ASAP7_75t_L g6540 ( 
.A(n_4881),
.B(n_4883),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_4759),
.Y(n_6541)
);

INVx2_ASAP7_75t_L g6542 ( 
.A(n_4641),
.Y(n_6542)
);

BUFx2_ASAP7_75t_L g6543 ( 
.A(n_4598),
.Y(n_6543)
);

OR2x6_ASAP7_75t_L g6544 ( 
.A(n_5240),
.B(n_5401),
.Y(n_6544)
);

INVx1_ASAP7_75t_L g6545 ( 
.A(n_4778),
.Y(n_6545)
);

INVx2_ASAP7_75t_L g6546 ( 
.A(n_4659),
.Y(n_6546)
);

BUFx8_ASAP7_75t_SL g6547 ( 
.A(n_5281),
.Y(n_6547)
);

INVx3_ASAP7_75t_L g6548 ( 
.A(n_4731),
.Y(n_6548)
);

CKINVDCx5p33_ASAP7_75t_R g6549 ( 
.A(n_5019),
.Y(n_6549)
);

AOI21xp5_ASAP7_75t_L g6550 ( 
.A1(n_5240),
.A2(n_5401),
.B(n_5334),
.Y(n_6550)
);

AOI22xp33_ASAP7_75t_L g6551 ( 
.A1(n_4884),
.A2(n_4894),
.B1(n_4899),
.B2(n_4889),
.Y(n_6551)
);

NOR2xp33_ASAP7_75t_L g6552 ( 
.A(n_4889),
.B(n_4894),
.Y(n_6552)
);

O2A1O1Ixp33_ASAP7_75t_L g6553 ( 
.A1(n_4899),
.A2(n_4909),
.B(n_4924),
.C(n_4910),
.Y(n_6553)
);

OAI22xp33_ASAP7_75t_L g6554 ( 
.A1(n_4909),
.A2(n_4924),
.B1(n_4925),
.B2(n_4910),
.Y(n_6554)
);

AOI21xp5_ASAP7_75t_L g6555 ( 
.A1(n_5331),
.A2(n_5385),
.B(n_5335),
.Y(n_6555)
);

NOR2xp33_ASAP7_75t_SL g6556 ( 
.A(n_5681),
.B(n_4542),
.Y(n_6556)
);

HB1xp67_ASAP7_75t_L g6557 ( 
.A(n_5924),
.Y(n_6557)
);

INVx4_ASAP7_75t_L g6558 ( 
.A(n_5528),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_6511),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6511),
.Y(n_6560)
);

AOI22xp5_ASAP7_75t_L g6561 ( 
.A1(n_5863),
.A2(n_5092),
.B1(n_5157),
.B2(n_4913),
.Y(n_6561)
);

INVx2_ASAP7_75t_L g6562 ( 
.A(n_6511),
.Y(n_6562)
);

INVx2_ASAP7_75t_L g6563 ( 
.A(n_6511),
.Y(n_6563)
);

AOI22xp33_ASAP7_75t_L g6564 ( 
.A1(n_5485),
.A2(n_5300),
.B1(n_4930),
.B2(n_4931),
.Y(n_6564)
);

OR2x6_ASAP7_75t_L g6565 ( 
.A(n_5960),
.B(n_6035),
.Y(n_6565)
);

INVx3_ASAP7_75t_L g6566 ( 
.A(n_5604),
.Y(n_6566)
);

INVx2_ASAP7_75t_L g6567 ( 
.A(n_6511),
.Y(n_6567)
);

NOR2xp33_ASAP7_75t_SL g6568 ( 
.A(n_5681),
.B(n_4588),
.Y(n_6568)
);

INVx1_ASAP7_75t_L g6569 ( 
.A(n_6511),
.Y(n_6569)
);

OR2x6_ASAP7_75t_L g6570 ( 
.A(n_5960),
.B(n_5426),
.Y(n_6570)
);

INVx2_ASAP7_75t_L g6571 ( 
.A(n_6511),
.Y(n_6571)
);

INVx1_ASAP7_75t_L g6572 ( 
.A(n_6511),
.Y(n_6572)
);

INVxp67_ASAP7_75t_SL g6573 ( 
.A(n_5924),
.Y(n_6573)
);

AOI21x1_ASAP7_75t_L g6574 ( 
.A1(n_5874),
.A2(n_4801),
.B(n_4800),
.Y(n_6574)
);

INVx5_ASAP7_75t_L g6575 ( 
.A(n_5559),
.Y(n_6575)
);

OR2x6_ASAP7_75t_L g6576 ( 
.A(n_5960),
.B(n_5426),
.Y(n_6576)
);

AND2x2_ASAP7_75t_L g6577 ( 
.A(n_5765),
.B(n_4696),
.Y(n_6577)
);

INVx1_ASAP7_75t_L g6578 ( 
.A(n_5472),
.Y(n_6578)
);

INVx2_ASAP7_75t_L g6579 ( 
.A(n_5470),
.Y(n_6579)
);

BUFx2_ASAP7_75t_L g6580 ( 
.A(n_6190),
.Y(n_6580)
);

INVx2_ASAP7_75t_SL g6581 ( 
.A(n_5604),
.Y(n_6581)
);

INVx2_ASAP7_75t_L g6582 ( 
.A(n_5470),
.Y(n_6582)
);

BUFx2_ASAP7_75t_L g6583 ( 
.A(n_6190),
.Y(n_6583)
);

INVx1_ASAP7_75t_L g6584 ( 
.A(n_5472),
.Y(n_6584)
);

NAND2xp5_ASAP7_75t_L g6585 ( 
.A(n_5900),
.B(n_5111),
.Y(n_6585)
);

CKINVDCx11_ASAP7_75t_R g6586 ( 
.A(n_5538),
.Y(n_6586)
);

INVx1_ASAP7_75t_SL g6587 ( 
.A(n_5829),
.Y(n_6587)
);

OAI22xp5_ASAP7_75t_L g6588 ( 
.A1(n_5901),
.A2(n_4930),
.B1(n_4931),
.B2(n_4925),
.Y(n_6588)
);

INVx1_ASAP7_75t_L g6589 ( 
.A(n_5480),
.Y(n_6589)
);

INVxp67_ASAP7_75t_L g6590 ( 
.A(n_5965),
.Y(n_6590)
);

BUFx6f_ASAP7_75t_L g6591 ( 
.A(n_5559),
.Y(n_6591)
);

BUFx12f_ASAP7_75t_L g6592 ( 
.A(n_5878),
.Y(n_6592)
);

BUFx2_ASAP7_75t_L g6593 ( 
.A(n_6190),
.Y(n_6593)
);

INVx1_ASAP7_75t_L g6594 ( 
.A(n_5480),
.Y(n_6594)
);

INVx2_ASAP7_75t_SL g6595 ( 
.A(n_5604),
.Y(n_6595)
);

NAND2xp5_ASAP7_75t_SL g6596 ( 
.A(n_6200),
.B(n_5143),
.Y(n_6596)
);

INVx1_ASAP7_75t_SL g6597 ( 
.A(n_5829),
.Y(n_6597)
);

INVx2_ASAP7_75t_L g6598 ( 
.A(n_5470),
.Y(n_6598)
);

OR2x2_ASAP7_75t_L g6599 ( 
.A(n_6078),
.B(n_4933),
.Y(n_6599)
);

NOR2xp67_ASAP7_75t_L g6600 ( 
.A(n_6417),
.B(n_4747),
.Y(n_6600)
);

INVx3_ASAP7_75t_L g6601 ( 
.A(n_5604),
.Y(n_6601)
);

INVx3_ASAP7_75t_L g6602 ( 
.A(n_5604),
.Y(n_6602)
);

CKINVDCx20_ASAP7_75t_R g6603 ( 
.A(n_6018),
.Y(n_6603)
);

BUFx6f_ASAP7_75t_L g6604 ( 
.A(n_5559),
.Y(n_6604)
);

BUFx12f_ASAP7_75t_L g6605 ( 
.A(n_5894),
.Y(n_6605)
);

CKINVDCx5p33_ASAP7_75t_R g6606 ( 
.A(n_6018),
.Y(n_6606)
);

AOI22xp5_ASAP7_75t_L g6607 ( 
.A1(n_5863),
.A2(n_5157),
.B1(n_4913),
.B2(n_4951),
.Y(n_6607)
);

AND2x2_ASAP7_75t_L g6608 ( 
.A(n_5765),
.B(n_4696),
.Y(n_6608)
);

NAND2xp5_ASAP7_75t_L g6609 ( 
.A(n_5900),
.B(n_4800),
.Y(n_6609)
);

CKINVDCx11_ASAP7_75t_R g6610 ( 
.A(n_5538),
.Y(n_6610)
);

AOI21xp33_ASAP7_75t_L g6611 ( 
.A1(n_5898),
.A2(n_5911),
.B(n_5874),
.Y(n_6611)
);

HB1xp67_ASAP7_75t_L g6612 ( 
.A(n_5981),
.Y(n_6612)
);

INVx1_ASAP7_75t_L g6613 ( 
.A(n_5489),
.Y(n_6613)
);

BUFx6f_ASAP7_75t_L g6614 ( 
.A(n_5559),
.Y(n_6614)
);

OAI22xp33_ASAP7_75t_L g6615 ( 
.A1(n_5921),
.A2(n_4459),
.B1(n_5451),
.B2(n_4936),
.Y(n_6615)
);

BUFx6f_ASAP7_75t_L g6616 ( 
.A(n_5559),
.Y(n_6616)
);

INVx1_ASAP7_75t_SL g6617 ( 
.A(n_5829),
.Y(n_6617)
);

INVx1_ASAP7_75t_L g6618 ( 
.A(n_5489),
.Y(n_6618)
);

BUFx6f_ASAP7_75t_L g6619 ( 
.A(n_5559),
.Y(n_6619)
);

INVx2_ASAP7_75t_L g6620 ( 
.A(n_5477),
.Y(n_6620)
);

INVx1_ASAP7_75t_L g6621 ( 
.A(n_5498),
.Y(n_6621)
);

INVx1_ASAP7_75t_L g6622 ( 
.A(n_5498),
.Y(n_6622)
);

INVx1_ASAP7_75t_L g6623 ( 
.A(n_5510),
.Y(n_6623)
);

INVx3_ASAP7_75t_L g6624 ( 
.A(n_5611),
.Y(n_6624)
);

NAND2x1p5_ASAP7_75t_L g6625 ( 
.A(n_5471),
.B(n_4588),
.Y(n_6625)
);

OR2x6_ASAP7_75t_L g6626 ( 
.A(n_5960),
.B(n_5267),
.Y(n_6626)
);

NAND2xp5_ASAP7_75t_SL g6627 ( 
.A(n_6200),
.B(n_5143),
.Y(n_6627)
);

BUFx3_ASAP7_75t_L g6628 ( 
.A(n_5619),
.Y(n_6628)
);

NOR2xp33_ASAP7_75t_L g6629 ( 
.A(n_5795),
.B(n_5415),
.Y(n_6629)
);

NAND2xp5_ASAP7_75t_L g6630 ( 
.A(n_5906),
.B(n_5111),
.Y(n_6630)
);

NAND2xp5_ASAP7_75t_L g6631 ( 
.A(n_5906),
.B(n_5116),
.Y(n_6631)
);

INVx1_ASAP7_75t_SL g6632 ( 
.A(n_5832),
.Y(n_6632)
);

INVx1_ASAP7_75t_L g6633 ( 
.A(n_5510),
.Y(n_6633)
);

NAND2xp5_ASAP7_75t_L g6634 ( 
.A(n_5524),
.B(n_5116),
.Y(n_6634)
);

BUFx6f_ASAP7_75t_L g6635 ( 
.A(n_5559),
.Y(n_6635)
);

INVx2_ASAP7_75t_SL g6636 ( 
.A(n_5611),
.Y(n_6636)
);

AOI22xp33_ASAP7_75t_L g6637 ( 
.A1(n_5485),
.A2(n_5870),
.B1(n_5653),
.B2(n_5665),
.Y(n_6637)
);

INVx1_ASAP7_75t_SL g6638 ( 
.A(n_5832),
.Y(n_6638)
);

OAI21x1_ASAP7_75t_L g6639 ( 
.A1(n_6029),
.A2(n_4696),
.B(n_4800),
.Y(n_6639)
);

BUFx6f_ASAP7_75t_L g6640 ( 
.A(n_5559),
.Y(n_6640)
);

INVx2_ASAP7_75t_L g6641 ( 
.A(n_5477),
.Y(n_6641)
);

INVx1_ASAP7_75t_SL g6642 ( 
.A(n_5832),
.Y(n_6642)
);

INVx2_ASAP7_75t_L g6643 ( 
.A(n_5477),
.Y(n_6643)
);

BUFx6f_ASAP7_75t_L g6644 ( 
.A(n_5568),
.Y(n_6644)
);

BUFx6f_ASAP7_75t_L g6645 ( 
.A(n_5568),
.Y(n_6645)
);

INVx2_ASAP7_75t_L g6646 ( 
.A(n_5482),
.Y(n_6646)
);

INVx2_ASAP7_75t_L g6647 ( 
.A(n_5482),
.Y(n_6647)
);

NAND2xp5_ASAP7_75t_L g6648 ( 
.A(n_5524),
.B(n_4735),
.Y(n_6648)
);

CKINVDCx11_ASAP7_75t_R g6649 ( 
.A(n_5547),
.Y(n_6649)
);

INVx1_ASAP7_75t_L g6650 ( 
.A(n_5517),
.Y(n_6650)
);

INVx5_ASAP7_75t_L g6651 ( 
.A(n_5568),
.Y(n_6651)
);

BUFx6f_ASAP7_75t_L g6652 ( 
.A(n_5568),
.Y(n_6652)
);

INVx5_ASAP7_75t_L g6653 ( 
.A(n_5568),
.Y(n_6653)
);

AND2x2_ASAP7_75t_L g6654 ( 
.A(n_5765),
.B(n_4696),
.Y(n_6654)
);

AND2x6_ASAP7_75t_L g6655 ( 
.A(n_6083),
.B(n_4442),
.Y(n_6655)
);

CKINVDCx20_ASAP7_75t_R g6656 ( 
.A(n_5547),
.Y(n_6656)
);

NAND2xp5_ASAP7_75t_L g6657 ( 
.A(n_6033),
.B(n_4982),
.Y(n_6657)
);

AOI22xp33_ASAP7_75t_L g6658 ( 
.A1(n_5870),
.A2(n_5300),
.B1(n_4936),
.B2(n_4940),
.Y(n_6658)
);

AOI21xp5_ASAP7_75t_L g6659 ( 
.A1(n_5493),
.A2(n_5385),
.B(n_5389),
.Y(n_6659)
);

OAI22xp5_ASAP7_75t_L g6660 ( 
.A1(n_5901),
.A2(n_4940),
.B1(n_4959),
.B2(n_4934),
.Y(n_6660)
);

NAND2xp5_ASAP7_75t_L g6661 ( 
.A(n_5576),
.B(n_4800),
.Y(n_6661)
);

BUFx3_ASAP7_75t_L g6662 ( 
.A(n_5619),
.Y(n_6662)
);

BUFx6f_ASAP7_75t_L g6663 ( 
.A(n_5568),
.Y(n_6663)
);

INVx1_ASAP7_75t_L g6664 ( 
.A(n_5517),
.Y(n_6664)
);

OR2x6_ASAP7_75t_SL g6665 ( 
.A(n_6111),
.B(n_5219),
.Y(n_6665)
);

OR2x6_ASAP7_75t_L g6666 ( 
.A(n_5960),
.B(n_5267),
.Y(n_6666)
);

BUFx2_ASAP7_75t_L g6667 ( 
.A(n_6190),
.Y(n_6667)
);

OR2x6_ASAP7_75t_L g6668 ( 
.A(n_6035),
.B(n_6249),
.Y(n_6668)
);

BUFx2_ASAP7_75t_L g6669 ( 
.A(n_6190),
.Y(n_6669)
);

HB1xp67_ASAP7_75t_L g6670 ( 
.A(n_5981),
.Y(n_6670)
);

INVx1_ASAP7_75t_L g6671 ( 
.A(n_5532),
.Y(n_6671)
);

AOI21xp5_ASAP7_75t_L g6672 ( 
.A1(n_5493),
.A2(n_5390),
.B(n_5389),
.Y(n_6672)
);

BUFx6f_ASAP7_75t_L g6673 ( 
.A(n_5568),
.Y(n_6673)
);

INVx2_ASAP7_75t_L g6674 ( 
.A(n_5482),
.Y(n_6674)
);

NAND2xp5_ASAP7_75t_L g6675 ( 
.A(n_5576),
.B(n_4801),
.Y(n_6675)
);

AND2x2_ASAP7_75t_L g6676 ( 
.A(n_5765),
.B(n_4696),
.Y(n_6676)
);

AOI22xp5_ASAP7_75t_L g6677 ( 
.A1(n_5868),
.A2(n_4914),
.B1(n_4971),
.B2(n_4951),
.Y(n_6677)
);

OAI22xp5_ASAP7_75t_L g6678 ( 
.A1(n_5921),
.A2(n_4959),
.B1(n_4961),
.B2(n_4934),
.Y(n_6678)
);

CKINVDCx5p33_ASAP7_75t_R g6679 ( 
.A(n_5860),
.Y(n_6679)
);

AOI22xp33_ASAP7_75t_L g6680 ( 
.A1(n_5653),
.A2(n_5300),
.B1(n_4968),
.B2(n_4978),
.Y(n_6680)
);

CKINVDCx8_ASAP7_75t_R g6681 ( 
.A(n_5509),
.Y(n_6681)
);

NAND2x1p5_ASAP7_75t_L g6682 ( 
.A(n_5471),
.B(n_4588),
.Y(n_6682)
);

INVx1_ASAP7_75t_L g6683 ( 
.A(n_5532),
.Y(n_6683)
);

INVx1_ASAP7_75t_SL g6684 ( 
.A(n_6518),
.Y(n_6684)
);

AND2x2_ASAP7_75t_L g6685 ( 
.A(n_5765),
.B(n_4692),
.Y(n_6685)
);

INVx1_ASAP7_75t_L g6686 ( 
.A(n_5483),
.Y(n_6686)
);

NOR2xp33_ASAP7_75t_L g6687 ( 
.A(n_5795),
.B(n_5415),
.Y(n_6687)
);

INVx2_ASAP7_75t_SL g6688 ( 
.A(n_5611),
.Y(n_6688)
);

AOI21xp5_ASAP7_75t_L g6689 ( 
.A1(n_5494),
.A2(n_5390),
.B(n_5389),
.Y(n_6689)
);

CKINVDCx6p67_ASAP7_75t_R g6690 ( 
.A(n_6205),
.Y(n_6690)
);

INVx2_ASAP7_75t_SL g6691 ( 
.A(n_5611),
.Y(n_6691)
);

BUFx12f_ASAP7_75t_L g6692 ( 
.A(n_5648),
.Y(n_6692)
);

INVx2_ASAP7_75t_L g6693 ( 
.A(n_5483),
.Y(n_6693)
);

INVx2_ASAP7_75t_SL g6694 ( 
.A(n_5611),
.Y(n_6694)
);

CKINVDCx8_ASAP7_75t_R g6695 ( 
.A(n_5509),
.Y(n_6695)
);

CKINVDCx8_ASAP7_75t_R g6696 ( 
.A(n_5521),
.Y(n_6696)
);

AND2x2_ASAP7_75t_L g6697 ( 
.A(n_5765),
.B(n_4692),
.Y(n_6697)
);

CKINVDCx5p33_ASAP7_75t_R g6698 ( 
.A(n_5860),
.Y(n_6698)
);

INVx4_ASAP7_75t_L g6699 ( 
.A(n_5528),
.Y(n_6699)
);

A2O1A1Ixp33_ASAP7_75t_L g6700 ( 
.A1(n_5876),
.A2(n_5352),
.B(n_5451),
.C(n_4583),
.Y(n_6700)
);

INVx2_ASAP7_75t_L g6701 ( 
.A(n_5483),
.Y(n_6701)
);

NAND3xp33_ASAP7_75t_L g6702 ( 
.A(n_5876),
.B(n_5912),
.C(n_5892),
.Y(n_6702)
);

NAND2xp5_ASAP7_75t_SL g6703 ( 
.A(n_5932),
.B(n_4746),
.Y(n_6703)
);

OAI21xp33_ASAP7_75t_L g6704 ( 
.A1(n_5499),
.A2(n_4968),
.B(n_4961),
.Y(n_6704)
);

BUFx12f_ASAP7_75t_L g6705 ( 
.A(n_5648),
.Y(n_6705)
);

INVx2_ASAP7_75t_SL g6706 ( 
.A(n_5649),
.Y(n_6706)
);

INVx3_ASAP7_75t_L g6707 ( 
.A(n_5649),
.Y(n_6707)
);

INVx1_ASAP7_75t_L g6708 ( 
.A(n_5542),
.Y(n_6708)
);

NAND2xp5_ASAP7_75t_L g6709 ( 
.A(n_6184),
.B(n_4801),
.Y(n_6709)
);

INVxp67_ASAP7_75t_L g6710 ( 
.A(n_5965),
.Y(n_6710)
);

NAND2xp5_ASAP7_75t_SL g6711 ( 
.A(n_5932),
.B(n_4746),
.Y(n_6711)
);

INVx1_ASAP7_75t_L g6712 ( 
.A(n_5542),
.Y(n_6712)
);

INVx4_ASAP7_75t_L g6713 ( 
.A(n_5528),
.Y(n_6713)
);

O2A1O1Ixp33_ASAP7_75t_L g6714 ( 
.A1(n_5911),
.A2(n_5384),
.B(n_4970),
.C(n_4969),
.Y(n_6714)
);

INVx2_ASAP7_75t_L g6715 ( 
.A(n_5513),
.Y(n_6715)
);

CKINVDCx20_ASAP7_75t_R g6716 ( 
.A(n_5914),
.Y(n_6716)
);

BUFx3_ASAP7_75t_L g6717 ( 
.A(n_5619),
.Y(n_6717)
);

BUFx3_ASAP7_75t_L g6718 ( 
.A(n_5619),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_5542),
.Y(n_6719)
);

INVx2_ASAP7_75t_L g6720 ( 
.A(n_5513),
.Y(n_6720)
);

INVx2_ASAP7_75t_L g6721 ( 
.A(n_5513),
.Y(n_6721)
);

HB1xp67_ASAP7_75t_L g6722 ( 
.A(n_5982),
.Y(n_6722)
);

INVx3_ASAP7_75t_L g6723 ( 
.A(n_5649),
.Y(n_6723)
);

AOI21xp5_ASAP7_75t_L g6724 ( 
.A1(n_6221),
.A2(n_6222),
.B(n_5502),
.Y(n_6724)
);

NAND2xp5_ASAP7_75t_L g6725 ( 
.A(n_6184),
.B(n_4801),
.Y(n_6725)
);

INVx5_ASAP7_75t_L g6726 ( 
.A(n_5570),
.Y(n_6726)
);

INVx4_ASAP7_75t_L g6727 ( 
.A(n_5528),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_5742),
.B(n_4941),
.Y(n_6728)
);

BUFx8_ASAP7_75t_L g6729 ( 
.A(n_6138),
.Y(n_6729)
);

OR2x6_ASAP7_75t_L g6730 ( 
.A(n_6035),
.B(n_5267),
.Y(n_6730)
);

AOI21xp5_ASAP7_75t_L g6731 ( 
.A1(n_6221),
.A2(n_6222),
.B(n_5502),
.Y(n_6731)
);

AOI22xp33_ASAP7_75t_L g6732 ( 
.A1(n_5665),
.A2(n_5300),
.B1(n_4989),
.B2(n_4991),
.Y(n_6732)
);

OR2x2_ASAP7_75t_L g6733 ( 
.A(n_6078),
.B(n_4942),
.Y(n_6733)
);

INVx1_ASAP7_75t_L g6734 ( 
.A(n_5537),
.Y(n_6734)
);

INVx3_ASAP7_75t_L g6735 ( 
.A(n_5649),
.Y(n_6735)
);

INVx1_ASAP7_75t_L g6736 ( 
.A(n_5537),
.Y(n_6736)
);

NAND2xp5_ASAP7_75t_L g6737 ( 
.A(n_5742),
.B(n_4942),
.Y(n_6737)
);

INVx2_ASAP7_75t_L g6738 ( 
.A(n_5526),
.Y(n_6738)
);

AOI22xp33_ASAP7_75t_L g6739 ( 
.A1(n_5844),
.A2(n_4989),
.B1(n_4991),
.B2(n_4978),
.Y(n_6739)
);

BUFx3_ASAP7_75t_L g6740 ( 
.A(n_5619),
.Y(n_6740)
);

HB1xp67_ASAP7_75t_L g6741 ( 
.A(n_5982),
.Y(n_6741)
);

INVxp67_ASAP7_75t_SL g6742 ( 
.A(n_5500),
.Y(n_6742)
);

INVx2_ASAP7_75t_L g6743 ( 
.A(n_5526),
.Y(n_6743)
);

INVx2_ASAP7_75t_L g6744 ( 
.A(n_5526),
.Y(n_6744)
);

AOI21xp5_ASAP7_75t_L g6745 ( 
.A1(n_6001),
.A2(n_4664),
.B(n_5433),
.Y(n_6745)
);

CKINVDCx5p33_ASAP7_75t_R g6746 ( 
.A(n_6415),
.Y(n_6746)
);

INVx1_ASAP7_75t_L g6747 ( 
.A(n_5668),
.Y(n_6747)
);

BUFx2_ASAP7_75t_L g6748 ( 
.A(n_6190),
.Y(n_6748)
);

OAI21xp33_ASAP7_75t_SL g6749 ( 
.A1(n_5848),
.A2(n_5352),
.B(n_4971),
.Y(n_6749)
);

BUFx3_ASAP7_75t_L g6750 ( 
.A(n_5864),
.Y(n_6750)
);

AND2x2_ASAP7_75t_L g6751 ( 
.A(n_5765),
.B(n_4692),
.Y(n_6751)
);

NAND2xp5_ASAP7_75t_L g6752 ( 
.A(n_6033),
.B(n_4982),
.Y(n_6752)
);

INVx1_ASAP7_75t_L g6753 ( 
.A(n_5668),
.Y(n_6753)
);

O2A1O1Ixp33_ASAP7_75t_L g6754 ( 
.A1(n_5898),
.A2(n_5384),
.B(n_5001),
.C(n_5007),
.Y(n_6754)
);

CKINVDCx20_ASAP7_75t_R g6755 ( 
.A(n_5914),
.Y(n_6755)
);

AND2x2_ASAP7_75t_L g6756 ( 
.A(n_5765),
.B(n_4692),
.Y(n_6756)
);

INVx1_ASAP7_75t_L g6757 ( 
.A(n_5668),
.Y(n_6757)
);

NAND2xp5_ASAP7_75t_L g6758 ( 
.A(n_6055),
.B(n_4984),
.Y(n_6758)
);

BUFx3_ASAP7_75t_L g6759 ( 
.A(n_5864),
.Y(n_6759)
);

CKINVDCx5p33_ASAP7_75t_R g6760 ( 
.A(n_6415),
.Y(n_6760)
);

NAND2xp5_ASAP7_75t_L g6761 ( 
.A(n_6170),
.B(n_4942),
.Y(n_6761)
);

INVx1_ASAP7_75t_SL g6762 ( 
.A(n_6518),
.Y(n_6762)
);

BUFx2_ASAP7_75t_L g6763 ( 
.A(n_6190),
.Y(n_6763)
);

BUFx2_ASAP7_75t_L g6764 ( 
.A(n_6190),
.Y(n_6764)
);

NOR2xp33_ASAP7_75t_L g6765 ( 
.A(n_5962),
.B(n_5451),
.Y(n_6765)
);

HB1xp67_ASAP7_75t_L g6766 ( 
.A(n_5500),
.Y(n_6766)
);

BUFx12f_ASAP7_75t_L g6767 ( 
.A(n_5733),
.Y(n_6767)
);

NAND2xp5_ASAP7_75t_L g6768 ( 
.A(n_6055),
.B(n_4984),
.Y(n_6768)
);

INVx3_ASAP7_75t_L g6769 ( 
.A(n_5649),
.Y(n_6769)
);

NAND2xp5_ASAP7_75t_L g6770 ( 
.A(n_5891),
.B(n_5041),
.Y(n_6770)
);

INVx1_ASAP7_75t_SL g6771 ( 
.A(n_5917),
.Y(n_6771)
);

INVx3_ASAP7_75t_SL g6772 ( 
.A(n_6303),
.Y(n_6772)
);

HB1xp67_ASAP7_75t_L g6773 ( 
.A(n_5512),
.Y(n_6773)
);

INVx3_ASAP7_75t_L g6774 ( 
.A(n_5679),
.Y(n_6774)
);

AOI21xp5_ASAP7_75t_L g6775 ( 
.A1(n_6001),
.A2(n_6367),
.B(n_6362),
.Y(n_6775)
);

INVx2_ASAP7_75t_L g6776 ( 
.A(n_5527),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_5773),
.Y(n_6777)
);

AOI22xp33_ASAP7_75t_L g6778 ( 
.A1(n_5844),
.A2(n_5001),
.B1(n_5007),
.B2(n_4994),
.Y(n_6778)
);

NOR2xp33_ASAP7_75t_L g6779 ( 
.A(n_5962),
.B(n_5284),
.Y(n_6779)
);

BUFx2_ASAP7_75t_L g6780 ( 
.A(n_6365),
.Y(n_6780)
);

INVx1_ASAP7_75t_L g6781 ( 
.A(n_5773),
.Y(n_6781)
);

NOR2xp33_ASAP7_75t_L g6782 ( 
.A(n_5908),
.B(n_5284),
.Y(n_6782)
);

NOR2xp33_ASAP7_75t_L g6783 ( 
.A(n_5908),
.B(n_5287),
.Y(n_6783)
);

NOR2xp33_ASAP7_75t_L g6784 ( 
.A(n_5854),
.B(n_5287),
.Y(n_6784)
);

INVx3_ASAP7_75t_L g6785 ( 
.A(n_5679),
.Y(n_6785)
);

HB1xp67_ASAP7_75t_L g6786 ( 
.A(n_5512),
.Y(n_6786)
);

CKINVDCx20_ASAP7_75t_R g6787 ( 
.A(n_5952),
.Y(n_6787)
);

NOR2xp33_ASAP7_75t_L g6788 ( 
.A(n_5854),
.B(n_5867),
.Y(n_6788)
);

INVx1_ASAP7_75t_L g6789 ( 
.A(n_5593),
.Y(n_6789)
);

INVx2_ASAP7_75t_SL g6790 ( 
.A(n_5679),
.Y(n_6790)
);

INVx1_ASAP7_75t_SL g6791 ( 
.A(n_5917),
.Y(n_6791)
);

BUFx5_ASAP7_75t_L g6792 ( 
.A(n_5717),
.Y(n_6792)
);

NAND2xp5_ASAP7_75t_L g6793 ( 
.A(n_5891),
.B(n_5041),
.Y(n_6793)
);

INVx3_ASAP7_75t_L g6794 ( 
.A(n_5679),
.Y(n_6794)
);

BUFx12f_ASAP7_75t_L g6795 ( 
.A(n_5733),
.Y(n_6795)
);

AOI22xp5_ASAP7_75t_L g6796 ( 
.A1(n_5868),
.A2(n_4914),
.B1(n_5044),
.B2(n_5012),
.Y(n_6796)
);

AOI22xp5_ASAP7_75t_L g6797 ( 
.A1(n_5835),
.A2(n_5044),
.B1(n_5049),
.B2(n_5012),
.Y(n_6797)
);

AOI22xp5_ASAP7_75t_L g6798 ( 
.A1(n_5835),
.A2(n_5053),
.B1(n_5056),
.B2(n_5049),
.Y(n_6798)
);

NAND2xp5_ASAP7_75t_L g6799 ( 
.A(n_5896),
.B(n_5047),
.Y(n_6799)
);

O2A1O1Ixp5_ASAP7_75t_L g6800 ( 
.A1(n_5890),
.A2(n_4606),
.B(n_4860),
.C(n_4741),
.Y(n_6800)
);

INVx2_ASAP7_75t_L g6801 ( 
.A(n_5527),
.Y(n_6801)
);

CKINVDCx11_ASAP7_75t_R g6802 ( 
.A(n_5952),
.Y(n_6802)
);

INVx2_ASAP7_75t_SL g6803 ( 
.A(n_5679),
.Y(n_6803)
);

BUFx12f_ASAP7_75t_L g6804 ( 
.A(n_5847),
.Y(n_6804)
);

BUFx2_ASAP7_75t_L g6805 ( 
.A(n_6365),
.Y(n_6805)
);

BUFx8_ASAP7_75t_L g6806 ( 
.A(n_6138),
.Y(n_6806)
);

NAND2xp5_ASAP7_75t_L g6807 ( 
.A(n_5896),
.B(n_5047),
.Y(n_6807)
);

INVx1_ASAP7_75t_L g6808 ( 
.A(n_5593),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_5593),
.Y(n_6809)
);

INVx2_ASAP7_75t_SL g6810 ( 
.A(n_5685),
.Y(n_6810)
);

BUFx3_ASAP7_75t_L g6811 ( 
.A(n_5864),
.Y(n_6811)
);

BUFx2_ASAP7_75t_L g6812 ( 
.A(n_6365),
.Y(n_6812)
);

HB1xp67_ASAP7_75t_L g6813 ( 
.A(n_6356),
.Y(n_6813)
);

INVx1_ASAP7_75t_L g6814 ( 
.A(n_5595),
.Y(n_6814)
);

AOI22xp5_ASAP7_75t_L g6815 ( 
.A1(n_5922),
.A2(n_5056),
.B1(n_5058),
.B2(n_5053),
.Y(n_6815)
);

NOR2xp33_ASAP7_75t_L g6816 ( 
.A(n_5867),
.B(n_5289),
.Y(n_6816)
);

INVx1_ASAP7_75t_L g6817 ( 
.A(n_5574),
.Y(n_6817)
);

NAND2xp5_ASAP7_75t_L g6818 ( 
.A(n_6170),
.B(n_4955),
.Y(n_6818)
);

HB1xp67_ASAP7_75t_L g6819 ( 
.A(n_6356),
.Y(n_6819)
);

NAND2xp5_ASAP7_75t_L g6820 ( 
.A(n_6170),
.B(n_4955),
.Y(n_6820)
);

OR2x6_ASAP7_75t_L g6821 ( 
.A(n_6035),
.B(n_5267),
.Y(n_6821)
);

INVx1_ASAP7_75t_L g6822 ( 
.A(n_5582),
.Y(n_6822)
);

AOI22xp33_ASAP7_75t_L g6823 ( 
.A1(n_5836),
.A2(n_4994),
.B1(n_5011),
.B2(n_5219),
.Y(n_6823)
);

AOI221xp5_ASAP7_75t_L g6824 ( 
.A1(n_5836),
.A2(n_5011),
.B1(n_5289),
.B2(n_5293),
.C(n_5290),
.Y(n_6824)
);

AOI21xp5_ASAP7_75t_L g6825 ( 
.A1(n_6362),
.A2(n_5436),
.B(n_5433),
.Y(n_6825)
);

NAND2xp5_ASAP7_75t_L g6826 ( 
.A(n_6276),
.B(n_5073),
.Y(n_6826)
);

NAND2xp33_ASAP7_75t_L g6827 ( 
.A(n_5721),
.B(n_5267),
.Y(n_6827)
);

INVx6_ASAP7_75t_L g6828 ( 
.A(n_6461),
.Y(n_6828)
);

INVx1_ASAP7_75t_L g6829 ( 
.A(n_5582),
.Y(n_6829)
);

NAND3xp33_ASAP7_75t_L g6830 ( 
.A(n_5912),
.B(n_5437),
.C(n_5436),
.Y(n_6830)
);

NAND2xp5_ASAP7_75t_L g6831 ( 
.A(n_6276),
.B(n_5073),
.Y(n_6831)
);

AOI211xp5_ASAP7_75t_L g6832 ( 
.A1(n_5893),
.A2(n_5078),
.B(n_5097),
.C(n_5058),
.Y(n_6832)
);

AOI221xp5_ASAP7_75t_L g6833 ( 
.A1(n_6111),
.A2(n_5892),
.B1(n_5893),
.B2(n_5499),
.C(n_5910),
.Y(n_6833)
);

BUFx2_ASAP7_75t_L g6834 ( 
.A(n_6365),
.Y(n_6834)
);

NAND2xp5_ASAP7_75t_L g6835 ( 
.A(n_6284),
.B(n_5106),
.Y(n_6835)
);

CKINVDCx20_ASAP7_75t_R g6836 ( 
.A(n_5629),
.Y(n_6836)
);

NAND2x1_ASAP7_75t_L g6837 ( 
.A(n_5551),
.B(n_4512),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6284),
.B(n_5106),
.Y(n_6838)
);

INVx3_ASAP7_75t_L g6839 ( 
.A(n_5685),
.Y(n_6839)
);

AOI22xp5_ASAP7_75t_L g6840 ( 
.A1(n_5922),
.A2(n_5078),
.B1(n_5117),
.B2(n_5097),
.Y(n_6840)
);

OAI21xp5_ASAP7_75t_L g6841 ( 
.A1(n_5848),
.A2(n_5440),
.B(n_5437),
.Y(n_6841)
);

INVx1_ASAP7_75t_L g6842 ( 
.A(n_5554),
.Y(n_6842)
);

INVx3_ASAP7_75t_L g6843 ( 
.A(n_5685),
.Y(n_6843)
);

INVx1_ASAP7_75t_L g6844 ( 
.A(n_5554),
.Y(n_6844)
);

OAI21x1_ASAP7_75t_L g6845 ( 
.A1(n_6029),
.A2(n_4743),
.B(n_4747),
.Y(n_6845)
);

NOR2xp33_ASAP7_75t_L g6846 ( 
.A(n_5913),
.B(n_5290),
.Y(n_6846)
);

BUFx2_ASAP7_75t_L g6847 ( 
.A(n_6365),
.Y(n_6847)
);

AOI22xp5_ASAP7_75t_L g6848 ( 
.A1(n_5910),
.A2(n_5935),
.B1(n_5889),
.B2(n_5967),
.Y(n_6848)
);

INVx1_ASAP7_75t_L g6849 ( 
.A(n_5562),
.Y(n_6849)
);

NAND2xp5_ASAP7_75t_L g6850 ( 
.A(n_6298),
.B(n_6232),
.Y(n_6850)
);

INVx1_ASAP7_75t_L g6851 ( 
.A(n_5562),
.Y(n_6851)
);

NOR2xp33_ASAP7_75t_SL g6852 ( 
.A(n_5933),
.B(n_4588),
.Y(n_6852)
);

INVx1_ASAP7_75t_L g6853 ( 
.A(n_5562),
.Y(n_6853)
);

NOR2xp33_ASAP7_75t_L g6854 ( 
.A(n_5913),
.B(n_5293),
.Y(n_6854)
);

BUFx2_ASAP7_75t_L g6855 ( 
.A(n_6365),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_5663),
.Y(n_6856)
);

CKINVDCx5p33_ASAP7_75t_R g6857 ( 
.A(n_6547),
.Y(n_6857)
);

CKINVDCx20_ASAP7_75t_R g6858 ( 
.A(n_5629),
.Y(n_6858)
);

INVx3_ASAP7_75t_L g6859 ( 
.A(n_5685),
.Y(n_6859)
);

NAND2xp5_ASAP7_75t_L g6860 ( 
.A(n_5917),
.B(n_4955),
.Y(n_6860)
);

OR2x6_ASAP7_75t_SL g6861 ( 
.A(n_5511),
.B(n_5350),
.Y(n_6861)
);

AOI222xp33_ASAP7_75t_L g6862 ( 
.A1(n_6050),
.A2(n_4481),
.B1(n_4639),
.B2(n_4935),
.C1(n_4927),
.C2(n_4905),
.Y(n_6862)
);

NAND2xp5_ASAP7_75t_L g6863 ( 
.A(n_5978),
.B(n_6039),
.Y(n_6863)
);

AOI21xp5_ASAP7_75t_L g6864 ( 
.A1(n_6367),
.A2(n_5448),
.B(n_5440),
.Y(n_6864)
);

INVx1_ASAP7_75t_L g6865 ( 
.A(n_5703),
.Y(n_6865)
);

AND2x2_ASAP7_75t_SL g6866 ( 
.A(n_5697),
.B(n_5352),
.Y(n_6866)
);

NOR2xp33_ASAP7_75t_SL g6867 ( 
.A(n_5933),
.B(n_4588),
.Y(n_6867)
);

NAND2xp5_ASAP7_75t_L g6868 ( 
.A(n_6298),
.B(n_5118),
.Y(n_6868)
);

BUFx8_ASAP7_75t_L g6869 ( 
.A(n_6138),
.Y(n_6869)
);

INVx1_ASAP7_75t_L g6870 ( 
.A(n_5703),
.Y(n_6870)
);

AOI22xp33_ASAP7_75t_L g6871 ( 
.A1(n_5643),
.A2(n_5463),
.B1(n_5357),
.B2(n_5065),
.Y(n_6871)
);

OAI21x1_ASAP7_75t_L g6872 ( 
.A1(n_6029),
.A2(n_4811),
.B(n_4747),
.Y(n_6872)
);

INVx2_ASAP7_75t_SL g6873 ( 
.A(n_5685),
.Y(n_6873)
);

BUFx12f_ASAP7_75t_L g6874 ( 
.A(n_5847),
.Y(n_6874)
);

INVx4_ASAP7_75t_L g6875 ( 
.A(n_5528),
.Y(n_6875)
);

NAND2xp5_ASAP7_75t_L g6876 ( 
.A(n_6232),
.B(n_5118),
.Y(n_6876)
);

INVxp67_ASAP7_75t_L g6877 ( 
.A(n_5971),
.Y(n_6877)
);

INVx4_ASAP7_75t_L g6878 ( 
.A(n_5528),
.Y(n_6878)
);

A2O1A1Ixp33_ASAP7_75t_SL g6879 ( 
.A1(n_5535),
.A2(n_5462),
.B(n_5450),
.C(n_4811),
.Y(n_6879)
);

AO21x2_ASAP7_75t_L g6880 ( 
.A1(n_6233),
.A2(n_5462),
.B(n_5450),
.Y(n_6880)
);

INVxp67_ASAP7_75t_SL g6881 ( 
.A(n_6385),
.Y(n_6881)
);

INVxp67_ASAP7_75t_L g6882 ( 
.A(n_5971),
.Y(n_6882)
);

AOI21xp5_ASAP7_75t_L g6883 ( 
.A1(n_6024),
.A2(n_5342),
.B(n_4937),
.Y(n_6883)
);

HB1xp67_ASAP7_75t_L g6884 ( 
.A(n_6385),
.Y(n_6884)
);

INVx3_ASAP7_75t_L g6885 ( 
.A(n_5691),
.Y(n_6885)
);

OR2x2_ASAP7_75t_L g6886 ( 
.A(n_6058),
.B(n_4811),
.Y(n_6886)
);

CKINVDCx5p33_ASAP7_75t_R g6887 ( 
.A(n_6547),
.Y(n_6887)
);

AOI21xp5_ASAP7_75t_L g6888 ( 
.A1(n_6024),
.A2(n_5342),
.B(n_4937),
.Y(n_6888)
);

AOI22xp33_ASAP7_75t_L g6889 ( 
.A1(n_5643),
.A2(n_5463),
.B1(n_5357),
.B2(n_5065),
.Y(n_6889)
);

INVxp67_ASAP7_75t_SL g6890 ( 
.A(n_6403),
.Y(n_6890)
);

A2O1A1Ixp33_ASAP7_75t_L g6891 ( 
.A1(n_5956),
.A2(n_4860),
.B(n_5082),
.C(n_4937),
.Y(n_6891)
);

BUFx2_ASAP7_75t_L g6892 ( 
.A(n_6365),
.Y(n_6892)
);

CKINVDCx5p33_ASAP7_75t_R g6893 ( 
.A(n_5875),
.Y(n_6893)
);

INVx3_ASAP7_75t_SL g6894 ( 
.A(n_6303),
.Y(n_6894)
);

INVx4_ASAP7_75t_L g6895 ( 
.A(n_5528),
.Y(n_6895)
);

INVx3_ASAP7_75t_L g6896 ( 
.A(n_5691),
.Y(n_6896)
);

NAND2xp5_ASAP7_75t_L g6897 ( 
.A(n_6056),
.B(n_5120),
.Y(n_6897)
);

INVx1_ASAP7_75t_SL g6898 ( 
.A(n_5978),
.Y(n_6898)
);

INVx2_ASAP7_75t_SL g6899 ( 
.A(n_5691),
.Y(n_6899)
);

NAND2xp5_ASAP7_75t_L g6900 ( 
.A(n_6056),
.B(n_5120),
.Y(n_6900)
);

BUFx2_ASAP7_75t_L g6901 ( 
.A(n_6365),
.Y(n_6901)
);

OR2x2_ASAP7_75t_L g6902 ( 
.A(n_6058),
.B(n_4811),
.Y(n_6902)
);

NAND2xp5_ASAP7_75t_L g6903 ( 
.A(n_6060),
.B(n_5833),
.Y(n_6903)
);

AOI22xp5_ASAP7_75t_L g6904 ( 
.A1(n_5935),
.A2(n_5117),
.B1(n_5121),
.B2(n_4431),
.Y(n_6904)
);

BUFx3_ASAP7_75t_L g6905 ( 
.A(n_5864),
.Y(n_6905)
);

BUFx3_ASAP7_75t_L g6906 ( 
.A(n_5864),
.Y(n_6906)
);

HB1xp67_ASAP7_75t_L g6907 ( 
.A(n_6403),
.Y(n_6907)
);

NAND2xp5_ASAP7_75t_L g6908 ( 
.A(n_6060),
.B(n_5137),
.Y(n_6908)
);

CKINVDCx5p33_ASAP7_75t_R g6909 ( 
.A(n_5875),
.Y(n_6909)
);

AOI21xp5_ASAP7_75t_L g6910 ( 
.A1(n_5530),
.A2(n_5342),
.B(n_4937),
.Y(n_6910)
);

NAND2xp5_ASAP7_75t_L g6911 ( 
.A(n_5833),
.B(n_5137),
.Y(n_6911)
);

BUFx3_ASAP7_75t_L g6912 ( 
.A(n_6127),
.Y(n_6912)
);

NAND2xp5_ASAP7_75t_L g6913 ( 
.A(n_5841),
.B(n_5152),
.Y(n_6913)
);

OAI22xp5_ASAP7_75t_L g6914 ( 
.A1(n_5721),
.A2(n_4459),
.B1(n_5121),
.B2(n_4937),
.Y(n_6914)
);

OR2x2_ASAP7_75t_SL g6915 ( 
.A(n_5602),
.B(n_5417),
.Y(n_6915)
);

INVx5_ASAP7_75t_L g6916 ( 
.A(n_5471),
.Y(n_6916)
);

BUFx2_ASAP7_75t_L g6917 ( 
.A(n_6450),
.Y(n_6917)
);

BUFx2_ASAP7_75t_L g6918 ( 
.A(n_6450),
.Y(n_6918)
);

CKINVDCx6p67_ASAP7_75t_R g6919 ( 
.A(n_6205),
.Y(n_6919)
);

INVx1_ASAP7_75t_SL g6920 ( 
.A(n_5978),
.Y(n_6920)
);

NAND2xp5_ASAP7_75t_SL g6921 ( 
.A(n_5889),
.B(n_4814),
.Y(n_6921)
);

INVx3_ASAP7_75t_SL g6922 ( 
.A(n_6303),
.Y(n_6922)
);

INVx5_ASAP7_75t_L g6923 ( 
.A(n_5471),
.Y(n_6923)
);

AOI21xp5_ASAP7_75t_L g6924 ( 
.A1(n_5530),
.A2(n_5342),
.B(n_5082),
.Y(n_6924)
);

INVxp67_ASAP7_75t_L g6925 ( 
.A(n_6135),
.Y(n_6925)
);

NOR4xp25_ASAP7_75t_L g6926 ( 
.A(n_5956),
.B(n_5181),
.C(n_5225),
.D(n_5164),
.Y(n_6926)
);

AND2x4_ASAP7_75t_L g6927 ( 
.A(n_6428),
.B(n_6429),
.Y(n_6927)
);

INVx1_ASAP7_75t_SL g6928 ( 
.A(n_6247),
.Y(n_6928)
);

OAI21x1_ASAP7_75t_SL g6929 ( 
.A1(n_5918),
.A2(n_4838),
.B(n_4834),
.Y(n_6929)
);

BUFx6f_ASAP7_75t_SL g6930 ( 
.A(n_5713),
.Y(n_6930)
);

AO32x2_ASAP7_75t_L g6931 ( 
.A1(n_5989),
.A2(n_4485),
.A3(n_4441),
.B1(n_4433),
.B2(n_4834),
.Y(n_6931)
);

NAND2xp5_ASAP7_75t_L g6932 ( 
.A(n_5841),
.B(n_5152),
.Y(n_6932)
);

NAND2xp5_ASAP7_75t_L g6933 ( 
.A(n_6380),
.B(n_5155),
.Y(n_6933)
);

INVx4_ASAP7_75t_L g6934 ( 
.A(n_5528),
.Y(n_6934)
);

NAND2xp5_ASAP7_75t_L g6935 ( 
.A(n_6380),
.B(n_5155),
.Y(n_6935)
);

AOI21xp5_ASAP7_75t_L g6936 ( 
.A1(n_6217),
.A2(n_6041),
.B(n_6038),
.Y(n_6936)
);

INVx3_ASAP7_75t_L g6937 ( 
.A(n_5691),
.Y(n_6937)
);

O2A1O1Ixp5_ASAP7_75t_L g6938 ( 
.A1(n_5890),
.A2(n_5082),
.B(n_5168),
.C(n_4860),
.Y(n_6938)
);

OR2x2_ASAP7_75t_L g6939 ( 
.A(n_6058),
.B(n_4823),
.Y(n_6939)
);

BUFx10_ASAP7_75t_L g6940 ( 
.A(n_6138),
.Y(n_6940)
);

BUFx3_ASAP7_75t_L g6941 ( 
.A(n_6127),
.Y(n_6941)
);

BUFx2_ASAP7_75t_SL g6942 ( 
.A(n_6127),
.Y(n_6942)
);

NAND2xp5_ASAP7_75t_SL g6943 ( 
.A(n_5970),
.B(n_4814),
.Y(n_6943)
);

NAND2xp5_ASAP7_75t_L g6944 ( 
.A(n_6039),
.B(n_4817),
.Y(n_6944)
);

BUFx10_ASAP7_75t_L g6945 ( 
.A(n_6138),
.Y(n_6945)
);

INVx4_ASAP7_75t_SL g6946 ( 
.A(n_5717),
.Y(n_6946)
);

O2A1O1Ixp33_ASAP7_75t_L g6947 ( 
.A1(n_5915),
.A2(n_5308),
.B(n_5337),
.C(n_5286),
.Y(n_6947)
);

INVx1_ASAP7_75t_L g6948 ( 
.A(n_5762),
.Y(n_6948)
);

AND2x2_ASAP7_75t_L g6949 ( 
.A(n_5766),
.B(n_5772),
.Y(n_6949)
);

AOI21xp5_ASAP7_75t_L g6950 ( 
.A1(n_6217),
.A2(n_5342),
.B(n_5168),
.Y(n_6950)
);

CKINVDCx5p33_ASAP7_75t_R g6951 ( 
.A(n_5977),
.Y(n_6951)
);

BUFx3_ASAP7_75t_L g6952 ( 
.A(n_6243),
.Y(n_6952)
);

INVx1_ASAP7_75t_SL g6953 ( 
.A(n_6247),
.Y(n_6953)
);

NOR2xp33_ASAP7_75t_L g6954 ( 
.A(n_5723),
.B(n_5164),
.Y(n_6954)
);

OR2x2_ASAP7_75t_SL g6955 ( 
.A(n_5602),
.B(n_5417),
.Y(n_6955)
);

AOI21xp5_ASAP7_75t_L g6956 ( 
.A1(n_6038),
.A2(n_5168),
.B(n_5082),
.Y(n_6956)
);

INVx1_ASAP7_75t_L g6957 ( 
.A(n_5763),
.Y(n_6957)
);

NAND2xp5_ASAP7_75t_L g6958 ( 
.A(n_6409),
.B(n_5188),
.Y(n_6958)
);

BUFx2_ASAP7_75t_SL g6959 ( 
.A(n_6243),
.Y(n_6959)
);

INVxp67_ASAP7_75t_L g6960 ( 
.A(n_6135),
.Y(n_6960)
);

BUFx3_ASAP7_75t_L g6961 ( 
.A(n_6243),
.Y(n_6961)
);

INVx2_ASAP7_75t_SL g6962 ( 
.A(n_5715),
.Y(n_6962)
);

INVx4_ASAP7_75t_L g6963 ( 
.A(n_5534),
.Y(n_6963)
);

INVx1_ASAP7_75t_SL g6964 ( 
.A(n_6247),
.Y(n_6964)
);

INVx4_ASAP7_75t_L g6965 ( 
.A(n_5534),
.Y(n_6965)
);

NAND2xp5_ASAP7_75t_L g6966 ( 
.A(n_6498),
.B(n_4400),
.Y(n_6966)
);

AND2x2_ASAP7_75t_L g6967 ( 
.A(n_5766),
.B(n_5772),
.Y(n_6967)
);

NAND2xp5_ASAP7_75t_L g6968 ( 
.A(n_6498),
.B(n_4400),
.Y(n_6968)
);

CKINVDCx5p33_ASAP7_75t_R g6969 ( 
.A(n_5977),
.Y(n_6969)
);

OAI22xp33_ASAP7_75t_L g6970 ( 
.A1(n_5840),
.A2(n_4459),
.B1(n_5064),
.B2(n_5149),
.Y(n_6970)
);

INVx1_ASAP7_75t_L g6971 ( 
.A(n_5764),
.Y(n_6971)
);

AND2x6_ASAP7_75t_L g6972 ( 
.A(n_6083),
.B(n_4442),
.Y(n_6972)
);

OR2x2_ASAP7_75t_L g6973 ( 
.A(n_6058),
.B(n_4826),
.Y(n_6973)
);

OR2x2_ASAP7_75t_L g6974 ( 
.A(n_6058),
.B(n_4826),
.Y(n_6974)
);

INVxp67_ASAP7_75t_SL g6975 ( 
.A(n_6448),
.Y(n_6975)
);

BUFx4f_ASAP7_75t_L g6976 ( 
.A(n_5662),
.Y(n_6976)
);

OR2x2_ASAP7_75t_L g6977 ( 
.A(n_6376),
.B(n_4826),
.Y(n_6977)
);

HB1xp67_ASAP7_75t_L g6978 ( 
.A(n_6448),
.Y(n_6978)
);

BUFx3_ASAP7_75t_L g6979 ( 
.A(n_6361),
.Y(n_6979)
);

INVxp67_ASAP7_75t_SL g6980 ( 
.A(n_6207),
.Y(n_6980)
);

OAI22xp5_ASAP7_75t_SL g6981 ( 
.A1(n_5871),
.A2(n_4459),
.B1(n_5096),
.B2(n_4993),
.Y(n_6981)
);

NAND2xp5_ASAP7_75t_L g6982 ( 
.A(n_6480),
.B(n_4418),
.Y(n_6982)
);

HB1xp67_ASAP7_75t_L g6983 ( 
.A(n_6062),
.Y(n_6983)
);

CKINVDCx16_ASAP7_75t_R g6984 ( 
.A(n_6135),
.Y(n_6984)
);

OA21x2_ASAP7_75t_L g6985 ( 
.A1(n_5861),
.A2(n_5042),
.B(n_5038),
.Y(n_6985)
);

BUFx3_ASAP7_75t_L g6986 ( 
.A(n_6361),
.Y(n_6986)
);

AOI21xp5_ASAP7_75t_L g6987 ( 
.A1(n_6041),
.A2(n_5168),
.B(n_5082),
.Y(n_6987)
);

NAND2xp5_ASAP7_75t_L g6988 ( 
.A(n_6480),
.B(n_4418),
.Y(n_6988)
);

AND2x2_ASAP7_75t_SL g6989 ( 
.A(n_5697),
.B(n_5311),
.Y(n_6989)
);

BUFx2_ASAP7_75t_L g6990 ( 
.A(n_6450),
.Y(n_6990)
);

AND2x2_ASAP7_75t_SL g6991 ( 
.A(n_5697),
.B(n_5311),
.Y(n_6991)
);

BUFx12f_ASAP7_75t_L g6992 ( 
.A(n_6116),
.Y(n_6992)
);

CKINVDCx8_ASAP7_75t_R g6993 ( 
.A(n_5521),
.Y(n_6993)
);

AOI22xp33_ASAP7_75t_L g6994 ( 
.A1(n_5925),
.A2(n_5065),
.B1(n_5420),
.B2(n_5255),
.Y(n_6994)
);

AOI22xp5_ASAP7_75t_L g6995 ( 
.A1(n_5967),
.A2(n_4431),
.B1(n_5420),
.B2(n_5148),
.Y(n_6995)
);

NAND2x1p5_ASAP7_75t_L g6996 ( 
.A(n_5487),
.B(n_4591),
.Y(n_6996)
);

AOI22xp33_ASAP7_75t_L g6997 ( 
.A1(n_5925),
.A2(n_5065),
.B1(n_5255),
.B2(n_5246),
.Y(n_6997)
);

BUFx3_ASAP7_75t_L g6998 ( 
.A(n_6361),
.Y(n_6998)
);

HB1xp67_ASAP7_75t_L g6999 ( 
.A(n_6062),
.Y(n_6999)
);

AO21x2_ASAP7_75t_L g7000 ( 
.A1(n_6233),
.A2(n_6263),
.B(n_6234),
.Y(n_7000)
);

NOR2xp33_ASAP7_75t_L g7001 ( 
.A(n_5723),
.B(n_5181),
.Y(n_7001)
);

INVx5_ASAP7_75t_L g7002 ( 
.A(n_5487),
.Y(n_7002)
);

NOR3xp33_ASAP7_75t_L g7003 ( 
.A(n_5861),
.B(n_4963),
.C(n_4672),
.Y(n_7003)
);

INVx2_ASAP7_75t_SL g7004 ( 
.A(n_5715),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_5700),
.Y(n_7005)
);

CKINVDCx8_ASAP7_75t_R g7006 ( 
.A(n_5872),
.Y(n_7006)
);

AOI22xp33_ASAP7_75t_L g7007 ( 
.A1(n_6050),
.A2(n_5065),
.B1(n_5349),
.B2(n_5246),
.Y(n_7007)
);

CKINVDCx5p33_ASAP7_75t_R g7008 ( 
.A(n_6116),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_5700),
.Y(n_7009)
);

OAI22xp5_ASAP7_75t_L g7010 ( 
.A1(n_5840),
.A2(n_5208),
.B1(n_5168),
.B2(n_5150),
.Y(n_7010)
);

AOI221x1_ASAP7_75t_L g7011 ( 
.A1(n_5940),
.A2(n_5405),
.B1(n_4854),
.B2(n_4832),
.C(n_4826),
.Y(n_7011)
);

OAI22x1_ASAP7_75t_L g7012 ( 
.A1(n_5961),
.A2(n_4497),
.B1(n_5018),
.B2(n_5013),
.Y(n_7012)
);

INVx2_ASAP7_75t_SL g7013 ( 
.A(n_5715),
.Y(n_7013)
);

BUFx12f_ASAP7_75t_L g7014 ( 
.A(n_6538),
.Y(n_7014)
);

BUFx8_ASAP7_75t_L g7015 ( 
.A(n_6364),
.Y(n_7015)
);

BUFx2_ASAP7_75t_L g7016 ( 
.A(n_6450),
.Y(n_7016)
);

NOR2x1_ASAP7_75t_L g7017 ( 
.A(n_6110),
.B(n_4832),
.Y(n_7017)
);

AOI22xp5_ASAP7_75t_L g7018 ( 
.A1(n_5929),
.A2(n_5953),
.B1(n_5834),
.B2(n_5928),
.Y(n_7018)
);

NAND2xp5_ASAP7_75t_L g7019 ( 
.A(n_6409),
.B(n_6427),
.Y(n_7019)
);

INVxp67_ASAP7_75t_L g7020 ( 
.A(n_5947),
.Y(n_7020)
);

NAND2xp5_ASAP7_75t_L g7021 ( 
.A(n_6427),
.B(n_6260),
.Y(n_7021)
);

INVx5_ASAP7_75t_L g7022 ( 
.A(n_6030),
.Y(n_7022)
);

NOR3xp33_ASAP7_75t_SL g7023 ( 
.A(n_5782),
.B(n_4944),
.C(n_4938),
.Y(n_7023)
);

NAND2xp5_ASAP7_75t_L g7024 ( 
.A(n_6260),
.B(n_5188),
.Y(n_7024)
);

BUFx6f_ASAP7_75t_L g7025 ( 
.A(n_6417),
.Y(n_7025)
);

AOI21xp5_ASAP7_75t_L g7026 ( 
.A1(n_6069),
.A2(n_5208),
.B(n_5325),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_5724),
.Y(n_7027)
);

AND2x4_ASAP7_75t_SL g7028 ( 
.A(n_5713),
.B(n_5948),
.Y(n_7028)
);

INVxp67_ASAP7_75t_L g7029 ( 
.A(n_5947),
.Y(n_7029)
);

AOI21xp33_ASAP7_75t_L g7030 ( 
.A1(n_5970),
.A2(n_5339),
.B(n_5325),
.Y(n_7030)
);

CKINVDCx20_ASAP7_75t_R g7031 ( 
.A(n_5712),
.Y(n_7031)
);

NAND2xp5_ASAP7_75t_SL g7032 ( 
.A(n_5519),
.B(n_5212),
.Y(n_7032)
);

AOI22xp33_ASAP7_75t_L g7033 ( 
.A1(n_6064),
.A2(n_5065),
.B1(n_5349),
.B2(n_5435),
.Y(n_7033)
);

AND2x2_ASAP7_75t_L g7034 ( 
.A(n_5784),
.B(n_6215),
.Y(n_7034)
);

NAND2x1p5_ASAP7_75t_L g7035 ( 
.A(n_5697),
.B(n_4591),
.Y(n_7035)
);

NOR2xp67_ASAP7_75t_SL g7036 ( 
.A(n_5927),
.B(n_4546),
.Y(n_7036)
);

INVx2_ASAP7_75t_SL g7037 ( 
.A(n_5727),
.Y(n_7037)
);

OAI22xp5_ASAP7_75t_L g7038 ( 
.A1(n_5953),
.A2(n_5895),
.B1(n_5824),
.B2(n_6216),
.Y(n_7038)
);

AND2x2_ASAP7_75t_SL g7039 ( 
.A(n_5697),
.B(n_5311),
.Y(n_7039)
);

AOI22xp33_ASAP7_75t_L g7040 ( 
.A1(n_6064),
.A2(n_5824),
.B1(n_6013),
.B2(n_5915),
.Y(n_7040)
);

AOI22xp33_ASAP7_75t_L g7041 ( 
.A1(n_6013),
.A2(n_5454),
.B1(n_5435),
.B2(n_5196),
.Y(n_7041)
);

AO21x1_ASAP7_75t_L g7042 ( 
.A1(n_6100),
.A2(n_5405),
.B(n_5004),
.Y(n_7042)
);

NAND2xp5_ASAP7_75t_SL g7043 ( 
.A(n_5519),
.B(n_5212),
.Y(n_7043)
);

OR2x2_ASAP7_75t_L g7044 ( 
.A(n_6376),
.B(n_4832),
.Y(n_7044)
);

INVx1_ASAP7_75t_SL g7045 ( 
.A(n_6297),
.Y(n_7045)
);

BUFx12f_ASAP7_75t_L g7046 ( 
.A(n_6538),
.Y(n_7046)
);

BUFx6f_ASAP7_75t_L g7047 ( 
.A(n_6417),
.Y(n_7047)
);

AOI22xp5_ASAP7_75t_L g7048 ( 
.A1(n_5929),
.A2(n_5148),
.B1(n_5252),
.B2(n_5150),
.Y(n_7048)
);

NAND2xp5_ASAP7_75t_L g7049 ( 
.A(n_6015),
.B(n_5209),
.Y(n_7049)
);

INVx4_ASAP7_75t_L g7050 ( 
.A(n_5534),
.Y(n_7050)
);

NAND2xp5_ASAP7_75t_L g7051 ( 
.A(n_6554),
.B(n_4418),
.Y(n_7051)
);

BUFx3_ASAP7_75t_L g7052 ( 
.A(n_6446),
.Y(n_7052)
);

NOR2xp33_ASAP7_75t_SL g7053 ( 
.A(n_6446),
.B(n_4591),
.Y(n_7053)
);

INVx1_ASAP7_75t_SL g7054 ( 
.A(n_6297),
.Y(n_7054)
);

INVx4_ASAP7_75t_L g7055 ( 
.A(n_5534),
.Y(n_7055)
);

AOI21xp5_ASAP7_75t_SL g7056 ( 
.A1(n_5674),
.A2(n_4457),
.B(n_4395),
.Y(n_7056)
);

INVx1_ASAP7_75t_L g7057 ( 
.A(n_5777),
.Y(n_7057)
);

BUFx2_ASAP7_75t_L g7058 ( 
.A(n_6450),
.Y(n_7058)
);

BUFx2_ASAP7_75t_L g7059 ( 
.A(n_6450),
.Y(n_7059)
);

BUFx6f_ASAP7_75t_L g7060 ( 
.A(n_6417),
.Y(n_7060)
);

BUFx3_ASAP7_75t_L g7061 ( 
.A(n_6446),
.Y(n_7061)
);

BUFx2_ASAP7_75t_L g7062 ( 
.A(n_6450),
.Y(n_7062)
);

NAND2xp5_ASAP7_75t_SL g7063 ( 
.A(n_5525),
.B(n_5212),
.Y(n_7063)
);

INVx4_ASAP7_75t_L g7064 ( 
.A(n_5534),
.Y(n_7064)
);

OAI22xp5_ASAP7_75t_L g7065 ( 
.A1(n_5895),
.A2(n_5208),
.B1(n_5156),
.B2(n_5149),
.Y(n_7065)
);

NAND2xp5_ASAP7_75t_SL g7066 ( 
.A(n_5525),
.B(n_5212),
.Y(n_7066)
);

NAND2xp5_ASAP7_75t_L g7067 ( 
.A(n_6554),
.B(n_4427),
.Y(n_7067)
);

AOI21xp33_ASAP7_75t_L g7068 ( 
.A1(n_5927),
.A2(n_5351),
.B(n_5339),
.Y(n_7068)
);

BUFx3_ASAP7_75t_L g7069 ( 
.A(n_5717),
.Y(n_7069)
);

AOI22xp33_ASAP7_75t_L g7070 ( 
.A1(n_5834),
.A2(n_5454),
.B1(n_5435),
.B2(n_5196),
.Y(n_7070)
);

OAI22xp5_ASAP7_75t_L g7071 ( 
.A1(n_6216),
.A2(n_5208),
.B1(n_5156),
.B2(n_4618),
.Y(n_7071)
);

INVx1_ASAP7_75t_SL g7072 ( 
.A(n_6297),
.Y(n_7072)
);

AOI22xp33_ASAP7_75t_L g7073 ( 
.A1(n_5543),
.A2(n_5454),
.B1(n_5114),
.B2(n_5148),
.Y(n_7073)
);

CKINVDCx11_ASAP7_75t_R g7074 ( 
.A(n_5712),
.Y(n_7074)
);

AOI21xp5_ASAP7_75t_L g7075 ( 
.A1(n_6069),
.A2(n_5208),
.B(n_5351),
.Y(n_7075)
);

NAND2xp5_ASAP7_75t_L g7076 ( 
.A(n_6015),
.B(n_5209),
.Y(n_7076)
);

INVx6_ASAP7_75t_L g7077 ( 
.A(n_6461),
.Y(n_7077)
);

OR2x2_ASAP7_75t_L g7078 ( 
.A(n_6376),
.B(n_4854),
.Y(n_7078)
);

BUFx6f_ASAP7_75t_L g7079 ( 
.A(n_6417),
.Y(n_7079)
);

NAND2xp5_ASAP7_75t_L g7080 ( 
.A(n_6021),
.B(n_4515),
.Y(n_7080)
);

BUFx2_ASAP7_75t_L g7081 ( 
.A(n_6458),
.Y(n_7081)
);

AND2x4_ASAP7_75t_SL g7082 ( 
.A(n_5713),
.B(n_4622),
.Y(n_7082)
);

INVx4_ASAP7_75t_L g7083 ( 
.A(n_5534),
.Y(n_7083)
);

NAND2xp5_ASAP7_75t_L g7084 ( 
.A(n_6021),
.B(n_4515),
.Y(n_7084)
);

BUFx2_ASAP7_75t_L g7085 ( 
.A(n_6458),
.Y(n_7085)
);

BUFx3_ASAP7_75t_L g7086 ( 
.A(n_5717),
.Y(n_7086)
);

BUFx2_ASAP7_75t_L g7087 ( 
.A(n_6458),
.Y(n_7087)
);

AOI22xp33_ASAP7_75t_L g7088 ( 
.A1(n_5543),
.A2(n_5114),
.B1(n_5337),
.B2(n_5308),
.Y(n_7088)
);

HB1xp67_ASAP7_75t_L g7089 ( 
.A(n_5596),
.Y(n_7089)
);

CKINVDCx20_ASAP7_75t_R g7090 ( 
.A(n_6529),
.Y(n_7090)
);

AOI22xp33_ASAP7_75t_SL g7091 ( 
.A1(n_5931),
.A2(n_4457),
.B1(n_4993),
.B2(n_4988),
.Y(n_7091)
);

A2O1A1Ixp33_ASAP7_75t_L g7092 ( 
.A1(n_6125),
.A2(n_5004),
.B(n_5458),
.C(n_5393),
.Y(n_7092)
);

INVx2_ASAP7_75t_SL g7093 ( 
.A(n_5732),
.Y(n_7093)
);

BUFx3_ASAP7_75t_L g7094 ( 
.A(n_5717),
.Y(n_7094)
);

INVx2_ASAP7_75t_SL g7095 ( 
.A(n_5732),
.Y(n_7095)
);

OAI21xp33_ASAP7_75t_L g7096 ( 
.A1(n_5928),
.A2(n_5225),
.B(n_5004),
.Y(n_7096)
);

AOI22xp5_ASAP7_75t_L g7097 ( 
.A1(n_5488),
.A2(n_5252),
.B1(n_4457),
.B2(n_5064),
.Y(n_7097)
);

AND2x6_ASAP7_75t_L g7098 ( 
.A(n_6083),
.B(n_4442),
.Y(n_7098)
);

BUFx2_ASAP7_75t_L g7099 ( 
.A(n_6458),
.Y(n_7099)
);

INVxp67_ASAP7_75t_L g7100 ( 
.A(n_6023),
.Y(n_7100)
);

CKINVDCx20_ASAP7_75t_R g7101 ( 
.A(n_6529),
.Y(n_7101)
);

AO21x1_ASAP7_75t_L g7102 ( 
.A1(n_6100),
.A2(n_5004),
.B(n_5356),
.Y(n_7102)
);

BUFx6f_ASAP7_75t_L g7103 ( 
.A(n_6417),
.Y(n_7103)
);

AOI22xp33_ASAP7_75t_SL g7104 ( 
.A1(n_5931),
.A2(n_4457),
.B1(n_4988),
.B2(n_4390),
.Y(n_7104)
);

AOI221xp5_ASAP7_75t_L g7105 ( 
.A1(n_5885),
.A2(n_5424),
.B1(n_5442),
.B2(n_5379),
.C(n_5360),
.Y(n_7105)
);

OAI22xp5_ASAP7_75t_L g7106 ( 
.A1(n_5888),
.A2(n_4618),
.B1(n_4729),
.B2(n_4591),
.Y(n_7106)
);

AOI221xp5_ASAP7_75t_L g7107 ( 
.A1(n_5885),
.A2(n_5424),
.B1(n_5442),
.B2(n_5379),
.C(n_5360),
.Y(n_7107)
);

CKINVDCx20_ASAP7_75t_R g7108 ( 
.A(n_6132),
.Y(n_7108)
);

AOI22xp33_ASAP7_75t_L g7109 ( 
.A1(n_5488),
.A2(n_5466),
.B1(n_5445),
.B2(n_4481),
.Y(n_7109)
);

AO22x1_ASAP7_75t_L g7110 ( 
.A1(n_6105),
.A2(n_4497),
.B1(n_5365),
.B2(n_4734),
.Y(n_7110)
);

NAND2xp5_ASAP7_75t_L g7111 ( 
.A(n_6150),
.B(n_4427),
.Y(n_7111)
);

OR2x2_ASAP7_75t_L g7112 ( 
.A(n_6376),
.B(n_4854),
.Y(n_7112)
);

CKINVDCx5p33_ASAP7_75t_R g7113 ( 
.A(n_6061),
.Y(n_7113)
);

AOI22xp5_ASAP7_75t_L g7114 ( 
.A1(n_6223),
.A2(n_5252),
.B1(n_4734),
.B2(n_5142),
.Y(n_7114)
);

AND2x2_ASAP7_75t_L g7115 ( 
.A(n_6228),
.B(n_6253),
.Y(n_7115)
);

INVx2_ASAP7_75t_SL g7116 ( 
.A(n_5736),
.Y(n_7116)
);

NAND2xp5_ASAP7_75t_L g7117 ( 
.A(n_5858),
.B(n_4985),
.Y(n_7117)
);

AOI22xp5_ASAP7_75t_L g7118 ( 
.A1(n_6223),
.A2(n_4734),
.B1(n_5142),
.B2(n_4512),
.Y(n_7118)
);

BUFx3_ASAP7_75t_L g7119 ( 
.A(n_5717),
.Y(n_7119)
);

BUFx2_ASAP7_75t_L g7120 ( 
.A(n_6458),
.Y(n_7120)
);

BUFx2_ASAP7_75t_L g7121 ( 
.A(n_6458),
.Y(n_7121)
);

BUFx3_ASAP7_75t_L g7122 ( 
.A(n_5717),
.Y(n_7122)
);

AOI22xp33_ASAP7_75t_L g7123 ( 
.A1(n_6113),
.A2(n_5466),
.B1(n_5445),
.B2(n_4639),
.Y(n_7123)
);

AND2x6_ASAP7_75t_L g7124 ( 
.A(n_6083),
.B(n_4442),
.Y(n_7124)
);

INVxp67_ASAP7_75t_L g7125 ( 
.A(n_6023),
.Y(n_7125)
);

NAND2xp5_ASAP7_75t_L g7126 ( 
.A(n_5858),
.B(n_4985),
.Y(n_7126)
);

BUFx6f_ASAP7_75t_L g7127 ( 
.A(n_6417),
.Y(n_7127)
);

INVx4_ASAP7_75t_L g7128 ( 
.A(n_5534),
.Y(n_7128)
);

OR2x2_ASAP7_75t_L g7129 ( 
.A(n_6376),
.B(n_6242),
.Y(n_7129)
);

NAND2xp5_ASAP7_75t_L g7130 ( 
.A(n_5862),
.B(n_4985),
.Y(n_7130)
);

NAND2xp5_ASAP7_75t_L g7131 ( 
.A(n_5862),
.B(n_4985),
.Y(n_7131)
);

OAI21xp33_ASAP7_75t_L g7132 ( 
.A1(n_5940),
.A2(n_5750),
.B(n_5936),
.Y(n_7132)
);

INVxp67_ASAP7_75t_L g7133 ( 
.A(n_6032),
.Y(n_7133)
);

AOI22xp33_ASAP7_75t_L g7134 ( 
.A1(n_6113),
.A2(n_4905),
.B1(n_4935),
.B2(n_4927),
.Y(n_7134)
);

BUFx12f_ASAP7_75t_L g7135 ( 
.A(n_6538),
.Y(n_7135)
);

INVx3_ASAP7_75t_L g7136 ( 
.A(n_6118),
.Y(n_7136)
);

AOI221xp5_ASAP7_75t_L g7137 ( 
.A1(n_5750),
.A2(n_4963),
.B1(n_5193),
.B2(n_4981),
.C(n_4672),
.Y(n_7137)
);

AND2x4_ASAP7_75t_L g7138 ( 
.A(n_6548),
.B(n_6011),
.Y(n_7138)
);

INVxp67_ASAP7_75t_L g7139 ( 
.A(n_6032),
.Y(n_7139)
);

INVx3_ASAP7_75t_SL g7140 ( 
.A(n_6417),
.Y(n_7140)
);

HB1xp67_ASAP7_75t_L g7141 ( 
.A(n_5596),
.Y(n_7141)
);

INVx5_ASAP7_75t_L g7142 ( 
.A(n_6030),
.Y(n_7142)
);

AOI221xp5_ASAP7_75t_L g7143 ( 
.A1(n_6144),
.A2(n_5193),
.B1(n_4981),
.B2(n_5439),
.C(n_5361),
.Y(n_7143)
);

CKINVDCx20_ASAP7_75t_R g7144 ( 
.A(n_6132),
.Y(n_7144)
);

AOI21xp5_ASAP7_75t_L g7145 ( 
.A1(n_6115),
.A2(n_5458),
.B(n_5393),
.Y(n_7145)
);

BUFx3_ASAP7_75t_L g7146 ( 
.A(n_5717),
.Y(n_7146)
);

A2O1A1Ixp33_ASAP7_75t_L g7147 ( 
.A1(n_6125),
.A2(n_5458),
.B(n_5393),
.C(n_4390),
.Y(n_7147)
);

AO21x1_ASAP7_75t_L g7148 ( 
.A1(n_5954),
.A2(n_5361),
.B(n_5358),
.Y(n_7148)
);

HB1xp67_ASAP7_75t_L g7149 ( 
.A(n_5614),
.Y(n_7149)
);

AOI22xp33_ASAP7_75t_L g7150 ( 
.A1(n_6002),
.A2(n_4442),
.B1(n_4390),
.B2(n_4440),
.Y(n_7150)
);

INVx3_ASAP7_75t_L g7151 ( 
.A(n_6118),
.Y(n_7151)
);

AOI22xp33_ASAP7_75t_L g7152 ( 
.A1(n_6002),
.A2(n_4442),
.B1(n_4390),
.B2(n_4440),
.Y(n_7152)
);

NAND2xp5_ASAP7_75t_L g7153 ( 
.A(n_5584),
.B(n_4990),
.Y(n_7153)
);

INVx2_ASAP7_75t_SL g7154 ( 
.A(n_5625),
.Y(n_7154)
);

INVx3_ASAP7_75t_L g7155 ( 
.A(n_6118),
.Y(n_7155)
);

INVx3_ASAP7_75t_L g7156 ( 
.A(n_6118),
.Y(n_7156)
);

INVx3_ASAP7_75t_L g7157 ( 
.A(n_6118),
.Y(n_7157)
);

A2O1A1Ixp33_ASAP7_75t_L g7158 ( 
.A1(n_5950),
.A2(n_4440),
.B(n_4395),
.C(n_4423),
.Y(n_7158)
);

INVx3_ASAP7_75t_L g7159 ( 
.A(n_6118),
.Y(n_7159)
);

AOI21xp33_ASAP7_75t_L g7160 ( 
.A1(n_5954),
.A2(n_6034),
.B(n_5491),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_L g7161 ( 
.A(n_5584),
.B(n_6000),
.Y(n_7161)
);

BUFx4f_ASAP7_75t_L g7162 ( 
.A(n_5662),
.Y(n_7162)
);

AOI22xp33_ASAP7_75t_L g7163 ( 
.A1(n_5988),
.A2(n_4442),
.B1(n_4440),
.B2(n_4395),
.Y(n_7163)
);

CKINVDCx8_ASAP7_75t_R g7164 ( 
.A(n_5872),
.Y(n_7164)
);

BUFx3_ASAP7_75t_L g7165 ( 
.A(n_5717),
.Y(n_7165)
);

AOI22xp33_ASAP7_75t_L g7166 ( 
.A1(n_5988),
.A2(n_4442),
.B1(n_4395),
.B2(n_4477),
.Y(n_7166)
);

AOI22xp33_ASAP7_75t_L g7167 ( 
.A1(n_5944),
.A2(n_6144),
.B1(n_5740),
.B2(n_5856),
.Y(n_7167)
);

AND2x2_ASAP7_75t_SL g7168 ( 
.A(n_5884),
.B(n_4423),
.Y(n_7168)
);

AOI22xp5_ASAP7_75t_L g7169 ( 
.A1(n_5944),
.A2(n_4512),
.B1(n_5142),
.B2(n_4734),
.Y(n_7169)
);

NAND2xp5_ASAP7_75t_L g7170 ( 
.A(n_6150),
.B(n_4427),
.Y(n_7170)
);

AOI222xp33_ASAP7_75t_L g7171 ( 
.A1(n_5567),
.A2(n_5481),
.B1(n_6224),
.B2(n_6202),
.C1(n_6386),
.C2(n_6155),
.Y(n_7171)
);

NAND2x1p5_ASAP7_75t_L g7172 ( 
.A(n_5884),
.B(n_4591),
.Y(n_7172)
);

AOI21xp5_ASAP7_75t_L g7173 ( 
.A1(n_6115),
.A2(n_4618),
.B(n_4591),
.Y(n_7173)
);

INVx3_ASAP7_75t_L g7174 ( 
.A(n_6118),
.Y(n_7174)
);

HB1xp67_ASAP7_75t_L g7175 ( 
.A(n_5614),
.Y(n_7175)
);

BUFx2_ASAP7_75t_L g7176 ( 
.A(n_6458),
.Y(n_7176)
);

AOI22xp33_ASAP7_75t_L g7177 ( 
.A1(n_5740),
.A2(n_5856),
.B1(n_6089),
.B2(n_5567),
.Y(n_7177)
);

INVx4_ASAP7_75t_L g7178 ( 
.A(n_5534),
.Y(n_7178)
);

INVx3_ASAP7_75t_SL g7179 ( 
.A(n_6464),
.Y(n_7179)
);

NOR2xp33_ASAP7_75t_L g7180 ( 
.A(n_5973),
.B(n_5439),
.Y(n_7180)
);

INVxp67_ASAP7_75t_SL g7181 ( 
.A(n_6207),
.Y(n_7181)
);

NAND2xp5_ASAP7_75t_SL g7182 ( 
.A(n_5973),
.B(n_5212),
.Y(n_7182)
);

AOI22xp33_ASAP7_75t_L g7183 ( 
.A1(n_5856),
.A2(n_4996),
.B1(n_5050),
.B2(n_4477),
.Y(n_7183)
);

INVx5_ASAP7_75t_L g7184 ( 
.A(n_6030),
.Y(n_7184)
);

O2A1O1Ixp5_ASAP7_75t_L g7185 ( 
.A1(n_6034),
.A2(n_4706),
.B(n_4837),
.C(n_4577),
.Y(n_7185)
);

INVx4_ASAP7_75t_L g7186 ( 
.A(n_5536),
.Y(n_7186)
);

NOR2xp33_ASAP7_75t_L g7187 ( 
.A(n_5535),
.B(n_5277),
.Y(n_7187)
);

CKINVDCx20_ASAP7_75t_R g7188 ( 
.A(n_6268),
.Y(n_7188)
);

AOI21xp33_ASAP7_75t_L g7189 ( 
.A1(n_5491),
.A2(n_5362),
.B(n_5358),
.Y(n_7189)
);

BUFx6f_ASAP7_75t_L g7190 ( 
.A(n_6464),
.Y(n_7190)
);

INVx2_ASAP7_75t_SL g7191 ( 
.A(n_5625),
.Y(n_7191)
);

AOI21xp5_ASAP7_75t_L g7192 ( 
.A1(n_6234),
.A2(n_4618),
.B(n_4591),
.Y(n_7192)
);

HB1xp67_ASAP7_75t_L g7193 ( 
.A(n_5640),
.Y(n_7193)
);

NAND2xp33_ASAP7_75t_L g7194 ( 
.A(n_5936),
.B(n_5350),
.Y(n_7194)
);

INVx5_ASAP7_75t_L g7195 ( 
.A(n_6030),
.Y(n_7195)
);

BUFx6f_ASAP7_75t_L g7196 ( 
.A(n_6464),
.Y(n_7196)
);

AOI22xp5_ASAP7_75t_L g7197 ( 
.A1(n_5871),
.A2(n_5142),
.B1(n_4734),
.B2(n_5277),
.Y(n_7197)
);

NOR2x1_ASAP7_75t_L g7198 ( 
.A(n_6110),
.B(n_5411),
.Y(n_7198)
);

BUFx6f_ASAP7_75t_L g7199 ( 
.A(n_6464),
.Y(n_7199)
);

BUFx6f_ASAP7_75t_L g7200 ( 
.A(n_6464),
.Y(n_7200)
);

AOI22xp33_ASAP7_75t_L g7201 ( 
.A1(n_6089),
.A2(n_5626),
.B1(n_6084),
.B2(n_5515),
.Y(n_7201)
);

INVx2_ASAP7_75t_SL g7202 ( 
.A(n_5625),
.Y(n_7202)
);

CKINVDCx11_ASAP7_75t_R g7203 ( 
.A(n_5505),
.Y(n_7203)
);

AND2x2_ASAP7_75t_SL g7204 ( 
.A(n_5884),
.B(n_4423),
.Y(n_7204)
);

OR2x2_ASAP7_75t_L g7205 ( 
.A(n_6376),
.B(n_4499),
.Y(n_7205)
);

CKINVDCx20_ASAP7_75t_R g7206 ( 
.A(n_6268),
.Y(n_7206)
);

AOI21xp5_ASAP7_75t_L g7207 ( 
.A1(n_6263),
.A2(n_4729),
.B(n_4618),
.Y(n_7207)
);

AOI21xp5_ASAP7_75t_L g7208 ( 
.A1(n_6274),
.A2(n_4729),
.B(n_4618),
.Y(n_7208)
);

BUFx6f_ASAP7_75t_L g7209 ( 
.A(n_6464),
.Y(n_7209)
);

OR2x2_ASAP7_75t_L g7210 ( 
.A(n_6376),
.B(n_4499),
.Y(n_7210)
);

NOR2xp33_ASAP7_75t_L g7211 ( 
.A(n_6531),
.B(n_5277),
.Y(n_7211)
);

BUFx8_ASAP7_75t_L g7212 ( 
.A(n_6364),
.Y(n_7212)
);

O2A1O1Ixp33_ASAP7_75t_L g7213 ( 
.A1(n_5803),
.A2(n_5413),
.B(n_5469),
.C(n_4765),
.Y(n_7213)
);

OAI21xp33_ASAP7_75t_L g7214 ( 
.A1(n_6395),
.A2(n_5371),
.B(n_5362),
.Y(n_7214)
);

NAND2xp5_ASAP7_75t_L g7215 ( 
.A(n_6153),
.B(n_4480),
.Y(n_7215)
);

BUFx8_ASAP7_75t_SL g7216 ( 
.A(n_5505),
.Y(n_7216)
);

HB1xp67_ASAP7_75t_L g7217 ( 
.A(n_5640),
.Y(n_7217)
);

AOI21xp5_ASAP7_75t_L g7218 ( 
.A1(n_6274),
.A2(n_4729),
.B(n_4618),
.Y(n_7218)
);

AOI21xp5_ASAP7_75t_L g7219 ( 
.A1(n_6275),
.A2(n_4767),
.B(n_4729),
.Y(n_7219)
);

AOI21xp5_ASAP7_75t_L g7220 ( 
.A1(n_6275),
.A2(n_6354),
.B(n_6209),
.Y(n_7220)
);

INVxp67_ASAP7_75t_L g7221 ( 
.A(n_6351),
.Y(n_7221)
);

HB1xp67_ASAP7_75t_L g7222 ( 
.A(n_5659),
.Y(n_7222)
);

AOI22xp5_ASAP7_75t_L g7223 ( 
.A1(n_5871),
.A2(n_5142),
.B1(n_4734),
.B2(n_5278),
.Y(n_7223)
);

AOI21xp33_ASAP7_75t_L g7224 ( 
.A1(n_5473),
.A2(n_5372),
.B(n_5371),
.Y(n_7224)
);

BUFx2_ASAP7_75t_L g7225 ( 
.A(n_5634),
.Y(n_7225)
);

OR2x6_ASAP7_75t_L g7226 ( 
.A(n_6350),
.B(n_4662),
.Y(n_7226)
);

INVx4_ASAP7_75t_L g7227 ( 
.A(n_5536),
.Y(n_7227)
);

BUFx6f_ASAP7_75t_L g7228 ( 
.A(n_6464),
.Y(n_7228)
);

AOI221xp5_ASAP7_75t_L g7229 ( 
.A1(n_5473),
.A2(n_5372),
.B1(n_5381),
.B2(n_5375),
.C(n_5373),
.Y(n_7229)
);

CKINVDCx11_ASAP7_75t_R g7230 ( 
.A(n_5505),
.Y(n_7230)
);

AOI21xp5_ASAP7_75t_L g7231 ( 
.A1(n_6354),
.A2(n_4767),
.B(n_4729),
.Y(n_7231)
);

AOI222xp33_ASAP7_75t_L g7232 ( 
.A1(n_5481),
.A2(n_4944),
.B1(n_4996),
.B2(n_5081),
.C1(n_5050),
.C2(n_4468),
.Y(n_7232)
);

BUFx8_ASAP7_75t_L g7233 ( 
.A(n_6364),
.Y(n_7233)
);

A2O1A1Ixp33_ASAP7_75t_L g7234 ( 
.A1(n_5950),
.A2(n_4833),
.B(n_4423),
.C(n_5413),
.Y(n_7234)
);

INVx4_ASAP7_75t_L g7235 ( 
.A(n_5536),
.Y(n_7235)
);

INVxp67_ASAP7_75t_SL g7236 ( 
.A(n_6207),
.Y(n_7236)
);

O2A1O1Ixp5_ASAP7_75t_L g7237 ( 
.A1(n_5803),
.A2(n_4706),
.B(n_4837),
.C(n_4577),
.Y(n_7237)
);

AOI21xp5_ASAP7_75t_L g7238 ( 
.A1(n_6209),
.A2(n_4767),
.B(n_4729),
.Y(n_7238)
);

NAND2xp5_ASAP7_75t_L g7239 ( 
.A(n_6047),
.B(n_4992),
.Y(n_7239)
);

BUFx6f_ASAP7_75t_L g7240 ( 
.A(n_6464),
.Y(n_7240)
);

INVxp67_ASAP7_75t_SL g7241 ( 
.A(n_6255),
.Y(n_7241)
);

INVx2_ASAP7_75t_SL g7242 ( 
.A(n_5634),
.Y(n_7242)
);

AOI21xp5_ASAP7_75t_L g7243 ( 
.A1(n_5780),
.A2(n_4767),
.B(n_4729),
.Y(n_7243)
);

NAND2xp33_ASAP7_75t_L g7244 ( 
.A(n_6061),
.B(n_4946),
.Y(n_7244)
);

NAND2x1p5_ASAP7_75t_L g7245 ( 
.A(n_5884),
.B(n_4729),
.Y(n_7245)
);

BUFx6f_ASAP7_75t_L g7246 ( 
.A(n_6468),
.Y(n_7246)
);

BUFx2_ASAP7_75t_L g7247 ( 
.A(n_5634),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_6047),
.B(n_4992),
.Y(n_7248)
);

HB1xp67_ASAP7_75t_L g7249 ( 
.A(n_5659),
.Y(n_7249)
);

OR2x2_ASAP7_75t_L g7250 ( 
.A(n_6376),
.B(n_4499),
.Y(n_7250)
);

AOI221xp5_ASAP7_75t_L g7251 ( 
.A1(n_5986),
.A2(n_5373),
.B1(n_5381),
.B2(n_5375),
.C(n_4765),
.Y(n_7251)
);

INVx2_ASAP7_75t_SL g7252 ( 
.A(n_5645),
.Y(n_7252)
);

NAND2xp5_ASAP7_75t_L g7253 ( 
.A(n_6153),
.B(n_4480),
.Y(n_7253)
);

BUFx2_ASAP7_75t_L g7254 ( 
.A(n_5667),
.Y(n_7254)
);

CKINVDCx6p67_ASAP7_75t_R g7255 ( 
.A(n_6205),
.Y(n_7255)
);

BUFx6f_ASAP7_75t_L g7256 ( 
.A(n_6468),
.Y(n_7256)
);

INVx2_ASAP7_75t_SL g7257 ( 
.A(n_5667),
.Y(n_7257)
);

OAI22xp5_ASAP7_75t_L g7258 ( 
.A1(n_5888),
.A2(n_4767),
.B1(n_4852),
.B2(n_4849),
.Y(n_7258)
);

CKINVDCx5p33_ASAP7_75t_R g7259 ( 
.A(n_6027),
.Y(n_7259)
);

INVx2_ASAP7_75t_SL g7260 ( 
.A(n_5667),
.Y(n_7260)
);

NAND2xp5_ASAP7_75t_L g7261 ( 
.A(n_6053),
.B(n_4992),
.Y(n_7261)
);

INVxp67_ASAP7_75t_SL g7262 ( 
.A(n_6255),
.Y(n_7262)
);

AO21x2_ASAP7_75t_L g7263 ( 
.A1(n_6555),
.A2(n_5051),
.B(n_4780),
.Y(n_7263)
);

BUFx6f_ASAP7_75t_L g7264 ( 
.A(n_6468),
.Y(n_7264)
);

INVx4_ASAP7_75t_L g7265 ( 
.A(n_5536),
.Y(n_7265)
);

INVx4_ASAP7_75t_L g7266 ( 
.A(n_5536),
.Y(n_7266)
);

NAND2xp5_ASAP7_75t_L g7267 ( 
.A(n_6053),
.B(n_4992),
.Y(n_7267)
);

HB1xp67_ASAP7_75t_L g7268 ( 
.A(n_5698),
.Y(n_7268)
);

NAND2xp5_ASAP7_75t_L g7269 ( 
.A(n_6054),
.B(n_4997),
.Y(n_7269)
);

BUFx6f_ASAP7_75t_L g7270 ( 
.A(n_6468),
.Y(n_7270)
);

OR2x2_ASAP7_75t_L g7271 ( 
.A(n_6242),
.B(n_4570),
.Y(n_7271)
);

AOI22xp33_ASAP7_75t_L g7272 ( 
.A1(n_5626),
.A2(n_4996),
.B1(n_5081),
.B2(n_5050),
.Y(n_7272)
);

NAND3xp33_ASAP7_75t_L g7273 ( 
.A(n_5848),
.B(n_5452),
.C(n_5404),
.Y(n_7273)
);

INVx3_ASAP7_75t_SL g7274 ( 
.A(n_6468),
.Y(n_7274)
);

NAND2xp5_ASAP7_75t_L g7275 ( 
.A(n_6159),
.B(n_4480),
.Y(n_7275)
);

BUFx6f_ASAP7_75t_L g7276 ( 
.A(n_6468),
.Y(n_7276)
);

HB1xp67_ASAP7_75t_L g7277 ( 
.A(n_5698),
.Y(n_7277)
);

NAND2xp5_ASAP7_75t_L g7278 ( 
.A(n_6159),
.B(n_4528),
.Y(n_7278)
);

NOR2xp33_ASAP7_75t_L g7279 ( 
.A(n_6531),
.B(n_5278),
.Y(n_7279)
);

BUFx3_ASAP7_75t_L g7280 ( 
.A(n_5717),
.Y(n_7280)
);

CKINVDCx5p33_ASAP7_75t_R g7281 ( 
.A(n_6052),
.Y(n_7281)
);

CKINVDCx8_ASAP7_75t_R g7282 ( 
.A(n_6137),
.Y(n_7282)
);

BUFx3_ASAP7_75t_L g7283 ( 
.A(n_5963),
.Y(n_7283)
);

CKINVDCx5p33_ASAP7_75t_R g7284 ( 
.A(n_5789),
.Y(n_7284)
);

INVx2_ASAP7_75t_SL g7285 ( 
.A(n_5688),
.Y(n_7285)
);

INVx1_ASAP7_75t_SL g7286 ( 
.A(n_6383),
.Y(n_7286)
);

NAND3xp33_ASAP7_75t_L g7287 ( 
.A(n_5799),
.B(n_5404),
.C(n_5397),
.Y(n_7287)
);

OAI22xp33_ASAP7_75t_L g7288 ( 
.A1(n_5871),
.A2(n_4849),
.B1(n_4852),
.B2(n_4767),
.Y(n_7288)
);

AOI21xp5_ASAP7_75t_L g7289 ( 
.A1(n_5780),
.A2(n_4849),
.B(n_4767),
.Y(n_7289)
);

NOR2xp33_ASAP7_75t_L g7290 ( 
.A(n_6485),
.B(n_5278),
.Y(n_7290)
);

AOI21xp5_ASAP7_75t_L g7291 ( 
.A1(n_5826),
.A2(n_4849),
.B(n_4767),
.Y(n_7291)
);

OAI22xp5_ASAP7_75t_L g7292 ( 
.A1(n_5888),
.A2(n_4767),
.B1(n_4852),
.B2(n_4849),
.Y(n_7292)
);

HB1xp67_ASAP7_75t_L g7293 ( 
.A(n_5728),
.Y(n_7293)
);

NAND2xp5_ASAP7_75t_L g7294 ( 
.A(n_6160),
.B(n_4528),
.Y(n_7294)
);

AOI22xp33_ASAP7_75t_SL g7295 ( 
.A1(n_5603),
.A2(n_4734),
.B1(n_5142),
.B2(n_4852),
.Y(n_7295)
);

AOI21xp5_ASAP7_75t_L g7296 ( 
.A1(n_5826),
.A2(n_4852),
.B(n_4849),
.Y(n_7296)
);

AOI21xp5_ASAP7_75t_L g7297 ( 
.A1(n_5838),
.A2(n_4852),
.B(n_4849),
.Y(n_7297)
);

INVx2_ASAP7_75t_SL g7298 ( 
.A(n_5688),
.Y(n_7298)
);

AOI22xp33_ASAP7_75t_L g7299 ( 
.A1(n_6084),
.A2(n_5050),
.B1(n_5081),
.B2(n_4468),
.Y(n_7299)
);

OR2x6_ASAP7_75t_SL g7300 ( 
.A(n_5511),
.B(n_4997),
.Y(n_7300)
);

OR2x2_ASAP7_75t_L g7301 ( 
.A(n_6242),
.B(n_4570),
.Y(n_7301)
);

AND2x2_ASAP7_75t_SL g7302 ( 
.A(n_5884),
.B(n_4833),
.Y(n_7302)
);

AOI22xp33_ASAP7_75t_L g7303 ( 
.A1(n_5515),
.A2(n_5081),
.B1(n_4468),
.B2(n_4734),
.Y(n_7303)
);

NAND2xp5_ASAP7_75t_L g7304 ( 
.A(n_6054),
.B(n_4997),
.Y(n_7304)
);

AOI21xp5_ASAP7_75t_L g7305 ( 
.A1(n_5838),
.A2(n_4852),
.B(n_4849),
.Y(n_7305)
);

O2A1O1Ixp33_ASAP7_75t_L g7306 ( 
.A1(n_5546),
.A2(n_5469),
.B(n_5397),
.C(n_5416),
.Y(n_7306)
);

NAND2xp5_ASAP7_75t_L g7307 ( 
.A(n_6057),
.B(n_4997),
.Y(n_7307)
);

NAND2x1p5_ASAP7_75t_L g7308 ( 
.A(n_5923),
.B(n_4849),
.Y(n_7308)
);

INVx4_ASAP7_75t_L g7309 ( 
.A(n_5536),
.Y(n_7309)
);

AOI21xp5_ASAP7_75t_SL g7310 ( 
.A1(n_5674),
.A2(n_5294),
.B(n_5288),
.Y(n_7310)
);

AOI21xp5_ASAP7_75t_L g7311 ( 
.A1(n_5850),
.A2(n_4866),
.B(n_4852),
.Y(n_7311)
);

CKINVDCx5p33_ASAP7_75t_R g7312 ( 
.A(n_5789),
.Y(n_7312)
);

AOI22xp5_ASAP7_75t_L g7313 ( 
.A1(n_6395),
.A2(n_5142),
.B1(n_4734),
.B2(n_5147),
.Y(n_7313)
);

CKINVDCx6p67_ASAP7_75t_R g7314 ( 
.A(n_6205),
.Y(n_7314)
);

A2O1A1Ixp33_ASAP7_75t_L g7315 ( 
.A1(n_6022),
.A2(n_4833),
.B(n_5294),
.C(n_5288),
.Y(n_7315)
);

NOR2xp67_ASAP7_75t_L g7316 ( 
.A(n_6468),
.B(n_5013),
.Y(n_7316)
);

NAND2xp5_ASAP7_75t_L g7317 ( 
.A(n_6057),
.B(n_6067),
.Y(n_7317)
);

NAND2xp5_ASAP7_75t_L g7318 ( 
.A(n_6067),
.B(n_5002),
.Y(n_7318)
);

NOR2xp33_ASAP7_75t_L g7319 ( 
.A(n_6485),
.B(n_5147),
.Y(n_7319)
);

BUFx6f_ASAP7_75t_L g7320 ( 
.A(n_5572),
.Y(n_7320)
);

NOR2xp67_ASAP7_75t_L g7321 ( 
.A(n_6270),
.B(n_5013),
.Y(n_7321)
);

BUFx6f_ASAP7_75t_L g7322 ( 
.A(n_5572),
.Y(n_7322)
);

INVx2_ASAP7_75t_SL g7323 ( 
.A(n_5688),
.Y(n_7323)
);

NAND2xp5_ASAP7_75t_L g7324 ( 
.A(n_6145),
.B(n_5002),
.Y(n_7324)
);

AOI21xp5_ASAP7_75t_L g7325 ( 
.A1(n_5850),
.A2(n_4866),
.B(n_4852),
.Y(n_7325)
);

NAND2xp5_ASAP7_75t_SL g7326 ( 
.A(n_6310),
.B(n_5212),
.Y(n_7326)
);

BUFx4f_ASAP7_75t_L g7327 ( 
.A(n_5662),
.Y(n_7327)
);

AOI22xp33_ASAP7_75t_L g7328 ( 
.A1(n_5918),
.A2(n_4468),
.B1(n_5142),
.B2(n_4734),
.Y(n_7328)
);

NAND3xp33_ASAP7_75t_L g7329 ( 
.A(n_5799),
.B(n_5516),
.C(n_5503),
.Y(n_7329)
);

INVx5_ASAP7_75t_L g7330 ( 
.A(n_6030),
.Y(n_7330)
);

AOI22xp33_ASAP7_75t_L g7331 ( 
.A1(n_5918),
.A2(n_5142),
.B1(n_4734),
.B2(n_5288),
.Y(n_7331)
);

NAND2xp5_ASAP7_75t_L g7332 ( 
.A(n_6145),
.B(n_5002),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_L g7333 ( 
.A(n_5601),
.B(n_5607),
.Y(n_7333)
);

INVxp67_ASAP7_75t_L g7334 ( 
.A(n_6351),
.Y(n_7334)
);

INVxp67_ASAP7_75t_SL g7335 ( 
.A(n_6229),
.Y(n_7335)
);

NAND2xp5_ASAP7_75t_L g7336 ( 
.A(n_5601),
.B(n_5002),
.Y(n_7336)
);

AOI22xp5_ASAP7_75t_L g7337 ( 
.A1(n_6173),
.A2(n_5142),
.B1(n_5147),
.B2(n_5317),
.Y(n_7337)
);

HB1xp67_ASAP7_75t_L g7338 ( 
.A(n_5728),
.Y(n_7338)
);

AOI22xp5_ASAP7_75t_L g7339 ( 
.A1(n_6173),
.A2(n_5142),
.B1(n_5147),
.B2(n_5317),
.Y(n_7339)
);

OAI21xp33_ASAP7_75t_L g7340 ( 
.A1(n_5799),
.A2(n_4722),
.B(n_4682),
.Y(n_7340)
);

OAI21xp33_ASAP7_75t_L g7341 ( 
.A1(n_5995),
.A2(n_4722),
.B(n_4682),
.Y(n_7341)
);

INVx2_ASAP7_75t_SL g7342 ( 
.A(n_5690),
.Y(n_7342)
);

INVx2_ASAP7_75t_SL g7343 ( 
.A(n_5946),
.Y(n_7343)
);

AND2x2_ASAP7_75t_L g7344 ( 
.A(n_5571),
.B(n_5580),
.Y(n_7344)
);

A2O1A1Ixp33_ASAP7_75t_L g7345 ( 
.A1(n_6022),
.A2(n_4833),
.B(n_5294),
.C(n_5288),
.Y(n_7345)
);

INVx5_ASAP7_75t_L g7346 ( 
.A(n_6030),
.Y(n_7346)
);

OR2x2_ASAP7_75t_L g7347 ( 
.A(n_6242),
.B(n_4589),
.Y(n_7347)
);

BUFx12f_ASAP7_75t_L g7348 ( 
.A(n_5529),
.Y(n_7348)
);

INVx2_ASAP7_75t_SL g7349 ( 
.A(n_5946),
.Y(n_7349)
);

BUFx6f_ASAP7_75t_L g7350 ( 
.A(n_5572),
.Y(n_7350)
);

BUFx12f_ASAP7_75t_L g7351 ( 
.A(n_5529),
.Y(n_7351)
);

CKINVDCx8_ASAP7_75t_R g7352 ( 
.A(n_6137),
.Y(n_7352)
);

NAND2xp33_ASAP7_75t_L g7353 ( 
.A(n_5490),
.B(n_4946),
.Y(n_7353)
);

AOI22xp5_ASAP7_75t_L g7354 ( 
.A1(n_6155),
.A2(n_5147),
.B1(n_5321),
.B2(n_5317),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_L g7355 ( 
.A(n_5607),
.B(n_5003),
.Y(n_7355)
);

AOI22xp33_ASAP7_75t_SL g7356 ( 
.A1(n_5603),
.A2(n_4866),
.B1(n_5028),
.B2(n_4952),
.Y(n_7356)
);

AOI21xp5_ASAP7_75t_L g7357 ( 
.A1(n_5852),
.A2(n_5934),
.B(n_5873),
.Y(n_7357)
);

NOR2xp33_ASAP7_75t_L g7358 ( 
.A(n_5938),
.B(n_5147),
.Y(n_7358)
);

NAND2xp5_ASAP7_75t_L g7359 ( 
.A(n_6071),
.B(n_5003),
.Y(n_7359)
);

NAND2xp5_ASAP7_75t_SL g7360 ( 
.A(n_6310),
.B(n_5231),
.Y(n_7360)
);

AOI22xp5_ASAP7_75t_L g7361 ( 
.A1(n_5672),
.A2(n_5321),
.B1(n_5322),
.B2(n_5317),
.Y(n_7361)
);

INVx4_ASAP7_75t_L g7362 ( 
.A(n_5536),
.Y(n_7362)
);

INVx1_ASAP7_75t_SL g7363 ( 
.A(n_6383),
.Y(n_7363)
);

BUFx6f_ASAP7_75t_L g7364 ( 
.A(n_5572),
.Y(n_7364)
);

BUFx3_ASAP7_75t_L g7365 ( 
.A(n_5963),
.Y(n_7365)
);

CKINVDCx5p33_ASAP7_75t_R g7366 ( 
.A(n_5789),
.Y(n_7366)
);

OAI21xp5_ASAP7_75t_L g7367 ( 
.A1(n_6117),
.A2(n_6308),
.B(n_5503),
.Y(n_7367)
);

HB1xp67_ASAP7_75t_L g7368 ( 
.A(n_5768),
.Y(n_7368)
);

BUFx3_ASAP7_75t_L g7369 ( 
.A(n_5963),
.Y(n_7369)
);

BUFx3_ASAP7_75t_L g7370 ( 
.A(n_5963),
.Y(n_7370)
);

NOR2x1_ASAP7_75t_L g7371 ( 
.A(n_6105),
.B(n_5411),
.Y(n_7371)
);

OAI22xp5_ASAP7_75t_L g7372 ( 
.A1(n_6043),
.A2(n_4866),
.B1(n_5028),
.B2(n_4952),
.Y(n_7372)
);

BUFx2_ASAP7_75t_L g7373 ( 
.A(n_5959),
.Y(n_7373)
);

AOI22xp5_ASAP7_75t_L g7374 ( 
.A1(n_5672),
.A2(n_5321),
.B1(n_5322),
.B2(n_5317),
.Y(n_7374)
);

AOI21xp5_ASAP7_75t_L g7375 ( 
.A1(n_5852),
.A2(n_5934),
.B(n_5873),
.Y(n_7375)
);

NOR2xp33_ASAP7_75t_SL g7376 ( 
.A(n_5662),
.B(n_4866),
.Y(n_7376)
);

A2O1A1Ixp33_ASAP7_75t_L g7377 ( 
.A1(n_6117),
.A2(n_5294),
.B(n_4952),
.C(n_5028),
.Y(n_7377)
);

BUFx3_ASAP7_75t_L g7378 ( 
.A(n_5963),
.Y(n_7378)
);

OR2x2_ASAP7_75t_L g7379 ( 
.A(n_6242),
.B(n_4589),
.Y(n_7379)
);

NOR2xp33_ASAP7_75t_L g7380 ( 
.A(n_5938),
.B(n_4723),
.Y(n_7380)
);

BUFx8_ASAP7_75t_SL g7381 ( 
.A(n_5529),
.Y(n_7381)
);

INVx1_ASAP7_75t_SL g7382 ( 
.A(n_6495),
.Y(n_7382)
);

BUFx2_ASAP7_75t_L g7383 ( 
.A(n_5959),
.Y(n_7383)
);

BUFx2_ASAP7_75t_SL g7384 ( 
.A(n_5963),
.Y(n_7384)
);

BUFx6f_ASAP7_75t_L g7385 ( 
.A(n_5666),
.Y(n_7385)
);

BUFx3_ASAP7_75t_L g7386 ( 
.A(n_5963),
.Y(n_7386)
);

NAND2xp5_ASAP7_75t_L g7387 ( 
.A(n_6160),
.B(n_4528),
.Y(n_7387)
);

INVx2_ASAP7_75t_SL g7388 ( 
.A(n_5946),
.Y(n_7388)
);

AOI21xp33_ASAP7_75t_L g7389 ( 
.A1(n_5546),
.A2(n_4601),
.B(n_4552),
.Y(n_7389)
);

AND2x2_ASAP7_75t_L g7390 ( 
.A(n_6226),
.B(n_4552),
.Y(n_7390)
);

BUFx6f_ASAP7_75t_SL g7391 ( 
.A(n_5713),
.Y(n_7391)
);

OAI22xp5_ASAP7_75t_SL g7392 ( 
.A1(n_6043),
.A2(n_4497),
.B1(n_4952),
.B2(n_4866),
.Y(n_7392)
);

AOI21xp5_ASAP7_75t_L g7393 ( 
.A1(n_5939),
.A2(n_5968),
.B(n_5951),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_6167),
.B(n_4592),
.Y(n_7394)
);

NAND2xp5_ASAP7_75t_L g7395 ( 
.A(n_6167),
.B(n_4592),
.Y(n_7395)
);

INVxp67_ASAP7_75t_SL g7396 ( 
.A(n_6229),
.Y(n_7396)
);

INVx4_ASAP7_75t_SL g7397 ( 
.A(n_5536),
.Y(n_7397)
);

INVx1_ASAP7_75t_SL g7398 ( 
.A(n_6495),
.Y(n_7398)
);

BUFx2_ASAP7_75t_L g7399 ( 
.A(n_5959),
.Y(n_7399)
);

HB1xp67_ASAP7_75t_L g7400 ( 
.A(n_5768),
.Y(n_7400)
);

AND2x2_ASAP7_75t_L g7401 ( 
.A(n_6199),
.B(n_4552),
.Y(n_7401)
);

NAND2xp5_ASAP7_75t_L g7402 ( 
.A(n_6071),
.B(n_5003),
.Y(n_7402)
);

BUFx3_ASAP7_75t_L g7403 ( 
.A(n_5963),
.Y(n_7403)
);

O2A1O1Ixp33_ASAP7_75t_L g7404 ( 
.A1(n_5475),
.A2(n_5416),
.B(n_4497),
.C(n_5453),
.Y(n_7404)
);

OR2x2_ASAP7_75t_L g7405 ( 
.A(n_6306),
.B(n_4597),
.Y(n_7405)
);

HB1xp67_ASAP7_75t_L g7406 ( 
.A(n_5776),
.Y(n_7406)
);

NAND2x1p5_ASAP7_75t_L g7407 ( 
.A(n_5923),
.B(n_4866),
.Y(n_7407)
);

NOR2x1_ASAP7_75t_L g7408 ( 
.A(n_6270),
.B(n_4597),
.Y(n_7408)
);

NAND2xp5_ASAP7_75t_SL g7409 ( 
.A(n_5964),
.B(n_5231),
.Y(n_7409)
);

AOI22xp33_ASAP7_75t_SL g7410 ( 
.A1(n_5603),
.A2(n_4866),
.B1(n_5028),
.B2(n_4952),
.Y(n_7410)
);

INVx2_ASAP7_75t_SL g7411 ( 
.A(n_5946),
.Y(n_7411)
);

BUFx3_ASAP7_75t_L g7412 ( 
.A(n_5975),
.Y(n_7412)
);

INVx1_ASAP7_75t_SL g7413 ( 
.A(n_6530),
.Y(n_7413)
);

INVx2_ASAP7_75t_SL g7414 ( 
.A(n_5946),
.Y(n_7414)
);

OAI22xp5_ASAP7_75t_L g7415 ( 
.A1(n_6095),
.A2(n_6388),
.B1(n_6410),
.B2(n_6331),
.Y(n_7415)
);

BUFx2_ASAP7_75t_L g7416 ( 
.A(n_5959),
.Y(n_7416)
);

NAND2xp5_ASAP7_75t_L g7417 ( 
.A(n_5843),
.B(n_5855),
.Y(n_7417)
);

AOI21xp5_ASAP7_75t_L g7418 ( 
.A1(n_5939),
.A2(n_4952),
.B(n_4866),
.Y(n_7418)
);

NOR2xp33_ASAP7_75t_L g7419 ( 
.A(n_5843),
.B(n_4733),
.Y(n_7419)
);

INVx2_ASAP7_75t_SL g7420 ( 
.A(n_5666),
.Y(n_7420)
);

BUFx6f_ASAP7_75t_L g7421 ( 
.A(n_5666),
.Y(n_7421)
);

BUFx6f_ASAP7_75t_L g7422 ( 
.A(n_5666),
.Y(n_7422)
);

BUFx2_ASAP7_75t_L g7423 ( 
.A(n_5975),
.Y(n_7423)
);

O2A1O1Ixp33_ASAP7_75t_L g7424 ( 
.A1(n_5475),
.A2(n_5453),
.B(n_4945),
.C(n_5113),
.Y(n_7424)
);

NAND2xp5_ASAP7_75t_L g7425 ( 
.A(n_5855),
.B(n_5006),
.Y(n_7425)
);

INVx2_ASAP7_75t_SL g7426 ( 
.A(n_5673),
.Y(n_7426)
);

INVx4_ASAP7_75t_L g7427 ( 
.A(n_5548),
.Y(n_7427)
);

INVx2_ASAP7_75t_SL g7428 ( 
.A(n_5673),
.Y(n_7428)
);

AOI21xp5_ASAP7_75t_L g7429 ( 
.A1(n_5951),
.A2(n_5028),
.B(n_4952),
.Y(n_7429)
);

BUFx3_ASAP7_75t_L g7430 ( 
.A(n_5975),
.Y(n_7430)
);

AOI22xp33_ASAP7_75t_L g7431 ( 
.A1(n_5738),
.A2(n_5317),
.B1(n_5322),
.B2(n_5321),
.Y(n_7431)
);

INVxp67_ASAP7_75t_SL g7432 ( 
.A(n_5819),
.Y(n_7432)
);

CKINVDCx5p33_ASAP7_75t_R g7433 ( 
.A(n_5825),
.Y(n_7433)
);

OAI22xp5_ASAP7_75t_L g7434 ( 
.A1(n_6095),
.A2(n_5028),
.B1(n_4952),
.B2(n_4858),
.Y(n_7434)
);

OR2x2_ASAP7_75t_L g7435 ( 
.A(n_6306),
.B(n_4552),
.Y(n_7435)
);

INVx6_ASAP7_75t_L g7436 ( 
.A(n_6461),
.Y(n_7436)
);

OAI22xp5_ASAP7_75t_L g7437 ( 
.A1(n_6331),
.A2(n_5028),
.B1(n_4952),
.B2(n_4858),
.Y(n_7437)
);

BUFx3_ASAP7_75t_L g7438 ( 
.A(n_5975),
.Y(n_7438)
);

BUFx3_ASAP7_75t_L g7439 ( 
.A(n_5975),
.Y(n_7439)
);

INVx2_ASAP7_75t_SL g7440 ( 
.A(n_5673),
.Y(n_7440)
);

AOI22xp33_ASAP7_75t_L g7441 ( 
.A1(n_5738),
.A2(n_5321),
.B1(n_5366),
.B2(n_5322),
.Y(n_7441)
);

OA21x2_ASAP7_75t_L g7442 ( 
.A1(n_6555),
.A2(n_4780),
.B(n_4779),
.Y(n_7442)
);

INVx2_ASAP7_75t_SL g7443 ( 
.A(n_5673),
.Y(n_7443)
);

NAND2xp5_ASAP7_75t_L g7444 ( 
.A(n_6264),
.B(n_5016),
.Y(n_7444)
);

NAND2xp5_ASAP7_75t_L g7445 ( 
.A(n_6264),
.B(n_5016),
.Y(n_7445)
);

INVx4_ASAP7_75t_L g7446 ( 
.A(n_5548),
.Y(n_7446)
);

NAND2xp5_ASAP7_75t_L g7447 ( 
.A(n_6176),
.B(n_4592),
.Y(n_7447)
);

AOI22xp5_ASAP7_75t_L g7448 ( 
.A1(n_5490),
.A2(n_5322),
.B1(n_5366),
.B2(n_5321),
.Y(n_7448)
);

O2A1O1Ixp33_ASAP7_75t_SL g7449 ( 
.A1(n_5704),
.A2(n_4945),
.B(n_5113),
.C(n_4903),
.Y(n_7449)
);

BUFx6f_ASAP7_75t_L g7450 ( 
.A(n_5739),
.Y(n_7450)
);

AOI21xp5_ASAP7_75t_L g7451 ( 
.A1(n_5968),
.A2(n_5028),
.B(n_5391),
.Y(n_7451)
);

AOI21xp5_ASAP7_75t_L g7452 ( 
.A1(n_5974),
.A2(n_5028),
.B(n_5391),
.Y(n_7452)
);

HB1xp67_ASAP7_75t_L g7453 ( 
.A(n_5776),
.Y(n_7453)
);

AND2x2_ASAP7_75t_L g7454 ( 
.A(n_6265),
.B(n_4552),
.Y(n_7454)
);

BUFx6f_ASAP7_75t_L g7455 ( 
.A(n_5739),
.Y(n_7455)
);

O2A1O1Ixp33_ASAP7_75t_L g7456 ( 
.A1(n_5565),
.A2(n_4945),
.B(n_5113),
.C(n_4903),
.Y(n_7456)
);

OR2x2_ASAP7_75t_L g7457 ( 
.A(n_6306),
.B(n_4552),
.Y(n_7457)
);

AOI22xp33_ASAP7_75t_L g7458 ( 
.A1(n_5550),
.A2(n_5322),
.B1(n_5366),
.B2(n_4598),
.Y(n_7458)
);

BUFx2_ASAP7_75t_L g7459 ( 
.A(n_5975),
.Y(n_7459)
);

NOR2xp33_ASAP7_75t_L g7460 ( 
.A(n_5986),
.B(n_4733),
.Y(n_7460)
);

BUFx12f_ASAP7_75t_L g7461 ( 
.A(n_5646),
.Y(n_7461)
);

BUFx2_ASAP7_75t_L g7462 ( 
.A(n_5975),
.Y(n_7462)
);

BUFx8_ASAP7_75t_L g7463 ( 
.A(n_5548),
.Y(n_7463)
);

BUFx6f_ASAP7_75t_L g7464 ( 
.A(n_5739),
.Y(n_7464)
);

CKINVDCx5p33_ASAP7_75t_R g7465 ( 
.A(n_5825),
.Y(n_7465)
);

BUFx2_ASAP7_75t_L g7466 ( 
.A(n_5975),
.Y(n_7466)
);

CKINVDCx5p33_ASAP7_75t_R g7467 ( 
.A(n_5825),
.Y(n_7467)
);

AOI222xp33_ASAP7_75t_L g7468 ( 
.A1(n_6224),
.A2(n_5105),
.B1(n_5128),
.B2(n_5179),
.C1(n_5055),
.C2(n_4820),
.Y(n_7468)
);

INVx2_ASAP7_75t_SL g7469 ( 
.A(n_5739),
.Y(n_7469)
);

BUFx3_ASAP7_75t_L g7470 ( 
.A(n_5979),
.Y(n_7470)
);

NAND2xp5_ASAP7_75t_L g7471 ( 
.A(n_6176),
.B(n_4628),
.Y(n_7471)
);

AOI21xp5_ASAP7_75t_L g7472 ( 
.A1(n_5974),
.A2(n_5391),
.B(n_4609),
.Y(n_7472)
);

INVxp67_ASAP7_75t_SL g7473 ( 
.A(n_5819),
.Y(n_7473)
);

AOI22xp5_ASAP7_75t_L g7474 ( 
.A1(n_5957),
.A2(n_5366),
.B1(n_5163),
.B2(n_5160),
.Y(n_7474)
);

AND2x2_ASAP7_75t_L g7475 ( 
.A(n_6177),
.B(n_4601),
.Y(n_7475)
);

BUFx3_ASAP7_75t_L g7476 ( 
.A(n_5979),
.Y(n_7476)
);

AOI22xp5_ASAP7_75t_L g7477 ( 
.A1(n_5957),
.A2(n_5366),
.B1(n_5163),
.B2(n_5160),
.Y(n_7477)
);

BUFx2_ASAP7_75t_L g7478 ( 
.A(n_5979),
.Y(n_7478)
);

BUFx6f_ASAP7_75t_SL g7479 ( 
.A(n_5948),
.Y(n_7479)
);

OAI22xp5_ASAP7_75t_L g7480 ( 
.A1(n_6388),
.A2(n_6473),
.B1(n_6551),
.B2(n_6410),
.Y(n_7480)
);

BUFx2_ASAP7_75t_L g7481 ( 
.A(n_5979),
.Y(n_7481)
);

INVx1_ASAP7_75t_SL g7482 ( 
.A(n_6530),
.Y(n_7482)
);

AOI21xp5_ASAP7_75t_L g7483 ( 
.A1(n_5976),
.A2(n_5391),
.B(n_4609),
.Y(n_7483)
);

BUFx12f_ASAP7_75t_L g7484 ( 
.A(n_5646),
.Y(n_7484)
);

BUFx2_ASAP7_75t_L g7485 ( 
.A(n_5979),
.Y(n_7485)
);

NOR2x1_ASAP7_75t_R g7486 ( 
.A(n_6147),
.B(n_5165),
.Y(n_7486)
);

OAI22xp5_ASAP7_75t_L g7487 ( 
.A1(n_6473),
.A2(n_4858),
.B1(n_4896),
.B2(n_4892),
.Y(n_7487)
);

AOI22xp5_ASAP7_75t_L g7488 ( 
.A1(n_6202),
.A2(n_5366),
.B1(n_5163),
.B2(n_5160),
.Y(n_7488)
);

AOI21xp5_ASAP7_75t_L g7489 ( 
.A1(n_5976),
.A2(n_5391),
.B(n_4609),
.Y(n_7489)
);

AOI22xp33_ASAP7_75t_L g7490 ( 
.A1(n_5550),
.A2(n_5633),
.B1(n_6183),
.B2(n_5995),
.Y(n_7490)
);

AOI21xp5_ASAP7_75t_L g7491 ( 
.A1(n_5999),
.A2(n_5391),
.B(n_4609),
.Y(n_7491)
);

BUFx6f_ASAP7_75t_L g7492 ( 
.A(n_5548),
.Y(n_7492)
);

INVx1_ASAP7_75t_SL g7493 ( 
.A(n_5958),
.Y(n_7493)
);

CKINVDCx20_ASAP7_75t_R g7494 ( 
.A(n_6271),
.Y(n_7494)
);

NOR2xp33_ASAP7_75t_L g7495 ( 
.A(n_6204),
.B(n_4739),
.Y(n_7495)
);

INVx5_ASAP7_75t_L g7496 ( 
.A(n_6030),
.Y(n_7496)
);

INVx6_ASAP7_75t_L g7497 ( 
.A(n_6461),
.Y(n_7497)
);

AOI21xp5_ASAP7_75t_L g7498 ( 
.A1(n_5999),
.A2(n_5391),
.B(n_4609),
.Y(n_7498)
);

OAI221xp5_ASAP7_75t_L g7499 ( 
.A1(n_5516),
.A2(n_4837),
.B1(n_4983),
.B2(n_4706),
.C(n_4577),
.Y(n_7499)
);

NAND2xp5_ASAP7_75t_L g7500 ( 
.A(n_5755),
.B(n_5017),
.Y(n_7500)
);

OR2x6_ASAP7_75t_SL g7501 ( 
.A(n_6130),
.B(n_5017),
.Y(n_7501)
);

AOI21xp5_ASAP7_75t_L g7502 ( 
.A1(n_6007),
.A2(n_5391),
.B(n_4609),
.Y(n_7502)
);

BUFx3_ASAP7_75t_L g7503 ( 
.A(n_5979),
.Y(n_7503)
);

OAI22xp5_ASAP7_75t_L g7504 ( 
.A1(n_6551),
.A2(n_4858),
.B1(n_4896),
.B2(n_4892),
.Y(n_7504)
);

INVx4_ASAP7_75t_L g7505 ( 
.A(n_5548),
.Y(n_7505)
);

NAND2xp5_ASAP7_75t_SL g7506 ( 
.A(n_5964),
.B(n_5231),
.Y(n_7506)
);

AOI21xp5_ASAP7_75t_L g7507 ( 
.A1(n_6007),
.A2(n_5391),
.B(n_4609),
.Y(n_7507)
);

OR2x2_ASAP7_75t_L g7508 ( 
.A(n_6306),
.B(n_4601),
.Y(n_7508)
);

NOR2xp33_ASAP7_75t_L g7509 ( 
.A(n_6204),
.B(n_4799),
.Y(n_7509)
);

INVx3_ASAP7_75t_SL g7510 ( 
.A(n_5579),
.Y(n_7510)
);

INVx1_ASAP7_75t_SL g7511 ( 
.A(n_5958),
.Y(n_7511)
);

O2A1O1Ixp5_ASAP7_75t_L g7512 ( 
.A1(n_6081),
.A2(n_4706),
.B(n_4837),
.C(n_4577),
.Y(n_7512)
);

A2O1A1Ixp33_ASAP7_75t_L g7513 ( 
.A1(n_5544),
.A2(n_5476),
.B(n_6129),
.C(n_6257),
.Y(n_7513)
);

AND2x2_ASAP7_75t_L g7514 ( 
.A(n_6199),
.B(n_4601),
.Y(n_7514)
);

INVx2_ASAP7_75t_SL g7515 ( 
.A(n_5587),
.Y(n_7515)
);

BUFx6f_ASAP7_75t_L g7516 ( 
.A(n_5548),
.Y(n_7516)
);

BUFx12f_ASAP7_75t_L g7517 ( 
.A(n_5646),
.Y(n_7517)
);

NAND2xp5_ASAP7_75t_L g7518 ( 
.A(n_5699),
.B(n_5021),
.Y(n_7518)
);

NOR2xp33_ASAP7_75t_L g7519 ( 
.A(n_6230),
.B(n_5417),
.Y(n_7519)
);

AOI22xp5_ASAP7_75t_L g7520 ( 
.A1(n_6183),
.A2(n_5231),
.B1(n_4769),
.B2(n_4598),
.Y(n_7520)
);

CKINVDCx5p33_ASAP7_75t_R g7521 ( 
.A(n_5845),
.Y(n_7521)
);

A2O1A1Ixp33_ASAP7_75t_L g7522 ( 
.A1(n_5544),
.A2(n_5376),
.B(n_4901),
.C(n_4911),
.Y(n_7522)
);

AOI22xp33_ASAP7_75t_L g7523 ( 
.A1(n_5633),
.A2(n_4598),
.B1(n_5417),
.B2(n_4892),
.Y(n_7523)
);

OAI22xp5_ASAP7_75t_L g7524 ( 
.A1(n_6309),
.A2(n_4858),
.B1(n_4896),
.B2(n_4892),
.Y(n_7524)
);

BUFx6f_ASAP7_75t_L g7525 ( 
.A(n_5548),
.Y(n_7525)
);

AND2x4_ASAP7_75t_L g7526 ( 
.A(n_6131),
.B(n_4392),
.Y(n_7526)
);

NOR2x1_ASAP7_75t_R g7527 ( 
.A(n_6188),
.B(n_6189),
.Y(n_7527)
);

AOI21xp5_ASAP7_75t_L g7528 ( 
.A1(n_6291),
.A2(n_4609),
.B(n_4601),
.Y(n_7528)
);

AOI21xp5_ASAP7_75t_L g7529 ( 
.A1(n_6291),
.A2(n_4624),
.B(n_4601),
.Y(n_7529)
);

BUFx6f_ASAP7_75t_L g7530 ( 
.A(n_5548),
.Y(n_7530)
);

AOI21xp5_ASAP7_75t_L g7531 ( 
.A1(n_6302),
.A2(n_4624),
.B(n_4601),
.Y(n_7531)
);

AOI21xp5_ASAP7_75t_L g7532 ( 
.A1(n_6302),
.A2(n_4624),
.B(n_4601),
.Y(n_7532)
);

BUFx2_ASAP7_75t_L g7533 ( 
.A(n_5979),
.Y(n_7533)
);

NAND2xp5_ASAP7_75t_L g7534 ( 
.A(n_6180),
.B(n_4628),
.Y(n_7534)
);

NAND2xp5_ASAP7_75t_L g7535 ( 
.A(n_6180),
.B(n_4628),
.Y(n_7535)
);

AND2x2_ASAP7_75t_L g7536 ( 
.A(n_6212),
.B(n_4624),
.Y(n_7536)
);

NOR2xp33_ASAP7_75t_L g7537 ( 
.A(n_6230),
.B(n_5417),
.Y(n_7537)
);

BUFx6f_ASAP7_75t_L g7538 ( 
.A(n_5557),
.Y(n_7538)
);

BUFx2_ASAP7_75t_L g7539 ( 
.A(n_5979),
.Y(n_7539)
);

AOI22xp33_ASAP7_75t_L g7540 ( 
.A1(n_5761),
.A2(n_4598),
.B1(n_5417),
.B2(n_4892),
.Y(n_7540)
);

AOI22xp33_ASAP7_75t_L g7541 ( 
.A1(n_5761),
.A2(n_4598),
.B1(n_5417),
.B2(n_4892),
.Y(n_7541)
);

CKINVDCx5p33_ASAP7_75t_R g7542 ( 
.A(n_5845),
.Y(n_7542)
);

NOR2xp33_ASAP7_75t_L g7543 ( 
.A(n_6235),
.B(n_5231),
.Y(n_7543)
);

NOR2xp33_ASAP7_75t_L g7544 ( 
.A(n_6235),
.B(n_5231),
.Y(n_7544)
);

AND2x2_ASAP7_75t_L g7545 ( 
.A(n_6212),
.B(n_4624),
.Y(n_7545)
);

AOI21xp5_ASAP7_75t_L g7546 ( 
.A1(n_6305),
.A2(n_4629),
.B(n_4624),
.Y(n_7546)
);

BUFx3_ASAP7_75t_L g7547 ( 
.A(n_5980),
.Y(n_7547)
);

NAND2xp5_ASAP7_75t_L g7548 ( 
.A(n_6387),
.B(n_4645),
.Y(n_7548)
);

BUFx3_ASAP7_75t_L g7549 ( 
.A(n_5980),
.Y(n_7549)
);

HB1xp67_ASAP7_75t_L g7550 ( 
.A(n_5983),
.Y(n_7550)
);

INVx5_ASAP7_75t_L g7551 ( 
.A(n_6312),
.Y(n_7551)
);

BUFx6f_ASAP7_75t_SL g7552 ( 
.A(n_5948),
.Y(n_7552)
);

BUFx6f_ASAP7_75t_L g7553 ( 
.A(n_5557),
.Y(n_7553)
);

BUFx12f_ASAP7_75t_L g7554 ( 
.A(n_5845),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_L g7555 ( 
.A(n_6387),
.B(n_4645),
.Y(n_7555)
);

AOI21xp5_ASAP7_75t_SL g7556 ( 
.A1(n_5704),
.A2(n_5138),
.B(n_4903),
.Y(n_7556)
);

AOI22xp5_ASAP7_75t_L g7557 ( 
.A1(n_5518),
.A2(n_4769),
.B1(n_5179),
.B2(n_4577),
.Y(n_7557)
);

CKINVDCx8_ASAP7_75t_R g7558 ( 
.A(n_6162),
.Y(n_7558)
);

NAND2xp5_ASAP7_75t_L g7559 ( 
.A(n_5699),
.B(n_5021),
.Y(n_7559)
);

BUFx2_ASAP7_75t_L g7560 ( 
.A(n_5980),
.Y(n_7560)
);

INVx2_ASAP7_75t_SL g7561 ( 
.A(n_5587),
.Y(n_7561)
);

OAI22xp5_ASAP7_75t_L g7562 ( 
.A1(n_6309),
.A2(n_4892),
.B1(n_4896),
.B2(n_4858),
.Y(n_7562)
);

AOI21xp5_ASAP7_75t_L g7563 ( 
.A1(n_6305),
.A2(n_4629),
.B(n_4624),
.Y(n_7563)
);

CKINVDCx5p33_ASAP7_75t_R g7564 ( 
.A(n_5849),
.Y(n_7564)
);

BUFx6f_ASAP7_75t_L g7565 ( 
.A(n_5557),
.Y(n_7565)
);

BUFx6f_ASAP7_75t_L g7566 ( 
.A(n_5557),
.Y(n_7566)
);

HB1xp67_ASAP7_75t_L g7567 ( 
.A(n_5983),
.Y(n_7567)
);

INVx2_ASAP7_75t_SL g7568 ( 
.A(n_5587),
.Y(n_7568)
);

BUFx3_ASAP7_75t_L g7569 ( 
.A(n_5980),
.Y(n_7569)
);

INVx5_ASAP7_75t_L g7570 ( 
.A(n_6312),
.Y(n_7570)
);

AND2x2_ASAP7_75t_L g7571 ( 
.A(n_6226),
.B(n_4624),
.Y(n_7571)
);

AOI21xp5_ASAP7_75t_L g7572 ( 
.A1(n_6318),
.A2(n_4694),
.B(n_4629),
.Y(n_7572)
);

AND2x2_ASAP7_75t_L g7573 ( 
.A(n_6226),
.B(n_4629),
.Y(n_7573)
);

OAI22xp5_ASAP7_75t_L g7574 ( 
.A1(n_6386),
.A2(n_4892),
.B1(n_4896),
.B2(n_4858),
.Y(n_7574)
);

AOI22xp5_ASAP7_75t_L g7575 ( 
.A1(n_5518),
.A2(n_4769),
.B1(n_5179),
.B2(n_4837),
.Y(n_7575)
);

AND2x2_ASAP7_75t_L g7576 ( 
.A(n_6265),
.B(n_4629),
.Y(n_7576)
);

AO21x2_ASAP7_75t_L g7577 ( 
.A1(n_6535),
.A2(n_4781),
.B(n_4779),
.Y(n_7577)
);

NAND2x2_ASAP7_75t_L g7578 ( 
.A(n_6225),
.B(n_4843),
.Y(n_7578)
);

INVx1_ASAP7_75t_SL g7579 ( 
.A(n_5958),
.Y(n_7579)
);

INVx2_ASAP7_75t_SL g7580 ( 
.A(n_5587),
.Y(n_7580)
);

HB1xp67_ASAP7_75t_L g7581 ( 
.A(n_5984),
.Y(n_7581)
);

BUFx2_ASAP7_75t_L g7582 ( 
.A(n_5980),
.Y(n_7582)
);

BUFx2_ASAP7_75t_L g7583 ( 
.A(n_5980),
.Y(n_7583)
);

AND2x6_ASAP7_75t_L g7584 ( 
.A(n_6083),
.B(n_4858),
.Y(n_7584)
);

INVx1_ASAP7_75t_SL g7585 ( 
.A(n_5972),
.Y(n_7585)
);

BUFx6f_ASAP7_75t_L g7586 ( 
.A(n_5557),
.Y(n_7586)
);

NAND2xp5_ASAP7_75t_L g7587 ( 
.A(n_5744),
.B(n_5018),
.Y(n_7587)
);

NAND2xp5_ASAP7_75t_L g7588 ( 
.A(n_5744),
.B(n_5018),
.Y(n_7588)
);

NOR2xp33_ASAP7_75t_L g7589 ( 
.A(n_6281),
.B(n_4869),
.Y(n_7589)
);

AND2x2_ASAP7_75t_SL g7590 ( 
.A(n_6068),
.B(n_4896),
.Y(n_7590)
);

NAND2xp5_ASAP7_75t_L g7591 ( 
.A(n_6299),
.B(n_4781),
.Y(n_7591)
);

INVx1_ASAP7_75t_SL g7592 ( 
.A(n_5972),
.Y(n_7592)
);

NOR2xp33_ASAP7_75t_L g7593 ( 
.A(n_6281),
.B(n_4869),
.Y(n_7593)
);

OAI222xp33_ASAP7_75t_L g7594 ( 
.A1(n_5484),
.A2(n_4706),
.B1(n_4983),
.B2(n_4986),
.C1(n_5057),
.C2(n_5136),
.Y(n_7594)
);

NAND2xp5_ASAP7_75t_L g7595 ( 
.A(n_6299),
.B(n_4789),
.Y(n_7595)
);

BUFx8_ASAP7_75t_L g7596 ( 
.A(n_5557),
.Y(n_7596)
);

INVx2_ASAP7_75t_L g7597 ( 
.A(n_6134),
.Y(n_7597)
);

INVx2_ASAP7_75t_L g7598 ( 
.A(n_6171),
.Y(n_7598)
);

NAND2xp5_ASAP7_75t_SL g7599 ( 
.A(n_6094),
.B(n_4896),
.Y(n_7599)
);

CKINVDCx11_ASAP7_75t_R g7600 ( 
.A(n_5849),
.Y(n_7600)
);

AOI21xp5_ASAP7_75t_SL g7601 ( 
.A1(n_5575),
.A2(n_5186),
.B(n_5138),
.Y(n_7601)
);

AND2x4_ASAP7_75t_L g7602 ( 
.A(n_6131),
.B(n_4392),
.Y(n_7602)
);

AOI22xp5_ASAP7_75t_L g7603 ( 
.A1(n_5636),
.A2(n_4769),
.B1(n_4986),
.B2(n_4983),
.Y(n_7603)
);

OR2x2_ASAP7_75t_L g7604 ( 
.A(n_6306),
.B(n_4629),
.Y(n_7604)
);

OAI21x1_ASAP7_75t_SL g7605 ( 
.A1(n_7042),
.A2(n_5821),
.B(n_5823),
.Y(n_7605)
);

INVxp33_ASAP7_75t_SL g7606 ( 
.A(n_7527),
.Y(n_7606)
);

O2A1O1Ixp33_ASAP7_75t_SL g7607 ( 
.A1(n_6611),
.A2(n_6257),
.B(n_6508),
.C(n_6271),
.Y(n_7607)
);

BUFx2_ASAP7_75t_L g7608 ( 
.A(n_6931),
.Y(n_7608)
);

NAND2x1p5_ASAP7_75t_L g7609 ( 
.A(n_6866),
.B(n_5775),
.Y(n_7609)
);

INVx3_ASAP7_75t_L g7610 ( 
.A(n_6927),
.Y(n_7610)
);

OAI21x1_ASAP7_75t_L g7611 ( 
.A1(n_7192),
.A2(n_7208),
.B(n_7207),
.Y(n_7611)
);

INVx1_ASAP7_75t_L g7612 ( 
.A(n_6621),
.Y(n_7612)
);

BUFx3_ASAP7_75t_L g7613 ( 
.A(n_6915),
.Y(n_7613)
);

BUFx6f_ASAP7_75t_L g7614 ( 
.A(n_7025),
.Y(n_7614)
);

NAND2xp5_ASAP7_75t_L g7615 ( 
.A(n_7021),
.B(n_6494),
.Y(n_7615)
);

NAND2x1_ASAP7_75t_L g7616 ( 
.A(n_7310),
.B(n_5980),
.Y(n_7616)
);

BUFx3_ASAP7_75t_L g7617 ( 
.A(n_6915),
.Y(n_7617)
);

INVx2_ASAP7_75t_L g7618 ( 
.A(n_6931),
.Y(n_7618)
);

OA21x2_ASAP7_75t_L g7619 ( 
.A1(n_6936),
.A2(n_7220),
.B(n_7528),
.Y(n_7619)
);

INVx2_ASAP7_75t_L g7620 ( 
.A(n_6931),
.Y(n_7620)
);

OAI21xp5_ASAP7_75t_L g7621 ( 
.A1(n_6702),
.A2(n_6094),
.B(n_6142),
.Y(n_7621)
);

INVx3_ASAP7_75t_L g7622 ( 
.A(n_6927),
.Y(n_7622)
);

AOI22xp5_ASAP7_75t_L g7623 ( 
.A1(n_7132),
.A2(n_6280),
.B1(n_6051),
.B2(n_5943),
.Y(n_7623)
);

INVx1_ASAP7_75t_L g7624 ( 
.A(n_6621),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_6621),
.Y(n_7625)
);

OR2x2_ASAP7_75t_L g7626 ( 
.A(n_6559),
.B(n_6528),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_6622),
.Y(n_7627)
);

AO21x1_ASAP7_75t_L g7628 ( 
.A1(n_6980),
.A2(n_6087),
.B(n_6120),
.Y(n_7628)
);

INVx2_ASAP7_75t_L g7629 ( 
.A(n_6931),
.Y(n_7629)
);

INVx4_ASAP7_75t_L g7630 ( 
.A(n_6692),
.Y(n_7630)
);

AOI22xp33_ASAP7_75t_L g7631 ( 
.A1(n_6637),
.A2(n_7132),
.B1(n_6833),
.B2(n_6702),
.Y(n_7631)
);

INVx3_ASAP7_75t_L g7632 ( 
.A(n_6927),
.Y(n_7632)
);

AOI22xp5_ASAP7_75t_L g7633 ( 
.A1(n_7132),
.A2(n_6637),
.B1(n_6848),
.B2(n_6833),
.Y(n_7633)
);

AOI22xp33_ASAP7_75t_SL g7634 ( 
.A1(n_6702),
.A2(n_5603),
.B1(n_6108),
.B2(n_6068),
.Y(n_7634)
);

INVx1_ASAP7_75t_L g7635 ( 
.A(n_6622),
.Y(n_7635)
);

OAI22xp5_ASAP7_75t_L g7636 ( 
.A1(n_6848),
.A2(n_5943),
.B1(n_6006),
.B2(n_5484),
.Y(n_7636)
);

INVx2_ASAP7_75t_L g7637 ( 
.A(n_6931),
.Y(n_7637)
);

INVx2_ASAP7_75t_L g7638 ( 
.A(n_6931),
.Y(n_7638)
);

INVx2_ASAP7_75t_L g7639 ( 
.A(n_6931),
.Y(n_7639)
);

CKINVDCx8_ASAP7_75t_R g7640 ( 
.A(n_6679),
.Y(n_7640)
);

OAI21xp5_ASAP7_75t_L g7641 ( 
.A1(n_6611),
.A2(n_6142),
.B(n_5694),
.Y(n_7641)
);

AND2x2_ASAP7_75t_L g7642 ( 
.A(n_6580),
.B(n_6583),
.Y(n_7642)
);

BUFx3_ASAP7_75t_L g7643 ( 
.A(n_6915),
.Y(n_7643)
);

OAI21x1_ASAP7_75t_L g7644 ( 
.A1(n_7218),
.A2(n_6353),
.B(n_6460),
.Y(n_7644)
);

OAI21x1_ASAP7_75t_L g7645 ( 
.A1(n_7218),
.A2(n_6353),
.B(n_6460),
.Y(n_7645)
);

CKINVDCx6p67_ASAP7_75t_R g7646 ( 
.A(n_6692),
.Y(n_7646)
);

INVx2_ASAP7_75t_L g7647 ( 
.A(n_6931),
.Y(n_7647)
);

INVx1_ASAP7_75t_L g7648 ( 
.A(n_6622),
.Y(n_7648)
);

NOR2xp33_ASAP7_75t_L g7649 ( 
.A(n_6788),
.B(n_6300),
.Y(n_7649)
);

AOI22xp33_ASAP7_75t_L g7650 ( 
.A1(n_6848),
.A2(n_6006),
.B1(n_5997),
.B2(n_6003),
.Y(n_7650)
);

CKINVDCx8_ASAP7_75t_R g7651 ( 
.A(n_6679),
.Y(n_7651)
);

AOI22xp33_ASAP7_75t_SL g7652 ( 
.A1(n_7038),
.A2(n_5603),
.B1(n_6108),
.B2(n_6068),
.Y(n_7652)
);

NAND2xp33_ASAP7_75t_R g7653 ( 
.A(n_7023),
.B(n_6066),
.Y(n_7653)
);

AO21x2_ASAP7_75t_L g7654 ( 
.A1(n_7148),
.A2(n_6227),
.B(n_6208),
.Y(n_7654)
);

INVx2_ASAP7_75t_L g7655 ( 
.A(n_6931),
.Y(n_7655)
);

INVx1_ASAP7_75t_L g7656 ( 
.A(n_6623),
.Y(n_7656)
);

AO31x2_ASAP7_75t_L g7657 ( 
.A1(n_7148),
.A2(n_7011),
.A3(n_7102),
.B(n_7042),
.Y(n_7657)
);

AO31x2_ASAP7_75t_L g7658 ( 
.A1(n_7148),
.A2(n_6097),
.A3(n_6211),
.B(n_6044),
.Y(n_7658)
);

AND3x1_ASAP7_75t_L g7659 ( 
.A(n_7023),
.B(n_6788),
.C(n_7096),
.Y(n_7659)
);

OAI21x1_ASAP7_75t_L g7660 ( 
.A1(n_7219),
.A2(n_6522),
.B(n_6460),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_6623),
.Y(n_7661)
);

AND2x2_ASAP7_75t_L g7662 ( 
.A(n_6580),
.B(n_6025),
.Y(n_7662)
);

AND2x4_ASAP7_75t_L g7663 ( 
.A(n_7316),
.B(n_5823),
.Y(n_7663)
);

NOR2xp33_ASAP7_75t_L g7664 ( 
.A(n_6954),
.B(n_6300),
.Y(n_7664)
);

AOI22xp33_ASAP7_75t_L g7665 ( 
.A1(n_7040),
.A2(n_5997),
.B1(n_6003),
.B2(n_5591),
.Y(n_7665)
);

AND2x2_ASAP7_75t_L g7666 ( 
.A(n_6580),
.B(n_6025),
.Y(n_7666)
);

INVx1_ASAP7_75t_L g7667 ( 
.A(n_6623),
.Y(n_7667)
);

INVxp67_ASAP7_75t_L g7668 ( 
.A(n_6665),
.Y(n_7668)
);

BUFx2_ASAP7_75t_L g7669 ( 
.A(n_6931),
.Y(n_7669)
);

INVx2_ASAP7_75t_L g7670 ( 
.A(n_6559),
.Y(n_7670)
);

NAND2x1p5_ASAP7_75t_L g7671 ( 
.A(n_6866),
.B(n_5775),
.Y(n_7671)
);

O2A1O1Ixp33_ASAP7_75t_L g7672 ( 
.A1(n_6611),
.A2(n_5565),
.B(n_5575),
.C(n_5545),
.Y(n_7672)
);

AOI21xp5_ASAP7_75t_SL g7673 ( 
.A1(n_6700),
.A2(n_5730),
.B(n_6288),
.Y(n_7673)
);

INVx3_ASAP7_75t_L g7674 ( 
.A(n_6927),
.Y(n_7674)
);

A2O1A1Ixp33_ASAP7_75t_L g7675 ( 
.A1(n_7096),
.A2(n_5476),
.B(n_6129),
.C(n_6120),
.Y(n_7675)
);

OAI21x1_ASAP7_75t_L g7676 ( 
.A1(n_6639),
.A2(n_7483),
.B(n_7472),
.Y(n_7676)
);

BUFx2_ASAP7_75t_L g7677 ( 
.A(n_7501),
.Y(n_7677)
);

AOI22xp33_ASAP7_75t_L g7678 ( 
.A1(n_7040),
.A2(n_5591),
.B1(n_5702),
.B2(n_5641),
.Y(n_7678)
);

INVx2_ASAP7_75t_L g7679 ( 
.A(n_6559),
.Y(n_7679)
);

AOI22xp33_ASAP7_75t_SL g7680 ( 
.A1(n_7038),
.A2(n_5603),
.B1(n_6108),
.B2(n_6068),
.Y(n_7680)
);

NAND3xp33_ASAP7_75t_L g7681 ( 
.A(n_7329),
.B(n_5506),
.C(n_5486),
.Y(n_7681)
);

INVx2_ASAP7_75t_L g7682 ( 
.A(n_6559),
.Y(n_7682)
);

AO21x2_ASAP7_75t_L g7683 ( 
.A1(n_7148),
.A2(n_6227),
.B(n_6208),
.Y(n_7683)
);

NAND2xp5_ASAP7_75t_L g7684 ( 
.A(n_7021),
.B(n_6609),
.Y(n_7684)
);

O2A1O1Ixp33_ASAP7_75t_SL g7685 ( 
.A1(n_6700),
.A2(n_6508),
.B(n_5822),
.C(n_6289),
.Y(n_7685)
);

OA21x2_ASAP7_75t_L g7686 ( 
.A1(n_6936),
.A2(n_7220),
.B(n_7528),
.Y(n_7686)
);

AOI22xp33_ASAP7_75t_L g7687 ( 
.A1(n_7038),
.A2(n_5702),
.B1(n_5641),
.B2(n_5656),
.Y(n_7687)
);

AOI222xp33_ASAP7_75t_L g7688 ( 
.A1(n_6678),
.A2(n_6328),
.B1(n_6339),
.B2(n_6423),
.C1(n_6407),
.C2(n_6295),
.Y(n_7688)
);

NOR2xp33_ASAP7_75t_L g7689 ( 
.A(n_6954),
.B(n_6327),
.Y(n_7689)
);

INVx1_ASAP7_75t_L g7690 ( 
.A(n_6633),
.Y(n_7690)
);

AOI22xp33_ASAP7_75t_L g7691 ( 
.A1(n_7171),
.A2(n_5656),
.B1(n_5636),
.B2(n_5600),
.Y(n_7691)
);

OAI21x1_ASAP7_75t_L g7692 ( 
.A1(n_6639),
.A2(n_6285),
.B(n_6272),
.Y(n_7692)
);

NOR2x1_ASAP7_75t_L g7693 ( 
.A(n_7601),
.B(n_6130),
.Y(n_7693)
);

OAI21x1_ASAP7_75t_L g7694 ( 
.A1(n_6639),
.A2(n_7483),
.B(n_7472),
.Y(n_7694)
);

NOR2xp33_ASAP7_75t_L g7695 ( 
.A(n_7001),
.B(n_6327),
.Y(n_7695)
);

BUFx2_ASAP7_75t_L g7696 ( 
.A(n_7501),
.Y(n_7696)
);

OAI22xp5_ASAP7_75t_L g7697 ( 
.A1(n_7018),
.A2(n_5822),
.B1(n_6108),
.B2(n_5624),
.Y(n_7697)
);

BUFx3_ASAP7_75t_L g7698 ( 
.A(n_6955),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_6633),
.Y(n_7699)
);

AO21x2_ASAP7_75t_L g7700 ( 
.A1(n_6980),
.A2(n_6494),
.B(n_5661),
.Y(n_7700)
);

OAI21x1_ASAP7_75t_L g7701 ( 
.A1(n_7489),
.A2(n_6272),
.B(n_6535),
.Y(n_7701)
);

BUFx2_ASAP7_75t_L g7702 ( 
.A(n_7501),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_6633),
.Y(n_7703)
);

BUFx12f_ASAP7_75t_L g7704 ( 
.A(n_7203),
.Y(n_7704)
);

AOI21xp5_ASAP7_75t_L g7705 ( 
.A1(n_6724),
.A2(n_6391),
.B(n_6390),
.Y(n_7705)
);

AND2x2_ASAP7_75t_L g7706 ( 
.A(n_6583),
.B(n_6044),
.Y(n_7706)
);

AOI21xp5_ASAP7_75t_L g7707 ( 
.A1(n_6724),
.A2(n_6391),
.B(n_6390),
.Y(n_7707)
);

INVx3_ASAP7_75t_L g7708 ( 
.A(n_6927),
.Y(n_7708)
);

OAI21xp5_ASAP7_75t_L g7709 ( 
.A1(n_7513),
.A2(n_5694),
.B(n_6288),
.Y(n_7709)
);

OAI21x1_ASAP7_75t_L g7710 ( 
.A1(n_7489),
.A2(n_6272),
.B(n_6536),
.Y(n_7710)
);

AND2x4_ASAP7_75t_L g7711 ( 
.A(n_7316),
.B(n_6131),
.Y(n_7711)
);

OAI21x1_ASAP7_75t_L g7712 ( 
.A1(n_7491),
.A2(n_6550),
.B(n_6536),
.Y(n_7712)
);

AOI22xp5_ASAP7_75t_L g7713 ( 
.A1(n_7018),
.A2(n_6280),
.B1(n_6051),
.B2(n_5589),
.Y(n_7713)
);

INVx1_ASAP7_75t_L g7714 ( 
.A(n_6650),
.Y(n_7714)
);

NAND2xp5_ASAP7_75t_L g7715 ( 
.A(n_6609),
.B(n_5788),
.Y(n_7715)
);

HB1xp67_ASAP7_75t_L g7716 ( 
.A(n_6557),
.Y(n_7716)
);

AO21x2_ASAP7_75t_L g7717 ( 
.A1(n_7181),
.A2(n_5661),
.B(n_5621),
.Y(n_7717)
);

OAI22xp5_ASAP7_75t_L g7718 ( 
.A1(n_7018),
.A2(n_5624),
.B1(n_6098),
.B2(n_6080),
.Y(n_7718)
);

A2O1A1Ixp33_ASAP7_75t_L g7719 ( 
.A1(n_7096),
.A2(n_6141),
.B(n_6289),
.C(n_5812),
.Y(n_7719)
);

INVx2_ASAP7_75t_SL g7720 ( 
.A(n_7025),
.Y(n_7720)
);

AOI21x1_ASAP7_75t_L g7721 ( 
.A1(n_6574),
.A2(n_5594),
.B(n_6211),
.Y(n_7721)
);

INVx2_ASAP7_75t_L g7722 ( 
.A(n_6562),
.Y(n_7722)
);

OAI21x1_ASAP7_75t_L g7723 ( 
.A1(n_7491),
.A2(n_6550),
.B(n_6500),
.Y(n_7723)
);

OA21x2_ASAP7_75t_L g7724 ( 
.A1(n_7529),
.A2(n_6075),
.B(n_6065),
.Y(n_7724)
);

INVx1_ASAP7_75t_L g7725 ( 
.A(n_6650),
.Y(n_7725)
);

INVx1_ASAP7_75t_L g7726 ( 
.A(n_6650),
.Y(n_7726)
);

HB1xp67_ASAP7_75t_L g7727 ( 
.A(n_6557),
.Y(n_7727)
);

BUFx2_ASAP7_75t_L g7728 ( 
.A(n_7501),
.Y(n_7728)
);

OAI22xp5_ASAP7_75t_L g7729 ( 
.A1(n_6904),
.A2(n_6080),
.B1(n_6124),
.B2(n_6098),
.Y(n_7729)
);

OAI21x1_ASAP7_75t_L g7730 ( 
.A1(n_7498),
.A2(n_6500),
.B(n_6492),
.Y(n_7730)
);

CKINVDCx5p33_ASAP7_75t_R g7731 ( 
.A(n_6802),
.Y(n_7731)
);

OAI21x1_ASAP7_75t_L g7732 ( 
.A1(n_7498),
.A2(n_6492),
.B(n_5670),
.Y(n_7732)
);

NOR2xp33_ASAP7_75t_L g7733 ( 
.A(n_7001),
.B(n_5725),
.Y(n_7733)
);

AND2x2_ASAP7_75t_L g7734 ( 
.A(n_6583),
.B(n_6065),
.Y(n_7734)
);

INVx1_ASAP7_75t_L g7735 ( 
.A(n_6664),
.Y(n_7735)
);

OR2x2_ASAP7_75t_L g7736 ( 
.A(n_6562),
.B(n_6528),
.Y(n_7736)
);

AO21x2_ASAP7_75t_L g7737 ( 
.A1(n_7181),
.A2(n_5621),
.B(n_6081),
.Y(n_7737)
);

OAI21x1_ASAP7_75t_SL g7738 ( 
.A1(n_7042),
.A2(n_5821),
.B(n_5786),
.Y(n_7738)
);

OAI21x1_ASAP7_75t_SL g7739 ( 
.A1(n_7042),
.A2(n_5821),
.B(n_5786),
.Y(n_7739)
);

INVx1_ASAP7_75t_L g7740 ( 
.A(n_6664),
.Y(n_7740)
);

OAI21x1_ASAP7_75t_L g7741 ( 
.A1(n_7502),
.A2(n_5670),
.B(n_5585),
.Y(n_7741)
);

INVx2_ASAP7_75t_L g7742 ( 
.A(n_6562),
.Y(n_7742)
);

INVx1_ASAP7_75t_L g7743 ( 
.A(n_6664),
.Y(n_7743)
);

AND2x4_ASAP7_75t_L g7744 ( 
.A(n_7316),
.B(n_6152),
.Y(n_7744)
);

OAI21x1_ASAP7_75t_L g7745 ( 
.A1(n_7502),
.A2(n_5670),
.B(n_5585),
.Y(n_7745)
);

BUFx2_ASAP7_75t_SL g7746 ( 
.A(n_7558),
.Y(n_7746)
);

OAI21x1_ASAP7_75t_SL g7747 ( 
.A1(n_7102),
.A2(n_5758),
.B(n_5798),
.Y(n_7747)
);

AOI222xp33_ASAP7_75t_L g7748 ( 
.A1(n_6678),
.A2(n_6407),
.B1(n_6328),
.B2(n_6423),
.C1(n_6339),
.C2(n_6295),
.Y(n_7748)
);

A2O1A1Ixp33_ASAP7_75t_L g7749 ( 
.A1(n_7513),
.A2(n_6141),
.B(n_5812),
.C(n_6106),
.Y(n_7749)
);

AO21x2_ASAP7_75t_L g7750 ( 
.A1(n_7236),
.A2(n_6238),
.B(n_6251),
.Y(n_7750)
);

INVx2_ASAP7_75t_L g7751 ( 
.A(n_6562),
.Y(n_7751)
);

AO31x2_ASAP7_75t_L g7752 ( 
.A1(n_7102),
.A2(n_6321),
.A3(n_6501),
.B(n_6238),
.Y(n_7752)
);

OAI21x1_ASAP7_75t_L g7753 ( 
.A1(n_7507),
.A2(n_5783),
.B(n_6445),
.Y(n_7753)
);

INVxp67_ASAP7_75t_L g7754 ( 
.A(n_6665),
.Y(n_7754)
);

INVx2_ASAP7_75t_SL g7755 ( 
.A(n_7025),
.Y(n_7755)
);

AOI21xp33_ASAP7_75t_SL g7756 ( 
.A1(n_6746),
.A2(n_5782),
.B(n_6262),
.Y(n_7756)
);

INVx1_ASAP7_75t_L g7757 ( 
.A(n_6671),
.Y(n_7757)
);

BUFx2_ASAP7_75t_L g7758 ( 
.A(n_6955),
.Y(n_7758)
);

AOI22xp33_ASAP7_75t_L g7759 ( 
.A1(n_7171),
.A2(n_5600),
.B1(n_5590),
.B2(n_5675),
.Y(n_7759)
);

INVx2_ASAP7_75t_L g7760 ( 
.A(n_6563),
.Y(n_7760)
);

INVx6_ASAP7_75t_L g7761 ( 
.A(n_7015),
.Y(n_7761)
);

HB1xp67_ASAP7_75t_L g7762 ( 
.A(n_6612),
.Y(n_7762)
);

AOI221xp5_ASAP7_75t_L g7763 ( 
.A1(n_7480),
.A2(n_6484),
.B1(n_6489),
.B2(n_6444),
.C(n_6436),
.Y(n_7763)
);

NOR2xp33_ASAP7_75t_SL g7764 ( 
.A(n_6866),
.B(n_5497),
.Y(n_7764)
);

AOI22xp5_ASAP7_75t_L g7765 ( 
.A1(n_7194),
.A2(n_5589),
.B1(n_6124),
.B2(n_5655),
.Y(n_7765)
);

NAND2xp5_ASAP7_75t_L g7766 ( 
.A(n_6609),
.B(n_5788),
.Y(n_7766)
);

INVx2_ASAP7_75t_SL g7767 ( 
.A(n_7025),
.Y(n_7767)
);

OAI21x1_ASAP7_75t_L g7768 ( 
.A1(n_7507),
.A2(n_5783),
.B(n_6445),
.Y(n_7768)
);

OR2x6_ASAP7_75t_L g7769 ( 
.A(n_6837),
.B(n_6399),
.Y(n_7769)
);

BUFx2_ASAP7_75t_SL g7770 ( 
.A(n_7558),
.Y(n_7770)
);

AO21x1_ASAP7_75t_L g7771 ( 
.A1(n_7236),
.A2(n_6087),
.B(n_5749),
.Y(n_7771)
);

NAND2x1p5_ASAP7_75t_L g7772 ( 
.A(n_6866),
.B(n_5775),
.Y(n_7772)
);

INVx1_ASAP7_75t_L g7773 ( 
.A(n_6671),
.Y(n_7773)
);

INVx1_ASAP7_75t_L g7774 ( 
.A(n_6671),
.Y(n_7774)
);

OAI21x1_ASAP7_75t_L g7775 ( 
.A1(n_7238),
.A2(n_6872),
.B(n_6845),
.Y(n_7775)
);

NAND2xp5_ASAP7_75t_L g7776 ( 
.A(n_6771),
.B(n_5788),
.Y(n_7776)
);

AND2x4_ASAP7_75t_L g7777 ( 
.A(n_6946),
.B(n_6152),
.Y(n_7777)
);

AOI22xp33_ASAP7_75t_SL g7778 ( 
.A1(n_6866),
.A2(n_5961),
.B1(n_6083),
.B2(n_6262),
.Y(n_7778)
);

OAI21x1_ASAP7_75t_SL g7779 ( 
.A1(n_7102),
.A2(n_5758),
.B(n_5798),
.Y(n_7779)
);

OAI21x1_ASAP7_75t_L g7780 ( 
.A1(n_7238),
.A2(n_5783),
.B(n_6445),
.Y(n_7780)
);

AO31x2_ASAP7_75t_L g7781 ( 
.A1(n_7012),
.A2(n_6501),
.A3(n_6408),
.B(n_6251),
.Y(n_7781)
);

AND2x2_ASAP7_75t_L g7782 ( 
.A(n_6593),
.B(n_5790),
.Y(n_7782)
);

AOI21xp5_ASAP7_75t_L g7783 ( 
.A1(n_6731),
.A2(n_6419),
.B(n_6402),
.Y(n_7783)
);

INVx3_ASAP7_75t_L g7784 ( 
.A(n_6927),
.Y(n_7784)
);

INVx1_ASAP7_75t_L g7785 ( 
.A(n_6683),
.Y(n_7785)
);

AOI21x1_ASAP7_75t_L g7786 ( 
.A1(n_6574),
.A2(n_5594),
.B(n_6411),
.Y(n_7786)
);

AND2x4_ASAP7_75t_L g7787 ( 
.A(n_6946),
.B(n_6152),
.Y(n_7787)
);

INVx3_ASAP7_75t_SL g7788 ( 
.A(n_6893),
.Y(n_7788)
);

AND2x4_ASAP7_75t_L g7789 ( 
.A(n_6946),
.B(n_6152),
.Y(n_7789)
);

OAI21xp5_ASAP7_75t_L g7790 ( 
.A1(n_7329),
.A2(n_5533),
.B(n_5730),
.Y(n_7790)
);

OAI21x1_ASAP7_75t_L g7791 ( 
.A1(n_6845),
.A2(n_6462),
.B(n_5606),
.Y(n_7791)
);

OAI21x1_ASAP7_75t_SL g7792 ( 
.A1(n_6947),
.A2(n_5749),
.B(n_5514),
.Y(n_7792)
);

CKINVDCx16_ASAP7_75t_R g7793 ( 
.A(n_6692),
.Y(n_7793)
);

AND2x4_ASAP7_75t_L g7794 ( 
.A(n_6946),
.B(n_7022),
.Y(n_7794)
);

NAND2xp5_ASAP7_75t_L g7795 ( 
.A(n_6771),
.B(n_6402),
.Y(n_7795)
);

INVx1_ASAP7_75t_L g7796 ( 
.A(n_6683),
.Y(n_7796)
);

NAND2xp5_ASAP7_75t_L g7797 ( 
.A(n_6771),
.B(n_6419),
.Y(n_7797)
);

OR2x6_ASAP7_75t_L g7798 ( 
.A(n_6837),
.B(n_6399),
.Y(n_7798)
);

OAI22xp5_ASAP7_75t_L g7799 ( 
.A1(n_6904),
.A2(n_5558),
.B1(n_5635),
.B2(n_5507),
.Y(n_7799)
);

AO21x2_ASAP7_75t_L g7800 ( 
.A1(n_7160),
.A2(n_6418),
.B(n_6374),
.Y(n_7800)
);

OAI21x1_ASAP7_75t_L g7801 ( 
.A1(n_6845),
.A2(n_6462),
.B(n_5606),
.Y(n_7801)
);

AO21x1_ASAP7_75t_L g7802 ( 
.A1(n_6852),
.A2(n_6269),
.B(n_5726),
.Y(n_7802)
);

BUFx12f_ASAP7_75t_L g7803 ( 
.A(n_7203),
.Y(n_7803)
);

OA21x2_ASAP7_75t_L g7804 ( 
.A1(n_7529),
.A2(n_7532),
.B(n_7531),
.Y(n_7804)
);

INVx2_ASAP7_75t_L g7805 ( 
.A(n_6563),
.Y(n_7805)
);

INVx1_ASAP7_75t_L g7806 ( 
.A(n_6683),
.Y(n_7806)
);

OAI21x1_ASAP7_75t_L g7807 ( 
.A1(n_6845),
.A2(n_6462),
.B(n_5615),
.Y(n_7807)
);

AOI22xp33_ASAP7_75t_L g7808 ( 
.A1(n_7171),
.A2(n_5590),
.B1(n_5675),
.B2(n_5745),
.Y(n_7808)
);

AOI21xp33_ASAP7_75t_L g7809 ( 
.A1(n_7329),
.A2(n_5990),
.B(n_5508),
.Y(n_7809)
);

OAI21x1_ASAP7_75t_L g7810 ( 
.A1(n_6872),
.A2(n_5598),
.B(n_6269),
.Y(n_7810)
);

OR2x6_ASAP7_75t_L g7811 ( 
.A(n_6837),
.B(n_6399),
.Y(n_7811)
);

OAI21xp5_ASAP7_75t_L g7812 ( 
.A1(n_6731),
.A2(n_5533),
.B(n_6408),
.Y(n_7812)
);

OAI21xp5_ASAP7_75t_L g7813 ( 
.A1(n_7367),
.A2(n_5708),
.B(n_5710),
.Y(n_7813)
);

BUFx6f_ASAP7_75t_L g7814 ( 
.A(n_7025),
.Y(n_7814)
);

A2O1A1Ixp33_ASAP7_75t_L g7815 ( 
.A1(n_7194),
.A2(n_5650),
.B(n_6282),
.C(n_6360),
.Y(n_7815)
);

OAI21x1_ASAP7_75t_L g7816 ( 
.A1(n_6872),
.A2(n_5796),
.B(n_5771),
.Y(n_7816)
);

OAI21x1_ASAP7_75t_L g7817 ( 
.A1(n_7451),
.A2(n_5796),
.B(n_5771),
.Y(n_7817)
);

OAI21x1_ASAP7_75t_L g7818 ( 
.A1(n_7451),
.A2(n_5814),
.B(n_5802),
.Y(n_7818)
);

NOR2xp33_ASAP7_75t_SL g7819 ( 
.A(n_7282),
.B(n_7352),
.Y(n_7819)
);

INVx1_ASAP7_75t_L g7820 ( 
.A(n_6578),
.Y(n_7820)
);

A2O1A1Ixp33_ASAP7_75t_L g7821 ( 
.A1(n_7367),
.A2(n_5650),
.B(n_6282),
.C(n_6258),
.Y(n_7821)
);

AOI22xp5_ASAP7_75t_L g7822 ( 
.A1(n_6678),
.A2(n_6827),
.B1(n_6904),
.B2(n_6588),
.Y(n_7822)
);

AO21x2_ASAP7_75t_L g7823 ( 
.A1(n_7160),
.A2(n_6418),
.B(n_6374),
.Y(n_7823)
);

INVx1_ASAP7_75t_L g7824 ( 
.A(n_6578),
.Y(n_7824)
);

NAND2x1p5_ASAP7_75t_L g7825 ( 
.A(n_6916),
.B(n_5775),
.Y(n_7825)
);

AOI21xp5_ASAP7_75t_L g7826 ( 
.A1(n_7367),
.A2(n_6426),
.B(n_6425),
.Y(n_7826)
);

OAI21x1_ASAP7_75t_L g7827 ( 
.A1(n_7452),
.A2(n_5814),
.B(n_5802),
.Y(n_7827)
);

BUFx2_ASAP7_75t_SL g7828 ( 
.A(n_7558),
.Y(n_7828)
);

OAI21x1_ASAP7_75t_SL g7829 ( 
.A1(n_6947),
.A2(n_5514),
.B(n_5990),
.Y(n_7829)
);

INVx1_ASAP7_75t_L g7830 ( 
.A(n_6578),
.Y(n_7830)
);

AND2x4_ASAP7_75t_SL g7831 ( 
.A(n_6940),
.B(n_5948),
.Y(n_7831)
);

AO21x2_ASAP7_75t_L g7832 ( 
.A1(n_7160),
.A2(n_6426),
.B(n_6425),
.Y(n_7832)
);

OAI21x1_ASAP7_75t_L g7833 ( 
.A1(n_7452),
.A2(n_5820),
.B(n_6491),
.Y(n_7833)
);

AOI21xp5_ASAP7_75t_L g7834 ( 
.A1(n_6672),
.A2(n_6478),
.B(n_6452),
.Y(n_7834)
);

OAI22xp33_ASAP7_75t_L g7835 ( 
.A1(n_6561),
.A2(n_5507),
.B1(n_5497),
.B2(n_5743),
.Y(n_7835)
);

OAI21x1_ASAP7_75t_L g7836 ( 
.A1(n_7173),
.A2(n_5820),
.B(n_6491),
.Y(n_7836)
);

INVxp67_ASAP7_75t_SL g7837 ( 
.A(n_7321),
.Y(n_7837)
);

XNOR2xp5_ASAP7_75t_L g7838 ( 
.A(n_7108),
.B(n_6436),
.Y(n_7838)
);

NAND2xp5_ASAP7_75t_L g7839 ( 
.A(n_6791),
.B(n_6452),
.Y(n_7839)
);

AND2x4_ASAP7_75t_L g7840 ( 
.A(n_6946),
.B(n_6152),
.Y(n_7840)
);

OAI21x1_ASAP7_75t_SL g7841 ( 
.A1(n_7213),
.A2(n_5514),
.B(n_5708),
.Y(n_7841)
);

OA21x2_ASAP7_75t_L g7842 ( 
.A1(n_7531),
.A2(n_6324),
.B(n_6478),
.Y(n_7842)
);

OA21x2_ASAP7_75t_L g7843 ( 
.A1(n_7532),
.A2(n_6324),
.B(n_5682),
.Y(n_7843)
);

NOR2xp67_ASAP7_75t_L g7844 ( 
.A(n_7022),
.B(n_5531),
.Y(n_7844)
);

INVx2_ASAP7_75t_SL g7845 ( 
.A(n_7025),
.Y(n_7845)
);

INVx1_ASAP7_75t_L g7846 ( 
.A(n_6584),
.Y(n_7846)
);

AO221x2_ASAP7_75t_L g7847 ( 
.A1(n_6615),
.A2(n_5555),
.B1(n_6501),
.B2(n_5678),
.C(n_6484),
.Y(n_7847)
);

INVx1_ASAP7_75t_L g7848 ( 
.A(n_6584),
.Y(n_7848)
);

OR2x2_ASAP7_75t_L g7849 ( 
.A(n_6563),
.B(n_6537),
.Y(n_7849)
);

INVx1_ASAP7_75t_L g7850 ( 
.A(n_6584),
.Y(n_7850)
);

INVx1_ASAP7_75t_L g7851 ( 
.A(n_6589),
.Y(n_7851)
);

OA21x2_ASAP7_75t_L g7852 ( 
.A1(n_7546),
.A2(n_5682),
.B(n_6431),
.Y(n_7852)
);

INVx2_ASAP7_75t_L g7853 ( 
.A(n_6563),
.Y(n_7853)
);

INVx1_ASAP7_75t_L g7854 ( 
.A(n_6589),
.Y(n_7854)
);

AOI22xp5_ASAP7_75t_L g7855 ( 
.A1(n_6827),
.A2(n_5655),
.B1(n_5664),
.B2(n_5651),
.Y(n_7855)
);

OAI21xp5_ASAP7_75t_L g7856 ( 
.A1(n_6926),
.A2(n_5731),
.B(n_5710),
.Y(n_7856)
);

INVx2_ASAP7_75t_SL g7857 ( 
.A(n_7025),
.Y(n_7857)
);

OAI22xp5_ASAP7_75t_L g7858 ( 
.A1(n_6797),
.A2(n_6798),
.B1(n_6561),
.B2(n_6778),
.Y(n_7858)
);

OAI21xp5_ASAP7_75t_L g7859 ( 
.A1(n_6926),
.A2(n_7167),
.B(n_7201),
.Y(n_7859)
);

AND2x4_ASAP7_75t_L g7860 ( 
.A(n_6946),
.B(n_6169),
.Y(n_7860)
);

AOI22xp33_ASAP7_75t_L g7861 ( 
.A1(n_7415),
.A2(n_5748),
.B1(n_5753),
.B2(n_5745),
.Y(n_7861)
);

AOI221x1_ASAP7_75t_L g7862 ( 
.A1(n_7068),
.A2(n_5555),
.B1(n_5545),
.B2(n_5751),
.C(n_5729),
.Y(n_7862)
);

OA21x2_ASAP7_75t_L g7863 ( 
.A1(n_7546),
.A2(n_6437),
.B(n_6431),
.Y(n_7863)
);

NOR2x1_ASAP7_75t_SL g7864 ( 
.A(n_6942),
.B(n_5551),
.Y(n_7864)
);

OAI21xp5_ASAP7_75t_L g7865 ( 
.A1(n_6926),
.A2(n_5731),
.B(n_5631),
.Y(n_7865)
);

NAND2xp5_ASAP7_75t_L g7866 ( 
.A(n_6791),
.B(n_6466),
.Y(n_7866)
);

BUFx10_ASAP7_75t_L g7867 ( 
.A(n_6828),
.Y(n_7867)
);

OR2x2_ASAP7_75t_L g7868 ( 
.A(n_6567),
.B(n_6537),
.Y(n_7868)
);

BUFx3_ASAP7_75t_L g7869 ( 
.A(n_6955),
.Y(n_7869)
);

HB1xp67_ASAP7_75t_L g7870 ( 
.A(n_6612),
.Y(n_7870)
);

INVx2_ASAP7_75t_L g7871 ( 
.A(n_6567),
.Y(n_7871)
);

INVx6_ASAP7_75t_SL g7872 ( 
.A(n_6565),
.Y(n_7872)
);

INVx1_ASAP7_75t_L g7873 ( 
.A(n_6589),
.Y(n_7873)
);

OAI21x1_ASAP7_75t_SL g7874 ( 
.A1(n_7213),
.A2(n_6283),
.B(n_6258),
.Y(n_7874)
);

AND2x2_ASAP7_75t_L g7875 ( 
.A(n_6593),
.B(n_5790),
.Y(n_7875)
);

AO21x2_ASAP7_75t_L g7876 ( 
.A1(n_6775),
.A2(n_5508),
.B(n_5495),
.Y(n_7876)
);

INVx2_ASAP7_75t_L g7877 ( 
.A(n_6567),
.Y(n_7877)
);

INVx1_ASAP7_75t_L g7878 ( 
.A(n_6594),
.Y(n_7878)
);

O2A1O1Ixp33_ASAP7_75t_SL g7879 ( 
.A1(n_7090),
.A2(n_5779),
.B(n_5805),
.C(n_5756),
.Y(n_7879)
);

INVx1_ASAP7_75t_L g7880 ( 
.A(n_6594),
.Y(n_7880)
);

NAND2x1p5_ASAP7_75t_L g7881 ( 
.A(n_6916),
.B(n_5775),
.Y(n_7881)
);

INVx3_ASAP7_75t_L g7882 ( 
.A(n_7025),
.Y(n_7882)
);

INVx1_ASAP7_75t_L g7883 ( 
.A(n_6594),
.Y(n_7883)
);

O2A1O1Ixp5_ASAP7_75t_L g7884 ( 
.A1(n_7036),
.A2(n_6443),
.B(n_6487),
.C(n_6437),
.Y(n_7884)
);

INVx2_ASAP7_75t_L g7885 ( 
.A(n_6567),
.Y(n_7885)
);

OR2x2_ASAP7_75t_L g7886 ( 
.A(n_6571),
.B(n_6466),
.Y(n_7886)
);

INVx1_ASAP7_75t_L g7887 ( 
.A(n_6613),
.Y(n_7887)
);

OAI21x1_ASAP7_75t_L g7888 ( 
.A1(n_7563),
.A2(n_5492),
.B(n_6206),
.Y(n_7888)
);

BUFx6f_ASAP7_75t_L g7889 ( 
.A(n_7025),
.Y(n_7889)
);

OAI221xp5_ASAP7_75t_L g7890 ( 
.A1(n_7201),
.A2(n_5486),
.B1(n_5558),
.B2(n_5635),
.C(n_5566),
.Y(n_7890)
);

INVx1_ASAP7_75t_L g7891 ( 
.A(n_6613),
.Y(n_7891)
);

AND2x2_ASAP7_75t_L g7892 ( 
.A(n_6593),
.B(n_5790),
.Y(n_7892)
);

INVx1_ASAP7_75t_L g7893 ( 
.A(n_6613),
.Y(n_7893)
);

BUFx6f_ASAP7_75t_L g7894 ( 
.A(n_7047),
.Y(n_7894)
);

AO21x2_ASAP7_75t_L g7895 ( 
.A1(n_6775),
.A2(n_5495),
.B(n_6443),
.Y(n_7895)
);

INVx1_ASAP7_75t_L g7896 ( 
.A(n_6618),
.Y(n_7896)
);

INVx2_ASAP7_75t_L g7897 ( 
.A(n_6571),
.Y(n_7897)
);

AND2x4_ASAP7_75t_L g7898 ( 
.A(n_6946),
.B(n_6169),
.Y(n_7898)
);

OAI21x1_ASAP7_75t_L g7899 ( 
.A1(n_7563),
.A2(n_6330),
.B(n_6206),
.Y(n_7899)
);

AND2x2_ASAP7_75t_L g7900 ( 
.A(n_6667),
.B(n_5801),
.Y(n_7900)
);

AND2x2_ASAP7_75t_L g7901 ( 
.A(n_6667),
.B(n_6669),
.Y(n_7901)
);

BUFx3_ASAP7_75t_L g7902 ( 
.A(n_6692),
.Y(n_7902)
);

OAI21x1_ASAP7_75t_L g7903 ( 
.A1(n_7572),
.A2(n_6330),
.B(n_6206),
.Y(n_7903)
);

INVx2_ASAP7_75t_L g7904 ( 
.A(n_6571),
.Y(n_7904)
);

OAI21xp5_ASAP7_75t_L g7905 ( 
.A1(n_7167),
.A2(n_5631),
.B(n_5756),
.Y(n_7905)
);

OA21x2_ASAP7_75t_L g7906 ( 
.A1(n_7572),
.A2(n_6488),
.B(n_6487),
.Y(n_7906)
);

AOI21xp33_ASAP7_75t_L g7907 ( 
.A1(n_7415),
.A2(n_6037),
.B(n_6010),
.Y(n_7907)
);

NOR2xp67_ASAP7_75t_L g7908 ( 
.A(n_7022),
.B(n_5531),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_6618),
.Y(n_7909)
);

INVx1_ASAP7_75t_L g7910 ( 
.A(n_6618),
.Y(n_7910)
);

AND2x2_ASAP7_75t_L g7911 ( 
.A(n_6667),
.B(n_5801),
.Y(n_7911)
);

OAI21x1_ASAP7_75t_L g7912 ( 
.A1(n_7231),
.A2(n_6330),
.B(n_6122),
.Y(n_7912)
);

INVx2_ASAP7_75t_L g7913 ( 
.A(n_6571),
.Y(n_7913)
);

AOI21xp5_ASAP7_75t_L g7914 ( 
.A1(n_6672),
.A2(n_6164),
.B(n_6312),
.Y(n_7914)
);

INVx1_ASAP7_75t_L g7915 ( 
.A(n_6670),
.Y(n_7915)
);

AND2x4_ASAP7_75t_L g7916 ( 
.A(n_6946),
.B(n_6169),
.Y(n_7916)
);

INVx1_ASAP7_75t_L g7917 ( 
.A(n_6670),
.Y(n_7917)
);

INVx2_ASAP7_75t_SL g7918 ( 
.A(n_7047),
.Y(n_7918)
);

INVxp67_ASAP7_75t_SL g7919 ( 
.A(n_7321),
.Y(n_7919)
);

OAI21x1_ASAP7_75t_L g7920 ( 
.A1(n_7231),
.A2(n_6330),
.B(n_6122),
.Y(n_7920)
);

NAND2xp5_ASAP7_75t_L g7921 ( 
.A(n_6791),
.B(n_6475),
.Y(n_7921)
);

AND2x4_ASAP7_75t_L g7922 ( 
.A(n_7022),
.B(n_6169),
.Y(n_7922)
);

AOI22xp33_ASAP7_75t_L g7923 ( 
.A1(n_7415),
.A2(n_5748),
.B1(n_5753),
.B2(n_6148),
.Y(n_7923)
);

AND2x4_ASAP7_75t_L g7924 ( 
.A(n_7022),
.B(n_6169),
.Y(n_7924)
);

AND2x4_ASAP7_75t_L g7925 ( 
.A(n_7022),
.B(n_6201),
.Y(n_7925)
);

AOI21xp5_ASAP7_75t_L g7926 ( 
.A1(n_6689),
.A2(n_6659),
.B(n_6852),
.Y(n_7926)
);

OAI21x1_ASAP7_75t_L g7927 ( 
.A1(n_7243),
.A2(n_5830),
.B(n_5759),
.Y(n_7927)
);

INVx1_ASAP7_75t_L g7928 ( 
.A(n_6722),
.Y(n_7928)
);

INVx1_ASAP7_75t_L g7929 ( 
.A(n_6722),
.Y(n_7929)
);

OA21x2_ASAP7_75t_L g7930 ( 
.A1(n_7357),
.A2(n_6533),
.B(n_6488),
.Y(n_7930)
);

AOI22xp33_ASAP7_75t_L g7931 ( 
.A1(n_7490),
.A2(n_6151),
.B1(n_6154),
.B2(n_6148),
.Y(n_7931)
);

OAI21x1_ASAP7_75t_L g7932 ( 
.A1(n_7243),
.A2(n_7291),
.B(n_7289),
.Y(n_7932)
);

INVx2_ASAP7_75t_L g7933 ( 
.A(n_6579),
.Y(n_7933)
);

INVx1_ASAP7_75t_L g7934 ( 
.A(n_6741),
.Y(n_7934)
);

INVx1_ASAP7_75t_L g7935 ( 
.A(n_6741),
.Y(n_7935)
);

BUFx2_ASAP7_75t_L g7936 ( 
.A(n_7584),
.Y(n_7936)
);

OAI21x1_ASAP7_75t_L g7937 ( 
.A1(n_7289),
.A2(n_5830),
.B(n_5759),
.Y(n_7937)
);

AOI22xp33_ASAP7_75t_SL g7938 ( 
.A1(n_6852),
.A2(n_6867),
.B1(n_6660),
.B2(n_6588),
.Y(n_7938)
);

AND2x4_ASAP7_75t_L g7939 ( 
.A(n_7022),
.B(n_6201),
.Y(n_7939)
);

AND2x2_ASAP7_75t_L g7940 ( 
.A(n_6669),
.B(n_5801),
.Y(n_7940)
);

OA21x2_ASAP7_75t_L g7941 ( 
.A1(n_7357),
.A2(n_6533),
.B(n_5828),
.Y(n_7941)
);

NAND2x1p5_ASAP7_75t_L g7942 ( 
.A(n_6916),
.B(n_5775),
.Y(n_7942)
);

BUFx3_ASAP7_75t_L g7943 ( 
.A(n_6705),
.Y(n_7943)
);

AND2x4_ASAP7_75t_L g7944 ( 
.A(n_7022),
.B(n_6201),
.Y(n_7944)
);

INVx2_ASAP7_75t_L g7945 ( 
.A(n_7597),
.Y(n_7945)
);

INVx2_ASAP7_75t_L g7946 ( 
.A(n_7597),
.Y(n_7946)
);

OAI21x1_ASAP7_75t_L g7947 ( 
.A1(n_7291),
.A2(n_5754),
.B(n_5747),
.Y(n_7947)
);

OAI21x1_ASAP7_75t_L g7948 ( 
.A1(n_7296),
.A2(n_5754),
.B(n_5747),
.Y(n_7948)
);

NAND2x1p5_ASAP7_75t_L g7949 ( 
.A(n_6916),
.B(n_5775),
.Y(n_7949)
);

NAND2xp5_ASAP7_75t_L g7950 ( 
.A(n_6898),
.B(n_6475),
.Y(n_7950)
);

OA21x2_ASAP7_75t_L g7951 ( 
.A1(n_7375),
.A2(n_5828),
.B(n_5808),
.Y(n_7951)
);

OAI211xp5_ASAP7_75t_SL g7952 ( 
.A1(n_6824),
.A2(n_6195),
.B(n_6213),
.C(n_6010),
.Y(n_7952)
);

INVx3_ASAP7_75t_L g7953 ( 
.A(n_7047),
.Y(n_7953)
);

HB1xp67_ASAP7_75t_L g7954 ( 
.A(n_6766),
.Y(n_7954)
);

OAI21x1_ASAP7_75t_L g7955 ( 
.A1(n_7296),
.A2(n_7305),
.B(n_7297),
.Y(n_7955)
);

INVx2_ASAP7_75t_SL g7956 ( 
.A(n_7047),
.Y(n_7956)
);

INVx1_ASAP7_75t_L g7957 ( 
.A(n_6766),
.Y(n_7957)
);

AND2x4_ASAP7_75t_L g7958 ( 
.A(n_7022),
.B(n_6201),
.Y(n_7958)
);

AND2x2_ASAP7_75t_L g7959 ( 
.A(n_6669),
.B(n_5808),
.Y(n_7959)
);

AOI21xp33_ASAP7_75t_SL g7960 ( 
.A1(n_6746),
.A2(n_6377),
.B(n_5807),
.Y(n_7960)
);

OAI21x1_ASAP7_75t_L g7961 ( 
.A1(n_7297),
.A2(n_5577),
.B(n_5746),
.Y(n_7961)
);

AOI22xp33_ASAP7_75t_L g7962 ( 
.A1(n_7490),
.A2(n_6154),
.B1(n_6161),
.B2(n_6151),
.Y(n_7962)
);

AO21x2_ASAP7_75t_L g7963 ( 
.A1(n_7389),
.A2(n_5581),
.B(n_6172),
.Y(n_7963)
);

AOI221x1_ASAP7_75t_L g7964 ( 
.A1(n_7068),
.A2(n_5555),
.B1(n_5751),
.B2(n_5729),
.C(n_5779),
.Y(n_7964)
);

INVx1_ASAP7_75t_L g7965 ( 
.A(n_6773),
.Y(n_7965)
);

OR2x2_ASAP7_75t_L g7966 ( 
.A(n_6560),
.B(n_6483),
.Y(n_7966)
);

AO31x2_ASAP7_75t_L g7967 ( 
.A1(n_7012),
.A2(n_6490),
.A3(n_6502),
.B(n_6394),
.Y(n_7967)
);

OA21x2_ASAP7_75t_L g7968 ( 
.A1(n_7375),
.A2(n_5828),
.B(n_5808),
.Y(n_7968)
);

OR2x6_ASAP7_75t_L g7969 ( 
.A(n_6565),
.B(n_6668),
.Y(n_7969)
);

O2A1O1Ixp33_ASAP7_75t_L g7970 ( 
.A1(n_6754),
.A2(n_5899),
.B(n_5707),
.C(n_5651),
.Y(n_7970)
);

OAI21x1_ASAP7_75t_L g7971 ( 
.A1(n_7305),
.A2(n_7325),
.B(n_7311),
.Y(n_7971)
);

INVx3_ASAP7_75t_L g7972 ( 
.A(n_7047),
.Y(n_7972)
);

INVx2_ASAP7_75t_L g7973 ( 
.A(n_6579),
.Y(n_7973)
);

BUFx3_ASAP7_75t_L g7974 ( 
.A(n_6705),
.Y(n_7974)
);

INVx2_ASAP7_75t_L g7975 ( 
.A(n_6579),
.Y(n_7975)
);

INVx1_ASAP7_75t_L g7976 ( 
.A(n_6773),
.Y(n_7976)
);

BUFx2_ASAP7_75t_R g7977 ( 
.A(n_7216),
.Y(n_7977)
);

AND2x2_ASAP7_75t_L g7978 ( 
.A(n_6748),
.B(n_5853),
.Y(n_7978)
);

AO21x2_ASAP7_75t_L g7979 ( 
.A1(n_7389),
.A2(n_5581),
.B(n_6172),
.Y(n_7979)
);

OA21x2_ASAP7_75t_L g7980 ( 
.A1(n_7393),
.A2(n_5857),
.B(n_5853),
.Y(n_7980)
);

O2A1O1Ixp33_ASAP7_75t_L g7981 ( 
.A1(n_6754),
.A2(n_5899),
.B(n_5707),
.C(n_5664),
.Y(n_7981)
);

INVx2_ASAP7_75t_L g7982 ( 
.A(n_6579),
.Y(n_7982)
);

OAI21x1_ASAP7_75t_L g7983 ( 
.A1(n_7311),
.A2(n_5577),
.B(n_5746),
.Y(n_7983)
);

OAI22xp33_ASAP7_75t_L g7984 ( 
.A1(n_6561),
.A2(n_5743),
.B1(n_6377),
.B2(n_5686),
.Y(n_7984)
);

INVx1_ASAP7_75t_SL g7985 ( 
.A(n_7286),
.Y(n_7985)
);

BUFx3_ASAP7_75t_L g7986 ( 
.A(n_6705),
.Y(n_7986)
);

OA21x2_ASAP7_75t_L g7987 ( 
.A1(n_7393),
.A2(n_5857),
.B(n_5853),
.Y(n_7987)
);

AND2x2_ASAP7_75t_L g7988 ( 
.A(n_6748),
.B(n_5857),
.Y(n_7988)
);

AOI21xp5_ASAP7_75t_L g7989 ( 
.A1(n_6689),
.A2(n_6164),
.B(n_6312),
.Y(n_7989)
);

INVx2_ASAP7_75t_L g7990 ( 
.A(n_7597),
.Y(n_7990)
);

OA21x2_ASAP7_75t_L g7991 ( 
.A1(n_6825),
.A2(n_5887),
.B(n_5880),
.Y(n_7991)
);

INVx1_ASAP7_75t_L g7992 ( 
.A(n_6786),
.Y(n_7992)
);

OAI21x1_ASAP7_75t_SL g7993 ( 
.A1(n_6797),
.A2(n_6283),
.B(n_6304),
.Y(n_7993)
);

OAI21x1_ASAP7_75t_L g7994 ( 
.A1(n_7325),
.A2(n_5577),
.B(n_5746),
.Y(n_7994)
);

OAI21x1_ASAP7_75t_L g7995 ( 
.A1(n_7418),
.A2(n_5577),
.B(n_5746),
.Y(n_7995)
);

INVx1_ASAP7_75t_L g7996 ( 
.A(n_6786),
.Y(n_7996)
);

INVx1_ASAP7_75t_L g7997 ( 
.A(n_6813),
.Y(n_7997)
);

OR2x2_ASAP7_75t_L g7998 ( 
.A(n_6560),
.B(n_6483),
.Y(n_7998)
);

NOR2xp33_ASAP7_75t_L g7999 ( 
.A(n_7020),
.B(n_5725),
.Y(n_7999)
);

OAI21x1_ASAP7_75t_L g8000 ( 
.A1(n_7418),
.A2(n_6004),
.B(n_5969),
.Y(n_8000)
);

INVx1_ASAP7_75t_L g8001 ( 
.A(n_6813),
.Y(n_8001)
);

OR2x6_ASAP7_75t_L g8002 ( 
.A(n_6565),
.B(n_6399),
.Y(n_8002)
);

AOI22xp33_ASAP7_75t_SL g8003 ( 
.A1(n_6867),
.A2(n_6444),
.B1(n_6505),
.B2(n_6489),
.Y(n_8003)
);

AOI21x1_ASAP7_75t_L g8004 ( 
.A1(n_6574),
.A2(n_6411),
.B(n_5859),
.Y(n_8004)
);

AOI22xp33_ASAP7_75t_L g8005 ( 
.A1(n_6739),
.A2(n_6178),
.B1(n_6179),
.B2(n_6161),
.Y(n_8005)
);

AO31x2_ASAP7_75t_L g8006 ( 
.A1(n_7012),
.A2(n_6490),
.A3(n_6502),
.B(n_6394),
.Y(n_8006)
);

OAI21x1_ASAP7_75t_L g8007 ( 
.A1(n_7429),
.A2(n_6004),
.B(n_5969),
.Y(n_8007)
);

INVx1_ASAP7_75t_L g8008 ( 
.A(n_6819),
.Y(n_8008)
);

OAI21xp33_ASAP7_75t_SL g8009 ( 
.A1(n_6596),
.A2(n_6479),
.B(n_5793),
.Y(n_8009)
);

BUFx2_ASAP7_75t_L g8010 ( 
.A(n_7584),
.Y(n_8010)
);

OA21x2_ASAP7_75t_L g8011 ( 
.A1(n_6825),
.A2(n_6864),
.B(n_6569),
.Y(n_8011)
);

AO21x2_ASAP7_75t_L g8012 ( 
.A1(n_7389),
.A2(n_6239),
.B(n_6220),
.Y(n_8012)
);

BUFx2_ASAP7_75t_SL g8013 ( 
.A(n_7558),
.Y(n_8013)
);

OAI22xp33_ASAP7_75t_L g8014 ( 
.A1(n_6797),
.A2(n_5686),
.B1(n_5722),
.B2(n_6085),
.Y(n_8014)
);

AOI21xp5_ASAP7_75t_L g8015 ( 
.A1(n_6659),
.A2(n_6164),
.B(n_6312),
.Y(n_8015)
);

NAND2xp5_ASAP7_75t_L g8016 ( 
.A(n_6898),
.B(n_6532),
.Y(n_8016)
);

NOR2xp67_ASAP7_75t_L g8017 ( 
.A(n_7022),
.B(n_5531),
.Y(n_8017)
);

NOR2xp33_ASAP7_75t_SL g8018 ( 
.A(n_7282),
.B(n_5859),
.Y(n_8018)
);

AOI21xp5_ASAP7_75t_L g8019 ( 
.A1(n_6867),
.A2(n_6164),
.B(n_6312),
.Y(n_8019)
);

BUFx6f_ASAP7_75t_L g8020 ( 
.A(n_7047),
.Y(n_8020)
);

CKINVDCx9p33_ASAP7_75t_R g8021 ( 
.A(n_7180),
.Y(n_8021)
);

INVx1_ASAP7_75t_SL g8022 ( 
.A(n_7286),
.Y(n_8022)
);

INVx2_ASAP7_75t_SL g8023 ( 
.A(n_7047),
.Y(n_8023)
);

AOI22xp33_ASAP7_75t_L g8024 ( 
.A1(n_6739),
.A2(n_6179),
.B1(n_6267),
.B2(n_6178),
.Y(n_8024)
);

INVx1_ASAP7_75t_L g8025 ( 
.A(n_6819),
.Y(n_8025)
);

CKINVDCx11_ASAP7_75t_R g8026 ( 
.A(n_6603),
.Y(n_8026)
);

INVx2_ASAP7_75t_L g8027 ( 
.A(n_6582),
.Y(n_8027)
);

INVx1_ASAP7_75t_L g8028 ( 
.A(n_6884),
.Y(n_8028)
);

OR2x2_ASAP7_75t_L g8029 ( 
.A(n_6560),
.B(n_6532),
.Y(n_8029)
);

NAND2x1p5_ASAP7_75t_L g8030 ( 
.A(n_6916),
.B(n_5775),
.Y(n_8030)
);

OR2x6_ASAP7_75t_L g8031 ( 
.A(n_6565),
.B(n_6433),
.Y(n_8031)
);

INVx2_ASAP7_75t_L g8032 ( 
.A(n_7597),
.Y(n_8032)
);

NAND2xp5_ASAP7_75t_L g8033 ( 
.A(n_6898),
.B(n_5767),
.Y(n_8033)
);

INVx1_ASAP7_75t_L g8034 ( 
.A(n_6884),
.Y(n_8034)
);

NAND2xp5_ASAP7_75t_L g8035 ( 
.A(n_6920),
.B(n_5767),
.Y(n_8035)
);

INVx2_ASAP7_75t_L g8036 ( 
.A(n_7598),
.Y(n_8036)
);

INVx2_ASAP7_75t_L g8037 ( 
.A(n_7598),
.Y(n_8037)
);

INVx2_ASAP7_75t_L g8038 ( 
.A(n_7598),
.Y(n_8038)
);

A2O1A1Ixp33_ASAP7_75t_L g8039 ( 
.A1(n_6798),
.A2(n_6282),
.B(n_6323),
.C(n_6304),
.Y(n_8039)
);

INVx1_ASAP7_75t_L g8040 ( 
.A(n_6907),
.Y(n_8040)
);

INVx2_ASAP7_75t_L g8041 ( 
.A(n_7598),
.Y(n_8041)
);

INVx4_ASAP7_75t_L g8042 ( 
.A(n_6705),
.Y(n_8042)
);

NAND2x1p5_ASAP7_75t_L g8043 ( 
.A(n_6916),
.B(n_5923),
.Y(n_8043)
);

O2A1O1Ixp33_ASAP7_75t_L g8044 ( 
.A1(n_7480),
.A2(n_5899),
.B(n_5687),
.C(n_5805),
.Y(n_8044)
);

INVx1_ASAP7_75t_L g8045 ( 
.A(n_6907),
.Y(n_8045)
);

NAND2xp5_ASAP7_75t_L g8046 ( 
.A(n_6920),
.B(n_5839),
.Y(n_8046)
);

OAI21xp5_ASAP7_75t_L g8047 ( 
.A1(n_6749),
.A2(n_5678),
.B(n_6323),
.Y(n_8047)
);

INVx1_ASAP7_75t_L g8048 ( 
.A(n_6978),
.Y(n_8048)
);

OAI21xp5_ASAP7_75t_L g8049 ( 
.A1(n_6749),
.A2(n_6360),
.B(n_6355),
.Y(n_8049)
);

AO21x2_ASAP7_75t_L g8050 ( 
.A1(n_7000),
.A2(n_6239),
.B(n_6220),
.Y(n_8050)
);

INVx6_ASAP7_75t_L g8051 ( 
.A(n_7015),
.Y(n_8051)
);

BUFx10_ASAP7_75t_L g8052 ( 
.A(n_6828),
.Y(n_8052)
);

NOR2x1_ASAP7_75t_SL g8053 ( 
.A(n_6942),
.B(n_6959),
.Y(n_8053)
);

OAI21x1_ASAP7_75t_SL g8054 ( 
.A1(n_6798),
.A2(n_6366),
.B(n_6355),
.Y(n_8054)
);

AOI221xp5_ASAP7_75t_SL g8055 ( 
.A1(n_7480),
.A2(n_6510),
.B1(n_6505),
.B2(n_6553),
.C(n_6372),
.Y(n_8055)
);

INVx2_ASAP7_75t_L g8056 ( 
.A(n_6582),
.Y(n_8056)
);

AOI21x1_ASAP7_75t_L g8057 ( 
.A1(n_6600),
.A2(n_6486),
.B(n_6292),
.Y(n_8057)
);

HB1xp67_ASAP7_75t_L g8058 ( 
.A(n_6978),
.Y(n_8058)
);

INVx2_ASAP7_75t_L g8059 ( 
.A(n_6582),
.Y(n_8059)
);

A2O1A1Ixp33_ASAP7_75t_L g8060 ( 
.A1(n_6832),
.A2(n_6372),
.B(n_6396),
.C(n_6366),
.Y(n_8060)
);

INVx1_ASAP7_75t_L g8061 ( 
.A(n_7089),
.Y(n_8061)
);

INVx2_ASAP7_75t_L g8062 ( 
.A(n_6582),
.Y(n_8062)
);

OAI21x1_ASAP7_75t_L g8063 ( 
.A1(n_7026),
.A2(n_7075),
.B(n_7185),
.Y(n_8063)
);

OAI21x1_ASAP7_75t_L g8064 ( 
.A1(n_7185),
.A2(n_6036),
.B(n_5719),
.Y(n_8064)
);

NAND2xp5_ASAP7_75t_L g8065 ( 
.A(n_6920),
.B(n_5839),
.Y(n_8065)
);

NAND2x1p5_ASAP7_75t_L g8066 ( 
.A(n_6916),
.B(n_5923),
.Y(n_8066)
);

INVx1_ASAP7_75t_L g8067 ( 
.A(n_7089),
.Y(n_8067)
);

AO21x2_ASAP7_75t_L g8068 ( 
.A1(n_7000),
.A2(n_6451),
.B(n_4790),
.Y(n_8068)
);

OA21x2_ASAP7_75t_L g8069 ( 
.A1(n_6569),
.A2(n_5887),
.B(n_5880),
.Y(n_8069)
);

AND2x2_ASAP7_75t_L g8070 ( 
.A(n_6748),
.B(n_5880),
.Y(n_8070)
);

INVx1_ASAP7_75t_L g8071 ( 
.A(n_7141),
.Y(n_8071)
);

AND2x2_ASAP7_75t_L g8072 ( 
.A(n_6763),
.B(n_5887),
.Y(n_8072)
);

INVx2_ASAP7_75t_L g8073 ( 
.A(n_6598),
.Y(n_8073)
);

INVx2_ASAP7_75t_L g8074 ( 
.A(n_6598),
.Y(n_8074)
);

AO21x2_ASAP7_75t_L g8075 ( 
.A1(n_7000),
.A2(n_6451),
.B(n_4790),
.Y(n_8075)
);

NOR2xp67_ASAP7_75t_L g8076 ( 
.A(n_7142),
.B(n_7184),
.Y(n_8076)
);

INVx2_ASAP7_75t_L g8077 ( 
.A(n_6598),
.Y(n_8077)
);

NOR2xp33_ASAP7_75t_SL g8078 ( 
.A(n_7282),
.B(n_6486),
.Y(n_8078)
);

OAI21x1_ASAP7_75t_L g8079 ( 
.A1(n_6625),
.A2(n_6076),
.B(n_6019),
.Y(n_8079)
);

OAI21x1_ASAP7_75t_L g8080 ( 
.A1(n_6625),
.A2(n_6076),
.B(n_6019),
.Y(n_8080)
);

AOI21xp5_ASAP7_75t_L g8081 ( 
.A1(n_7377),
.A2(n_6164),
.B(n_6312),
.Y(n_8081)
);

OAI21xp5_ASAP7_75t_L g8082 ( 
.A1(n_6749),
.A2(n_6414),
.B(n_6396),
.Y(n_8082)
);

NOR2xp33_ASAP7_75t_L g8083 ( 
.A(n_7020),
.B(n_5726),
.Y(n_8083)
);

AOI22xp33_ASAP7_75t_L g8084 ( 
.A1(n_6778),
.A2(n_6267),
.B1(n_6371),
.B2(n_6325),
.Y(n_8084)
);

INVx1_ASAP7_75t_L g8085 ( 
.A(n_7141),
.Y(n_8085)
);

NOR2xp33_ASAP7_75t_L g8086 ( 
.A(n_7029),
.B(n_6139),
.Y(n_8086)
);

INVx2_ASAP7_75t_L g8087 ( 
.A(n_6598),
.Y(n_8087)
);

OAI21xp5_ASAP7_75t_L g8088 ( 
.A1(n_7177),
.A2(n_6424),
.B(n_6414),
.Y(n_8088)
);

INVx2_ASAP7_75t_L g8089 ( 
.A(n_6620),
.Y(n_8089)
);

INVx2_ASAP7_75t_L g8090 ( 
.A(n_6620),
.Y(n_8090)
);

A2O1A1Ixp33_ASAP7_75t_L g8091 ( 
.A1(n_6832),
.A2(n_6424),
.B(n_6514),
.C(n_6509),
.Y(n_8091)
);

INVx1_ASAP7_75t_L g8092 ( 
.A(n_7149),
.Y(n_8092)
);

OAI21x1_ASAP7_75t_L g8093 ( 
.A1(n_6625),
.A2(n_6076),
.B(n_6019),
.Y(n_8093)
);

AND2x2_ASAP7_75t_L g8094 ( 
.A(n_6763),
.B(n_5916),
.Y(n_8094)
);

INVx2_ASAP7_75t_L g8095 ( 
.A(n_6620),
.Y(n_8095)
);

AOI21xp5_ASAP7_75t_L g8096 ( 
.A1(n_7377),
.A2(n_6164),
.B(n_6496),
.Y(n_8096)
);

INVx1_ASAP7_75t_L g8097 ( 
.A(n_7149),
.Y(n_8097)
);

AND2x2_ASAP7_75t_L g8098 ( 
.A(n_6763),
.B(n_5916),
.Y(n_8098)
);

OAI21x1_ASAP7_75t_L g8099 ( 
.A1(n_6625),
.A2(n_6104),
.B(n_6076),
.Y(n_8099)
);

OAI21x1_ASAP7_75t_L g8100 ( 
.A1(n_6682),
.A2(n_6104),
.B(n_6076),
.Y(n_8100)
);

INVx1_ASAP7_75t_L g8101 ( 
.A(n_7175),
.Y(n_8101)
);

INVx1_ASAP7_75t_SL g8102 ( 
.A(n_7286),
.Y(n_8102)
);

INVx2_ASAP7_75t_L g8103 ( 
.A(n_6620),
.Y(n_8103)
);

OAI21xp5_ASAP7_75t_L g8104 ( 
.A1(n_7177),
.A2(n_6514),
.B(n_6509),
.Y(n_8104)
);

OAI21x1_ASAP7_75t_SL g8105 ( 
.A1(n_6914),
.A2(n_6553),
.B(n_6213),
.Y(n_8105)
);

INVx1_ASAP7_75t_L g8106 ( 
.A(n_7175),
.Y(n_8106)
);

INVx1_ASAP7_75t_L g8107 ( 
.A(n_7193),
.Y(n_8107)
);

OAI21x1_ASAP7_75t_SL g8108 ( 
.A1(n_6914),
.A2(n_7456),
.B(n_7145),
.Y(n_8108)
);

AO31x2_ASAP7_75t_L g8109 ( 
.A1(n_7012),
.A2(n_6490),
.A3(n_6502),
.B(n_6394),
.Y(n_8109)
);

INVx1_ASAP7_75t_L g8110 ( 
.A(n_7193),
.Y(n_8110)
);

OA21x2_ASAP7_75t_L g8111 ( 
.A1(n_6569),
.A2(n_5926),
.B(n_5916),
.Y(n_8111)
);

INVx1_ASAP7_75t_L g8112 ( 
.A(n_7217),
.Y(n_8112)
);

CKINVDCx6p67_ASAP7_75t_R g8113 ( 
.A(n_6767),
.Y(n_8113)
);

INVx1_ASAP7_75t_L g8114 ( 
.A(n_7217),
.Y(n_8114)
);

AND2x4_ASAP7_75t_L g8115 ( 
.A(n_7142),
.B(n_6201),
.Y(n_8115)
);

AOI22xp33_ASAP7_75t_L g8116 ( 
.A1(n_6588),
.A2(n_6660),
.B1(n_6824),
.B2(n_7353),
.Y(n_8116)
);

CKINVDCx20_ASAP7_75t_R g8117 ( 
.A(n_6603),
.Y(n_8117)
);

AND2x2_ASAP7_75t_L g8118 ( 
.A(n_6764),
.B(n_5926),
.Y(n_8118)
);

INVx1_ASAP7_75t_L g8119 ( 
.A(n_7222),
.Y(n_8119)
);

OAI22xp5_ASAP7_75t_L g8120 ( 
.A1(n_6815),
.A2(n_5566),
.B1(n_6371),
.B2(n_6325),
.Y(n_8120)
);

INVx1_ASAP7_75t_L g8121 ( 
.A(n_7222),
.Y(n_8121)
);

OAI211xp5_ASAP7_75t_SL g8122 ( 
.A1(n_7123),
.A2(n_6195),
.B(n_6037),
.C(n_6091),
.Y(n_8122)
);

AO21x2_ASAP7_75t_L g8123 ( 
.A1(n_7000),
.A2(n_4789),
.B(n_5716),
.Y(n_8123)
);

INVx1_ASAP7_75t_L g8124 ( 
.A(n_7249),
.Y(n_8124)
);

NAND2xp5_ASAP7_75t_L g8125 ( 
.A(n_6863),
.B(n_5877),
.Y(n_8125)
);

INVx1_ASAP7_75t_L g8126 ( 
.A(n_7249),
.Y(n_8126)
);

INVx2_ASAP7_75t_L g8127 ( 
.A(n_6641),
.Y(n_8127)
);

AOI22xp33_ASAP7_75t_L g8128 ( 
.A1(n_6660),
.A2(n_6389),
.B1(n_6441),
.B2(n_6412),
.Y(n_8128)
);

AO21x2_ASAP7_75t_L g8129 ( 
.A1(n_7000),
.A2(n_5718),
.B(n_5716),
.Y(n_8129)
);

OAI21xp5_ASAP7_75t_L g8130 ( 
.A1(n_7068),
.A2(n_5693),
.B(n_5689),
.Y(n_8130)
);

OAI21xp5_ASAP7_75t_L g8131 ( 
.A1(n_6850),
.A2(n_6840),
.B(n_6815),
.Y(n_8131)
);

CKINVDCx5p33_ASAP7_75t_R g8132 ( 
.A(n_6802),
.Y(n_8132)
);

O2A1O1Ixp33_ASAP7_75t_L g8133 ( 
.A1(n_6714),
.A2(n_5899),
.B(n_5687),
.C(n_6510),
.Y(n_8133)
);

AOI22xp5_ASAP7_75t_L g8134 ( 
.A1(n_6815),
.A2(n_6412),
.B1(n_6441),
.B2(n_6389),
.Y(n_8134)
);

NAND2xp5_ASAP7_75t_L g8135 ( 
.A(n_6863),
.B(n_5877),
.Y(n_8135)
);

OAI22xp5_ASAP7_75t_L g8136 ( 
.A1(n_6840),
.A2(n_6456),
.B1(n_6463),
.B2(n_6457),
.Y(n_8136)
);

OR2x2_ASAP7_75t_L g8137 ( 
.A(n_6572),
.B(n_6526),
.Y(n_8137)
);

AND2x2_ASAP7_75t_L g8138 ( 
.A(n_6764),
.B(n_5926),
.Y(n_8138)
);

INVx3_ASAP7_75t_L g8139 ( 
.A(n_7047),
.Y(n_8139)
);

NAND2x1p5_ASAP7_75t_L g8140 ( 
.A(n_6916),
.B(n_5923),
.Y(n_8140)
);

BUFx3_ASAP7_75t_L g8141 ( 
.A(n_6767),
.Y(n_8141)
);

INVx1_ASAP7_75t_L g8142 ( 
.A(n_7268),
.Y(n_8142)
);

BUFx2_ASAP7_75t_L g8143 ( 
.A(n_7584),
.Y(n_8143)
);

OAI21x1_ASAP7_75t_SL g8144 ( 
.A1(n_6914),
.A2(n_5693),
.B(n_5689),
.Y(n_8144)
);

INVx1_ASAP7_75t_L g8145 ( 
.A(n_7268),
.Y(n_8145)
);

NAND2xp5_ASAP7_75t_L g8146 ( 
.A(n_6863),
.B(n_5945),
.Y(n_8146)
);

CKINVDCx11_ASAP7_75t_R g8147 ( 
.A(n_7074),
.Y(n_8147)
);

OR2x6_ASAP7_75t_L g8148 ( 
.A(n_6565),
.B(n_6433),
.Y(n_8148)
);

AO21x2_ASAP7_75t_L g8149 ( 
.A1(n_7000),
.A2(n_5718),
.B(n_5781),
.Y(n_8149)
);

OR2x2_ASAP7_75t_L g8150 ( 
.A(n_6572),
.B(n_6526),
.Y(n_8150)
);

NAND3xp33_ASAP7_75t_L g8151 ( 
.A(n_7105),
.B(n_6091),
.C(n_6059),
.Y(n_8151)
);

AND2x2_ASAP7_75t_L g8152 ( 
.A(n_6764),
.B(n_5949),
.Y(n_8152)
);

BUFx3_ASAP7_75t_L g8153 ( 
.A(n_6767),
.Y(n_8153)
);

INVx2_ASAP7_75t_L g8154 ( 
.A(n_6641),
.Y(n_8154)
);

NAND2xp33_ASAP7_75t_L g8155 ( 
.A(n_6698),
.B(n_6340),
.Y(n_8155)
);

NOR2xp33_ASAP7_75t_L g8156 ( 
.A(n_7029),
.B(n_6139),
.Y(n_8156)
);

AO21x2_ASAP7_75t_L g8157 ( 
.A1(n_6841),
.A2(n_5785),
.B(n_5781),
.Y(n_8157)
);

INVx3_ASAP7_75t_L g8158 ( 
.A(n_7047),
.Y(n_8158)
);

AO32x2_ASAP7_75t_L g8159 ( 
.A1(n_7154),
.A2(n_5994),
.A3(n_6017),
.B1(n_5991),
.B2(n_5989),
.Y(n_8159)
);

AND2x4_ASAP7_75t_L g8160 ( 
.A(n_7142),
.B(n_6294),
.Y(n_8160)
);

CKINVDCx8_ASAP7_75t_R g8161 ( 
.A(n_6698),
.Y(n_8161)
);

AND2x2_ASAP7_75t_L g8162 ( 
.A(n_6780),
.B(n_5949),
.Y(n_8162)
);

OAI21xp5_ASAP7_75t_L g8163 ( 
.A1(n_6850),
.A2(n_5774),
.B(n_5722),
.Y(n_8163)
);

AOI22xp33_ASAP7_75t_L g8164 ( 
.A1(n_7353),
.A2(n_6456),
.B1(n_6463),
.B2(n_6457),
.Y(n_8164)
);

BUFx3_ASAP7_75t_L g8165 ( 
.A(n_6767),
.Y(n_8165)
);

A2O1A1Ixp33_ASAP7_75t_L g8166 ( 
.A1(n_6832),
.A2(n_6493),
.B(n_6540),
.C(n_6525),
.Y(n_8166)
);

INVx1_ASAP7_75t_L g8167 ( 
.A(n_7277),
.Y(n_8167)
);

BUFx6f_ASAP7_75t_L g8168 ( 
.A(n_7060),
.Y(n_8168)
);

NOR2xp33_ASAP7_75t_L g8169 ( 
.A(n_6779),
.B(n_6192),
.Y(n_8169)
);

BUFx2_ASAP7_75t_L g8170 ( 
.A(n_7584),
.Y(n_8170)
);

INVx2_ASAP7_75t_L g8171 ( 
.A(n_6641),
.Y(n_8171)
);

INVx1_ASAP7_75t_L g8172 ( 
.A(n_7277),
.Y(n_8172)
);

INVx1_ASAP7_75t_L g8173 ( 
.A(n_7293),
.Y(n_8173)
);

NAND2xp5_ASAP7_75t_L g8174 ( 
.A(n_7161),
.B(n_5945),
.Y(n_8174)
);

BUFx6f_ASAP7_75t_L g8175 ( 
.A(n_7060),
.Y(n_8175)
);

INVx1_ASAP7_75t_L g8176 ( 
.A(n_7293),
.Y(n_8176)
);

AOI22xp33_ASAP7_75t_L g8177 ( 
.A1(n_6823),
.A2(n_6493),
.B1(n_6540),
.B2(n_6525),
.Y(n_8177)
);

INVx1_ASAP7_75t_L g8178 ( 
.A(n_7338),
.Y(n_8178)
);

OA21x2_ASAP7_75t_L g8179 ( 
.A1(n_6572),
.A2(n_5949),
.B(n_6322),
.Y(n_8179)
);

NOR2xp33_ASAP7_75t_L g8180 ( 
.A(n_6779),
.B(n_6192),
.Y(n_8180)
);

OAI22xp5_ASAP7_75t_L g8181 ( 
.A1(n_6840),
.A2(n_6552),
.B1(n_6198),
.B2(n_6516),
.Y(n_8181)
);

NOR2x1_ASAP7_75t_R g8182 ( 
.A(n_6795),
.B(n_5849),
.Y(n_8182)
);

OA21x2_ASAP7_75t_L g8183 ( 
.A1(n_6780),
.A2(n_6346),
.B(n_6322),
.Y(n_8183)
);

INVx6_ASAP7_75t_SL g8184 ( 
.A(n_6565),
.Y(n_8184)
);

NOR2xp67_ASAP7_75t_L g8185 ( 
.A(n_7142),
.B(n_5592),
.Y(n_8185)
);

NAND2xp5_ASAP7_75t_L g8186 ( 
.A(n_7161),
.B(n_6020),
.Y(n_8186)
);

NOR2xp33_ASAP7_75t_L g8187 ( 
.A(n_6903),
.B(n_7100),
.Y(n_8187)
);

INVx1_ASAP7_75t_L g8188 ( 
.A(n_7338),
.Y(n_8188)
);

NAND2xp5_ASAP7_75t_L g8189 ( 
.A(n_7333),
.B(n_6020),
.Y(n_8189)
);

AND2x4_ASAP7_75t_L g8190 ( 
.A(n_7142),
.B(n_6294),
.Y(n_8190)
);

BUFx2_ASAP7_75t_L g8191 ( 
.A(n_7584),
.Y(n_8191)
);

AO21x2_ASAP7_75t_L g8192 ( 
.A1(n_6841),
.A2(n_5785),
.B(n_6469),
.Y(n_8192)
);

BUFx2_ASAP7_75t_L g8193 ( 
.A(n_7584),
.Y(n_8193)
);

OA21x2_ASAP7_75t_L g8194 ( 
.A1(n_6780),
.A2(n_6347),
.B(n_6346),
.Y(n_8194)
);

BUFx3_ASAP7_75t_L g8195 ( 
.A(n_6795),
.Y(n_8195)
);

INVx1_ASAP7_75t_L g8196 ( 
.A(n_7368),
.Y(n_8196)
);

OAI221xp5_ASAP7_75t_L g8197 ( 
.A1(n_7134),
.A2(n_6250),
.B1(n_6198),
.B2(n_5774),
.C(n_6552),
.Y(n_8197)
);

AOI21xp33_ASAP7_75t_L g8198 ( 
.A1(n_7214),
.A2(n_6059),
.B(n_5741),
.Y(n_8198)
);

OR2x2_ASAP7_75t_L g8199 ( 
.A(n_6805),
.B(n_6812),
.Y(n_8199)
);

NAND2xp5_ASAP7_75t_L g8200 ( 
.A(n_7333),
.B(n_6031),
.Y(n_8200)
);

INVx1_ASAP7_75t_L g8201 ( 
.A(n_7368),
.Y(n_8201)
);

INVx4_ASAP7_75t_SL g8202 ( 
.A(n_6655),
.Y(n_8202)
);

AOI21xp5_ASAP7_75t_L g8203 ( 
.A1(n_6556),
.A2(n_6164),
.B(n_6496),
.Y(n_8203)
);

INVx2_ASAP7_75t_SL g8204 ( 
.A(n_7060),
.Y(n_8204)
);

A2O1A1Ixp33_ASAP7_75t_L g8205 ( 
.A1(n_7036),
.A2(n_6507),
.B(n_6516),
.C(n_5797),
.Y(n_8205)
);

OA21x2_ASAP7_75t_L g8206 ( 
.A1(n_6805),
.A2(n_6352),
.B(n_6347),
.Y(n_8206)
);

BUFx6f_ASAP7_75t_L g8207 ( 
.A(n_7060),
.Y(n_8207)
);

BUFx4f_ASAP7_75t_SL g8208 ( 
.A(n_6795),
.Y(n_8208)
);

INVx1_ASAP7_75t_L g8209 ( 
.A(n_7400),
.Y(n_8209)
);

OA21x2_ASAP7_75t_L g8210 ( 
.A1(n_6805),
.A2(n_6404),
.B(n_6352),
.Y(n_8210)
);

INVx1_ASAP7_75t_L g8211 ( 
.A(n_7400),
.Y(n_8211)
);

INVx2_ASAP7_75t_L g8212 ( 
.A(n_6641),
.Y(n_8212)
);

OAI22xp5_ASAP7_75t_SL g8213 ( 
.A1(n_6984),
.A2(n_6194),
.B1(n_6316),
.B2(n_6248),
.Y(n_8213)
);

INVx2_ASAP7_75t_L g8214 ( 
.A(n_6643),
.Y(n_8214)
);

AND2x4_ASAP7_75t_L g8215 ( 
.A(n_7142),
.B(n_6294),
.Y(n_8215)
);

INVx1_ASAP7_75t_L g8216 ( 
.A(n_7406),
.Y(n_8216)
);

NAND2x1p5_ASAP7_75t_L g8217 ( 
.A(n_6916),
.B(n_5923),
.Y(n_8217)
);

INVx1_ASAP7_75t_L g8218 ( 
.A(n_7406),
.Y(n_8218)
);

AOI22xp33_ASAP7_75t_L g8219 ( 
.A1(n_6823),
.A2(n_5787),
.B1(n_5948),
.B2(n_5617),
.Y(n_8219)
);

AOI21xp33_ASAP7_75t_L g8220 ( 
.A1(n_7214),
.A2(n_5741),
.B(n_5737),
.Y(n_8220)
);

OAI221xp5_ASAP7_75t_L g8221 ( 
.A1(n_7134),
.A2(n_6250),
.B1(n_5737),
.B2(n_5735),
.C(n_5787),
.Y(n_8221)
);

AOI21xp5_ASAP7_75t_L g8222 ( 
.A1(n_6556),
.A2(n_6539),
.B(n_6496),
.Y(n_8222)
);

OR2x2_ASAP7_75t_L g8223 ( 
.A(n_6812),
.B(n_6031),
.Y(n_8223)
);

INVx1_ASAP7_75t_L g8224 ( 
.A(n_7453),
.Y(n_8224)
);

AO21x2_ASAP7_75t_L g8225 ( 
.A1(n_6841),
.A2(n_6470),
.B(n_6469),
.Y(n_8225)
);

BUFx3_ASAP7_75t_L g8226 ( 
.A(n_6795),
.Y(n_8226)
);

INVx1_ASAP7_75t_L g8227 ( 
.A(n_7453),
.Y(n_8227)
);

O2A1O1Ixp33_ASAP7_75t_L g8228 ( 
.A1(n_6714),
.A2(n_5714),
.B(n_5792),
.C(n_5813),
.Y(n_8228)
);

OAI21xp5_ASAP7_75t_L g8229 ( 
.A1(n_7123),
.A2(n_5617),
.B(n_5714),
.Y(n_8229)
);

INVx1_ASAP7_75t_L g8230 ( 
.A(n_6573),
.Y(n_8230)
);

OAI21x1_ASAP7_75t_L g8231 ( 
.A1(n_6996),
.A2(n_7407),
.B(n_7308),
.Y(n_8231)
);

NAND2xp5_ASAP7_75t_L g8232 ( 
.A(n_6590),
.B(n_6046),
.Y(n_8232)
);

AOI22xp33_ASAP7_75t_L g8233 ( 
.A1(n_6704),
.A2(n_5797),
.B1(n_5735),
.B2(n_6049),
.Y(n_8233)
);

A2O1A1Ixp33_ASAP7_75t_SL g8234 ( 
.A1(n_7036),
.A2(n_7460),
.B(n_7003),
.C(n_7180),
.Y(n_8234)
);

AND2x4_ASAP7_75t_L g8235 ( 
.A(n_7142),
.B(n_6294),
.Y(n_8235)
);

NAND2x1p5_ASAP7_75t_L g8236 ( 
.A(n_6916),
.B(n_6923),
.Y(n_8236)
);

OAI21x1_ASAP7_75t_L g8237 ( 
.A1(n_7308),
.A2(n_6335),
.B(n_6334),
.Y(n_8237)
);

OR2x6_ASAP7_75t_L g8238 ( 
.A(n_6565),
.B(n_6433),
.Y(n_8238)
);

OA21x2_ASAP7_75t_L g8239 ( 
.A1(n_6812),
.A2(n_6421),
.B(n_6404),
.Y(n_8239)
);

AO21x2_ASAP7_75t_L g8240 ( 
.A1(n_7189),
.A2(n_6472),
.B(n_6470),
.Y(n_8240)
);

BUFx3_ASAP7_75t_L g8241 ( 
.A(n_6804),
.Y(n_8241)
);

BUFx2_ASAP7_75t_L g8242 ( 
.A(n_7584),
.Y(n_8242)
);

A2O1A1Ixp33_ASAP7_75t_L g8243 ( 
.A1(n_6677),
.A2(n_6507),
.B(n_6512),
.C(n_6503),
.Y(n_8243)
);

INVx1_ASAP7_75t_L g8244 ( 
.A(n_6573),
.Y(n_8244)
);

BUFx2_ASAP7_75t_L g8245 ( 
.A(n_7584),
.Y(n_8245)
);

OAI21xp5_ASAP7_75t_L g8246 ( 
.A1(n_7166),
.A2(n_7251),
.B(n_7404),
.Y(n_8246)
);

OA21x2_ASAP7_75t_L g8247 ( 
.A1(n_6834),
.A2(n_6421),
.B(n_6503),
.Y(n_8247)
);

INVx2_ASAP7_75t_L g8248 ( 
.A(n_6643),
.Y(n_8248)
);

AO21x2_ASAP7_75t_L g8249 ( 
.A1(n_7189),
.A2(n_6474),
.B(n_6472),
.Y(n_8249)
);

CKINVDCx5p33_ASAP7_75t_R g8250 ( 
.A(n_6586),
.Y(n_8250)
);

CKINVDCx8_ASAP7_75t_R g8251 ( 
.A(n_6760),
.Y(n_8251)
);

AO21x2_ASAP7_75t_L g8252 ( 
.A1(n_7189),
.A2(n_6482),
.B(n_6474),
.Y(n_8252)
);

AO21x2_ASAP7_75t_L g8253 ( 
.A1(n_6879),
.A2(n_6497),
.B(n_6482),
.Y(n_8253)
);

INVx3_ASAP7_75t_L g8254 ( 
.A(n_7060),
.Y(n_8254)
);

BUFx12f_ASAP7_75t_L g8255 ( 
.A(n_7230),
.Y(n_8255)
);

OAI21xp5_ASAP7_75t_L g8256 ( 
.A1(n_7166),
.A2(n_5792),
.B(n_5778),
.Y(n_8256)
);

CKINVDCx5p33_ASAP7_75t_R g8257 ( 
.A(n_6586),
.Y(n_8257)
);

OAI21x1_ASAP7_75t_L g8258 ( 
.A1(n_7308),
.A2(n_6335),
.B(n_6334),
.Y(n_8258)
);

HB1xp67_ASAP7_75t_L g8259 ( 
.A(n_7550),
.Y(n_8259)
);

OAI21x1_ASAP7_75t_L g8260 ( 
.A1(n_7308),
.A2(n_6359),
.B(n_6335),
.Y(n_8260)
);

INVx2_ASAP7_75t_L g8261 ( 
.A(n_6643),
.Y(n_8261)
);

OAI21x1_ASAP7_75t_L g8262 ( 
.A1(n_7308),
.A2(n_6359),
.B(n_6335),
.Y(n_8262)
);

CKINVDCx11_ASAP7_75t_R g8263 ( 
.A(n_7074),
.Y(n_8263)
);

NOR2xp33_ASAP7_75t_L g8264 ( 
.A(n_6903),
.B(n_5496),
.Y(n_8264)
);

A2O1A1Ixp33_ASAP7_75t_L g8265 ( 
.A1(n_6677),
.A2(n_6512),
.B(n_6517),
.C(n_6503),
.Y(n_8265)
);

INVx1_ASAP7_75t_L g8266 ( 
.A(n_6742),
.Y(n_8266)
);

OAI21x1_ASAP7_75t_L g8267 ( 
.A1(n_7407),
.A2(n_6359),
.B(n_6335),
.Y(n_8267)
);

OR2x2_ASAP7_75t_L g8268 ( 
.A(n_6834),
.B(n_6046),
.Y(n_8268)
);

INVx3_ASAP7_75t_L g8269 ( 
.A(n_7060),
.Y(n_8269)
);

AOI22xp33_ASAP7_75t_L g8270 ( 
.A1(n_6704),
.A2(n_6049),
.B1(n_6126),
.B2(n_5599),
.Y(n_8270)
);

INVx4_ASAP7_75t_L g8271 ( 
.A(n_6804),
.Y(n_8271)
);

A2O1A1Ixp33_ASAP7_75t_L g8272 ( 
.A1(n_6677),
.A2(n_6519),
.B(n_6543),
.C(n_6517),
.Y(n_8272)
);

NAND2xp5_ASAP7_75t_SL g8273 ( 
.A(n_6984),
.B(n_6479),
.Y(n_8273)
);

O2A1O1Ixp33_ASAP7_75t_L g8274 ( 
.A1(n_7224),
.A2(n_5813),
.B(n_6340),
.C(n_5522),
.Y(n_8274)
);

O2A1O1Ixp33_ASAP7_75t_SL g8275 ( 
.A1(n_7090),
.A2(n_7101),
.B(n_6891),
.C(n_7092),
.Y(n_8275)
);

NAND2xp5_ASAP7_75t_L g8276 ( 
.A(n_6590),
.B(n_6063),
.Y(n_8276)
);

OAI22xp33_ASAP7_75t_L g8277 ( 
.A1(n_6796),
.A2(n_6085),
.B1(n_6398),
.B2(n_5644),
.Y(n_8277)
);

INVx2_ASAP7_75t_L g8278 ( 
.A(n_6643),
.Y(n_8278)
);

BUFx4_ASAP7_75t_SL g8279 ( 
.A(n_7101),
.Y(n_8279)
);

OAI21x1_ASAP7_75t_L g8280 ( 
.A1(n_7407),
.A2(n_6902),
.B(n_6886),
.Y(n_8280)
);

CKINVDCx5p33_ASAP7_75t_R g8281 ( 
.A(n_6610),
.Y(n_8281)
);

OAI22xp33_ASAP7_75t_L g8282 ( 
.A1(n_6796),
.A2(n_6085),
.B1(n_6398),
.B2(n_5644),
.Y(n_8282)
);

NAND2xp5_ASAP7_75t_L g8283 ( 
.A(n_6710),
.B(n_6063),
.Y(n_8283)
);

OAI21x1_ASAP7_75t_SL g8284 ( 
.A1(n_7456),
.A2(n_5623),
.B(n_5605),
.Y(n_8284)
);

INVx2_ASAP7_75t_L g8285 ( 
.A(n_6646),
.Y(n_8285)
);

INVx1_ASAP7_75t_L g8286 ( 
.A(n_6742),
.Y(n_8286)
);

INVx2_ASAP7_75t_L g8287 ( 
.A(n_6646),
.Y(n_8287)
);

AOI22x1_ASAP7_75t_L g8288 ( 
.A1(n_6862),
.A2(n_7232),
.B1(n_6984),
.B2(n_6874),
.Y(n_8288)
);

INVx1_ASAP7_75t_L g8289 ( 
.A(n_6881),
.Y(n_8289)
);

AND2x4_ASAP7_75t_L g8290 ( 
.A(n_7142),
.B(n_6294),
.Y(n_8290)
);

AND2x4_ASAP7_75t_SL g8291 ( 
.A(n_6940),
.B(n_5557),
.Y(n_8291)
);

BUFx3_ASAP7_75t_L g8292 ( 
.A(n_6804),
.Y(n_8292)
);

OAI21x1_ASAP7_75t_L g8293 ( 
.A1(n_7407),
.A2(n_6902),
.B(n_6886),
.Y(n_8293)
);

INVx1_ASAP7_75t_L g8294 ( 
.A(n_6881),
.Y(n_8294)
);

INVx1_ASAP7_75t_L g8295 ( 
.A(n_6890),
.Y(n_8295)
);

INVx2_ASAP7_75t_L g8296 ( 
.A(n_6646),
.Y(n_8296)
);

INVx2_ASAP7_75t_L g8297 ( 
.A(n_6646),
.Y(n_8297)
);

AOI22xp33_ASAP7_75t_L g8298 ( 
.A1(n_6704),
.A2(n_6126),
.B1(n_5599),
.B2(n_5557),
.Y(n_8298)
);

INVx1_ASAP7_75t_L g8299 ( 
.A(n_6890),
.Y(n_8299)
);

NOR2xp67_ASAP7_75t_SL g8300 ( 
.A(n_7056),
.B(n_5937),
.Y(n_8300)
);

CKINVDCx6p67_ASAP7_75t_R g8301 ( 
.A(n_6804),
.Y(n_8301)
);

INVx1_ASAP7_75t_L g8302 ( 
.A(n_6975),
.Y(n_8302)
);

AOI221xp5_ASAP7_75t_L g8303 ( 
.A1(n_7224),
.A2(n_6442),
.B1(n_6440),
.B2(n_5769),
.C(n_5778),
.Y(n_8303)
);

OA21x2_ASAP7_75t_L g8304 ( 
.A1(n_6847),
.A2(n_6519),
.B(n_6543),
.Y(n_8304)
);

INVx1_ASAP7_75t_L g8305 ( 
.A(n_6975),
.Y(n_8305)
);

INVx1_ASAP7_75t_SL g8306 ( 
.A(n_7363),
.Y(n_8306)
);

OA21x2_ASAP7_75t_L g8307 ( 
.A1(n_6847),
.A2(n_6543),
.B(n_5556),
.Y(n_8307)
);

INVx2_ASAP7_75t_L g8308 ( 
.A(n_6647),
.Y(n_8308)
);

AND2x2_ASAP7_75t_L g8309 ( 
.A(n_6847),
.B(n_6237),
.Y(n_8309)
);

AOI21xp33_ASAP7_75t_L g8310 ( 
.A1(n_7214),
.A2(n_6266),
.B(n_6077),
.Y(n_8310)
);

OAI221xp5_ASAP7_75t_L g8311 ( 
.A1(n_7088),
.A2(n_5809),
.B1(n_5810),
.B2(n_5818),
.C(n_5806),
.Y(n_8311)
);

NAND3xp33_ASAP7_75t_L g8312 ( 
.A(n_7105),
.B(n_5818),
.C(n_5769),
.Y(n_8312)
);

HB1xp67_ASAP7_75t_L g8313 ( 
.A(n_7550),
.Y(n_8313)
);

A2O1A1Ixp33_ASAP7_75t_L g8314 ( 
.A1(n_6796),
.A2(n_6520),
.B(n_6523),
.C(n_5806),
.Y(n_8314)
);

HB1xp67_ASAP7_75t_L g8315 ( 
.A(n_7567),
.Y(n_8315)
);

CKINVDCx6p67_ASAP7_75t_R g8316 ( 
.A(n_6874),
.Y(n_8316)
);

OA21x2_ASAP7_75t_L g8317 ( 
.A1(n_6855),
.A2(n_5556),
.B(n_5553),
.Y(n_8317)
);

INVx1_ASAP7_75t_L g8318 ( 
.A(n_7567),
.Y(n_8318)
);

INVx5_ASAP7_75t_L g8319 ( 
.A(n_7060),
.Y(n_8319)
);

BUFx3_ASAP7_75t_L g8320 ( 
.A(n_6874),
.Y(n_8320)
);

OR2x2_ASAP7_75t_L g8321 ( 
.A(n_6855),
.B(n_6077),
.Y(n_8321)
);

OAI21xp5_ASAP7_75t_L g8322 ( 
.A1(n_7251),
.A2(n_5809),
.B(n_5810),
.Y(n_8322)
);

NOR2x1_ASAP7_75t_SL g8323 ( 
.A(n_6942),
.B(n_5551),
.Y(n_8323)
);

A2O1A1Ixp33_ASAP7_75t_L g8324 ( 
.A1(n_6607),
.A2(n_6520),
.B(n_6523),
.C(n_6479),
.Y(n_8324)
);

AND2x2_ASAP7_75t_L g8325 ( 
.A(n_6855),
.B(n_6237),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7581),
.Y(n_8326)
);

NAND2xp5_ASAP7_75t_L g8327 ( 
.A(n_6710),
.B(n_6266),
.Y(n_8327)
);

INVx1_ASAP7_75t_L g8328 ( 
.A(n_7581),
.Y(n_8328)
);

INVxp33_ASAP7_75t_L g8329 ( 
.A(n_7527),
.Y(n_8329)
);

AOI22xp5_ASAP7_75t_L g8330 ( 
.A1(n_6995),
.A2(n_5800),
.B1(n_6479),
.B2(n_6085),
.Y(n_8330)
);

INVx1_ASAP7_75t_L g8331 ( 
.A(n_6686),
.Y(n_8331)
);

INVx1_ASAP7_75t_L g8332 ( 
.A(n_6686),
.Y(n_8332)
);

AND2x2_ASAP7_75t_L g8333 ( 
.A(n_6892),
.B(n_6901),
.Y(n_8333)
);

INVx1_ASAP7_75t_L g8334 ( 
.A(n_6686),
.Y(n_8334)
);

CKINVDCx16_ASAP7_75t_R g8335 ( 
.A(n_6874),
.Y(n_8335)
);

NAND2xp5_ASAP7_75t_L g8336 ( 
.A(n_6877),
.B(n_6174),
.Y(n_8336)
);

AOI22xp5_ASAP7_75t_L g8337 ( 
.A1(n_6995),
.A2(n_5800),
.B1(n_5644),
.B2(n_5692),
.Y(n_8337)
);

NAND2xp5_ASAP7_75t_SL g8338 ( 
.A(n_7282),
.B(n_5980),
.Y(n_8338)
);

OAI21xp5_ASAP7_75t_L g8339 ( 
.A1(n_7404),
.A2(n_5637),
.B(n_5630),
.Y(n_8339)
);

AND2x4_ASAP7_75t_L g8340 ( 
.A(n_7142),
.B(n_6373),
.Y(n_8340)
);

NAND2x1_ASAP7_75t_L g8341 ( 
.A(n_7556),
.B(n_5985),
.Y(n_8341)
);

OAI21x1_ASAP7_75t_L g8342 ( 
.A1(n_6939),
.A2(n_6974),
.B(n_6973),
.Y(n_8342)
);

AOI221xp5_ASAP7_75t_L g8343 ( 
.A1(n_7224),
.A2(n_6854),
.B1(n_6846),
.B2(n_7107),
.C(n_6816),
.Y(n_8343)
);

NOR4xp25_ASAP7_75t_L g8344 ( 
.A(n_7273),
.B(n_5522),
.C(n_5523),
.D(n_5496),
.Y(n_8344)
);

AOI22xp33_ASAP7_75t_L g8345 ( 
.A1(n_6564),
.A2(n_5579),
.B1(n_6107),
.B2(n_5692),
.Y(n_8345)
);

OAI22xp33_ASAP7_75t_L g8346 ( 
.A1(n_6607),
.A2(n_5579),
.B1(n_6107),
.B2(n_5692),
.Y(n_8346)
);

INVx2_ASAP7_75t_L g8347 ( 
.A(n_6647),
.Y(n_8347)
);

OAI21x1_ASAP7_75t_L g8348 ( 
.A1(n_6973),
.A2(n_6974),
.B(n_7017),
.Y(n_8348)
);

OA21x2_ASAP7_75t_L g8349 ( 
.A1(n_6892),
.A2(n_5560),
.B(n_5553),
.Y(n_8349)
);

OA21x2_ASAP7_75t_L g8350 ( 
.A1(n_6892),
.A2(n_5561),
.B(n_5560),
.Y(n_8350)
);

INVx1_ASAP7_75t_SL g8351 ( 
.A(n_7363),
.Y(n_8351)
);

NOR2xp33_ASAP7_75t_L g8352 ( 
.A(n_7100),
.B(n_5523),
.Y(n_8352)
);

OR2x2_ASAP7_75t_L g8353 ( 
.A(n_6901),
.B(n_5552),
.Y(n_8353)
);

BUFx2_ASAP7_75t_L g8354 ( 
.A(n_7584),
.Y(n_8354)
);

INVx2_ASAP7_75t_L g8355 ( 
.A(n_6647),
.Y(n_8355)
);

NOR2xp67_ASAP7_75t_L g8356 ( 
.A(n_7142),
.B(n_5592),
.Y(n_8356)
);

INVx5_ASAP7_75t_SL g8357 ( 
.A(n_6690),
.Y(n_8357)
);

AOI22xp33_ASAP7_75t_L g8358 ( 
.A1(n_6564),
.A2(n_6107),
.B1(n_6136),
.B2(n_5551),
.Y(n_8358)
);

AO21x2_ASAP7_75t_L g8359 ( 
.A1(n_6879),
.A2(n_5479),
.B(n_5478),
.Y(n_8359)
);

INVx1_ASAP7_75t_L g8360 ( 
.A(n_6708),
.Y(n_8360)
);

AOI22xp5_ASAP7_75t_L g8361 ( 
.A1(n_6995),
.A2(n_6136),
.B1(n_5551),
.B2(n_5955),
.Y(n_8361)
);

AOI22xp33_ASAP7_75t_L g8362 ( 
.A1(n_6732),
.A2(n_6136),
.B1(n_5551),
.B2(n_5479),
.Y(n_8362)
);

OAI21xp5_ASAP7_75t_L g8363 ( 
.A1(n_6830),
.A2(n_6607),
.B(n_6732),
.Y(n_8363)
);

AOI22xp5_ASAP7_75t_L g8364 ( 
.A1(n_6615),
.A2(n_5551),
.B1(n_5955),
.B2(n_5105),
.Y(n_8364)
);

AOI21xp5_ASAP7_75t_L g8365 ( 
.A1(n_6556),
.A2(n_6539),
.B(n_6496),
.Y(n_8365)
);

OAI21xp5_ASAP7_75t_L g8366 ( 
.A1(n_6830),
.A2(n_5637),
.B(n_5630),
.Y(n_8366)
);

AO21x2_ASAP7_75t_L g8367 ( 
.A1(n_7030),
.A2(n_5479),
.B(n_5478),
.Y(n_8367)
);

OAI22x1_ASAP7_75t_L g8368 ( 
.A1(n_6925),
.A2(n_5616),
.B1(n_5669),
.B2(n_5592),
.Y(n_8368)
);

HB1xp67_ASAP7_75t_L g8369 ( 
.A(n_6587),
.Y(n_8369)
);

OAI22xp5_ASAP7_75t_L g8370 ( 
.A1(n_6665),
.A2(n_6442),
.B1(n_6440),
.B2(n_5616),
.Y(n_8370)
);

NOR2x1_ASAP7_75t_SL g8371 ( 
.A(n_6959),
.B(n_5985),
.Y(n_8371)
);

AOI22xp33_ASAP7_75t_L g8372 ( 
.A1(n_6816),
.A2(n_5479),
.B1(n_5478),
.B2(n_5520),
.Y(n_8372)
);

OAI21xp5_ASAP7_75t_L g8373 ( 
.A1(n_6830),
.A2(n_5479),
.B(n_5478),
.Y(n_8373)
);

BUFx3_ASAP7_75t_L g8374 ( 
.A(n_6992),
.Y(n_8374)
);

NAND2xp5_ASAP7_75t_L g8375 ( 
.A(n_6877),
.B(n_6174),
.Y(n_8375)
);

INVx2_ASAP7_75t_L g8376 ( 
.A(n_6647),
.Y(n_8376)
);

NAND2xp5_ASAP7_75t_L g8377 ( 
.A(n_6882),
.B(n_6174),
.Y(n_8377)
);

AOI21xp5_ASAP7_75t_L g8378 ( 
.A1(n_6568),
.A2(n_6539),
.B(n_6496),
.Y(n_8378)
);

INVx4_ASAP7_75t_L g8379 ( 
.A(n_6992),
.Y(n_8379)
);

NAND2xp5_ASAP7_75t_L g8380 ( 
.A(n_6882),
.B(n_6203),
.Y(n_8380)
);

AOI21xp5_ASAP7_75t_L g8381 ( 
.A1(n_6568),
.A2(n_6539),
.B(n_6496),
.Y(n_8381)
);

NAND2xp5_ASAP7_75t_L g8382 ( 
.A(n_6585),
.B(n_6203),
.Y(n_8382)
);

NAND2xp5_ASAP7_75t_SL g8383 ( 
.A(n_7352),
.B(n_5985),
.Y(n_8383)
);

INVx2_ASAP7_75t_L g8384 ( 
.A(n_6674),
.Y(n_8384)
);

INVx1_ASAP7_75t_L g8385 ( 
.A(n_6708),
.Y(n_8385)
);

AO21x2_ASAP7_75t_L g8386 ( 
.A1(n_7030),
.A2(n_5478),
.B(n_5561),
.Y(n_8386)
);

INVx1_ASAP7_75t_L g8387 ( 
.A(n_6708),
.Y(n_8387)
);

INVx2_ASAP7_75t_L g8388 ( 
.A(n_6674),
.Y(n_8388)
);

AOI221xp5_ASAP7_75t_L g8389 ( 
.A1(n_6846),
.A2(n_5706),
.B1(n_5709),
.B2(n_5660),
.C(n_5654),
.Y(n_8389)
);

AND2x2_ASAP7_75t_L g8390 ( 
.A(n_6901),
.B(n_6237),
.Y(n_8390)
);

AOI21xp5_ASAP7_75t_L g8391 ( 
.A1(n_6568),
.A2(n_6539),
.B(n_6496),
.Y(n_8391)
);

INVx6_ASAP7_75t_L g8392 ( 
.A(n_7015),
.Y(n_8392)
);

NAND2xp5_ASAP7_75t_L g8393 ( 
.A(n_6585),
.B(n_6203),
.Y(n_8393)
);

AO222x2_ASAP7_75t_L g8394 ( 
.A1(n_6862),
.A2(n_5881),
.B1(n_5851),
.B2(n_5520),
.C1(n_5549),
.C2(n_5608),
.Y(n_8394)
);

OAI21xp5_ASAP7_75t_L g8395 ( 
.A1(n_7273),
.A2(n_5660),
.B(n_5654),
.Y(n_8395)
);

NAND2x1p5_ASAP7_75t_L g8396 ( 
.A(n_6923),
.B(n_5923),
.Y(n_8396)
);

INVx2_ASAP7_75t_L g8397 ( 
.A(n_6674),
.Y(n_8397)
);

OAI21x1_ASAP7_75t_L g8398 ( 
.A1(n_6883),
.A2(n_6888),
.B(n_7129),
.Y(n_8398)
);

AOI221x1_ASAP7_75t_L g8399 ( 
.A1(n_7273),
.A2(n_6465),
.B1(n_5998),
.B2(n_6008),
.C(n_5987),
.Y(n_8399)
);

OAI21x1_ASAP7_75t_SL g8400 ( 
.A1(n_6950),
.A2(n_5623),
.B(n_5605),
.Y(n_8400)
);

OAI21x1_ASAP7_75t_SL g8401 ( 
.A1(n_6950),
.A2(n_5623),
.B(n_5605),
.Y(n_8401)
);

INVx2_ASAP7_75t_L g8402 ( 
.A(n_6674),
.Y(n_8402)
);

INVx2_ASAP7_75t_L g8403 ( 
.A(n_6693),
.Y(n_8403)
);

INVx1_ASAP7_75t_L g8404 ( 
.A(n_6712),
.Y(n_8404)
);

INVx1_ASAP7_75t_L g8405 ( 
.A(n_6712),
.Y(n_8405)
);

OAI21x1_ASAP7_75t_L g8406 ( 
.A1(n_7129),
.A2(n_6279),
.B(n_6261),
.Y(n_8406)
);

INVx2_ASAP7_75t_L g8407 ( 
.A(n_6693),
.Y(n_8407)
);

INVx1_ASAP7_75t_L g8408 ( 
.A(n_6712),
.Y(n_8408)
);

AND2x4_ASAP7_75t_L g8409 ( 
.A(n_7184),
.B(n_7195),
.Y(n_8409)
);

AND2x2_ASAP7_75t_L g8410 ( 
.A(n_6577),
.B(n_6301),
.Y(n_8410)
);

NAND2xp5_ASAP7_75t_L g8411 ( 
.A(n_6630),
.B(n_5552),
.Y(n_8411)
);

NAND2xp5_ASAP7_75t_L g8412 ( 
.A(n_6630),
.B(n_5909),
.Y(n_8412)
);

NOR2xp33_ASAP7_75t_L g8413 ( 
.A(n_7125),
.B(n_5879),
.Y(n_8413)
);

INVxp67_ASAP7_75t_SL g8414 ( 
.A(n_7321),
.Y(n_8414)
);

HB1xp67_ASAP7_75t_L g8415 ( 
.A(n_6587),
.Y(n_8415)
);

OA21x2_ASAP7_75t_L g8416 ( 
.A1(n_7129),
.A2(n_6608),
.B(n_6577),
.Y(n_8416)
);

INVx1_ASAP7_75t_SL g8417 ( 
.A(n_7363),
.Y(n_8417)
);

INVx1_ASAP7_75t_L g8418 ( 
.A(n_6719),
.Y(n_8418)
);

INVx1_ASAP7_75t_L g8419 ( 
.A(n_6719),
.Y(n_8419)
);

OA21x2_ASAP7_75t_L g8420 ( 
.A1(n_7129),
.A2(n_6608),
.B(n_6577),
.Y(n_8420)
);

AOI21x1_ASAP7_75t_L g8421 ( 
.A1(n_6600),
.A2(n_6292),
.B(n_6449),
.Y(n_8421)
);

OAI21x1_ASAP7_75t_L g8422 ( 
.A1(n_7435),
.A2(n_6286),
.B(n_6279),
.Y(n_8422)
);

INVx2_ASAP7_75t_L g8423 ( 
.A(n_6693),
.Y(n_8423)
);

INVx1_ASAP7_75t_L g8424 ( 
.A(n_6719),
.Y(n_8424)
);

AOI21xp5_ASAP7_75t_L g8425 ( 
.A1(n_7449),
.A2(n_6544),
.B(n_6539),
.Y(n_8425)
);

NAND2xp33_ASAP7_75t_L g8426 ( 
.A(n_6760),
.B(n_6340),
.Y(n_8426)
);

INVx1_ASAP7_75t_L g8427 ( 
.A(n_6734),
.Y(n_8427)
);

OAI21x1_ASAP7_75t_L g8428 ( 
.A1(n_7435),
.A2(n_6293),
.B(n_6286),
.Y(n_8428)
);

NAND2x1p5_ASAP7_75t_L g8429 ( 
.A(n_6923),
.B(n_5923),
.Y(n_8429)
);

AOI22xp5_ASAP7_75t_L g8430 ( 
.A1(n_6658),
.A2(n_5955),
.B1(n_5677),
.B2(n_5658),
.Y(n_8430)
);

OAI21x1_ASAP7_75t_L g8431 ( 
.A1(n_7435),
.A2(n_6293),
.B(n_6286),
.Y(n_8431)
);

AOI21x1_ASAP7_75t_L g8432 ( 
.A1(n_6600),
.A2(n_6449),
.B(n_5680),
.Y(n_8432)
);

INVx3_ASAP7_75t_L g8433 ( 
.A(n_7060),
.Y(n_8433)
);

NAND2xp33_ASAP7_75t_L g8434 ( 
.A(n_6857),
.B(n_6340),
.Y(n_8434)
);

OAI21x1_ASAP7_75t_L g8435 ( 
.A1(n_7435),
.A2(n_6296),
.B(n_6293),
.Y(n_8435)
);

INVx2_ASAP7_75t_L g8436 ( 
.A(n_6693),
.Y(n_8436)
);

OAI21x1_ASAP7_75t_L g8437 ( 
.A1(n_7457),
.A2(n_6315),
.B(n_6296),
.Y(n_8437)
);

AND2x2_ASAP7_75t_L g8438 ( 
.A(n_6577),
.B(n_6301),
.Y(n_8438)
);

OAI21xp5_ASAP7_75t_L g8439 ( 
.A1(n_7229),
.A2(n_5709),
.B(n_5706),
.Y(n_8439)
);

INVx2_ASAP7_75t_L g8440 ( 
.A(n_6701),
.Y(n_8440)
);

OR2x2_ASAP7_75t_L g8441 ( 
.A(n_6587),
.B(n_6597),
.Y(n_8441)
);

OAI21x1_ASAP7_75t_L g8442 ( 
.A1(n_7457),
.A2(n_7604),
.B(n_7508),
.Y(n_8442)
);

AND2x4_ASAP7_75t_L g8443 ( 
.A(n_7184),
.B(n_6373),
.Y(n_8443)
);

INVx1_ASAP7_75t_L g8444 ( 
.A(n_6734),
.Y(n_8444)
);

INVx2_ASAP7_75t_SL g8445 ( 
.A(n_7060),
.Y(n_8445)
);

OAI21x1_ASAP7_75t_L g8446 ( 
.A1(n_7457),
.A2(n_6315),
.B(n_6296),
.Y(n_8446)
);

OAI21x1_ASAP7_75t_L g8447 ( 
.A1(n_7457),
.A2(n_7604),
.B(n_7508),
.Y(n_8447)
);

BUFx3_ASAP7_75t_L g8448 ( 
.A(n_6992),
.Y(n_8448)
);

INVx2_ASAP7_75t_L g8449 ( 
.A(n_6701),
.Y(n_8449)
);

NAND2xp5_ASAP7_75t_L g8450 ( 
.A(n_6631),
.B(n_5909),
.Y(n_8450)
);

NOR2xp67_ASAP7_75t_L g8451 ( 
.A(n_7184),
.B(n_5669),
.Y(n_8451)
);

INVx4_ASAP7_75t_L g8452 ( 
.A(n_6992),
.Y(n_8452)
);

AO21x2_ASAP7_75t_L g8453 ( 
.A1(n_7030),
.A2(n_5564),
.B(n_5563),
.Y(n_8453)
);

INVx6_ASAP7_75t_L g8454 ( 
.A(n_7015),
.Y(n_8454)
);

AOI21xp33_ASAP7_75t_SL g8455 ( 
.A1(n_6857),
.A2(n_5541),
.B(n_5474),
.Y(n_8455)
);

OAI21x1_ASAP7_75t_L g8456 ( 
.A1(n_7508),
.A2(n_6317),
.B(n_6315),
.Y(n_8456)
);

BUFx3_ASAP7_75t_L g8457 ( 
.A(n_6655),
.Y(n_8457)
);

NAND2xp5_ASAP7_75t_L g8458 ( 
.A(n_6631),
.B(n_6103),
.Y(n_8458)
);

NAND2xp5_ASAP7_75t_SL g8459 ( 
.A(n_7352),
.B(n_5985),
.Y(n_8459)
);

CKINVDCx20_ASAP7_75t_R g8460 ( 
.A(n_6716),
.Y(n_8460)
);

BUFx2_ASAP7_75t_L g8461 ( 
.A(n_7584),
.Y(n_8461)
);

O2A1O1Ixp33_ASAP7_75t_SL g8462 ( 
.A1(n_6891),
.A2(n_5827),
.B(n_5883),
.C(n_5811),
.Y(n_8462)
);

OAI21xp5_ASAP7_75t_L g8463 ( 
.A1(n_7229),
.A2(n_6092),
.B(n_5793),
.Y(n_8463)
);

NAND2xp5_ASAP7_75t_L g8464 ( 
.A(n_7125),
.B(n_6103),
.Y(n_8464)
);

OAI21xp5_ASAP7_75t_L g8465 ( 
.A1(n_6680),
.A2(n_6092),
.B(n_6182),
.Y(n_8465)
);

O2A1O1Ixp33_ASAP7_75t_L g8466 ( 
.A1(n_6596),
.A2(n_6465),
.B(n_5620),
.C(n_5622),
.Y(n_8466)
);

AOI21xp5_ASAP7_75t_L g8467 ( 
.A1(n_7449),
.A2(n_6544),
.B(n_6539),
.Y(n_8467)
);

AOI221xp5_ASAP7_75t_L g8468 ( 
.A1(n_6854),
.A2(n_5622),
.B1(n_5620),
.B2(n_5618),
.C(n_6182),
.Y(n_8468)
);

AO21x2_ASAP7_75t_L g8469 ( 
.A1(n_6709),
.A2(n_5564),
.B(n_5563),
.Y(n_8469)
);

NAND2xp5_ASAP7_75t_L g8470 ( 
.A(n_7133),
.B(n_6187),
.Y(n_8470)
);

OR2x6_ASAP7_75t_SL g8471 ( 
.A(n_7113),
.B(n_6893),
.Y(n_8471)
);

OAI21x1_ASAP7_75t_L g8472 ( 
.A1(n_7604),
.A2(n_7437),
.B(n_6929),
.Y(n_8472)
);

OAI221xp5_ASAP7_75t_L g8473 ( 
.A1(n_7088),
.A2(n_5987),
.B1(n_6008),
.B2(n_5998),
.C(n_5985),
.Y(n_8473)
);

OAI22xp33_ASAP7_75t_L g8474 ( 
.A1(n_6665),
.A2(n_4896),
.B1(n_4915),
.B2(n_4908),
.Y(n_8474)
);

AOI21xp5_ASAP7_75t_L g8475 ( 
.A1(n_7147),
.A2(n_6544),
.B(n_5869),
.Y(n_8475)
);

A2O1A1Ixp33_ASAP7_75t_L g8476 ( 
.A1(n_7107),
.A2(n_5985),
.B(n_5998),
.C(n_5987),
.Y(n_8476)
);

OAI21x1_ASAP7_75t_L g8477 ( 
.A1(n_7437),
.A2(n_6345),
.B(n_6332),
.Y(n_8477)
);

OAI21x1_ASAP7_75t_L g8478 ( 
.A1(n_7437),
.A2(n_6345),
.B(n_6332),
.Y(n_8478)
);

NOR2xp67_ASAP7_75t_SL g8479 ( 
.A(n_7352),
.B(n_5937),
.Y(n_8479)
);

AO31x2_ASAP7_75t_L g8480 ( 
.A1(n_7574),
.A2(n_6319),
.A3(n_6326),
.B(n_6307),
.Y(n_8480)
);

BUFx4f_ASAP7_75t_SL g8481 ( 
.A(n_6716),
.Y(n_8481)
);

BUFx3_ASAP7_75t_L g8482 ( 
.A(n_6655),
.Y(n_8482)
);

NAND2xp5_ASAP7_75t_L g8483 ( 
.A(n_7133),
.B(n_6187),
.Y(n_8483)
);

INVxp67_ASAP7_75t_L g8484 ( 
.A(n_7241),
.Y(n_8484)
);

AO21x2_ASAP7_75t_L g8485 ( 
.A1(n_6709),
.A2(n_5573),
.B(n_5569),
.Y(n_8485)
);

A2O1A1Ixp33_ASAP7_75t_L g8486 ( 
.A1(n_7092),
.A2(n_5985),
.B(n_5998),
.C(n_5987),
.Y(n_8486)
);

CKINVDCx11_ASAP7_75t_R g8487 ( 
.A(n_6610),
.Y(n_8487)
);

CKINVDCx20_ASAP7_75t_R g8488 ( 
.A(n_6755),
.Y(n_8488)
);

INVx2_ASAP7_75t_L g8489 ( 
.A(n_6701),
.Y(n_8489)
);

BUFx3_ASAP7_75t_L g8490 ( 
.A(n_6655),
.Y(n_8490)
);

NAND2xp5_ASAP7_75t_L g8491 ( 
.A(n_7139),
.B(n_6245),
.Y(n_8491)
);

OAI22xp5_ASAP7_75t_L g8492 ( 
.A1(n_6627),
.A2(n_6121),
.B1(n_6175),
.B2(n_6163),
.Y(n_8492)
);

AND2x2_ASAP7_75t_L g8493 ( 
.A(n_6608),
.B(n_6301),
.Y(n_8493)
);

AND2x2_ASAP7_75t_L g8494 ( 
.A(n_6608),
.B(n_6343),
.Y(n_8494)
);

INVx1_ASAP7_75t_L g8495 ( 
.A(n_6734),
.Y(n_8495)
);

OAI21x1_ASAP7_75t_L g8496 ( 
.A1(n_6977),
.A2(n_6363),
.B(n_6357),
.Y(n_8496)
);

CKINVDCx8_ASAP7_75t_R g8497 ( 
.A(n_6887),
.Y(n_8497)
);

OAI21x1_ASAP7_75t_L g8498 ( 
.A1(n_6977),
.A2(n_6392),
.B(n_6363),
.Y(n_8498)
);

NAND2xp5_ASAP7_75t_L g8499 ( 
.A(n_7139),
.B(n_6245),
.Y(n_8499)
);

AO31x2_ASAP7_75t_L g8500 ( 
.A1(n_7574),
.A2(n_6319),
.A3(n_6326),
.B(n_6307),
.Y(n_8500)
);

OAI21x1_ASAP7_75t_L g8501 ( 
.A1(n_6977),
.A2(n_6397),
.B(n_6392),
.Y(n_8501)
);

OAI21x1_ASAP7_75t_L g8502 ( 
.A1(n_6977),
.A2(n_6397),
.B(n_6392),
.Y(n_8502)
);

OAI21x1_ASAP7_75t_L g8503 ( 
.A1(n_7044),
.A2(n_7112),
.B(n_7078),
.Y(n_8503)
);

INVx2_ASAP7_75t_L g8504 ( 
.A(n_6701),
.Y(n_8504)
);

INVxp33_ASAP7_75t_L g8505 ( 
.A(n_7527),
.Y(n_8505)
);

OAI21x1_ASAP7_75t_L g8506 ( 
.A1(n_7044),
.A2(n_6400),
.B(n_6397),
.Y(n_8506)
);

AOI21xp5_ASAP7_75t_L g8507 ( 
.A1(n_7147),
.A2(n_6544),
.B(n_5869),
.Y(n_8507)
);

INVx2_ASAP7_75t_L g8508 ( 
.A(n_6715),
.Y(n_8508)
);

INVxp67_ASAP7_75t_L g8509 ( 
.A(n_7241),
.Y(n_8509)
);

OAI21x1_ASAP7_75t_L g8510 ( 
.A1(n_7044),
.A2(n_6405),
.B(n_6400),
.Y(n_8510)
);

AND2x4_ASAP7_75t_L g8511 ( 
.A(n_7184),
.B(n_6373),
.Y(n_8511)
);

AO31x2_ASAP7_75t_L g8512 ( 
.A1(n_7574),
.A2(n_7372),
.A3(n_7504),
.B(n_7487),
.Y(n_8512)
);

HB1xp67_ASAP7_75t_L g8513 ( 
.A(n_6597),
.Y(n_8513)
);

CKINVDCx5p33_ASAP7_75t_R g8514 ( 
.A(n_6649),
.Y(n_8514)
);

INVx1_ASAP7_75t_L g8515 ( 
.A(n_6736),
.Y(n_8515)
);

A2O1A1Ixp33_ASAP7_75t_L g8516 ( 
.A1(n_6627),
.A2(n_5985),
.B(n_5998),
.C(n_5987),
.Y(n_8516)
);

INVx4_ASAP7_75t_SL g8517 ( 
.A(n_6655),
.Y(n_8517)
);

INVx3_ASAP7_75t_L g8518 ( 
.A(n_7079),
.Y(n_8518)
);

OR2x2_ASAP7_75t_L g8519 ( 
.A(n_6597),
.B(n_6381),
.Y(n_8519)
);

OAI21x1_ASAP7_75t_L g8520 ( 
.A1(n_7044),
.A2(n_6405),
.B(n_6400),
.Y(n_8520)
);

INVx1_ASAP7_75t_L g8521 ( 
.A(n_6736),
.Y(n_8521)
);

OAI21x1_ASAP7_75t_L g8522 ( 
.A1(n_7078),
.A2(n_7112),
.B(n_6987),
.Y(n_8522)
);

INVx2_ASAP7_75t_SL g8523 ( 
.A(n_7079),
.Y(n_8523)
);

OAI21xp5_ASAP7_75t_L g8524 ( 
.A1(n_6680),
.A2(n_6471),
.B(n_6381),
.Y(n_8524)
);

CKINVDCx5p33_ASAP7_75t_R g8525 ( 
.A(n_6649),
.Y(n_8525)
);

INVx1_ASAP7_75t_L g8526 ( 
.A(n_6736),
.Y(n_8526)
);

AOI21xp5_ASAP7_75t_L g8527 ( 
.A1(n_7408),
.A2(n_6544),
.B(n_5869),
.Y(n_8527)
);

INVx3_ASAP7_75t_L g8528 ( 
.A(n_7079),
.Y(n_8528)
);

AOI21xp5_ASAP7_75t_L g8529 ( 
.A1(n_7408),
.A2(n_6544),
.B(n_5869),
.Y(n_8529)
);

AOI22xp33_ASAP7_75t_L g8530 ( 
.A1(n_6658),
.A2(n_5539),
.B1(n_5549),
.B2(n_5520),
.Y(n_8530)
);

AOI22xp5_ASAP7_75t_L g8531 ( 
.A1(n_6862),
.A2(n_5677),
.B1(n_5658),
.B2(n_5549),
.Y(n_8531)
);

OAI21xp5_ASAP7_75t_L g8532 ( 
.A1(n_7163),
.A2(n_6515),
.B(n_6471),
.Y(n_8532)
);

BUFx4f_ASAP7_75t_L g8533 ( 
.A(n_7348),
.Y(n_8533)
);

AOI22xp5_ASAP7_75t_L g8534 ( 
.A1(n_7065),
.A2(n_5658),
.B1(n_5677),
.B2(n_5583),
.Y(n_8534)
);

OAI21x1_ASAP7_75t_L g8535 ( 
.A1(n_7078),
.A2(n_6406),
.B(n_6405),
.Y(n_8535)
);

NAND2xp5_ASAP7_75t_L g8536 ( 
.A(n_6944),
.B(n_6515),
.Y(n_8536)
);

AO21x2_ASAP7_75t_L g8537 ( 
.A1(n_6709),
.A2(n_5573),
.B(n_5569),
.Y(n_8537)
);

O2A1O1Ixp33_ASAP7_75t_L g8538 ( 
.A1(n_7424),
.A2(n_5618),
.B(n_5815),
.C(n_5794),
.Y(n_8538)
);

INVx1_ASAP7_75t_L g8539 ( 
.A(n_6747),
.Y(n_8539)
);

OAI21xp5_ASAP7_75t_L g8540 ( 
.A1(n_7163),
.A2(n_5671),
.B(n_5669),
.Y(n_8540)
);

AOI22xp33_ASAP7_75t_L g8541 ( 
.A1(n_6782),
.A2(n_5583),
.B1(n_5608),
.B2(n_5539),
.Y(n_8541)
);

INVx3_ASAP7_75t_SL g8542 ( 
.A(n_6909),
.Y(n_8542)
);

OAI21x1_ASAP7_75t_L g8543 ( 
.A1(n_7078),
.A2(n_6420),
.B(n_6406),
.Y(n_8543)
);

INVx3_ASAP7_75t_L g8544 ( 
.A(n_7079),
.Y(n_8544)
);

OAI21xp5_ASAP7_75t_L g8545 ( 
.A1(n_7424),
.A2(n_5705),
.B(n_5671),
.Y(n_8545)
);

OAI21x1_ASAP7_75t_L g8546 ( 
.A1(n_7112),
.A2(n_6987),
.B(n_6956),
.Y(n_8546)
);

BUFx10_ASAP7_75t_L g8547 ( 
.A(n_6828),
.Y(n_8547)
);

OAI21x1_ASAP7_75t_L g8548 ( 
.A1(n_7112),
.A2(n_6420),
.B(n_6406),
.Y(n_8548)
);

NAND2x1p5_ASAP7_75t_L g8549 ( 
.A(n_6923),
.B(n_5930),
.Y(n_8549)
);

NAND2xp5_ASAP7_75t_L g8550 ( 
.A(n_6944),
.B(n_5811),
.Y(n_8550)
);

NOR3xp33_ASAP7_75t_L g8551 ( 
.A(n_7137),
.B(n_5623),
.C(n_5605),
.Y(n_8551)
);

O2A1O1Ixp33_ASAP7_75t_SL g8552 ( 
.A1(n_7522),
.A2(n_5883),
.B(n_5827),
.C(n_6073),
.Y(n_8552)
);

OAI21x1_ASAP7_75t_L g8553 ( 
.A1(n_7442),
.A2(n_6430),
.B(n_6422),
.Y(n_8553)
);

CKINVDCx16_ASAP7_75t_R g8554 ( 
.A(n_6836),
.Y(n_8554)
);

OR2x2_ASAP7_75t_L g8555 ( 
.A(n_6617),
.B(n_6314),
.Y(n_8555)
);

BUFx3_ASAP7_75t_L g8556 ( 
.A(n_6655),
.Y(n_8556)
);

OAI21x1_ASAP7_75t_L g8557 ( 
.A1(n_7442),
.A2(n_6430),
.B(n_6422),
.Y(n_8557)
);

OAI21x1_ASAP7_75t_L g8558 ( 
.A1(n_7442),
.A2(n_6438),
.B(n_6430),
.Y(n_8558)
);

INVx1_ASAP7_75t_L g8559 ( 
.A(n_6747),
.Y(n_8559)
);

INVx2_ASAP7_75t_L g8560 ( 
.A(n_6715),
.Y(n_8560)
);

AOI21x1_ASAP7_75t_L g8561 ( 
.A1(n_7599),
.A2(n_5680),
.B(n_6307),
.Y(n_8561)
);

INVxp67_ASAP7_75t_L g8562 ( 
.A(n_7262),
.Y(n_8562)
);

OAI22xp33_ASAP7_75t_L g8563 ( 
.A1(n_7048),
.A2(n_4908),
.B1(n_4919),
.B2(n_4915),
.Y(n_8563)
);

OAI21x1_ASAP7_75t_L g8564 ( 
.A1(n_7442),
.A2(n_6447),
.B(n_6438),
.Y(n_8564)
);

AOI22xp33_ASAP7_75t_L g8565 ( 
.A1(n_6782),
.A2(n_5583),
.B1(n_5608),
.B2(n_5539),
.Y(n_8565)
);

OAI21x1_ASAP7_75t_L g8566 ( 
.A1(n_7442),
.A2(n_7372),
.B(n_7172),
.Y(n_8566)
);

INVxp67_ASAP7_75t_L g8567 ( 
.A(n_7262),
.Y(n_8567)
);

OA21x2_ASAP7_75t_L g8568 ( 
.A1(n_6654),
.A2(n_5586),
.B(n_5578),
.Y(n_8568)
);

OAI21x1_ASAP7_75t_L g8569 ( 
.A1(n_7442),
.A2(n_6447),
.B(n_6438),
.Y(n_8569)
);

AO21x2_ASAP7_75t_L g8570 ( 
.A1(n_6725),
.A2(n_6880),
.B(n_7577),
.Y(n_8570)
);

INVx2_ASAP7_75t_L g8571 ( 
.A(n_6715),
.Y(n_8571)
);

AO21x2_ASAP7_75t_L g8572 ( 
.A1(n_6725),
.A2(n_5586),
.B(n_5578),
.Y(n_8572)
);

AOI22xp33_ASAP7_75t_L g8573 ( 
.A1(n_6783),
.A2(n_5609),
.B1(n_5647),
.B2(n_5632),
.Y(n_8573)
);

OAI21x1_ASAP7_75t_L g8574 ( 
.A1(n_7442),
.A2(n_6454),
.B(n_6447),
.Y(n_8574)
);

INVx1_ASAP7_75t_L g8575 ( 
.A(n_6747),
.Y(n_8575)
);

NAND2xp5_ASAP7_75t_L g8576 ( 
.A(n_6944),
.B(n_5984),
.Y(n_8576)
);

OAI21x1_ASAP7_75t_L g8577 ( 
.A1(n_7372),
.A2(n_6467),
.B(n_6454),
.Y(n_8577)
);

INVx2_ASAP7_75t_L g8578 ( 
.A(n_6715),
.Y(n_8578)
);

BUFx3_ASAP7_75t_L g8579 ( 
.A(n_6655),
.Y(n_8579)
);

AO21x2_ASAP7_75t_L g8580 ( 
.A1(n_6725),
.A2(n_5610),
.B(n_5597),
.Y(n_8580)
);

INVx1_ASAP7_75t_L g8581 ( 
.A(n_6753),
.Y(n_8581)
);

BUFx12f_ASAP7_75t_L g8582 ( 
.A(n_7600),
.Y(n_8582)
);

INVx2_ASAP7_75t_SL g8583 ( 
.A(n_7079),
.Y(n_8583)
);

AOI21x1_ASAP7_75t_L g8584 ( 
.A1(n_7599),
.A2(n_6326),
.B(n_6319),
.Y(n_8584)
);

A2O1A1Ixp33_ASAP7_75t_L g8585 ( 
.A1(n_6800),
.A2(n_5998),
.B(n_6008),
.C(n_5987),
.Y(n_8585)
);

OA21x2_ASAP7_75t_L g8586 ( 
.A1(n_6654),
.A2(n_5610),
.B(n_5597),
.Y(n_8586)
);

INVx1_ASAP7_75t_L g8587 ( 
.A(n_6753),
.Y(n_8587)
);

INVx1_ASAP7_75t_L g8588 ( 
.A(n_6753),
.Y(n_8588)
);

INVx3_ASAP7_75t_L g8589 ( 
.A(n_7079),
.Y(n_8589)
);

AOI22xp33_ASAP7_75t_L g8590 ( 
.A1(n_6783),
.A2(n_5609),
.B1(n_5647),
.B2(n_5632),
.Y(n_8590)
);

AOI221xp5_ASAP7_75t_L g8591 ( 
.A1(n_6784),
.A2(n_7137),
.B1(n_7143),
.B2(n_6629),
.C(n_6687),
.Y(n_8591)
);

OAI21xp5_ASAP7_75t_L g8592 ( 
.A1(n_6997),
.A2(n_5705),
.B(n_5671),
.Y(n_8592)
);

OAI21x1_ASAP7_75t_L g8593 ( 
.A1(n_7035),
.A2(n_7245),
.B(n_7172),
.Y(n_8593)
);

OAI22xp5_ASAP7_75t_L g8594 ( 
.A1(n_6871),
.A2(n_6121),
.B1(n_6175),
.B2(n_6163),
.Y(n_8594)
);

OA21x2_ASAP7_75t_L g8595 ( 
.A1(n_6654),
.A2(n_5628),
.B(n_5613),
.Y(n_8595)
);

OAI22xp5_ASAP7_75t_L g8596 ( 
.A1(n_6871),
.A2(n_6121),
.B1(n_6175),
.B2(n_6163),
.Y(n_8596)
);

NAND2xp5_ASAP7_75t_L g8597 ( 
.A(n_7324),
.B(n_5996),
.Y(n_8597)
);

OAI21xp5_ASAP7_75t_L g8598 ( 
.A1(n_6997),
.A2(n_5760),
.B(n_5705),
.Y(n_8598)
);

INVx1_ASAP7_75t_L g8599 ( 
.A(n_6757),
.Y(n_8599)
);

AO21x1_ASAP7_75t_L g8600 ( 
.A1(n_7003),
.A2(n_6545),
.B(n_6541),
.Y(n_8600)
);

OAI211xp5_ASAP7_75t_L g8601 ( 
.A1(n_7143),
.A2(n_5794),
.B(n_5816),
.C(n_5815),
.Y(n_8601)
);

INVx1_ASAP7_75t_L g8602 ( 
.A(n_6757),
.Y(n_8602)
);

BUFx2_ASAP7_75t_L g8603 ( 
.A(n_7584),
.Y(n_8603)
);

INVx2_ASAP7_75t_L g8604 ( 
.A(n_6720),
.Y(n_8604)
);

AND2x2_ASAP7_75t_L g8605 ( 
.A(n_6654),
.B(n_6343),
.Y(n_8605)
);

OA21x2_ASAP7_75t_L g8606 ( 
.A1(n_6676),
.A2(n_5628),
.B(n_5613),
.Y(n_8606)
);

AOI221xp5_ASAP7_75t_L g8607 ( 
.A1(n_6784),
.A2(n_5816),
.B1(n_6074),
.B2(n_6086),
.C(n_6073),
.Y(n_8607)
);

NAND2x1p5_ASAP7_75t_L g8608 ( 
.A(n_6923),
.B(n_5930),
.Y(n_8608)
);

AO31x2_ASAP7_75t_L g8609 ( 
.A1(n_7487),
.A2(n_6382),
.A3(n_6337),
.B(n_6348),
.Y(n_8609)
);

OAI21xp5_ASAP7_75t_L g8610 ( 
.A1(n_6994),
.A2(n_5760),
.B(n_6121),
.Y(n_8610)
);

INVx1_ASAP7_75t_L g8611 ( 
.A(n_6757),
.Y(n_8611)
);

AOI22xp33_ASAP7_75t_L g8612 ( 
.A1(n_7232),
.A2(n_5609),
.B1(n_5647),
.B2(n_5632),
.Y(n_8612)
);

O2A1O1Ixp33_ASAP7_75t_L g8613 ( 
.A1(n_6703),
.A2(n_5186),
.B(n_5203),
.C(n_5138),
.Y(n_8613)
);

OR2x6_ASAP7_75t_L g8614 ( 
.A(n_6565),
.B(n_6433),
.Y(n_8614)
);

INVx2_ASAP7_75t_L g8615 ( 
.A(n_6720),
.Y(n_8615)
);

AOI21xp5_ASAP7_75t_L g8616 ( 
.A1(n_7408),
.A2(n_6544),
.B(n_5869),
.Y(n_8616)
);

OAI21xp5_ASAP7_75t_L g8617 ( 
.A1(n_6994),
.A2(n_5760),
.B(n_6121),
.Y(n_8617)
);

BUFx6f_ASAP7_75t_L g8618 ( 
.A(n_7079),
.Y(n_8618)
);

AOI21xp5_ASAP7_75t_L g8619 ( 
.A1(n_6976),
.A2(n_5869),
.B(n_5588),
.Y(n_8619)
);

INVx2_ASAP7_75t_L g8620 ( 
.A(n_6720),
.Y(n_8620)
);

AOI21xp5_ASAP7_75t_L g8621 ( 
.A1(n_6976),
.A2(n_5869),
.B(n_5588),
.Y(n_8621)
);

OA21x2_ASAP7_75t_L g8622 ( 
.A1(n_6676),
.A2(n_5642),
.B(n_5638),
.Y(n_8622)
);

AO31x2_ASAP7_75t_L g8623 ( 
.A1(n_7487),
.A2(n_6337),
.A3(n_6348),
.B(n_6333),
.Y(n_8623)
);

O2A1O1Ixp33_ASAP7_75t_SL g8624 ( 
.A1(n_7522),
.A2(n_6086),
.B(n_6090),
.C(n_6074),
.Y(n_8624)
);

AND2x4_ASAP7_75t_L g8625 ( 
.A(n_7184),
.B(n_6373),
.Y(n_8625)
);

NAND2xp5_ASAP7_75t_L g8626 ( 
.A(n_7324),
.B(n_5996),
.Y(n_8626)
);

INVx1_ASAP7_75t_L g8627 ( 
.A(n_6777),
.Y(n_8627)
);

AOI21xp5_ASAP7_75t_L g8628 ( 
.A1(n_6976),
.A2(n_5588),
.B(n_6175),
.Y(n_8628)
);

AOI22xp33_ASAP7_75t_L g8629 ( 
.A1(n_7232),
.A2(n_6687),
.B1(n_6629),
.B2(n_7065),
.Y(n_8629)
);

INVx2_ASAP7_75t_L g8630 ( 
.A(n_6720),
.Y(n_8630)
);

AO32x2_ASAP7_75t_L g8631 ( 
.A1(n_7154),
.A2(n_5994),
.A3(n_6017),
.B1(n_5991),
.B2(n_5989),
.Y(n_8631)
);

BUFx12f_ASAP7_75t_L g8632 ( 
.A(n_7230),
.Y(n_8632)
);

BUFx6f_ASAP7_75t_L g8633 ( 
.A(n_7079),
.Y(n_8633)
);

NOR2xp67_ASAP7_75t_L g8634 ( 
.A(n_7184),
.B(n_5501),
.Y(n_8634)
);

HB1xp67_ASAP7_75t_L g8635 ( 
.A(n_6617),
.Y(n_8635)
);

AOI21xp5_ASAP7_75t_L g8636 ( 
.A1(n_6976),
.A2(n_5588),
.B(n_6481),
.Y(n_8636)
);

INVx2_ASAP7_75t_L g8637 ( 
.A(n_6721),
.Y(n_8637)
);

INVx1_ASAP7_75t_L g8638 ( 
.A(n_6777),
.Y(n_8638)
);

AOI22xp33_ASAP7_75t_L g8639 ( 
.A1(n_7065),
.A2(n_6093),
.B1(n_6042),
.B2(n_5998),
.Y(n_8639)
);

HB1xp67_ASAP7_75t_L g8640 ( 
.A(n_6617),
.Y(n_8640)
);

INVx5_ASAP7_75t_L g8641 ( 
.A(n_7079),
.Y(n_8641)
);

BUFx6f_ASAP7_75t_L g8642 ( 
.A(n_7103),
.Y(n_8642)
);

HB1xp67_ASAP7_75t_L g8643 ( 
.A(n_6632),
.Y(n_8643)
);

BUFx6f_ASAP7_75t_L g8644 ( 
.A(n_7103),
.Y(n_8644)
);

INVx1_ASAP7_75t_L g8645 ( 
.A(n_6777),
.Y(n_8645)
);

INVx1_ASAP7_75t_SL g8646 ( 
.A(n_7382),
.Y(n_8646)
);

AOI221xp5_ASAP7_75t_L g8647 ( 
.A1(n_7279),
.A2(n_7211),
.B1(n_6703),
.B2(n_6711),
.C(n_6960),
.Y(n_8647)
);

NAND2xp5_ASAP7_75t_SL g8648 ( 
.A(n_7590),
.B(n_5987),
.Y(n_8648)
);

INVx6_ASAP7_75t_L g8649 ( 
.A(n_7015),
.Y(n_8649)
);

HB1xp67_ASAP7_75t_L g8650 ( 
.A(n_6632),
.Y(n_8650)
);

NAND2xp5_ASAP7_75t_L g8651 ( 
.A(n_7332),
.B(n_6005),
.Y(n_8651)
);

INVx3_ASAP7_75t_L g8652 ( 
.A(n_7103),
.Y(n_8652)
);

OR2x2_ASAP7_75t_L g8653 ( 
.A(n_6632),
.B(n_6638),
.Y(n_8653)
);

INVx2_ASAP7_75t_L g8654 ( 
.A(n_6721),
.Y(n_8654)
);

OAI21x1_ASAP7_75t_L g8655 ( 
.A1(n_7172),
.A2(n_7245),
.B(n_7512),
.Y(n_8655)
);

OAI21x1_ASAP7_75t_SL g8656 ( 
.A1(n_7306),
.A2(n_5623),
.B(n_5605),
.Y(n_8656)
);

AOI22xp5_ASAP7_75t_L g8657 ( 
.A1(n_7041),
.A2(n_4769),
.B1(n_5652),
.B2(n_5627),
.Y(n_8657)
);

HB1xp67_ASAP7_75t_L g8658 ( 
.A(n_6638),
.Y(n_8658)
);

INVx2_ASAP7_75t_L g8659 ( 
.A(n_6721),
.Y(n_8659)
);

OAI221xp5_ASAP7_75t_L g8660 ( 
.A1(n_7041),
.A2(n_6008),
.B1(n_6012),
.B2(n_5998),
.C(n_5987),
.Y(n_8660)
);

INVx1_ASAP7_75t_L g8661 ( 
.A(n_6781),
.Y(n_8661)
);

NOR2xp33_ASAP7_75t_L g8662 ( 
.A(n_7417),
.B(n_5882),
.Y(n_8662)
);

AO21x1_ASAP7_75t_L g8663 ( 
.A1(n_7205),
.A2(n_6534),
.B(n_6527),
.Y(n_8663)
);

OAI21x1_ASAP7_75t_L g8664 ( 
.A1(n_7245),
.A2(n_7512),
.B(n_6737),
.Y(n_8664)
);

INVx2_ASAP7_75t_L g8665 ( 
.A(n_6721),
.Y(n_8665)
);

INVx3_ASAP7_75t_L g8666 ( 
.A(n_7103),
.Y(n_8666)
);

INVx1_ASAP7_75t_L g8667 ( 
.A(n_6781),
.Y(n_8667)
);

INVx1_ASAP7_75t_L g8668 ( 
.A(n_6781),
.Y(n_8668)
);

OAI22xp5_ASAP7_75t_L g8669 ( 
.A1(n_6889),
.A2(n_6163),
.B1(n_6214),
.B2(n_6175),
.Y(n_8669)
);

BUFx2_ASAP7_75t_R g8670 ( 
.A(n_7216),
.Y(n_8670)
);

OAI22xp33_ASAP7_75t_L g8671 ( 
.A1(n_7048),
.A2(n_4908),
.B1(n_4919),
.B2(n_4915),
.Y(n_8671)
);

INVx2_ASAP7_75t_L g8672 ( 
.A(n_6738),
.Y(n_8672)
);

AND2x4_ASAP7_75t_L g8673 ( 
.A(n_7184),
.B(n_7195),
.Y(n_8673)
);

O2A1O1Ixp33_ASAP7_75t_SL g8674 ( 
.A1(n_6836),
.A2(n_6101),
.B(n_6102),
.C(n_6090),
.Y(n_8674)
);

OAI21x1_ASAP7_75t_L g8675 ( 
.A1(n_6737),
.A2(n_6521),
.B(n_6513),
.Y(n_8675)
);

OAI21x1_ASAP7_75t_L g8676 ( 
.A1(n_6737),
.A2(n_6524),
.B(n_6521),
.Y(n_8676)
);

AND2x4_ASAP7_75t_L g8677 ( 
.A(n_7184),
.B(n_6373),
.Y(n_8677)
);

OAI21xp5_ASAP7_75t_L g8678 ( 
.A1(n_6711),
.A2(n_6214),
.B(n_6163),
.Y(n_8678)
);

NAND2xp5_ASAP7_75t_L g8679 ( 
.A(n_7332),
.B(n_6005),
.Y(n_8679)
);

AOI22xp33_ASAP7_75t_L g8680 ( 
.A1(n_6889),
.A2(n_6093),
.B1(n_6012),
.B2(n_6014),
.Y(n_8680)
);

OAI21x1_ASAP7_75t_L g8681 ( 
.A1(n_6728),
.A2(n_6524),
.B(n_6521),
.Y(n_8681)
);

INVx1_ASAP7_75t_L g8682 ( 
.A(n_6789),
.Y(n_8682)
);

NOR2x1_ASAP7_75t_R g8683 ( 
.A(n_7600),
.B(n_5851),
.Y(n_8683)
);

AOI221xp5_ASAP7_75t_L g8684 ( 
.A1(n_7211),
.A2(n_6109),
.B1(n_6112),
.B2(n_6102),
.C(n_6101),
.Y(n_8684)
);

CKINVDCx8_ASAP7_75t_R g8685 ( 
.A(n_6887),
.Y(n_8685)
);

OAI21x1_ASAP7_75t_L g8686 ( 
.A1(n_6728),
.A2(n_6542),
.B(n_6524),
.Y(n_8686)
);

NAND2x1p5_ASAP7_75t_L g8687 ( 
.A(n_6923),
.B(n_5930),
.Y(n_8687)
);

OAI21xp5_ASAP7_75t_L g8688 ( 
.A1(n_6943),
.A2(n_6252),
.B(n_6214),
.Y(n_8688)
);

AND2x4_ASAP7_75t_L g8689 ( 
.A(n_7184),
.B(n_6384),
.Y(n_8689)
);

NOR2xp67_ASAP7_75t_L g8690 ( 
.A(n_7195),
.B(n_5501),
.Y(n_8690)
);

OAI21x1_ASAP7_75t_L g8691 ( 
.A1(n_6728),
.A2(n_6546),
.B(n_6542),
.Y(n_8691)
);

NAND2xp5_ASAP7_75t_L g8692 ( 
.A(n_6634),
.B(n_6009),
.Y(n_8692)
);

OAI21x1_ASAP7_75t_L g8693 ( 
.A1(n_6985),
.A2(n_6546),
.B(n_6542),
.Y(n_8693)
);

AO31x2_ASAP7_75t_L g8694 ( 
.A1(n_7504),
.A2(n_6337),
.A3(n_6348),
.B(n_6333),
.Y(n_8694)
);

OAI21xp5_ASAP7_75t_L g8695 ( 
.A1(n_6943),
.A2(n_6252),
.B(n_6214),
.Y(n_8695)
);

INVx2_ASAP7_75t_L g8696 ( 
.A(n_6738),
.Y(n_8696)
);

INVx2_ASAP7_75t_L g8697 ( 
.A(n_6738),
.Y(n_8697)
);

AOI22xp33_ASAP7_75t_L g8698 ( 
.A1(n_7033),
.A2(n_6093),
.B1(n_6012),
.B2(n_6014),
.Y(n_8698)
);

NAND2xp5_ASAP7_75t_SL g8699 ( 
.A(n_7590),
.B(n_7356),
.Y(n_8699)
);

OAI21x1_ASAP7_75t_L g8700 ( 
.A1(n_6985),
.A2(n_6546),
.B(n_5757),
.Y(n_8700)
);

OAI21x1_ASAP7_75t_L g8701 ( 
.A1(n_6985),
.A2(n_5757),
.B(n_5752),
.Y(n_8701)
);

AND2x4_ASAP7_75t_L g8702 ( 
.A(n_7195),
.B(n_6384),
.Y(n_8702)
);

AND2x4_ASAP7_75t_L g8703 ( 
.A(n_7195),
.B(n_6384),
.Y(n_8703)
);

OAI21x1_ASAP7_75t_L g8704 ( 
.A1(n_6985),
.A2(n_5757),
.B(n_5752),
.Y(n_8704)
);

NOR2xp33_ASAP7_75t_L g8705 ( 
.A(n_7417),
.B(n_5879),
.Y(n_8705)
);

NAND3xp33_ASAP7_75t_L g8706 ( 
.A(n_7109),
.B(n_6012),
.C(n_6008),
.Y(n_8706)
);

HB1xp67_ASAP7_75t_L g8707 ( 
.A(n_6638),
.Y(n_8707)
);

AO31x2_ASAP7_75t_L g8708 ( 
.A1(n_7504),
.A2(n_6378),
.A3(n_6382),
.B(n_6333),
.Y(n_8708)
);

O2A1O1Ixp33_ASAP7_75t_L g8709 ( 
.A1(n_7158),
.A2(n_5203),
.B(n_5318),
.C(n_5186),
.Y(n_8709)
);

BUFx2_ASAP7_75t_L g8710 ( 
.A(n_7584),
.Y(n_8710)
);

INVx5_ASAP7_75t_L g8711 ( 
.A(n_7103),
.Y(n_8711)
);

CKINVDCx5p33_ASAP7_75t_R g8712 ( 
.A(n_6606),
.Y(n_8712)
);

AND2x2_ASAP7_75t_L g8713 ( 
.A(n_6676),
.B(n_6343),
.Y(n_8713)
);

OAI21x1_ASAP7_75t_L g8714 ( 
.A1(n_6985),
.A2(n_5757),
.B(n_5752),
.Y(n_8714)
);

INVx1_ASAP7_75t_L g8715 ( 
.A(n_6789),
.Y(n_8715)
);

OAI22xp5_ASAP7_75t_L g8716 ( 
.A1(n_7300),
.A2(n_6214),
.B1(n_6379),
.B2(n_6252),
.Y(n_8716)
);

INVx2_ASAP7_75t_L g8717 ( 
.A(n_6738),
.Y(n_8717)
);

AOI22xp33_ASAP7_75t_L g8718 ( 
.A1(n_7033),
.A2(n_6042),
.B1(n_6012),
.B2(n_6014),
.Y(n_8718)
);

AOI222xp33_ASAP7_75t_L g8719 ( 
.A1(n_7244),
.A2(n_5851),
.B1(n_5881),
.B2(n_5937),
.C1(n_6259),
.C2(n_6248),
.Y(n_8719)
);

INVx1_ASAP7_75t_L g8720 ( 
.A(n_6789),
.Y(n_8720)
);

OAI21x1_ASAP7_75t_L g8721 ( 
.A1(n_6985),
.A2(n_5757),
.B(n_5752),
.Y(n_8721)
);

OAI21xp5_ASAP7_75t_L g8722 ( 
.A1(n_6745),
.A2(n_6379),
.B(n_6252),
.Y(n_8722)
);

INVx2_ASAP7_75t_L g8723 ( 
.A(n_6743),
.Y(n_8723)
);

HB1xp67_ASAP7_75t_L g8724 ( 
.A(n_6642),
.Y(n_8724)
);

INVx2_ASAP7_75t_L g8725 ( 
.A(n_6743),
.Y(n_8725)
);

INVx1_ASAP7_75t_L g8726 ( 
.A(n_6808),
.Y(n_8726)
);

NAND2xp5_ASAP7_75t_L g8727 ( 
.A(n_6634),
.B(n_6009),
.Y(n_8727)
);

INVx1_ASAP7_75t_L g8728 ( 
.A(n_6808),
.Y(n_8728)
);

AND2x2_ASAP7_75t_L g8729 ( 
.A(n_6676),
.B(n_6349),
.Y(n_8729)
);

INVx2_ASAP7_75t_L g8730 ( 
.A(n_6743),
.Y(n_8730)
);

HB1xp67_ASAP7_75t_L g8731 ( 
.A(n_6642),
.Y(n_8731)
);

OAI22xp5_ASAP7_75t_L g8732 ( 
.A1(n_7300),
.A2(n_6252),
.B1(n_6481),
.B2(n_6379),
.Y(n_8732)
);

OAI21x1_ASAP7_75t_L g8733 ( 
.A1(n_6985),
.A2(n_5791),
.B(n_5752),
.Y(n_8733)
);

INVx1_ASAP7_75t_L g8734 ( 
.A(n_6808),
.Y(n_8734)
);

OAI21x1_ASAP7_75t_L g8735 ( 
.A1(n_7434),
.A2(n_5842),
.B(n_5791),
.Y(n_8735)
);

INVx2_ASAP7_75t_L g8736 ( 
.A(n_6743),
.Y(n_8736)
);

BUFx2_ASAP7_75t_L g8737 ( 
.A(n_7373),
.Y(n_8737)
);

NOR2x1_ASAP7_75t_SL g8738 ( 
.A(n_6959),
.B(n_6008),
.Y(n_8738)
);

CKINVDCx5p33_ASAP7_75t_R g8739 ( 
.A(n_6606),
.Y(n_8739)
);

NAND2x1p5_ASAP7_75t_L g8740 ( 
.A(n_6923),
.B(n_5930),
.Y(n_8740)
);

NAND2xp5_ASAP7_75t_L g8741 ( 
.A(n_7111),
.B(n_6016),
.Y(n_8741)
);

BUFx2_ASAP7_75t_L g8742 ( 
.A(n_7373),
.Y(n_8742)
);

NAND3xp33_ASAP7_75t_L g8743 ( 
.A(n_7109),
.B(n_6012),
.C(n_6008),
.Y(n_8743)
);

INVxp67_ASAP7_75t_L g8744 ( 
.A(n_7589),
.Y(n_8744)
);

CKINVDCx5p33_ASAP7_75t_R g8745 ( 
.A(n_6755),
.Y(n_8745)
);

INVx1_ASAP7_75t_L g8746 ( 
.A(n_6809),
.Y(n_8746)
);

AOI21xp33_ASAP7_75t_SL g8747 ( 
.A1(n_6909),
.A2(n_6434),
.B(n_6375),
.Y(n_8747)
);

BUFx6f_ASAP7_75t_L g8748 ( 
.A(n_7103),
.Y(n_8748)
);

OA21x2_ASAP7_75t_L g8749 ( 
.A1(n_6685),
.A2(n_6751),
.B(n_6697),
.Y(n_8749)
);

INVx2_ASAP7_75t_L g8750 ( 
.A(n_6744),
.Y(n_8750)
);

AOI21xp5_ASAP7_75t_L g8751 ( 
.A1(n_6976),
.A2(n_5588),
.B(n_6379),
.Y(n_8751)
);

OAI21x1_ASAP7_75t_SL g8752 ( 
.A1(n_7306),
.A2(n_6924),
.B(n_6910),
.Y(n_8752)
);

NAND2xp5_ASAP7_75t_L g8753 ( 
.A(n_7111),
.B(n_6016),
.Y(n_8753)
);

NAND2x1p5_ASAP7_75t_L g8754 ( 
.A(n_6923),
.B(n_5930),
.Y(n_8754)
);

OAI21xp5_ASAP7_75t_L g8755 ( 
.A1(n_6745),
.A2(n_6481),
.B(n_6379),
.Y(n_8755)
);

OAI21xp5_ASAP7_75t_L g8756 ( 
.A1(n_7007),
.A2(n_6481),
.B(n_6112),
.Y(n_8756)
);

AOI21x1_ASAP7_75t_L g8757 ( 
.A1(n_7110),
.A2(n_6382),
.B(n_6378),
.Y(n_8757)
);

OAI21xp5_ASAP7_75t_L g8758 ( 
.A1(n_7007),
.A2(n_6481),
.B(n_6114),
.Y(n_8758)
);

OA21x2_ASAP7_75t_L g8759 ( 
.A1(n_6685),
.A2(n_5683),
.B(n_5657),
.Y(n_8759)
);

AOI22xp33_ASAP7_75t_L g8760 ( 
.A1(n_7341),
.A2(n_6042),
.B1(n_6012),
.B2(n_6014),
.Y(n_8760)
);

NOR2x1_ASAP7_75t_R g8761 ( 
.A(n_7348),
.B(n_5881),
.Y(n_8761)
);

OAI21x1_ASAP7_75t_L g8762 ( 
.A1(n_7434),
.A2(n_7198),
.B(n_6924),
.Y(n_8762)
);

AO32x2_ASAP7_75t_L g8763 ( 
.A1(n_7154),
.A2(n_6017),
.A3(n_6096),
.B1(n_5994),
.B2(n_5991),
.Y(n_8763)
);

INVx1_ASAP7_75t_L g8764 ( 
.A(n_6809),
.Y(n_8764)
);

OAI21x1_ASAP7_75t_L g8765 ( 
.A1(n_7434),
.A2(n_5842),
.B(n_5791),
.Y(n_8765)
);

INVx2_ASAP7_75t_L g8766 ( 
.A(n_6744),
.Y(n_8766)
);

INVx1_ASAP7_75t_L g8767 ( 
.A(n_6809),
.Y(n_8767)
);

BUFx2_ASAP7_75t_L g8768 ( 
.A(n_7373),
.Y(n_8768)
);

AOI22xp33_ASAP7_75t_L g8769 ( 
.A1(n_7341),
.A2(n_6048),
.B1(n_6082),
.B2(n_6008),
.Y(n_8769)
);

NOR2xp33_ASAP7_75t_L g8770 ( 
.A(n_7279),
.B(n_5879),
.Y(n_8770)
);

INVx1_ASAP7_75t_L g8771 ( 
.A(n_6814),
.Y(n_8771)
);

NOR2xp33_ASAP7_75t_L g8772 ( 
.A(n_6966),
.B(n_5879),
.Y(n_8772)
);

OAI21x1_ASAP7_75t_SL g8773 ( 
.A1(n_6910),
.A2(n_7477),
.B(n_7474),
.Y(n_8773)
);

INVx1_ASAP7_75t_L g8774 ( 
.A(n_6814),
.Y(n_8774)
);

AOI22xp33_ASAP7_75t_L g8775 ( 
.A1(n_7341),
.A2(n_6088),
.B1(n_6014),
.B2(n_6026),
.Y(n_8775)
);

NOR2xp33_ASAP7_75t_L g8776 ( 
.A(n_6966),
.B(n_5879),
.Y(n_8776)
);

AND2x2_ASAP7_75t_L g8777 ( 
.A(n_6949),
.B(n_6349),
.Y(n_8777)
);

INVx1_ASAP7_75t_L g8778 ( 
.A(n_6814),
.Y(n_8778)
);

OAI21x1_ASAP7_75t_L g8779 ( 
.A1(n_7198),
.A2(n_5842),
.B(n_5791),
.Y(n_8779)
);

INVx1_ASAP7_75t_L g8780 ( 
.A(n_6817),
.Y(n_8780)
);

A2O1A1Ixp33_ASAP7_75t_L g8781 ( 
.A1(n_6800),
.A2(n_6014),
.B(n_6026),
.C(n_6012),
.Y(n_8781)
);

INVx2_ASAP7_75t_L g8782 ( 
.A(n_6744),
.Y(n_8782)
);

AND2x2_ASAP7_75t_L g8783 ( 
.A(n_6949),
.B(n_6967),
.Y(n_8783)
);

OAI21x1_ASAP7_75t_L g8784 ( 
.A1(n_7198),
.A2(n_5842),
.B(n_5791),
.Y(n_8784)
);

HB1xp67_ASAP7_75t_L g8785 ( 
.A(n_6642),
.Y(n_8785)
);

INVx1_ASAP7_75t_L g8786 ( 
.A(n_6817),
.Y(n_8786)
);

INVx1_ASAP7_75t_L g8787 ( 
.A(n_6817),
.Y(n_8787)
);

AOI221xp5_ASAP7_75t_L g8788 ( 
.A1(n_6925),
.A2(n_6128),
.B1(n_6146),
.B2(n_6114),
.C(n_6109),
.Y(n_8788)
);

NOR2xp33_ASAP7_75t_R g8789 ( 
.A(n_6951),
.B(n_5684),
.Y(n_8789)
);

OAI21x1_ASAP7_75t_SL g8790 ( 
.A1(n_7474),
.A2(n_5652),
.B(n_5627),
.Y(n_8790)
);

BUFx3_ASAP7_75t_L g8791 ( 
.A(n_6655),
.Y(n_8791)
);

OR2x6_ASAP7_75t_L g8792 ( 
.A(n_6668),
.B(n_6433),
.Y(n_8792)
);

AND2x2_ASAP7_75t_L g8793 ( 
.A(n_6949),
.B(n_6349),
.Y(n_8793)
);

AND2x2_ASAP7_75t_L g8794 ( 
.A(n_6949),
.B(n_6369),
.Y(n_8794)
);

INVx2_ASAP7_75t_L g8795 ( 
.A(n_6744),
.Y(n_8795)
);

HB1xp67_ASAP7_75t_L g8796 ( 
.A(n_7225),
.Y(n_8796)
);

NAND2xp5_ASAP7_75t_L g8797 ( 
.A(n_7111),
.B(n_6165),
.Y(n_8797)
);

INVx5_ASAP7_75t_L g8798 ( 
.A(n_7103),
.Y(n_8798)
);

OAI222xp33_ASAP7_75t_L g8799 ( 
.A1(n_7048),
.A2(n_6273),
.B1(n_6287),
.B2(n_6277),
.C1(n_5804),
.C2(n_5882),
.Y(n_8799)
);

OR2x2_ASAP7_75t_L g8800 ( 
.A(n_7205),
.B(n_6314),
.Y(n_8800)
);

OAI22xp5_ASAP7_75t_L g8801 ( 
.A1(n_7300),
.A2(n_4769),
.B1(n_6287),
.B2(n_6273),
.Y(n_8801)
);

AND2x2_ASAP7_75t_L g8802 ( 
.A(n_6967),
.B(n_6369),
.Y(n_8802)
);

OAI21x1_ASAP7_75t_L g8803 ( 
.A1(n_7371),
.A2(n_5865),
.B(n_5842),
.Y(n_8803)
);

OAI21x1_ASAP7_75t_L g8804 ( 
.A1(n_7371),
.A2(n_5902),
.B(n_5865),
.Y(n_8804)
);

HB1xp67_ASAP7_75t_L g8805 ( 
.A(n_7225),
.Y(n_8805)
);

AO32x2_ASAP7_75t_L g8806 ( 
.A1(n_7154),
.A2(n_6157),
.A3(n_6185),
.B1(n_6123),
.B2(n_6096),
.Y(n_8806)
);

INVxp67_ASAP7_75t_L g8807 ( 
.A(n_7589),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_6822),
.Y(n_8808)
);

OAI21xp5_ASAP7_75t_L g8809 ( 
.A1(n_7158),
.A2(n_6146),
.B(n_6128),
.Y(n_8809)
);

OAI21x1_ASAP7_75t_L g8810 ( 
.A1(n_7371),
.A2(n_5902),
.B(n_5865),
.Y(n_8810)
);

O2A1O1Ixp33_ASAP7_75t_L g8811 ( 
.A1(n_7182),
.A2(n_5318),
.B(n_5374),
.C(n_5203),
.Y(n_8811)
);

OAI21x1_ASAP7_75t_L g8812 ( 
.A1(n_7405),
.A2(n_5902),
.B(n_5865),
.Y(n_8812)
);

NOR2xp33_ASAP7_75t_L g8813 ( 
.A(n_6966),
.B(n_6968),
.Y(n_8813)
);

OAI21x1_ASAP7_75t_L g8814 ( 
.A1(n_7301),
.A2(n_5902),
.B(n_5865),
.Y(n_8814)
);

AOI21xp33_ASAP7_75t_L g8815 ( 
.A1(n_6684),
.A2(n_6762),
.B(n_6835),
.Y(n_8815)
);

OAI21xp5_ASAP7_75t_L g8816 ( 
.A1(n_6684),
.A2(n_6156),
.B(n_6149),
.Y(n_8816)
);

OR2x2_ASAP7_75t_L g8817 ( 
.A(n_7205),
.B(n_6329),
.Y(n_8817)
);

OR2x2_ASAP7_75t_L g8818 ( 
.A(n_7205),
.B(n_6329),
.Y(n_8818)
);

OAI21x1_ASAP7_75t_L g8819 ( 
.A1(n_7271),
.A2(n_5904),
.B(n_5902),
.Y(n_8819)
);

AOI22xp33_ASAP7_75t_L g8820 ( 
.A1(n_6765),
.A2(n_6088),
.B1(n_6026),
.B2(n_6042),
.Y(n_8820)
);

INVx1_ASAP7_75t_L g8821 ( 
.A(n_6822),
.Y(n_8821)
);

INVx3_ASAP7_75t_L g8822 ( 
.A(n_7103),
.Y(n_8822)
);

BUFx4f_ASAP7_75t_SL g8823 ( 
.A(n_6787),
.Y(n_8823)
);

INVxp67_ASAP7_75t_SL g8824 ( 
.A(n_7210),
.Y(n_8824)
);

NOR2xp33_ASAP7_75t_L g8825 ( 
.A(n_6968),
.B(n_6765),
.Y(n_8825)
);

OAI21x1_ASAP7_75t_L g8826 ( 
.A1(n_7347),
.A2(n_5907),
.B(n_5904),
.Y(n_8826)
);

INVx2_ASAP7_75t_SL g8827 ( 
.A(n_7103),
.Y(n_8827)
);

INVx1_ASAP7_75t_L g8828 ( 
.A(n_6822),
.Y(n_8828)
);

OAI21x1_ASAP7_75t_L g8829 ( 
.A1(n_7271),
.A2(n_5907),
.B(n_5904),
.Y(n_8829)
);

CKINVDCx9p33_ASAP7_75t_R g8830 ( 
.A(n_7460),
.Y(n_8830)
);

AND2x4_ASAP7_75t_L g8831 ( 
.A(n_7195),
.B(n_6384),
.Y(n_8831)
);

NAND2xp5_ASAP7_75t_L g8832 ( 
.A(n_7170),
.B(n_6165),
.Y(n_8832)
);

CKINVDCx11_ASAP7_75t_R g8833 ( 
.A(n_6787),
.Y(n_8833)
);

AOI22xp33_ASAP7_75t_L g8834 ( 
.A1(n_6921),
.A2(n_6088),
.B1(n_6026),
.B2(n_6042),
.Y(n_8834)
);

INVx1_ASAP7_75t_L g8835 ( 
.A(n_6829),
.Y(n_8835)
);

AO31x2_ASAP7_75t_L g8836 ( 
.A1(n_7524),
.A2(n_6378),
.A3(n_5992),
.B(n_6070),
.Y(n_8836)
);

NOR2x1_ASAP7_75t_SL g8837 ( 
.A(n_7226),
.B(n_6014),
.Y(n_8837)
);

A2O1A1Ixp33_ASAP7_75t_L g8838 ( 
.A1(n_6938),
.A2(n_6026),
.B(n_6042),
.C(n_6014),
.Y(n_8838)
);

O2A1O1Ixp33_ASAP7_75t_L g8839 ( 
.A1(n_7182),
.A2(n_5374),
.B(n_5318),
.C(n_6149),
.Y(n_8839)
);

NAND2xp5_ASAP7_75t_L g8840 ( 
.A(n_7170),
.B(n_6193),
.Y(n_8840)
);

OAI21x1_ASAP7_75t_L g8841 ( 
.A1(n_7271),
.A2(n_5907),
.B(n_5904),
.Y(n_8841)
);

OAI21xp5_ASAP7_75t_L g8842 ( 
.A1(n_6684),
.A2(n_6158),
.B(n_6156),
.Y(n_8842)
);

INVx1_ASAP7_75t_L g8843 ( 
.A(n_6829),
.Y(n_8843)
);

INVx1_ASAP7_75t_L g8844 ( 
.A(n_6829),
.Y(n_8844)
);

OAI21x1_ASAP7_75t_L g8845 ( 
.A1(n_7301),
.A2(n_5907),
.B(n_5904),
.Y(n_8845)
);

OA21x2_ASAP7_75t_L g8846 ( 
.A1(n_6685),
.A2(n_5701),
.B(n_5696),
.Y(n_8846)
);

INVx2_ASAP7_75t_L g8847 ( 
.A(n_6776),
.Y(n_8847)
);

OAI21x1_ASAP7_75t_L g8848 ( 
.A1(n_7301),
.A2(n_7347),
.B(n_7271),
.Y(n_8848)
);

BUFx3_ASAP7_75t_L g8849 ( 
.A(n_6655),
.Y(n_8849)
);

OAI222xp33_ASAP7_75t_L g8850 ( 
.A1(n_7326),
.A2(n_6273),
.B1(n_6287),
.B2(n_6277),
.C1(n_5804),
.C2(n_5882),
.Y(n_8850)
);

CKINVDCx6p67_ASAP7_75t_R g8851 ( 
.A(n_7348),
.Y(n_8851)
);

NAND2xp5_ASAP7_75t_SL g8852 ( 
.A(n_7590),
.B(n_6026),
.Y(n_8852)
);

OAI22xp5_ASAP7_75t_L g8853 ( 
.A1(n_7300),
.A2(n_4769),
.B1(n_4915),
.B2(n_4908),
.Y(n_8853)
);

INVx1_ASAP7_75t_L g8854 ( 
.A(n_6842),
.Y(n_8854)
);

HB1xp67_ASAP7_75t_L g8855 ( 
.A(n_7225),
.Y(n_8855)
);

AOI22xp33_ASAP7_75t_L g8856 ( 
.A1(n_6921),
.A2(n_6042),
.B1(n_6048),
.B2(n_6026),
.Y(n_8856)
);

INVx2_ASAP7_75t_R g8857 ( 
.A(n_7140),
.Y(n_8857)
);

AOI21x1_ASAP7_75t_L g8858 ( 
.A1(n_7110),
.A2(n_5992),
.B(n_5972),
.Y(n_8858)
);

OAI22x1_ASAP7_75t_L g8859 ( 
.A1(n_6960),
.A2(n_6191),
.B1(n_6079),
.B2(n_5992),
.Y(n_8859)
);

INVx1_ASAP7_75t_L g8860 ( 
.A(n_6842),
.Y(n_8860)
);

BUFx10_ASAP7_75t_L g8861 ( 
.A(n_6828),
.Y(n_8861)
);

AND2x4_ASAP7_75t_SL g8862 ( 
.A(n_6940),
.B(n_5831),
.Y(n_8862)
);

BUFx2_ASAP7_75t_L g8863 ( 
.A(n_7383),
.Y(n_8863)
);

CKINVDCx5p33_ASAP7_75t_R g8864 ( 
.A(n_7381),
.Y(n_8864)
);

INVx2_ASAP7_75t_L g8865 ( 
.A(n_6776),
.Y(n_8865)
);

INVx3_ASAP7_75t_L g8866 ( 
.A(n_7127),
.Y(n_8866)
);

INVxp33_ASAP7_75t_L g8867 ( 
.A(n_7486),
.Y(n_8867)
);

OR2x2_ASAP7_75t_L g8868 ( 
.A(n_7210),
.B(n_6336),
.Y(n_8868)
);

OAI21x1_ASAP7_75t_L g8869 ( 
.A1(n_7301),
.A2(n_5919),
.B(n_5907),
.Y(n_8869)
);

OAI21x1_ASAP7_75t_L g8870 ( 
.A1(n_7347),
.A2(n_5920),
.B(n_5919),
.Y(n_8870)
);

OAI21x1_ASAP7_75t_L g8871 ( 
.A1(n_7347),
.A2(n_5920),
.B(n_5919),
.Y(n_8871)
);

OAI21xp33_ASAP7_75t_SL g8872 ( 
.A1(n_7590),
.A2(n_6277),
.B(n_6123),
.Y(n_8872)
);

AND2x2_ASAP7_75t_L g8873 ( 
.A(n_6967),
.B(n_6369),
.Y(n_8873)
);

AND2x2_ASAP7_75t_L g8874 ( 
.A(n_6967),
.B(n_6435),
.Y(n_8874)
);

BUFx2_ASAP7_75t_L g8875 ( 
.A(n_7383),
.Y(n_8875)
);

INVx2_ASAP7_75t_SL g8876 ( 
.A(n_7127),
.Y(n_8876)
);

OAI21x1_ASAP7_75t_L g8877 ( 
.A1(n_7379),
.A2(n_7405),
.B(n_7258),
.Y(n_8877)
);

O2A1O1Ixp33_ASAP7_75t_SL g8878 ( 
.A1(n_6858),
.A2(n_6166),
.B(n_6181),
.C(n_6158),
.Y(n_8878)
);

AND2x2_ASAP7_75t_L g8879 ( 
.A(n_7034),
.B(n_6435),
.Y(n_8879)
);

OAI21x1_ASAP7_75t_L g8880 ( 
.A1(n_7379),
.A2(n_5920),
.B(n_5919),
.Y(n_8880)
);

OAI21x1_ASAP7_75t_L g8881 ( 
.A1(n_7379),
.A2(n_5920),
.B(n_5919),
.Y(n_8881)
);

AOI221xp5_ASAP7_75t_L g8882 ( 
.A1(n_7290),
.A2(n_6186),
.B1(n_6210),
.B2(n_6181),
.C(n_6166),
.Y(n_8882)
);

AOI22xp33_ASAP7_75t_SL g8883 ( 
.A1(n_7590),
.A2(n_6461),
.B1(n_6088),
.B2(n_6042),
.Y(n_8883)
);

NOR2xp33_ASAP7_75t_L g8884 ( 
.A(n_6968),
.B(n_5882),
.Y(n_8884)
);

OAI21x1_ASAP7_75t_L g8885 ( 
.A1(n_7379),
.A2(n_7405),
.B(n_7258),
.Y(n_8885)
);

OAI21xp5_ASAP7_75t_L g8886 ( 
.A1(n_6762),
.A2(n_6210),
.B(n_6186),
.Y(n_8886)
);

XOR2xp5_ASAP7_75t_L g8887 ( 
.A(n_7108),
.B(n_6549),
.Y(n_8887)
);

BUFx12f_ASAP7_75t_L g8888 ( 
.A(n_7284),
.Y(n_8888)
);

OA21x2_ASAP7_75t_L g8889 ( 
.A1(n_6685),
.A2(n_5701),
.B(n_5696),
.Y(n_8889)
);

OR2x6_ASAP7_75t_L g8890 ( 
.A(n_6668),
.B(n_6433),
.Y(n_8890)
);

O2A1O1Ixp5_ASAP7_75t_L g8891 ( 
.A1(n_7326),
.A2(n_5770),
.B(n_5817),
.C(n_5695),
.Y(n_8891)
);

BUFx12f_ASAP7_75t_L g8892 ( 
.A(n_7284),
.Y(n_8892)
);

OA21x2_ASAP7_75t_L g8893 ( 
.A1(n_6697),
.A2(n_5720),
.B(n_5711),
.Y(n_8893)
);

NAND2x1_ASAP7_75t_L g8894 ( 
.A(n_6655),
.B(n_6026),
.Y(n_8894)
);

AO31x2_ASAP7_75t_L g8895 ( 
.A1(n_7524),
.A2(n_6079),
.A3(n_6099),
.B(n_6070),
.Y(n_8895)
);

BUFx10_ASAP7_75t_L g8896 ( 
.A(n_6828),
.Y(n_8896)
);

AOI22xp33_ASAP7_75t_L g8897 ( 
.A1(n_7290),
.A2(n_6082),
.B1(n_6088),
.B2(n_6048),
.Y(n_8897)
);

OR2x6_ASAP7_75t_L g8898 ( 
.A(n_6668),
.B(n_6433),
.Y(n_8898)
);

OAI21xp5_ASAP7_75t_L g8899 ( 
.A1(n_6762),
.A2(n_6219),
.B(n_6218),
.Y(n_8899)
);

INVx2_ASAP7_75t_L g8900 ( 
.A(n_6776),
.Y(n_8900)
);

INVx8_ASAP7_75t_L g8901 ( 
.A(n_7014),
.Y(n_8901)
);

HB1xp67_ASAP7_75t_L g8902 ( 
.A(n_7247),
.Y(n_8902)
);

INVx2_ASAP7_75t_SL g8903 ( 
.A(n_7127),
.Y(n_8903)
);

OR2x2_ASAP7_75t_L g8904 ( 
.A(n_7210),
.B(n_7250),
.Y(n_8904)
);

NAND2xp5_ASAP7_75t_L g8905 ( 
.A(n_7170),
.B(n_6193),
.Y(n_8905)
);

INVx1_ASAP7_75t_L g8906 ( 
.A(n_6842),
.Y(n_8906)
);

INVxp67_ASAP7_75t_L g8907 ( 
.A(n_7593),
.Y(n_8907)
);

NAND2xp5_ASAP7_75t_L g8908 ( 
.A(n_6761),
.B(n_6256),
.Y(n_8908)
);

AND2x2_ASAP7_75t_SL g8909 ( 
.A(n_6976),
.B(n_6048),
.Y(n_8909)
);

AND2x4_ASAP7_75t_L g8910 ( 
.A(n_7195),
.B(n_6384),
.Y(n_8910)
);

BUFx12f_ASAP7_75t_L g8911 ( 
.A(n_7312),
.Y(n_8911)
);

INVx2_ASAP7_75t_SL g8912 ( 
.A(n_7127),
.Y(n_8912)
);

AOI22xp33_ASAP7_75t_SL g8913 ( 
.A1(n_7071),
.A2(n_6082),
.B1(n_6088),
.B2(n_6048),
.Y(n_8913)
);

OAI21x1_ASAP7_75t_SL g8914 ( 
.A1(n_7474),
.A2(n_5652),
.B(n_5627),
.Y(n_8914)
);

INVx1_ASAP7_75t_SL g8915 ( 
.A(n_7382),
.Y(n_8915)
);

NAND2xp5_ASAP7_75t_L g8916 ( 
.A(n_6761),
.B(n_6256),
.Y(n_8916)
);

CKINVDCx11_ASAP7_75t_R g8917 ( 
.A(n_6858),
.Y(n_8917)
);

AOI22xp33_ASAP7_75t_L g8918 ( 
.A1(n_7360),
.A2(n_6082),
.B1(n_6088),
.B2(n_6048),
.Y(n_8918)
);

AOI21xp5_ASAP7_75t_L g8919 ( 
.A1(n_7162),
.A2(n_7327),
.B(n_7376),
.Y(n_8919)
);

INVx2_ASAP7_75t_L g8920 ( 
.A(n_6776),
.Y(n_8920)
);

AND2x2_ASAP7_75t_L g8921 ( 
.A(n_7034),
.B(n_7115),
.Y(n_8921)
);

OA21x2_ASAP7_75t_L g8922 ( 
.A1(n_6697),
.A2(n_5720),
.B(n_5711),
.Y(n_8922)
);

INVx2_ASAP7_75t_L g8923 ( 
.A(n_6801),
.Y(n_8923)
);

NAND3xp33_ASAP7_75t_L g8924 ( 
.A(n_7299),
.B(n_6082),
.C(n_6048),
.Y(n_8924)
);

NAND2x1p5_ASAP7_75t_L g8925 ( 
.A(n_6923),
.B(n_5930),
.Y(n_8925)
);

OAI21x1_ASAP7_75t_L g8926 ( 
.A1(n_7405),
.A2(n_5941),
.B(n_5920),
.Y(n_8926)
);

INVx1_ASAP7_75t_L g8927 ( 
.A(n_6844),
.Y(n_8927)
);

OAI21x1_ASAP7_75t_L g8928 ( 
.A1(n_7106),
.A2(n_5941),
.B(n_5612),
.Y(n_8928)
);

OAI22xp5_ASAP7_75t_L g8929 ( 
.A1(n_7295),
.A2(n_4915),
.B1(n_4919),
.B2(n_4908),
.Y(n_8929)
);

INVx1_ASAP7_75t_L g8930 ( 
.A(n_6844),
.Y(n_8930)
);

NAND3xp33_ASAP7_75t_L g8931 ( 
.A(n_7299),
.B(n_7272),
.C(n_7070),
.Y(n_8931)
);

OAI21x1_ASAP7_75t_L g8932 ( 
.A1(n_7106),
.A2(n_5941),
.B(n_5612),
.Y(n_8932)
);

INVx1_ASAP7_75t_SL g8933 ( 
.A(n_7382),
.Y(n_8933)
);

OAI22xp5_ASAP7_75t_L g8934 ( 
.A1(n_7295),
.A2(n_4915),
.B1(n_4919),
.B2(n_4908),
.Y(n_8934)
);

INVx1_ASAP7_75t_L g8935 ( 
.A(n_6844),
.Y(n_8935)
);

INVx1_ASAP7_75t_L g8936 ( 
.A(n_6849),
.Y(n_8936)
);

CKINVDCx20_ASAP7_75t_R g8937 ( 
.A(n_7144),
.Y(n_8937)
);

CKINVDCx11_ASAP7_75t_R g8938 ( 
.A(n_7031),
.Y(n_8938)
);

BUFx2_ASAP7_75t_L g8939 ( 
.A(n_7383),
.Y(n_8939)
);

NAND2xp5_ASAP7_75t_L g8940 ( 
.A(n_6761),
.B(n_6342),
.Y(n_8940)
);

NOR2x1_ASAP7_75t_R g8941 ( 
.A(n_7348),
.B(n_6248),
.Y(n_8941)
);

AO32x2_ASAP7_75t_L g8942 ( 
.A1(n_7191),
.A2(n_6157),
.A3(n_6185),
.B1(n_6123),
.B2(n_6096),
.Y(n_8942)
);

OAI221xp5_ASAP7_75t_L g8943 ( 
.A1(n_7073),
.A2(n_6088),
.B1(n_6093),
.B2(n_6082),
.C(n_6048),
.Y(n_8943)
);

AOI21xp33_ASAP7_75t_L g8944 ( 
.A1(n_6835),
.A2(n_6868),
.B(n_6838),
.Y(n_8944)
);

INVx1_ASAP7_75t_L g8945 ( 
.A(n_6849),
.Y(n_8945)
);

OAI22xp5_ASAP7_75t_L g8946 ( 
.A1(n_7356),
.A2(n_4915),
.B1(n_4919),
.B2(n_4908),
.Y(n_8946)
);

BUFx6f_ASAP7_75t_L g8947 ( 
.A(n_7127),
.Y(n_8947)
);

OAI21xp5_ASAP7_75t_L g8948 ( 
.A1(n_7337),
.A2(n_6219),
.B(n_6218),
.Y(n_8948)
);

INVx1_ASAP7_75t_L g8949 ( 
.A(n_6849),
.Y(n_8949)
);

CKINVDCx20_ASAP7_75t_R g8950 ( 
.A(n_7144),
.Y(n_8950)
);

OAI21x1_ASAP7_75t_L g8951 ( 
.A1(n_7106),
.A2(n_5941),
.B(n_5612),
.Y(n_8951)
);

AND2x2_ASAP7_75t_L g8952 ( 
.A(n_7034),
.B(n_6435),
.Y(n_8952)
);

INVx2_ASAP7_75t_L g8953 ( 
.A(n_8759),
.Y(n_8953)
);

BUFx6f_ASAP7_75t_L g8954 ( 
.A(n_7803),
.Y(n_8954)
);

OR2x2_ASAP7_75t_L g8955 ( 
.A(n_7795),
.B(n_7215),
.Y(n_8955)
);

INVx1_ASAP7_75t_L g8956 ( 
.A(n_7820),
.Y(n_8956)
);

INVx2_ASAP7_75t_L g8957 ( 
.A(n_8759),
.Y(n_8957)
);

INVx1_ASAP7_75t_L g8958 ( 
.A(n_7820),
.Y(n_8958)
);

INVx6_ASAP7_75t_L g8959 ( 
.A(n_7704),
.Y(n_8959)
);

BUFx2_ASAP7_75t_L g8960 ( 
.A(n_7872),
.Y(n_8960)
);

INVx3_ASAP7_75t_L g8961 ( 
.A(n_7614),
.Y(n_8961)
);

OAI21x1_ASAP7_75t_L g8962 ( 
.A1(n_8566),
.A2(n_7292),
.B(n_7258),
.Y(n_8962)
);

AOI22xp33_ASAP7_75t_L g8963 ( 
.A1(n_7858),
.A2(n_7032),
.B1(n_7063),
.B2(n_7043),
.Y(n_8963)
);

INVx2_ASAP7_75t_L g8964 ( 
.A(n_8759),
.Y(n_8964)
);

CKINVDCx20_ASAP7_75t_R g8965 ( 
.A(n_8937),
.Y(n_8965)
);

NOR2x1_ASAP7_75t_SL g8966 ( 
.A(n_8273),
.B(n_7746),
.Y(n_8966)
);

INVxp33_ASAP7_75t_L g8967 ( 
.A(n_8789),
.Y(n_8967)
);

INVx1_ASAP7_75t_L g8968 ( 
.A(n_7824),
.Y(n_8968)
);

AOI222xp33_ASAP7_75t_L g8969 ( 
.A1(n_7631),
.A2(n_7360),
.B1(n_6981),
.B2(n_7244),
.C1(n_7010),
.C2(n_7073),
.Y(n_8969)
);

INVx1_ASAP7_75t_L g8970 ( 
.A(n_7824),
.Y(n_8970)
);

INVx1_ASAP7_75t_L g8971 ( 
.A(n_7830),
.Y(n_8971)
);

HB1xp67_ASAP7_75t_L g8972 ( 
.A(n_7716),
.Y(n_8972)
);

AND2x2_ASAP7_75t_L g8973 ( 
.A(n_7758),
.B(n_7343),
.Y(n_8973)
);

INVx3_ASAP7_75t_L g8974 ( 
.A(n_7614),
.Y(n_8974)
);

AOI22xp5_ASAP7_75t_L g8975 ( 
.A1(n_7633),
.A2(n_7010),
.B1(n_6981),
.B2(n_7071),
.Y(n_8975)
);

INVx1_ASAP7_75t_L g8976 ( 
.A(n_7830),
.Y(n_8976)
);

INVx2_ASAP7_75t_L g8977 ( 
.A(n_8759),
.Y(n_8977)
);

INVx1_ASAP7_75t_L g8978 ( 
.A(n_7846),
.Y(n_8978)
);

HB1xp67_ASAP7_75t_SL g8979 ( 
.A(n_7977),
.Y(n_8979)
);

INVx2_ASAP7_75t_L g8980 ( 
.A(n_8759),
.Y(n_8980)
);

OAI22xp33_ASAP7_75t_L g8981 ( 
.A1(n_7822),
.A2(n_6861),
.B1(n_7339),
.B2(n_7337),
.Y(n_8981)
);

INVxp33_ASAP7_75t_L g8982 ( 
.A(n_8789),
.Y(n_8982)
);

INVx1_ASAP7_75t_L g8983 ( 
.A(n_7846),
.Y(n_8983)
);

INVx1_ASAP7_75t_L g8984 ( 
.A(n_7848),
.Y(n_8984)
);

INVx1_ASAP7_75t_L g8985 ( 
.A(n_7848),
.Y(n_8985)
);

NAND2x1p5_ASAP7_75t_L g8986 ( 
.A(n_7693),
.B(n_6575),
.Y(n_8986)
);

INVx2_ASAP7_75t_L g8987 ( 
.A(n_8759),
.Y(n_8987)
);

AOI21xp5_ASAP7_75t_L g8988 ( 
.A1(n_7705),
.A2(n_7783),
.B(n_7707),
.Y(n_8988)
);

AOI22xp5_ASAP7_75t_L g8989 ( 
.A1(n_7633),
.A2(n_7010),
.B1(n_6981),
.B2(n_7071),
.Y(n_8989)
);

NAND2x1p5_ASAP7_75t_L g8990 ( 
.A(n_7693),
.B(n_6575),
.Y(n_8990)
);

HB1xp67_ASAP7_75t_L g8991 ( 
.A(n_7716),
.Y(n_8991)
);

INVx1_ASAP7_75t_L g8992 ( 
.A(n_7850),
.Y(n_8992)
);

INVx2_ASAP7_75t_L g8993 ( 
.A(n_8846),
.Y(n_8993)
);

INVx2_ASAP7_75t_L g8994 ( 
.A(n_8846),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_7850),
.Y(n_8995)
);

INVx2_ASAP7_75t_L g8996 ( 
.A(n_8846),
.Y(n_8996)
);

INVx3_ASAP7_75t_L g8997 ( 
.A(n_7614),
.Y(n_8997)
);

INVx4_ASAP7_75t_L g8998 ( 
.A(n_7704),
.Y(n_8998)
);

INVx1_ASAP7_75t_L g8999 ( 
.A(n_7851),
.Y(n_8999)
);

INVx1_ASAP7_75t_L g9000 ( 
.A(n_7851),
.Y(n_9000)
);

INVx1_ASAP7_75t_L g9001 ( 
.A(n_7854),
.Y(n_9001)
);

INVx1_ASAP7_75t_L g9002 ( 
.A(n_7854),
.Y(n_9002)
);

AOI22xp5_ASAP7_75t_L g9003 ( 
.A1(n_7631),
.A2(n_6970),
.B1(n_7319),
.B2(n_7337),
.Y(n_9003)
);

INVx2_ASAP7_75t_L g9004 ( 
.A(n_8846),
.Y(n_9004)
);

INVx2_ASAP7_75t_L g9005 ( 
.A(n_8846),
.Y(n_9005)
);

INVx2_ASAP7_75t_L g9006 ( 
.A(n_8846),
.Y(n_9006)
);

BUFx2_ASAP7_75t_L g9007 ( 
.A(n_7872),
.Y(n_9007)
);

AOI22xp33_ASAP7_75t_SL g9008 ( 
.A1(n_8288),
.A2(n_7392),
.B1(n_6991),
.B2(n_7039),
.Y(n_9008)
);

OAI22xp5_ASAP7_75t_L g9009 ( 
.A1(n_7691),
.A2(n_7759),
.B1(n_7808),
.B2(n_7678),
.Y(n_9009)
);

INVx2_ASAP7_75t_L g9010 ( 
.A(n_8889),
.Y(n_9010)
);

AND2x4_ASAP7_75t_L g9011 ( 
.A(n_8202),
.B(n_7195),
.Y(n_9011)
);

INVx1_ASAP7_75t_L g9012 ( 
.A(n_7873),
.Y(n_9012)
);

BUFx6f_ASAP7_75t_L g9013 ( 
.A(n_7704),
.Y(n_9013)
);

HB1xp67_ASAP7_75t_L g9014 ( 
.A(n_7727),
.Y(n_9014)
);

AND2x2_ASAP7_75t_L g9015 ( 
.A(n_7758),
.B(n_7343),
.Y(n_9015)
);

INVx2_ASAP7_75t_L g9016 ( 
.A(n_8889),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_7873),
.Y(n_9017)
);

INVx2_ASAP7_75t_L g9018 ( 
.A(n_8889),
.Y(n_9018)
);

OAI21x1_ASAP7_75t_L g9019 ( 
.A1(n_8566),
.A2(n_7292),
.B(n_7250),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_7878),
.Y(n_9020)
);

BUFx2_ASAP7_75t_SL g9021 ( 
.A(n_7640),
.Y(n_9021)
);

INVx1_ASAP7_75t_L g9022 ( 
.A(n_7878),
.Y(n_9022)
);

INVx2_ASAP7_75t_L g9023 ( 
.A(n_8889),
.Y(n_9023)
);

HB1xp67_ASAP7_75t_L g9024 ( 
.A(n_7727),
.Y(n_9024)
);

INVx1_ASAP7_75t_L g9025 ( 
.A(n_7880),
.Y(n_9025)
);

BUFx6f_ASAP7_75t_L g9026 ( 
.A(n_7704),
.Y(n_9026)
);

INVx1_ASAP7_75t_L g9027 ( 
.A(n_7880),
.Y(n_9027)
);

BUFx2_ASAP7_75t_R g9028 ( 
.A(n_8251),
.Y(n_9028)
);

INVx2_ASAP7_75t_SL g9029 ( 
.A(n_7902),
.Y(n_9029)
);

CKINVDCx5p33_ASAP7_75t_R g9030 ( 
.A(n_8026),
.Y(n_9030)
);

INVx1_ASAP7_75t_L g9031 ( 
.A(n_7883),
.Y(n_9031)
);

INVx1_ASAP7_75t_SL g9032 ( 
.A(n_8021),
.Y(n_9032)
);

BUFx6f_ASAP7_75t_L g9033 ( 
.A(n_7803),
.Y(n_9033)
);

NAND2xp5_ASAP7_75t_L g9034 ( 
.A(n_8813),
.B(n_7019),
.Y(n_9034)
);

CKINVDCx11_ASAP7_75t_R g9035 ( 
.A(n_8026),
.Y(n_9035)
);

INVx1_ASAP7_75t_L g9036 ( 
.A(n_7883),
.Y(n_9036)
);

AO21x2_ASAP7_75t_L g9037 ( 
.A1(n_7747),
.A2(n_7577),
.B(n_6675),
.Y(n_9037)
);

BUFx2_ASAP7_75t_L g9038 ( 
.A(n_7872),
.Y(n_9038)
);

HB1xp67_ASAP7_75t_L g9039 ( 
.A(n_7762),
.Y(n_9039)
);

OAI21x1_ASAP7_75t_L g9040 ( 
.A1(n_8566),
.A2(n_7292),
.B(n_7250),
.Y(n_9040)
);

INVx1_ASAP7_75t_L g9041 ( 
.A(n_7887),
.Y(n_9041)
);

AOI22xp33_ASAP7_75t_SL g9042 ( 
.A1(n_8288),
.A2(n_7392),
.B1(n_6991),
.B2(n_7039),
.Y(n_9042)
);

INVx1_ASAP7_75t_L g9043 ( 
.A(n_7887),
.Y(n_9043)
);

INVx6_ASAP7_75t_L g9044 ( 
.A(n_7803),
.Y(n_9044)
);

INVx1_ASAP7_75t_L g9045 ( 
.A(n_7891),
.Y(n_9045)
);

AOI22xp33_ASAP7_75t_L g9046 ( 
.A1(n_7858),
.A2(n_7043),
.B1(n_7063),
.B2(n_7032),
.Y(n_9046)
);

AND2x4_ASAP7_75t_L g9047 ( 
.A(n_8202),
.B(n_7195),
.Y(n_9047)
);

INVx1_ASAP7_75t_L g9048 ( 
.A(n_7891),
.Y(n_9048)
);

AOI222xp33_ASAP7_75t_L g9049 ( 
.A1(n_7678),
.A2(n_7392),
.B1(n_6970),
.B2(n_7272),
.C1(n_7188),
.C2(n_7206),
.Y(n_9049)
);

HB1xp67_ASAP7_75t_L g9050 ( 
.A(n_7762),
.Y(n_9050)
);

INVx2_ASAP7_75t_L g9051 ( 
.A(n_8889),
.Y(n_9051)
);

INVx1_ASAP7_75t_L g9052 ( 
.A(n_7893),
.Y(n_9052)
);

BUFx6f_ASAP7_75t_SL g9053 ( 
.A(n_7630),
.Y(n_9053)
);

BUFx6f_ASAP7_75t_SL g9054 ( 
.A(n_7630),
.Y(n_9054)
);

INVx1_ASAP7_75t_SL g9055 ( 
.A(n_8021),
.Y(n_9055)
);

INVx1_ASAP7_75t_L g9056 ( 
.A(n_7893),
.Y(n_9056)
);

INVx1_ASAP7_75t_L g9057 ( 
.A(n_7896),
.Y(n_9057)
);

INVx1_ASAP7_75t_L g9058 ( 
.A(n_7896),
.Y(n_9058)
);

OAI21xp5_ASAP7_75t_L g9059 ( 
.A1(n_7859),
.A2(n_7339),
.B(n_7319),
.Y(n_9059)
);

NAND2xp5_ASAP7_75t_L g9060 ( 
.A(n_8813),
.B(n_7019),
.Y(n_9060)
);

INVx1_ASAP7_75t_L g9061 ( 
.A(n_7909),
.Y(n_9061)
);

INVx2_ASAP7_75t_L g9062 ( 
.A(n_8889),
.Y(n_9062)
);

INVx2_ASAP7_75t_L g9063 ( 
.A(n_8893),
.Y(n_9063)
);

NAND2x1p5_ASAP7_75t_L g9064 ( 
.A(n_7616),
.B(n_6575),
.Y(n_9064)
);

INVx8_ASAP7_75t_L g9065 ( 
.A(n_7803),
.Y(n_9065)
);

CKINVDCx8_ASAP7_75t_R g9066 ( 
.A(n_7793),
.Y(n_9066)
);

OAI22xp5_ASAP7_75t_L g9067 ( 
.A1(n_7691),
.A2(n_6861),
.B1(n_7410),
.B2(n_7431),
.Y(n_9067)
);

INVx2_ASAP7_75t_SL g9068 ( 
.A(n_7902),
.Y(n_9068)
);

INVx1_ASAP7_75t_L g9069 ( 
.A(n_7909),
.Y(n_9069)
);

OR2x6_ASAP7_75t_L g9070 ( 
.A(n_7673),
.B(n_7110),
.Y(n_9070)
);

INVx2_ASAP7_75t_L g9071 ( 
.A(n_8893),
.Y(n_9071)
);

OA21x2_ASAP7_75t_L g9072 ( 
.A1(n_8399),
.A2(n_7334),
.B(n_7221),
.Y(n_9072)
);

AOI22xp33_ASAP7_75t_SL g9073 ( 
.A1(n_8288),
.A2(n_6991),
.B1(n_7039),
.B2(n_6989),
.Y(n_9073)
);

AOI21x1_ASAP7_75t_L g9074 ( 
.A1(n_8300),
.A2(n_6999),
.B(n_6983),
.Y(n_9074)
);

INVx1_ASAP7_75t_L g9075 ( 
.A(n_7910),
.Y(n_9075)
);

OAI22xp33_ASAP7_75t_L g9076 ( 
.A1(n_7822),
.A2(n_6861),
.B1(n_7339),
.B2(n_7313),
.Y(n_9076)
);

INVx2_ASAP7_75t_L g9077 ( 
.A(n_8893),
.Y(n_9077)
);

NAND2x1p5_ASAP7_75t_L g9078 ( 
.A(n_7616),
.B(n_6575),
.Y(n_9078)
);

AND2x2_ASAP7_75t_L g9079 ( 
.A(n_7758),
.B(n_7343),
.Y(n_9079)
);

INVx1_ASAP7_75t_L g9080 ( 
.A(n_7910),
.Y(n_9080)
);

CKINVDCx12_ASAP7_75t_R g9081 ( 
.A(n_8683),
.Y(n_9081)
);

INVx1_ASAP7_75t_L g9082 ( 
.A(n_7612),
.Y(n_9082)
);

INVx1_ASAP7_75t_L g9083 ( 
.A(n_7612),
.Y(n_9083)
);

INVx2_ASAP7_75t_L g9084 ( 
.A(n_8893),
.Y(n_9084)
);

INVx2_ASAP7_75t_L g9085 ( 
.A(n_8893),
.Y(n_9085)
);

BUFx6f_ASAP7_75t_L g9086 ( 
.A(n_8255),
.Y(n_9086)
);

AOI22xp33_ASAP7_75t_SL g9087 ( 
.A1(n_7764),
.A2(n_6991),
.B1(n_7039),
.B2(n_6989),
.Y(n_9087)
);

INVx1_ASAP7_75t_L g9088 ( 
.A(n_7624),
.Y(n_9088)
);

INVx2_ASAP7_75t_L g9089 ( 
.A(n_8893),
.Y(n_9089)
);

AO21x1_ASAP7_75t_SL g9090 ( 
.A1(n_8850),
.A2(n_7575),
.B(n_7557),
.Y(n_9090)
);

INVx1_ASAP7_75t_L g9091 ( 
.A(n_7624),
.Y(n_9091)
);

INVx1_ASAP7_75t_L g9092 ( 
.A(n_7625),
.Y(n_9092)
);

BUFx6f_ASAP7_75t_L g9093 ( 
.A(n_8255),
.Y(n_9093)
);

AOI22xp33_ASAP7_75t_L g9094 ( 
.A1(n_8647),
.A2(n_7859),
.B1(n_7847),
.B2(n_8131),
.Y(n_9094)
);

INVx1_ASAP7_75t_L g9095 ( 
.A(n_7625),
.Y(n_9095)
);

INVx3_ASAP7_75t_L g9096 ( 
.A(n_7614),
.Y(n_9096)
);

BUFx10_ASAP7_75t_L g9097 ( 
.A(n_8864),
.Y(n_9097)
);

INVx2_ASAP7_75t_L g9098 ( 
.A(n_8922),
.Y(n_9098)
);

INVx1_ASAP7_75t_L g9099 ( 
.A(n_7627),
.Y(n_9099)
);

INVx3_ASAP7_75t_L g9100 ( 
.A(n_7614),
.Y(n_9100)
);

INVx1_ASAP7_75t_L g9101 ( 
.A(n_7627),
.Y(n_9101)
);

INVx1_ASAP7_75t_L g9102 ( 
.A(n_7635),
.Y(n_9102)
);

BUFx2_ASAP7_75t_R g9103 ( 
.A(n_8251),
.Y(n_9103)
);

NOR2xp33_ASAP7_75t_L g9104 ( 
.A(n_7606),
.B(n_7351),
.Y(n_9104)
);

BUFx2_ASAP7_75t_R g9105 ( 
.A(n_8251),
.Y(n_9105)
);

CKINVDCx5p33_ASAP7_75t_R g9106 ( 
.A(n_8917),
.Y(n_9106)
);

INVx1_ASAP7_75t_L g9107 ( 
.A(n_7635),
.Y(n_9107)
);

INVx1_ASAP7_75t_L g9108 ( 
.A(n_7648),
.Y(n_9108)
);

BUFx12f_ASAP7_75t_L g9109 ( 
.A(n_8255),
.Y(n_9109)
);

HB1xp67_ASAP7_75t_L g9110 ( 
.A(n_7870),
.Y(n_9110)
);

AOI22xp33_ASAP7_75t_L g9111 ( 
.A1(n_8647),
.A2(n_7066),
.B1(n_6991),
.B2(n_7039),
.Y(n_9111)
);

AOI22xp33_ASAP7_75t_L g9112 ( 
.A1(n_7847),
.A2(n_7066),
.B1(n_6989),
.B2(n_7519),
.Y(n_9112)
);

INVx2_ASAP7_75t_L g9113 ( 
.A(n_8922),
.Y(n_9113)
);

AND2x2_ASAP7_75t_L g9114 ( 
.A(n_7613),
.B(n_7343),
.Y(n_9114)
);

INVx2_ASAP7_75t_SL g9115 ( 
.A(n_7902),
.Y(n_9115)
);

INVx1_ASAP7_75t_L g9116 ( 
.A(n_7648),
.Y(n_9116)
);

INVx1_ASAP7_75t_L g9117 ( 
.A(n_7656),
.Y(n_9117)
);

HB1xp67_ASAP7_75t_L g9118 ( 
.A(n_7870),
.Y(n_9118)
);

OAI21x1_ASAP7_75t_L g9119 ( 
.A1(n_8757),
.A2(n_7694),
.B(n_7676),
.Y(n_9119)
);

NAND2x1p5_ASAP7_75t_L g9120 ( 
.A(n_7616),
.B(n_6575),
.Y(n_9120)
);

INVx2_ASAP7_75t_L g9121 ( 
.A(n_8922),
.Y(n_9121)
);

AOI22xp33_ASAP7_75t_SL g9122 ( 
.A1(n_7764),
.A2(n_6989),
.B1(n_7206),
.B2(n_7188),
.Y(n_9122)
);

NAND2xp5_ASAP7_75t_L g9123 ( 
.A(n_7615),
.B(n_7317),
.Y(n_9123)
);

INVx3_ASAP7_75t_L g9124 ( 
.A(n_7614),
.Y(n_9124)
);

INVx1_ASAP7_75t_L g9125 ( 
.A(n_7656),
.Y(n_9125)
);

INVx2_ASAP7_75t_L g9126 ( 
.A(n_8922),
.Y(n_9126)
);

AND2x2_ASAP7_75t_L g9127 ( 
.A(n_7613),
.B(n_7617),
.Y(n_9127)
);

INVx3_ASAP7_75t_L g9128 ( 
.A(n_7614),
.Y(n_9128)
);

AOI22xp5_ASAP7_75t_L g9129 ( 
.A1(n_7636),
.A2(n_7431),
.B1(n_7441),
.B2(n_7523),
.Y(n_9129)
);

INVx2_ASAP7_75t_L g9130 ( 
.A(n_8922),
.Y(n_9130)
);

HB1xp67_ASAP7_75t_L g9131 ( 
.A(n_7954),
.Y(n_9131)
);

OAI22xp5_ASAP7_75t_L g9132 ( 
.A1(n_7759),
.A2(n_6861),
.B1(n_7410),
.B2(n_7441),
.Y(n_9132)
);

AOI22xp33_ASAP7_75t_L g9133 ( 
.A1(n_7847),
.A2(n_6989),
.B1(n_7537),
.B2(n_7519),
.Y(n_9133)
);

BUFx10_ASAP7_75t_L g9134 ( 
.A(n_8864),
.Y(n_9134)
);

INVx2_ASAP7_75t_L g9135 ( 
.A(n_8922),
.Y(n_9135)
);

AND2x4_ASAP7_75t_L g9136 ( 
.A(n_8202),
.B(n_7195),
.Y(n_9136)
);

INVx1_ASAP7_75t_L g9137 ( 
.A(n_7661),
.Y(n_9137)
);

INVx1_ASAP7_75t_L g9138 ( 
.A(n_7661),
.Y(n_9138)
);

INVx3_ASAP7_75t_L g9139 ( 
.A(n_7614),
.Y(n_9139)
);

NAND2xp5_ASAP7_75t_L g9140 ( 
.A(n_7615),
.B(n_7317),
.Y(n_9140)
);

INVx1_ASAP7_75t_L g9141 ( 
.A(n_7667),
.Y(n_9141)
);

INVx2_ASAP7_75t_L g9142 ( 
.A(n_8568),
.Y(n_9142)
);

AOI22xp33_ASAP7_75t_L g9143 ( 
.A1(n_7847),
.A2(n_7537),
.B1(n_6265),
.B2(n_6246),
.Y(n_9143)
);

INVx2_ASAP7_75t_L g9144 ( 
.A(n_8568),
.Y(n_9144)
);

AO21x2_ASAP7_75t_L g9145 ( 
.A1(n_7747),
.A2(n_7577),
.B(n_6675),
.Y(n_9145)
);

INVx2_ASAP7_75t_L g9146 ( 
.A(n_8568),
.Y(n_9146)
);

HB1xp67_ASAP7_75t_L g9147 ( 
.A(n_7954),
.Y(n_9147)
);

BUFx2_ASAP7_75t_L g9148 ( 
.A(n_7872),
.Y(n_9148)
);

INVx1_ASAP7_75t_L g9149 ( 
.A(n_7667),
.Y(n_9149)
);

INVx8_ASAP7_75t_L g9150 ( 
.A(n_8255),
.Y(n_9150)
);

AND2x2_ASAP7_75t_L g9151 ( 
.A(n_7613),
.B(n_7349),
.Y(n_9151)
);

BUFx6f_ASAP7_75t_L g9152 ( 
.A(n_8582),
.Y(n_9152)
);

INVx3_ASAP7_75t_L g9153 ( 
.A(n_7814),
.Y(n_9153)
);

INVx3_ASAP7_75t_L g9154 ( 
.A(n_7814),
.Y(n_9154)
);

INVx3_ASAP7_75t_L g9155 ( 
.A(n_7814),
.Y(n_9155)
);

INVx2_ASAP7_75t_SL g9156 ( 
.A(n_7902),
.Y(n_9156)
);

INVx1_ASAP7_75t_L g9157 ( 
.A(n_7690),
.Y(n_9157)
);

AOI22xp33_ASAP7_75t_L g9158 ( 
.A1(n_7847),
.A2(n_6265),
.B1(n_6246),
.B2(n_7162),
.Y(n_9158)
);

BUFx2_ASAP7_75t_L g9159 ( 
.A(n_7872),
.Y(n_9159)
);

INVx1_ASAP7_75t_L g9160 ( 
.A(n_7690),
.Y(n_9160)
);

BUFx2_ASAP7_75t_L g9161 ( 
.A(n_7872),
.Y(n_9161)
);

INVx1_ASAP7_75t_L g9162 ( 
.A(n_7703),
.Y(n_9162)
);

INVx2_ASAP7_75t_L g9163 ( 
.A(n_8568),
.Y(n_9163)
);

HB1xp67_ASAP7_75t_L g9164 ( 
.A(n_8058),
.Y(n_9164)
);

NAND2xp5_ASAP7_75t_L g9165 ( 
.A(n_8825),
.B(n_6657),
.Y(n_9165)
);

HB1xp67_ASAP7_75t_L g9166 ( 
.A(n_8058),
.Y(n_9166)
);

CKINVDCx20_ASAP7_75t_R g9167 ( 
.A(n_8937),
.Y(n_9167)
);

OA21x2_ASAP7_75t_L g9168 ( 
.A1(n_8399),
.A2(n_7334),
.B(n_7221),
.Y(n_9168)
);

INVx1_ASAP7_75t_L g9169 ( 
.A(n_7703),
.Y(n_9169)
);

OAI21x1_ASAP7_75t_L g9170 ( 
.A1(n_8757),
.A2(n_7250),
.B(n_7210),
.Y(n_9170)
);

INVx1_ASAP7_75t_L g9171 ( 
.A(n_7714),
.Y(n_9171)
);

HB1xp67_ASAP7_75t_L g9172 ( 
.A(n_8259),
.Y(n_9172)
);

INVx1_ASAP7_75t_L g9173 ( 
.A(n_7714),
.Y(n_9173)
);

CKINVDCx11_ASAP7_75t_R g9174 ( 
.A(n_8117),
.Y(n_9174)
);

INVx1_ASAP7_75t_L g9175 ( 
.A(n_7725),
.Y(n_9175)
);

INVx2_ASAP7_75t_L g9176 ( 
.A(n_8568),
.Y(n_9176)
);

INVx1_ASAP7_75t_L g9177 ( 
.A(n_7725),
.Y(n_9177)
);

INVx1_ASAP7_75t_L g9178 ( 
.A(n_7726),
.Y(n_9178)
);

OAI22x1_ASAP7_75t_L g9179 ( 
.A1(n_7838),
.A2(n_7113),
.B1(n_7575),
.B2(n_7557),
.Y(n_9179)
);

AO21x1_ASAP7_75t_L g9180 ( 
.A1(n_7837),
.A2(n_7562),
.B(n_7524),
.Y(n_9180)
);

INVxp67_ASAP7_75t_L g9181 ( 
.A(n_8086),
.Y(n_9181)
);

OAI21x1_ASAP7_75t_L g9182 ( 
.A1(n_8757),
.A2(n_7562),
.B(n_6601),
.Y(n_9182)
);

INVx3_ASAP7_75t_L g9183 ( 
.A(n_7814),
.Y(n_9183)
);

BUFx2_ASAP7_75t_L g9184 ( 
.A(n_8184),
.Y(n_9184)
);

CKINVDCx11_ASAP7_75t_R g9185 ( 
.A(n_8117),
.Y(n_9185)
);

INVx1_ASAP7_75t_L g9186 ( 
.A(n_7726),
.Y(n_9186)
);

AOI22xp33_ASAP7_75t_L g9187 ( 
.A1(n_7847),
.A2(n_6265),
.B1(n_6246),
.B2(n_7162),
.Y(n_9187)
);

INVx1_ASAP7_75t_L g9188 ( 
.A(n_7735),
.Y(n_9188)
);

INVx1_ASAP7_75t_L g9189 ( 
.A(n_7735),
.Y(n_9189)
);

INVx1_ASAP7_75t_L g9190 ( 
.A(n_7740),
.Y(n_9190)
);

BUFx2_ASAP7_75t_R g9191 ( 
.A(n_8497),
.Y(n_9191)
);

INVx2_ASAP7_75t_L g9192 ( 
.A(n_8568),
.Y(n_9192)
);

NOR2x1_ASAP7_75t_R g9193 ( 
.A(n_8582),
.B(n_7351),
.Y(n_9193)
);

INVx3_ASAP7_75t_L g9194 ( 
.A(n_7814),
.Y(n_9194)
);

INVx1_ASAP7_75t_L g9195 ( 
.A(n_7740),
.Y(n_9195)
);

BUFx10_ASAP7_75t_L g9196 ( 
.A(n_7731),
.Y(n_9196)
);

INVx1_ASAP7_75t_L g9197 ( 
.A(n_7743),
.Y(n_9197)
);

HB1xp67_ASAP7_75t_L g9198 ( 
.A(n_8259),
.Y(n_9198)
);

AND2x4_ASAP7_75t_L g9199 ( 
.A(n_8202),
.B(n_7330),
.Y(n_9199)
);

BUFx3_ASAP7_75t_L g9200 ( 
.A(n_8582),
.Y(n_9200)
);

OAI22xp33_ASAP7_75t_L g9201 ( 
.A1(n_7765),
.A2(n_7313),
.B1(n_7575),
.B2(n_7557),
.Y(n_9201)
);

INVxp67_ASAP7_75t_L g9202 ( 
.A(n_8086),
.Y(n_9202)
);

INVx2_ASAP7_75t_L g9203 ( 
.A(n_8586),
.Y(n_9203)
);

AND2x2_ASAP7_75t_L g9204 ( 
.A(n_7613),
.B(n_7349),
.Y(n_9204)
);

INVx1_ASAP7_75t_L g9205 ( 
.A(n_7699),
.Y(n_9205)
);

INVx6_ASAP7_75t_L g9206 ( 
.A(n_8582),
.Y(n_9206)
);

INVx1_ASAP7_75t_L g9207 ( 
.A(n_7699),
.Y(n_9207)
);

INVx1_ASAP7_75t_L g9208 ( 
.A(n_7743),
.Y(n_9208)
);

INVx1_ASAP7_75t_L g9209 ( 
.A(n_7773),
.Y(n_9209)
);

BUFx2_ASAP7_75t_SL g9210 ( 
.A(n_7640),
.Y(n_9210)
);

INVx1_ASAP7_75t_L g9211 ( 
.A(n_7773),
.Y(n_9211)
);

OAI22xp5_ASAP7_75t_L g9212 ( 
.A1(n_7808),
.A2(n_6695),
.B1(n_6696),
.B2(n_6681),
.Y(n_9212)
);

OAI22xp33_ASAP7_75t_L g9213 ( 
.A1(n_7765),
.A2(n_7313),
.B1(n_7114),
.B2(n_7118),
.Y(n_9213)
);

OAI22xp33_ASAP7_75t_L g9214 ( 
.A1(n_7855),
.A2(n_7114),
.B1(n_7118),
.B2(n_7097),
.Y(n_9214)
);

INVx1_ASAP7_75t_L g9215 ( 
.A(n_7774),
.Y(n_9215)
);

AND2x2_ASAP7_75t_L g9216 ( 
.A(n_7617),
.B(n_7349),
.Y(n_9216)
);

INVx1_ASAP7_75t_L g9217 ( 
.A(n_7774),
.Y(n_9217)
);

OAI21x1_ASAP7_75t_L g9218 ( 
.A1(n_7676),
.A2(n_7562),
.B(n_6601),
.Y(n_9218)
);

INVx1_ASAP7_75t_L g9219 ( 
.A(n_7785),
.Y(n_9219)
);

INVx1_ASAP7_75t_L g9220 ( 
.A(n_7785),
.Y(n_9220)
);

INVx2_ASAP7_75t_L g9221 ( 
.A(n_8586),
.Y(n_9221)
);

INVx1_ASAP7_75t_L g9222 ( 
.A(n_7796),
.Y(n_9222)
);

BUFx3_ASAP7_75t_L g9223 ( 
.A(n_8632),
.Y(n_9223)
);

OAI22xp33_ASAP7_75t_L g9224 ( 
.A1(n_7855),
.A2(n_7636),
.B1(n_7709),
.B2(n_7729),
.Y(n_9224)
);

NAND2xp5_ASAP7_75t_L g9225 ( 
.A(n_8825),
.B(n_8944),
.Y(n_9225)
);

AOI22xp33_ASAP7_75t_L g9226 ( 
.A1(n_8131),
.A2(n_6265),
.B1(n_6246),
.B2(n_7162),
.Y(n_9226)
);

AND2x4_ASAP7_75t_L g9227 ( 
.A(n_8202),
.B(n_7330),
.Y(n_9227)
);

AND2x2_ASAP7_75t_L g9228 ( 
.A(n_7617),
.B(n_7349),
.Y(n_9228)
);

INVx3_ASAP7_75t_L g9229 ( 
.A(n_7814),
.Y(n_9229)
);

INVx1_ASAP7_75t_L g9230 ( 
.A(n_7757),
.Y(n_9230)
);

INVx1_ASAP7_75t_L g9231 ( 
.A(n_7757),
.Y(n_9231)
);

INVx2_ASAP7_75t_L g9232 ( 
.A(n_8586),
.Y(n_9232)
);

INVx4_ASAP7_75t_SL g9233 ( 
.A(n_8208),
.Y(n_9233)
);

INVx2_ASAP7_75t_L g9234 ( 
.A(n_8586),
.Y(n_9234)
);

INVx1_ASAP7_75t_L g9235 ( 
.A(n_7796),
.Y(n_9235)
);

OAI21x1_ASAP7_75t_L g9236 ( 
.A1(n_7676),
.A2(n_7694),
.B(n_8735),
.Y(n_9236)
);

INVx2_ASAP7_75t_L g9237 ( 
.A(n_8586),
.Y(n_9237)
);

OAI22xp5_ASAP7_75t_L g9238 ( 
.A1(n_8116),
.A2(n_6695),
.B1(n_6696),
.B2(n_6681),
.Y(n_9238)
);

AO21x1_ASAP7_75t_SL g9239 ( 
.A1(n_8850),
.A2(n_7183),
.B(n_7594),
.Y(n_9239)
);

INVx2_ASAP7_75t_L g9240 ( 
.A(n_8586),
.Y(n_9240)
);

INVx2_ASAP7_75t_SL g9241 ( 
.A(n_7943),
.Y(n_9241)
);

CKINVDCx16_ASAP7_75t_R g9242 ( 
.A(n_8471),
.Y(n_9242)
);

BUFx12f_ASAP7_75t_L g9243 ( 
.A(n_8632),
.Y(n_9243)
);

INVx2_ASAP7_75t_L g9244 ( 
.A(n_8595),
.Y(n_9244)
);

INVx3_ASAP7_75t_L g9245 ( 
.A(n_7814),
.Y(n_9245)
);

INVx2_ASAP7_75t_L g9246 ( 
.A(n_8595),
.Y(n_9246)
);

AO21x2_ASAP7_75t_L g9247 ( 
.A1(n_7747),
.A2(n_7577),
.B(n_6675),
.Y(n_9247)
);

NAND2xp5_ASAP7_75t_L g9248 ( 
.A(n_8944),
.B(n_6657),
.Y(n_9248)
);

OAI22xp5_ASAP7_75t_L g9249 ( 
.A1(n_8116),
.A2(n_6695),
.B1(n_6696),
.B2(n_6681),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_7806),
.Y(n_9250)
);

INVx1_ASAP7_75t_L g9251 ( 
.A(n_7806),
.Y(n_9251)
);

INVx1_ASAP7_75t_L g9252 ( 
.A(n_8331),
.Y(n_9252)
);

OAI21x1_ASAP7_75t_L g9253 ( 
.A1(n_7694),
.A2(n_6601),
.B(n_6566),
.Y(n_9253)
);

AND2x4_ASAP7_75t_L g9254 ( 
.A(n_8202),
.B(n_7330),
.Y(n_9254)
);

OAI21x1_ASAP7_75t_SL g9255 ( 
.A1(n_8053),
.A2(n_7477),
.B(n_7183),
.Y(n_9255)
);

INVx2_ASAP7_75t_L g9256 ( 
.A(n_8595),
.Y(n_9256)
);

INVx4_ASAP7_75t_SL g9257 ( 
.A(n_8208),
.Y(n_9257)
);

INVx2_ASAP7_75t_L g9258 ( 
.A(n_8595),
.Y(n_9258)
);

INVx2_ASAP7_75t_L g9259 ( 
.A(n_8595),
.Y(n_9259)
);

HB1xp67_ASAP7_75t_L g9260 ( 
.A(n_8313),
.Y(n_9260)
);

AO21x1_ASAP7_75t_SL g9261 ( 
.A1(n_7709),
.A2(n_7594),
.B(n_7097),
.Y(n_9261)
);

INVx3_ASAP7_75t_L g9262 ( 
.A(n_7814),
.Y(n_9262)
);

INVx1_ASAP7_75t_L g9263 ( 
.A(n_8331),
.Y(n_9263)
);

CKINVDCx5p33_ASAP7_75t_R g9264 ( 
.A(n_8917),
.Y(n_9264)
);

INVx1_ASAP7_75t_L g9265 ( 
.A(n_8332),
.Y(n_9265)
);

INVx2_ASAP7_75t_L g9266 ( 
.A(n_8595),
.Y(n_9266)
);

CKINVDCx5p33_ASAP7_75t_R g9267 ( 
.A(n_8938),
.Y(n_9267)
);

OAI22xp33_ASAP7_75t_L g9268 ( 
.A1(n_7729),
.A2(n_7114),
.B1(n_7118),
.B2(n_7097),
.Y(n_9268)
);

AOI22xp33_ASAP7_75t_L g9269 ( 
.A1(n_8363),
.A2(n_6265),
.B1(n_7327),
.B2(n_7162),
.Y(n_9269)
);

INVx1_ASAP7_75t_L g9270 ( 
.A(n_8332),
.Y(n_9270)
);

AOI22xp33_ASAP7_75t_SL g9271 ( 
.A1(n_7812),
.A2(n_7494),
.B1(n_7204),
.B2(n_7302),
.Y(n_9271)
);

AOI21x1_ASAP7_75t_L g9272 ( 
.A1(n_8300),
.A2(n_6999),
.B(n_6983),
.Y(n_9272)
);

BUFx12f_ASAP7_75t_L g9273 ( 
.A(n_8632),
.Y(n_9273)
);

OAI21x1_ASAP7_75t_L g9274 ( 
.A1(n_8735),
.A2(n_6601),
.B(n_6566),
.Y(n_9274)
);

INVx6_ASAP7_75t_L g9275 ( 
.A(n_8632),
.Y(n_9275)
);

INVx2_ASAP7_75t_L g9276 ( 
.A(n_8606),
.Y(n_9276)
);

INVx3_ASAP7_75t_SL g9277 ( 
.A(n_7646),
.Y(n_9277)
);

OAI21x1_ASAP7_75t_L g9278 ( 
.A1(n_8735),
.A2(n_6601),
.B(n_6566),
.Y(n_9278)
);

AOI22xp33_ASAP7_75t_L g9279 ( 
.A1(n_8363),
.A2(n_7327),
.B1(n_7162),
.B2(n_7204),
.Y(n_9279)
);

INVx1_ASAP7_75t_L g9280 ( 
.A(n_8334),
.Y(n_9280)
);

HB1xp67_ASAP7_75t_L g9281 ( 
.A(n_8313),
.Y(n_9281)
);

AOI22xp33_ASAP7_75t_L g9282 ( 
.A1(n_8931),
.A2(n_7327),
.B1(n_7204),
.B2(n_7302),
.Y(n_9282)
);

AOI22xp33_ASAP7_75t_L g9283 ( 
.A1(n_8931),
.A2(n_7327),
.B1(n_7204),
.B2(n_7302),
.Y(n_9283)
);

INVx2_ASAP7_75t_L g9284 ( 
.A(n_8606),
.Y(n_9284)
);

INVx2_ASAP7_75t_L g9285 ( 
.A(n_8606),
.Y(n_9285)
);

OAI22xp33_ASAP7_75t_L g9286 ( 
.A1(n_7890),
.A2(n_8337),
.B1(n_7697),
.B2(n_7905),
.Y(n_9286)
);

OAI21x1_ASAP7_75t_L g9287 ( 
.A1(n_8765),
.A2(n_6601),
.B(n_6566),
.Y(n_9287)
);

CKINVDCx20_ASAP7_75t_R g9288 ( 
.A(n_8950),
.Y(n_9288)
);

BUFx3_ASAP7_75t_L g9289 ( 
.A(n_8471),
.Y(n_9289)
);

NAND2xp5_ASAP7_75t_L g9290 ( 
.A(n_8187),
.B(n_6752),
.Y(n_9290)
);

INVx1_ASAP7_75t_SL g9291 ( 
.A(n_8830),
.Y(n_9291)
);

AOI22xp33_ASAP7_75t_L g9292 ( 
.A1(n_7799),
.A2(n_7327),
.B1(n_7204),
.B2(n_7302),
.Y(n_9292)
);

HB1xp67_ASAP7_75t_L g9293 ( 
.A(n_8315),
.Y(n_9293)
);

AOI22xp33_ASAP7_75t_L g9294 ( 
.A1(n_7799),
.A2(n_7302),
.B1(n_7168),
.B2(n_7409),
.Y(n_9294)
);

CKINVDCx10_ASAP7_75t_R g9295 ( 
.A(n_7793),
.Y(n_9295)
);

INVx1_ASAP7_75t_L g9296 ( 
.A(n_8334),
.Y(n_9296)
);

INVx1_ASAP7_75t_L g9297 ( 
.A(n_8360),
.Y(n_9297)
);

INVx1_ASAP7_75t_SL g9298 ( 
.A(n_8830),
.Y(n_9298)
);

INVx3_ASAP7_75t_L g9299 ( 
.A(n_7889),
.Y(n_9299)
);

INVx3_ASAP7_75t_L g9300 ( 
.A(n_7889),
.Y(n_9300)
);

AND2x2_ASAP7_75t_L g9301 ( 
.A(n_7617),
.B(n_7388),
.Y(n_9301)
);

AOI22xp33_ASAP7_75t_L g9302 ( 
.A1(n_7665),
.A2(n_7168),
.B1(n_7506),
.B2(n_7409),
.Y(n_9302)
);

OAI21x1_ASAP7_75t_L g9303 ( 
.A1(n_8765),
.A2(n_6602),
.B(n_6566),
.Y(n_9303)
);

NAND2xp5_ASAP7_75t_L g9304 ( 
.A(n_8187),
.B(n_8169),
.Y(n_9304)
);

OAI22xp5_ASAP7_75t_L g9305 ( 
.A1(n_7687),
.A2(n_6695),
.B1(n_6696),
.B2(n_6681),
.Y(n_9305)
);

AO21x1_ASAP7_75t_L g9306 ( 
.A1(n_7837),
.A2(n_7473),
.B(n_7432),
.Y(n_9306)
);

AOI22xp33_ASAP7_75t_L g9307 ( 
.A1(n_7665),
.A2(n_7168),
.B1(n_7506),
.B2(n_7104),
.Y(n_9307)
);

AND2x2_ASAP7_75t_L g9308 ( 
.A(n_7643),
.B(n_7388),
.Y(n_9308)
);

INVx3_ASAP7_75t_L g9309 ( 
.A(n_7889),
.Y(n_9309)
);

OA21x2_ASAP7_75t_L g9310 ( 
.A1(n_8399),
.A2(n_6751),
.B(n_6697),
.Y(n_9310)
);

INVx1_ASAP7_75t_L g9311 ( 
.A(n_8360),
.Y(n_9311)
);

INVx1_ASAP7_75t_L g9312 ( 
.A(n_8385),
.Y(n_9312)
);

INVx1_ASAP7_75t_L g9313 ( 
.A(n_8385),
.Y(n_9313)
);

OA21x2_ASAP7_75t_L g9314 ( 
.A1(n_8701),
.A2(n_6756),
.B(n_6751),
.Y(n_9314)
);

CKINVDCx20_ASAP7_75t_R g9315 ( 
.A(n_8950),
.Y(n_9315)
);

BUFx3_ASAP7_75t_L g9316 ( 
.A(n_8471),
.Y(n_9316)
);

OA21x2_ASAP7_75t_L g9317 ( 
.A1(n_8701),
.A2(n_6756),
.B(n_6751),
.Y(n_9317)
);

INVx3_ASAP7_75t_L g9318 ( 
.A(n_7889),
.Y(n_9318)
);

AO21x2_ASAP7_75t_L g9319 ( 
.A1(n_7779),
.A2(n_7826),
.B(n_8570),
.Y(n_9319)
);

BUFx12f_ASAP7_75t_L g9320 ( 
.A(n_8147),
.Y(n_9320)
);

AOI22xp33_ASAP7_75t_SL g9321 ( 
.A1(n_7621),
.A2(n_8054),
.B1(n_8104),
.B2(n_8088),
.Y(n_9321)
);

INVx2_ASAP7_75t_L g9322 ( 
.A(n_8606),
.Y(n_9322)
);

OAI21x1_ASAP7_75t_L g9323 ( 
.A1(n_8765),
.A2(n_6602),
.B(n_6566),
.Y(n_9323)
);

AOI22xp33_ASAP7_75t_L g9324 ( 
.A1(n_7697),
.A2(n_7168),
.B1(n_7104),
.B2(n_7091),
.Y(n_9324)
);

BUFx3_ASAP7_75t_L g9325 ( 
.A(n_7646),
.Y(n_9325)
);

AOI22xp33_ASAP7_75t_SL g9326 ( 
.A1(n_7621),
.A2(n_7494),
.B1(n_7031),
.B2(n_7495),
.Y(n_9326)
);

HB1xp67_ASAP7_75t_L g9327 ( 
.A(n_8315),
.Y(n_9327)
);

OAI22xp5_ASAP7_75t_L g9328 ( 
.A1(n_7687),
.A2(n_7006),
.B1(n_7164),
.B2(n_6993),
.Y(n_9328)
);

INVx1_ASAP7_75t_L g9329 ( 
.A(n_8387),
.Y(n_9329)
);

INVx1_ASAP7_75t_L g9330 ( 
.A(n_8387),
.Y(n_9330)
);

AOI22xp33_ASAP7_75t_L g9331 ( 
.A1(n_7813),
.A2(n_7168),
.B1(n_7091),
.B2(n_6972),
.Y(n_9331)
);

OAI22xp5_ASAP7_75t_L g9332 ( 
.A1(n_7861),
.A2(n_7006),
.B1(n_7164),
.B2(n_6993),
.Y(n_9332)
);

OA21x2_ASAP7_75t_L g9333 ( 
.A1(n_8701),
.A2(n_6756),
.B(n_7399),
.Y(n_9333)
);

INVx2_ASAP7_75t_L g9334 ( 
.A(n_8606),
.Y(n_9334)
);

INVx1_ASAP7_75t_L g9335 ( 
.A(n_8404),
.Y(n_9335)
);

INVx2_ASAP7_75t_L g9336 ( 
.A(n_8606),
.Y(n_9336)
);

AND2x2_ASAP7_75t_L g9337 ( 
.A(n_7643),
.B(n_7388),
.Y(n_9337)
);

INVx1_ASAP7_75t_L g9338 ( 
.A(n_8404),
.Y(n_9338)
);

INVx1_ASAP7_75t_L g9339 ( 
.A(n_8405),
.Y(n_9339)
);

INVx2_ASAP7_75t_L g9340 ( 
.A(n_8622),
.Y(n_9340)
);

AOI22xp33_ASAP7_75t_SL g9341 ( 
.A1(n_8054),
.A2(n_7509),
.B1(n_7495),
.B2(n_7046),
.Y(n_9341)
);

INVx1_ASAP7_75t_L g9342 ( 
.A(n_8405),
.Y(n_9342)
);

AND2x2_ASAP7_75t_L g9343 ( 
.A(n_7643),
.B(n_7388),
.Y(n_9343)
);

HB1xp67_ASAP7_75t_L g9344 ( 
.A(n_8796),
.Y(n_9344)
);

OAI21xp33_ASAP7_75t_L g9345 ( 
.A1(n_7812),
.A2(n_7488),
.B(n_7458),
.Y(n_9345)
);

OAI21x1_ASAP7_75t_L g9346 ( 
.A1(n_8472),
.A2(n_6624),
.B(n_6602),
.Y(n_9346)
);

AO21x1_ASAP7_75t_L g9347 ( 
.A1(n_7919),
.A2(n_7473),
.B(n_7432),
.Y(n_9347)
);

INVx1_ASAP7_75t_L g9348 ( 
.A(n_8408),
.Y(n_9348)
);

OA21x2_ASAP7_75t_L g9349 ( 
.A1(n_8704),
.A2(n_6756),
.B(n_7399),
.Y(n_9349)
);

INVx1_ASAP7_75t_L g9350 ( 
.A(n_8408),
.Y(n_9350)
);

BUFx2_ASAP7_75t_L g9351 ( 
.A(n_8184),
.Y(n_9351)
);

INVx3_ASAP7_75t_L g9352 ( 
.A(n_7889),
.Y(n_9352)
);

AO21x2_ASAP7_75t_L g9353 ( 
.A1(n_7779),
.A2(n_7826),
.B(n_8570),
.Y(n_9353)
);

HB1xp67_ASAP7_75t_L g9354 ( 
.A(n_8796),
.Y(n_9354)
);

INVx2_ASAP7_75t_L g9355 ( 
.A(n_8622),
.Y(n_9355)
);

INVx2_ASAP7_75t_L g9356 ( 
.A(n_8622),
.Y(n_9356)
);

CKINVDCx20_ASAP7_75t_R g9357 ( 
.A(n_8460),
.Y(n_9357)
);

OAI22xp5_ASAP7_75t_L g9358 ( 
.A1(n_7861),
.A2(n_7006),
.B1(n_7164),
.B2(n_6993),
.Y(n_9358)
);

AOI22xp33_ASAP7_75t_SL g9359 ( 
.A1(n_7813),
.A2(n_7376),
.B1(n_7053),
.B2(n_7399),
.Y(n_9359)
);

INVx1_ASAP7_75t_L g9360 ( 
.A(n_8418),
.Y(n_9360)
);

INVx1_ASAP7_75t_L g9361 ( 
.A(n_8418),
.Y(n_9361)
);

INVx2_ASAP7_75t_L g9362 ( 
.A(n_8622),
.Y(n_9362)
);

INVx2_ASAP7_75t_L g9363 ( 
.A(n_8622),
.Y(n_9363)
);

INVx8_ASAP7_75t_L g9364 ( 
.A(n_8901),
.Y(n_9364)
);

AND2x2_ASAP7_75t_L g9365 ( 
.A(n_7643),
.B(n_7698),
.Y(n_9365)
);

INVx1_ASAP7_75t_L g9366 ( 
.A(n_8419),
.Y(n_9366)
);

INVx2_ASAP7_75t_L g9367 ( 
.A(n_8622),
.Y(n_9367)
);

INVx1_ASAP7_75t_L g9368 ( 
.A(n_8419),
.Y(n_9368)
);

INVx1_ASAP7_75t_L g9369 ( 
.A(n_8424),
.Y(n_9369)
);

CKINVDCx20_ASAP7_75t_R g9370 ( 
.A(n_8460),
.Y(n_9370)
);

AOI22xp33_ASAP7_75t_SL g9371 ( 
.A1(n_8054),
.A2(n_7509),
.B1(n_7046),
.B2(n_7135),
.Y(n_9371)
);

AOI21x1_ASAP7_75t_L g9372 ( 
.A1(n_8300),
.A2(n_7459),
.B(n_7423),
.Y(n_9372)
);

INVx2_ASAP7_75t_L g9373 ( 
.A(n_8496),
.Y(n_9373)
);

AOI22xp33_ASAP7_75t_L g9374 ( 
.A1(n_7984),
.A2(n_6972),
.B1(n_7098),
.B2(n_6655),
.Y(n_9374)
);

INVx2_ASAP7_75t_L g9375 ( 
.A(n_8496),
.Y(n_9375)
);

INVx2_ASAP7_75t_L g9376 ( 
.A(n_8496),
.Y(n_9376)
);

AOI22xp33_ASAP7_75t_SL g9377 ( 
.A1(n_7905),
.A2(n_7376),
.B1(n_7053),
.B2(n_7416),
.Y(n_9377)
);

BUFx3_ASAP7_75t_L g9378 ( 
.A(n_7646),
.Y(n_9378)
);

OR2x6_ASAP7_75t_L g9379 ( 
.A(n_7705),
.B(n_6828),
.Y(n_9379)
);

OAI22xp5_ASAP7_75t_L g9380 ( 
.A1(n_7634),
.A2(n_7006),
.B1(n_7164),
.B2(n_6993),
.Y(n_9380)
);

INVx1_ASAP7_75t_L g9381 ( 
.A(n_8424),
.Y(n_9381)
);

INVx1_ASAP7_75t_L g9382 ( 
.A(n_8427),
.Y(n_9382)
);

AOI22xp33_ASAP7_75t_L g9383 ( 
.A1(n_7984),
.A2(n_6972),
.B1(n_7098),
.B2(n_6655),
.Y(n_9383)
);

AOI21xp5_ASAP7_75t_L g9384 ( 
.A1(n_7707),
.A2(n_7053),
.B(n_7315),
.Y(n_9384)
);

NAND2x1p5_ASAP7_75t_L g9385 ( 
.A(n_8341),
.B(n_8319),
.Y(n_9385)
);

AOI22xp33_ASAP7_75t_SL g9386 ( 
.A1(n_8088),
.A2(n_7416),
.B1(n_7014),
.B2(n_7135),
.Y(n_9386)
);

BUFx6f_ASAP7_75t_L g9387 ( 
.A(n_7943),
.Y(n_9387)
);

OAI21x1_ASAP7_75t_L g9388 ( 
.A1(n_8472),
.A2(n_6624),
.B(n_6602),
.Y(n_9388)
);

HB1xp67_ASAP7_75t_L g9389 ( 
.A(n_8805),
.Y(n_9389)
);

INVx2_ASAP7_75t_SL g9390 ( 
.A(n_7943),
.Y(n_9390)
);

INVx2_ASAP7_75t_L g9391 ( 
.A(n_8498),
.Y(n_9391)
);

INVx2_ASAP7_75t_L g9392 ( 
.A(n_8498),
.Y(n_9392)
);

OA21x2_ASAP7_75t_L g9393 ( 
.A1(n_8704),
.A2(n_8721),
.B(n_8714),
.Y(n_9393)
);

OAI22xp5_ASAP7_75t_L g9394 ( 
.A1(n_7634),
.A2(n_7680),
.B1(n_7652),
.B2(n_7923),
.Y(n_9394)
);

INVx2_ASAP7_75t_L g9395 ( 
.A(n_8498),
.Y(n_9395)
);

INVx1_ASAP7_75t_L g9396 ( 
.A(n_8427),
.Y(n_9396)
);

INVx2_ASAP7_75t_L g9397 ( 
.A(n_8501),
.Y(n_9397)
);

INVx1_ASAP7_75t_L g9398 ( 
.A(n_8444),
.Y(n_9398)
);

OAI21xp5_ASAP7_75t_L g9399 ( 
.A1(n_8151),
.A2(n_6938),
.B(n_7315),
.Y(n_9399)
);

HB1xp67_ASAP7_75t_L g9400 ( 
.A(n_8805),
.Y(n_9400)
);

AOI22xp33_ASAP7_75t_L g9401 ( 
.A1(n_7681),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9401)
);

INVx2_ASAP7_75t_L g9402 ( 
.A(n_8501),
.Y(n_9402)
);

AOI22xp33_ASAP7_75t_L g9403 ( 
.A1(n_7681),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9403)
);

BUFx12f_ASAP7_75t_L g9404 ( 
.A(n_8147),
.Y(n_9404)
);

INVx2_ASAP7_75t_L g9405 ( 
.A(n_8501),
.Y(n_9405)
);

INVx1_ASAP7_75t_L g9406 ( 
.A(n_8444),
.Y(n_9406)
);

AND2x4_ASAP7_75t_L g9407 ( 
.A(n_8202),
.B(n_7330),
.Y(n_9407)
);

OAI22xp33_ASAP7_75t_L g9408 ( 
.A1(n_7890),
.A2(n_7477),
.B1(n_7197),
.B2(n_7223),
.Y(n_9408)
);

INVx1_ASAP7_75t_L g9409 ( 
.A(n_8495),
.Y(n_9409)
);

AO22x1_ASAP7_75t_L g9410 ( 
.A1(n_7606),
.A2(n_6969),
.B1(n_7008),
.B2(n_6951),
.Y(n_9410)
);

INVx1_ASAP7_75t_L g9411 ( 
.A(n_8495),
.Y(n_9411)
);

OR2x6_ASAP7_75t_L g9412 ( 
.A(n_7783),
.B(n_7856),
.Y(n_9412)
);

INVx2_ASAP7_75t_L g9413 ( 
.A(n_8502),
.Y(n_9413)
);

AND2x2_ASAP7_75t_L g9414 ( 
.A(n_7698),
.B(n_7411),
.Y(n_9414)
);

INVx1_ASAP7_75t_L g9415 ( 
.A(n_8515),
.Y(n_9415)
);

INVx4_ASAP7_75t_SL g9416 ( 
.A(n_7788),
.Y(n_9416)
);

INVx1_ASAP7_75t_L g9417 ( 
.A(n_8515),
.Y(n_9417)
);

AO21x1_ASAP7_75t_L g9418 ( 
.A1(n_7919),
.A2(n_6900),
.B(n_6897),
.Y(n_9418)
);

INVx1_ASAP7_75t_L g9419 ( 
.A(n_8521),
.Y(n_9419)
);

INVx1_ASAP7_75t_L g9420 ( 
.A(n_8521),
.Y(n_9420)
);

INVx1_ASAP7_75t_L g9421 ( 
.A(n_8526),
.Y(n_9421)
);

INVx1_ASAP7_75t_L g9422 ( 
.A(n_8526),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_8539),
.Y(n_9423)
);

INVx1_ASAP7_75t_L g9424 ( 
.A(n_8539),
.Y(n_9424)
);

INVx1_ASAP7_75t_L g9425 ( 
.A(n_8559),
.Y(n_9425)
);

INVx2_ASAP7_75t_L g9426 ( 
.A(n_8502),
.Y(n_9426)
);

INVx1_ASAP7_75t_L g9427 ( 
.A(n_8559),
.Y(n_9427)
);

CKINVDCx5p33_ASAP7_75t_R g9428 ( 
.A(n_8938),
.Y(n_9428)
);

INVx2_ASAP7_75t_L g9429 ( 
.A(n_8502),
.Y(n_9429)
);

INVx2_ASAP7_75t_L g9430 ( 
.A(n_8510),
.Y(n_9430)
);

OAI21x1_ASAP7_75t_L g9431 ( 
.A1(n_8472),
.A2(n_6624),
.B(n_6602),
.Y(n_9431)
);

INVx2_ASAP7_75t_L g9432 ( 
.A(n_8506),
.Y(n_9432)
);

NAND2xp5_ASAP7_75t_L g9433 ( 
.A(n_8169),
.B(n_6752),
.Y(n_9433)
);

INVx1_ASAP7_75t_L g9434 ( 
.A(n_8575),
.Y(n_9434)
);

OAI21x1_ASAP7_75t_L g9435 ( 
.A1(n_8704),
.A2(n_6624),
.B(n_6602),
.Y(n_9435)
);

INVxp67_ASAP7_75t_L g9436 ( 
.A(n_8156),
.Y(n_9436)
);

INVx1_ASAP7_75t_L g9437 ( 
.A(n_8575),
.Y(n_9437)
);

INVx3_ASAP7_75t_L g9438 ( 
.A(n_7889),
.Y(n_9438)
);

INVx1_ASAP7_75t_L g9439 ( 
.A(n_8581),
.Y(n_9439)
);

INVx2_ASAP7_75t_L g9440 ( 
.A(n_8506),
.Y(n_9440)
);

INVx2_ASAP7_75t_L g9441 ( 
.A(n_8506),
.Y(n_9441)
);

INVx1_ASAP7_75t_SL g9442 ( 
.A(n_8833),
.Y(n_9442)
);

AOI22xp33_ASAP7_75t_SL g9443 ( 
.A1(n_8104),
.A2(n_7416),
.B1(n_7014),
.B2(n_7135),
.Y(n_9443)
);

INVx1_ASAP7_75t_L g9444 ( 
.A(n_8581),
.Y(n_9444)
);

OAI21x1_ASAP7_75t_L g9445 ( 
.A1(n_8714),
.A2(n_6707),
.B(n_6624),
.Y(n_9445)
);

INVx4_ASAP7_75t_L g9446 ( 
.A(n_8113),
.Y(n_9446)
);

INVx1_ASAP7_75t_L g9447 ( 
.A(n_8587),
.Y(n_9447)
);

INVx1_ASAP7_75t_L g9448 ( 
.A(n_8587),
.Y(n_9448)
);

INVx3_ASAP7_75t_L g9449 ( 
.A(n_7889),
.Y(n_9449)
);

INVx1_ASAP7_75t_L g9450 ( 
.A(n_8588),
.Y(n_9450)
);

INVx2_ASAP7_75t_L g9451 ( 
.A(n_8520),
.Y(n_9451)
);

AND2x2_ASAP7_75t_L g9452 ( 
.A(n_7698),
.B(n_7411),
.Y(n_9452)
);

INVxp67_ASAP7_75t_L g9453 ( 
.A(n_8156),
.Y(n_9453)
);

INVx1_ASAP7_75t_L g9454 ( 
.A(n_8588),
.Y(n_9454)
);

OAI21xp5_ASAP7_75t_SL g9455 ( 
.A1(n_7778),
.A2(n_7468),
.B(n_7070),
.Y(n_9455)
);

INVx1_ASAP7_75t_L g9456 ( 
.A(n_8599),
.Y(n_9456)
);

INVx1_ASAP7_75t_L g9457 ( 
.A(n_8599),
.Y(n_9457)
);

BUFx3_ASAP7_75t_L g9458 ( 
.A(n_8113),
.Y(n_9458)
);

INVx1_ASAP7_75t_L g9459 ( 
.A(n_8602),
.Y(n_9459)
);

HB1xp67_ASAP7_75t_L g9460 ( 
.A(n_8855),
.Y(n_9460)
);

OAI21x1_ASAP7_75t_L g9461 ( 
.A1(n_8714),
.A2(n_6707),
.B(n_6624),
.Y(n_9461)
);

INVx1_ASAP7_75t_L g9462 ( 
.A(n_8602),
.Y(n_9462)
);

AOI22xp33_ASAP7_75t_SL g9463 ( 
.A1(n_8151),
.A2(n_7014),
.B1(n_7135),
.B2(n_7046),
.Y(n_9463)
);

AOI22xp5_ASAP7_75t_SL g9464 ( 
.A1(n_7838),
.A2(n_6656),
.B1(n_7008),
.B2(n_6969),
.Y(n_9464)
);

INVx2_ASAP7_75t_L g9465 ( 
.A(n_8510),
.Y(n_9465)
);

BUFx2_ASAP7_75t_L g9466 ( 
.A(n_8184),
.Y(n_9466)
);

CKINVDCx6p67_ASAP7_75t_R g9467 ( 
.A(n_7788),
.Y(n_9467)
);

INVx1_ASAP7_75t_L g9468 ( 
.A(n_8611),
.Y(n_9468)
);

AND2x2_ASAP7_75t_L g9469 ( 
.A(n_7698),
.B(n_7869),
.Y(n_9469)
);

BUFx2_ASAP7_75t_L g9470 ( 
.A(n_8184),
.Y(n_9470)
);

AOI22xp33_ASAP7_75t_SL g9471 ( 
.A1(n_7993),
.A2(n_7046),
.B1(n_7346),
.B2(n_7330),
.Y(n_9471)
);

INVx3_ASAP7_75t_L g9472 ( 
.A(n_7889),
.Y(n_9472)
);

CKINVDCx5p33_ASAP7_75t_R g9473 ( 
.A(n_8833),
.Y(n_9473)
);

INVx1_ASAP7_75t_L g9474 ( 
.A(n_8611),
.Y(n_9474)
);

BUFx8_ASAP7_75t_L g9475 ( 
.A(n_8888),
.Y(n_9475)
);

INVx2_ASAP7_75t_L g9476 ( 
.A(n_8510),
.Y(n_9476)
);

INVx2_ASAP7_75t_L g9477 ( 
.A(n_8520),
.Y(n_9477)
);

INVx2_ASAP7_75t_L g9478 ( 
.A(n_8520),
.Y(n_9478)
);

INVx2_ASAP7_75t_L g9479 ( 
.A(n_8543),
.Y(n_9479)
);

INVx1_ASAP7_75t_L g9480 ( 
.A(n_8627),
.Y(n_9480)
);

BUFx3_ASAP7_75t_L g9481 ( 
.A(n_8113),
.Y(n_9481)
);

HB1xp67_ASAP7_75t_L g9482 ( 
.A(n_8855),
.Y(n_9482)
);

INVx1_ASAP7_75t_L g9483 ( 
.A(n_8627),
.Y(n_9483)
);

HB1xp67_ASAP7_75t_L g9484 ( 
.A(n_8902),
.Y(n_9484)
);

NOR2x1_ASAP7_75t_R g9485 ( 
.A(n_8263),
.B(n_7351),
.Y(n_9485)
);

AO21x1_ASAP7_75t_L g9486 ( 
.A1(n_8414),
.A2(n_6900),
.B(n_6897),
.Y(n_9486)
);

INVx4_ASAP7_75t_L g9487 ( 
.A(n_8301),
.Y(n_9487)
);

INVx1_ASAP7_75t_L g9488 ( 
.A(n_8638),
.Y(n_9488)
);

CKINVDCx16_ASAP7_75t_R g9489 ( 
.A(n_8335),
.Y(n_9489)
);

INVx4_ASAP7_75t_L g9490 ( 
.A(n_8301),
.Y(n_9490)
);

NAND2x1p5_ASAP7_75t_L g9491 ( 
.A(n_8341),
.B(n_6575),
.Y(n_9491)
);

OAI22xp5_ASAP7_75t_L g9492 ( 
.A1(n_7652),
.A2(n_7523),
.B1(n_7152),
.B2(n_7150),
.Y(n_9492)
);

AOI22xp33_ASAP7_75t_L g9493 ( 
.A1(n_7680),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9493)
);

AOI21x1_ASAP7_75t_L g9494 ( 
.A1(n_7677),
.A2(n_7459),
.B(n_7423),
.Y(n_9494)
);

OAI22xp5_ASAP7_75t_L g9495 ( 
.A1(n_7923),
.A2(n_7838),
.B1(n_8091),
.B2(n_8060),
.Y(n_9495)
);

BUFx2_ASAP7_75t_L g9496 ( 
.A(n_8184),
.Y(n_9496)
);

BUFx10_ASAP7_75t_L g9497 ( 
.A(n_7731),
.Y(n_9497)
);

BUFx2_ASAP7_75t_L g9498 ( 
.A(n_8184),
.Y(n_9498)
);

AND2x2_ASAP7_75t_L g9499 ( 
.A(n_7869),
.B(n_7411),
.Y(n_9499)
);

AOI22xp5_ASAP7_75t_L g9500 ( 
.A1(n_7659),
.A2(n_7354),
.B1(n_7448),
.B2(n_7520),
.Y(n_9500)
);

BUFx6f_ASAP7_75t_L g9501 ( 
.A(n_7943),
.Y(n_9501)
);

INVx2_ASAP7_75t_L g9502 ( 
.A(n_8543),
.Y(n_9502)
);

INVx2_ASAP7_75t_L g9503 ( 
.A(n_8543),
.Y(n_9503)
);

HB1xp67_ASAP7_75t_L g9504 ( 
.A(n_8902),
.Y(n_9504)
);

INVx2_ASAP7_75t_L g9505 ( 
.A(n_8548),
.Y(n_9505)
);

INVx1_ASAP7_75t_L g9506 ( 
.A(n_8638),
.Y(n_9506)
);

BUFx3_ASAP7_75t_L g9507 ( 
.A(n_8301),
.Y(n_9507)
);

INVx2_ASAP7_75t_L g9508 ( 
.A(n_8535),
.Y(n_9508)
);

INVx2_ASAP7_75t_SL g9509 ( 
.A(n_7974),
.Y(n_9509)
);

BUFx4f_ASAP7_75t_L g9510 ( 
.A(n_8316),
.Y(n_9510)
);

AOI22xp33_ASAP7_75t_SL g9511 ( 
.A1(n_7993),
.A2(n_7330),
.B1(n_7496),
.B2(n_7346),
.Y(n_9511)
);

INVx2_ASAP7_75t_L g9512 ( 
.A(n_8535),
.Y(n_9512)
);

BUFx6f_ASAP7_75t_L g9513 ( 
.A(n_7974),
.Y(n_9513)
);

INVx2_ASAP7_75t_L g9514 ( 
.A(n_8535),
.Y(n_9514)
);

INVx2_ASAP7_75t_SL g9515 ( 
.A(n_7974),
.Y(n_9515)
);

HB1xp67_ASAP7_75t_L g9516 ( 
.A(n_8223),
.Y(n_9516)
);

BUFx6f_ASAP7_75t_L g9517 ( 
.A(n_7974),
.Y(n_9517)
);

INVx2_ASAP7_75t_L g9518 ( 
.A(n_8548),
.Y(n_9518)
);

HB1xp67_ASAP7_75t_L g9519 ( 
.A(n_8223),
.Y(n_9519)
);

AND2x4_ASAP7_75t_L g9520 ( 
.A(n_8517),
.B(n_7330),
.Y(n_9520)
);

INVx1_ASAP7_75t_L g9521 ( 
.A(n_8645),
.Y(n_9521)
);

INVx2_ASAP7_75t_L g9522 ( 
.A(n_8548),
.Y(n_9522)
);

HB1xp67_ASAP7_75t_L g9523 ( 
.A(n_8223),
.Y(n_9523)
);

AOI22xp33_ASAP7_75t_L g9524 ( 
.A1(n_8343),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9524)
);

INVx2_ASAP7_75t_L g9525 ( 
.A(n_8553),
.Y(n_9525)
);

INVx2_ASAP7_75t_L g9526 ( 
.A(n_8553),
.Y(n_9526)
);

AND2x4_ASAP7_75t_L g9527 ( 
.A(n_8517),
.B(n_7330),
.Y(n_9527)
);

OAI21x1_ASAP7_75t_L g9528 ( 
.A1(n_8721),
.A2(n_6723),
.B(n_6707),
.Y(n_9528)
);

INVx4_ASAP7_75t_L g9529 ( 
.A(n_8316),
.Y(n_9529)
);

INVx1_ASAP7_75t_L g9530 ( 
.A(n_8645),
.Y(n_9530)
);

INVx2_ASAP7_75t_L g9531 ( 
.A(n_8553),
.Y(n_9531)
);

AOI22xp33_ASAP7_75t_L g9532 ( 
.A1(n_8343),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9532)
);

INVx2_ASAP7_75t_L g9533 ( 
.A(n_8557),
.Y(n_9533)
);

INVx2_ASAP7_75t_L g9534 ( 
.A(n_8557),
.Y(n_9534)
);

INVx1_ASAP7_75t_L g9535 ( 
.A(n_8661),
.Y(n_9535)
);

OAI22xp33_ASAP7_75t_L g9536 ( 
.A1(n_8337),
.A2(n_7197),
.B1(n_7223),
.B2(n_7169),
.Y(n_9536)
);

AOI22x1_ASAP7_75t_L g9537 ( 
.A1(n_8335),
.A2(n_7366),
.B1(n_7433),
.B2(n_7312),
.Y(n_9537)
);

AOI22xp33_ASAP7_75t_L g9538 ( 
.A1(n_7835),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9538)
);

INVx1_ASAP7_75t_L g9539 ( 
.A(n_8661),
.Y(n_9539)
);

INVx1_ASAP7_75t_L g9540 ( 
.A(n_8667),
.Y(n_9540)
);

OAI22xp33_ASAP7_75t_L g9541 ( 
.A1(n_8330),
.A2(n_7197),
.B1(n_7223),
.B2(n_7169),
.Y(n_9541)
);

AND2x4_ASAP7_75t_L g9542 ( 
.A(n_8517),
.B(n_7330),
.Y(n_9542)
);

BUFx3_ASAP7_75t_L g9543 ( 
.A(n_8316),
.Y(n_9543)
);

OR2x6_ASAP7_75t_L g9544 ( 
.A(n_7856),
.B(n_6828),
.Y(n_9544)
);

INVxp33_ASAP7_75t_L g9545 ( 
.A(n_8683),
.Y(n_9545)
);

INVx1_ASAP7_75t_L g9546 ( 
.A(n_8667),
.Y(n_9546)
);

INVx1_ASAP7_75t_L g9547 ( 
.A(n_8668),
.Y(n_9547)
);

BUFx3_ASAP7_75t_L g9548 ( 
.A(n_7986),
.Y(n_9548)
);

NAND2x1p5_ASAP7_75t_L g9549 ( 
.A(n_8341),
.B(n_8319),
.Y(n_9549)
);

INVx1_ASAP7_75t_L g9550 ( 
.A(n_8668),
.Y(n_9550)
);

AOI22xp33_ASAP7_75t_L g9551 ( 
.A1(n_7835),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9551)
);

AO21x1_ASAP7_75t_L g9552 ( 
.A1(n_8414),
.A2(n_7049),
.B(n_6908),
.Y(n_9552)
);

INVx2_ASAP7_75t_L g9553 ( 
.A(n_8557),
.Y(n_9553)
);

INVx4_ASAP7_75t_L g9554 ( 
.A(n_7630),
.Y(n_9554)
);

INVx1_ASAP7_75t_L g9555 ( 
.A(n_8682),
.Y(n_9555)
);

INVx8_ASAP7_75t_L g9556 ( 
.A(n_8901),
.Y(n_9556)
);

OAI21x1_ASAP7_75t_SL g9557 ( 
.A1(n_8053),
.A2(n_7426),
.B(n_7420),
.Y(n_9557)
);

INVx2_ASAP7_75t_SL g9558 ( 
.A(n_7986),
.Y(n_9558)
);

INVx2_ASAP7_75t_L g9559 ( 
.A(n_8558),
.Y(n_9559)
);

AOI22xp33_ASAP7_75t_L g9560 ( 
.A1(n_8229),
.A2(n_7763),
.B1(n_7650),
.B2(n_8629),
.Y(n_9560)
);

AND2x2_ASAP7_75t_L g9561 ( 
.A(n_7869),
.B(n_7411),
.Y(n_9561)
);

INVx2_ASAP7_75t_SL g9562 ( 
.A(n_7986),
.Y(n_9562)
);

OAI22xp5_ASAP7_75t_L g9563 ( 
.A1(n_8060),
.A2(n_7152),
.B1(n_7150),
.B2(n_7520),
.Y(n_9563)
);

AO21x1_ASAP7_75t_SL g9564 ( 
.A1(n_8463),
.A2(n_7303),
.B(n_7169),
.Y(n_9564)
);

BUFx6f_ASAP7_75t_L g9565 ( 
.A(n_7986),
.Y(n_9565)
);

NAND2xp5_ASAP7_75t_L g9566 ( 
.A(n_8180),
.B(n_6758),
.Y(n_9566)
);

BUFx2_ASAP7_75t_R g9567 ( 
.A(n_8497),
.Y(n_9567)
);

INVx1_ASAP7_75t_L g9568 ( 
.A(n_8682),
.Y(n_9568)
);

NAND2xp5_ASAP7_75t_L g9569 ( 
.A(n_8180),
.B(n_6758),
.Y(n_9569)
);

BUFx6f_ASAP7_75t_L g9570 ( 
.A(n_8141),
.Y(n_9570)
);

INVx11_ASAP7_75t_L g9571 ( 
.A(n_8888),
.Y(n_9571)
);

BUFx2_ASAP7_75t_L g9572 ( 
.A(n_8009),
.Y(n_9572)
);

INVx1_ASAP7_75t_L g9573 ( 
.A(n_8715),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_8715),
.Y(n_9574)
);

INVx2_ASAP7_75t_L g9575 ( 
.A(n_8558),
.Y(n_9575)
);

AOI22xp33_ASAP7_75t_L g9576 ( 
.A1(n_8229),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9576)
);

OAI21x1_ASAP7_75t_L g9577 ( 
.A1(n_8721),
.A2(n_6723),
.B(n_6707),
.Y(n_9577)
);

OAI22xp33_ASAP7_75t_L g9578 ( 
.A1(n_8330),
.A2(n_7520),
.B1(n_7448),
.B2(n_7488),
.Y(n_9578)
);

INVx1_ASAP7_75t_L g9579 ( 
.A(n_8720),
.Y(n_9579)
);

INVx1_ASAP7_75t_L g9580 ( 
.A(n_8720),
.Y(n_9580)
);

INVx1_ASAP7_75t_L g9581 ( 
.A(n_8726),
.Y(n_9581)
);

INVx1_ASAP7_75t_L g9582 ( 
.A(n_8726),
.Y(n_9582)
);

NAND2xp5_ASAP7_75t_L g9583 ( 
.A(n_8055),
.B(n_6768),
.Y(n_9583)
);

INVx2_ASAP7_75t_L g9584 ( 
.A(n_8558),
.Y(n_9584)
);

INVx1_ASAP7_75t_L g9585 ( 
.A(n_8728),
.Y(n_9585)
);

BUFx6f_ASAP7_75t_L g9586 ( 
.A(n_8141),
.Y(n_9586)
);

INVx2_ASAP7_75t_L g9587 ( 
.A(n_8564),
.Y(n_9587)
);

AOI22xp33_ASAP7_75t_L g9588 ( 
.A1(n_7763),
.A2(n_6972),
.B1(n_7124),
.B2(n_7098),
.Y(n_9588)
);

INVx2_ASAP7_75t_L g9589 ( 
.A(n_8564),
.Y(n_9589)
);

OAI21x1_ASAP7_75t_L g9590 ( 
.A1(n_8733),
.A2(n_6723),
.B(n_6707),
.Y(n_9590)
);

INVx2_ASAP7_75t_L g9591 ( 
.A(n_8564),
.Y(n_9591)
);

BUFx2_ASAP7_75t_L g9592 ( 
.A(n_8009),
.Y(n_9592)
);

AOI21x1_ASAP7_75t_L g9593 ( 
.A1(n_7677),
.A2(n_7459),
.B(n_7423),
.Y(n_9593)
);

INVx1_ASAP7_75t_L g9594 ( 
.A(n_8728),
.Y(n_9594)
);

CKINVDCx20_ASAP7_75t_R g9595 ( 
.A(n_8488),
.Y(n_9595)
);

INVx4_ASAP7_75t_L g9596 ( 
.A(n_7630),
.Y(n_9596)
);

OR2x6_ASAP7_75t_L g9597 ( 
.A(n_7865),
.B(n_7077),
.Y(n_9597)
);

INVx1_ASAP7_75t_L g9598 ( 
.A(n_8734),
.Y(n_9598)
);

BUFx12f_ASAP7_75t_L g9599 ( 
.A(n_8263),
.Y(n_9599)
);

INVx2_ASAP7_75t_L g9600 ( 
.A(n_8569),
.Y(n_9600)
);

INVx1_ASAP7_75t_L g9601 ( 
.A(n_8734),
.Y(n_9601)
);

AOI22xp5_ASAP7_75t_L g9602 ( 
.A1(n_7659),
.A2(n_7354),
.B1(n_7448),
.B2(n_7458),
.Y(n_9602)
);

AOI22xp33_ASAP7_75t_L g9603 ( 
.A1(n_7650),
.A2(n_7098),
.B1(n_7124),
.B2(n_7543),
.Y(n_9603)
);

BUFx6f_ASAP7_75t_L g9604 ( 
.A(n_8141),
.Y(n_9604)
);

INVxp67_ASAP7_75t_L g9605 ( 
.A(n_7999),
.Y(n_9605)
);

BUFx3_ASAP7_75t_L g9606 ( 
.A(n_8141),
.Y(n_9606)
);

INVx1_ASAP7_75t_L g9607 ( 
.A(n_8746),
.Y(n_9607)
);

AND2x4_ASAP7_75t_L g9608 ( 
.A(n_8517),
.B(n_7330),
.Y(n_9608)
);

BUFx12f_ASAP7_75t_L g9609 ( 
.A(n_8487),
.Y(n_9609)
);

INVx1_ASAP7_75t_L g9610 ( 
.A(n_8746),
.Y(n_9610)
);

OAI22xp33_ASAP7_75t_L g9611 ( 
.A1(n_7964),
.A2(n_7488),
.B1(n_7354),
.B2(n_7374),
.Y(n_9611)
);

INVx1_ASAP7_75t_L g9612 ( 
.A(n_8764),
.Y(n_9612)
);

INVx1_ASAP7_75t_L g9613 ( 
.A(n_8764),
.Y(n_9613)
);

BUFx2_ASAP7_75t_L g9614 ( 
.A(n_7869),
.Y(n_9614)
);

OAI21x1_ASAP7_75t_L g9615 ( 
.A1(n_8733),
.A2(n_6723),
.B(n_6707),
.Y(n_9615)
);

AND2x2_ASAP7_75t_L g9616 ( 
.A(n_8309),
.B(n_7414),
.Y(n_9616)
);

AND2x2_ASAP7_75t_L g9617 ( 
.A(n_8309),
.B(n_7414),
.Y(n_9617)
);

CKINVDCx6p67_ASAP7_75t_R g9618 ( 
.A(n_7788),
.Y(n_9618)
);

AND2x4_ASAP7_75t_L g9619 ( 
.A(n_8517),
.B(n_7346),
.Y(n_9619)
);

INVx2_ASAP7_75t_L g9620 ( 
.A(n_8569),
.Y(n_9620)
);

OAI21x1_ASAP7_75t_SL g9621 ( 
.A1(n_8053),
.A2(n_7426),
.B(n_7420),
.Y(n_9621)
);

INVx2_ASAP7_75t_L g9622 ( 
.A(n_8569),
.Y(n_9622)
);

CKINVDCx20_ASAP7_75t_R g9623 ( 
.A(n_8488),
.Y(n_9623)
);

BUFx10_ASAP7_75t_L g9624 ( 
.A(n_8132),
.Y(n_9624)
);

AOI22xp33_ASAP7_75t_L g9625 ( 
.A1(n_8629),
.A2(n_7124),
.B1(n_7544),
.B2(n_7543),
.Y(n_9625)
);

INVx1_ASAP7_75t_L g9626 ( 
.A(n_8767),
.Y(n_9626)
);

CKINVDCx11_ASAP7_75t_R g9627 ( 
.A(n_8497),
.Y(n_9627)
);

INVx2_ASAP7_75t_L g9628 ( 
.A(n_8574),
.Y(n_9628)
);

AOI22xp33_ASAP7_75t_L g9629 ( 
.A1(n_7907),
.A2(n_7124),
.B1(n_7544),
.B2(n_7391),
.Y(n_9629)
);

INVx1_ASAP7_75t_L g9630 ( 
.A(n_8767),
.Y(n_9630)
);

INVx1_ASAP7_75t_L g9631 ( 
.A(n_8771),
.Y(n_9631)
);

BUFx6f_ASAP7_75t_L g9632 ( 
.A(n_8153),
.Y(n_9632)
);

INVx1_ASAP7_75t_L g9633 ( 
.A(n_8771),
.Y(n_9633)
);

OAI21x1_ASAP7_75t_SL g9634 ( 
.A1(n_8600),
.A2(n_7426),
.B(n_7420),
.Y(n_9634)
);

OA21x2_ASAP7_75t_L g9635 ( 
.A1(n_8733),
.A2(n_6918),
.B(n_6917),
.Y(n_9635)
);

AOI22xp33_ASAP7_75t_L g9636 ( 
.A1(n_7907),
.A2(n_7391),
.B1(n_7479),
.B2(n_6930),
.Y(n_9636)
);

AOI22xp33_ASAP7_75t_L g9637 ( 
.A1(n_8591),
.A2(n_7391),
.B1(n_7479),
.B2(n_6930),
.Y(n_9637)
);

OAI22xp5_ASAP7_75t_L g9638 ( 
.A1(n_8091),
.A2(n_7345),
.B1(n_7234),
.B2(n_7303),
.Y(n_9638)
);

AOI22xp33_ASAP7_75t_SL g9639 ( 
.A1(n_7993),
.A2(n_7346),
.B1(n_7551),
.B2(n_7496),
.Y(n_9639)
);

INVx1_ASAP7_75t_L g9640 ( 
.A(n_8774),
.Y(n_9640)
);

INVx2_ASAP7_75t_L g9641 ( 
.A(n_8574),
.Y(n_9641)
);

AOI22xp33_ASAP7_75t_L g9642 ( 
.A1(n_8591),
.A2(n_7391),
.B1(n_7479),
.B2(n_6930),
.Y(n_9642)
);

AOI21x1_ASAP7_75t_L g9643 ( 
.A1(n_7677),
.A2(n_7466),
.B(n_7462),
.Y(n_9643)
);

INVx1_ASAP7_75t_L g9644 ( 
.A(n_8774),
.Y(n_9644)
);

INVx1_ASAP7_75t_L g9645 ( 
.A(n_8778),
.Y(n_9645)
);

BUFx3_ASAP7_75t_L g9646 ( 
.A(n_8153),
.Y(n_9646)
);

INVx2_ASAP7_75t_L g9647 ( 
.A(n_8574),
.Y(n_9647)
);

NAND2xp5_ASAP7_75t_L g9648 ( 
.A(n_8055),
.B(n_6768),
.Y(n_9648)
);

CKINVDCx14_ASAP7_75t_R g9649 ( 
.A(n_8487),
.Y(n_9649)
);

INVx1_ASAP7_75t_L g9650 ( 
.A(n_8778),
.Y(n_9650)
);

CKINVDCx11_ASAP7_75t_R g9651 ( 
.A(n_8685),
.Y(n_9651)
);

AOI21x1_ASAP7_75t_L g9652 ( 
.A1(n_7696),
.A2(n_7728),
.B(n_7702),
.Y(n_9652)
);

OA21x2_ASAP7_75t_L g9653 ( 
.A1(n_8064),
.A2(n_6918),
.B(n_6917),
.Y(n_9653)
);

AOI22xp33_ASAP7_75t_L g9654 ( 
.A1(n_8246),
.A2(n_7391),
.B1(n_7479),
.B2(n_6930),
.Y(n_9654)
);

INVx2_ASAP7_75t_L g9655 ( 
.A(n_8693),
.Y(n_9655)
);

CKINVDCx5p33_ASAP7_75t_R g9656 ( 
.A(n_8279),
.Y(n_9656)
);

NAND2xp5_ASAP7_75t_L g9657 ( 
.A(n_8741),
.B(n_6908),
.Y(n_9657)
);

INVx1_ASAP7_75t_L g9658 ( 
.A(n_8780),
.Y(n_9658)
);

HB1xp67_ASAP7_75t_L g9659 ( 
.A(n_8268),
.Y(n_9659)
);

INVx1_ASAP7_75t_L g9660 ( 
.A(n_8780),
.Y(n_9660)
);

HB1xp67_ASAP7_75t_SL g9661 ( 
.A(n_7977),
.Y(n_9661)
);

AOI22xp33_ASAP7_75t_L g9662 ( 
.A1(n_8246),
.A2(n_7391),
.B1(n_7479),
.B2(n_6930),
.Y(n_9662)
);

BUFx2_ASAP7_75t_L g9663 ( 
.A(n_8872),
.Y(n_9663)
);

INVx11_ASAP7_75t_L g9664 ( 
.A(n_8888),
.Y(n_9664)
);

INVx3_ASAP7_75t_L g9665 ( 
.A(n_7894),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_8786),
.Y(n_9666)
);

OR2x2_ASAP7_75t_L g9667 ( 
.A(n_7795),
.B(n_7215),
.Y(n_9667)
);

AOI22xp33_ASAP7_75t_L g9668 ( 
.A1(n_8014),
.A2(n_7938),
.B1(n_8181),
.B2(n_7641),
.Y(n_9668)
);

INVx1_ASAP7_75t_L g9669 ( 
.A(n_8786),
.Y(n_9669)
);

INVx1_ASAP7_75t_L g9670 ( 
.A(n_8787),
.Y(n_9670)
);

INVx4_ASAP7_75t_L g9671 ( 
.A(n_7630),
.Y(n_9671)
);

INVx1_ASAP7_75t_L g9672 ( 
.A(n_8787),
.Y(n_9672)
);

OA21x2_ASAP7_75t_L g9673 ( 
.A1(n_8064),
.A2(n_6918),
.B(n_6917),
.Y(n_9673)
);

INVx3_ASAP7_75t_L g9674 ( 
.A(n_7894),
.Y(n_9674)
);

INVx1_ASAP7_75t_L g9675 ( 
.A(n_8808),
.Y(n_9675)
);

CKINVDCx11_ASAP7_75t_R g9676 ( 
.A(n_8685),
.Y(n_9676)
);

INVx2_ASAP7_75t_L g9677 ( 
.A(n_8693),
.Y(n_9677)
);

OR2x6_ASAP7_75t_L g9678 ( 
.A(n_7865),
.B(n_7077),
.Y(n_9678)
);

INVx8_ASAP7_75t_L g9679 ( 
.A(n_8901),
.Y(n_9679)
);

AOI22xp33_ASAP7_75t_SL g9680 ( 
.A1(n_8105),
.A2(n_7346),
.B1(n_7551),
.B2(n_7496),
.Y(n_9680)
);

BUFx4f_ASAP7_75t_SL g9681 ( 
.A(n_8888),
.Y(n_9681)
);

HB1xp67_ASAP7_75t_L g9682 ( 
.A(n_8268),
.Y(n_9682)
);

AOI22xp33_ASAP7_75t_SL g9683 ( 
.A1(n_8105),
.A2(n_7346),
.B1(n_7551),
.B2(n_7496),
.Y(n_9683)
);

INVx1_ASAP7_75t_L g9684 ( 
.A(n_8808),
.Y(n_9684)
);

INVx3_ASAP7_75t_L g9685 ( 
.A(n_7894),
.Y(n_9685)
);

INVx1_ASAP7_75t_L g9686 ( 
.A(n_8821),
.Y(n_9686)
);

HB1xp67_ASAP7_75t_L g9687 ( 
.A(n_8268),
.Y(n_9687)
);

INVx1_ASAP7_75t_L g9688 ( 
.A(n_8821),
.Y(n_9688)
);

AOI22xp33_ASAP7_75t_SL g9689 ( 
.A1(n_8105),
.A2(n_7346),
.B1(n_7551),
.B2(n_7496),
.Y(n_9689)
);

INVx1_ASAP7_75t_SL g9690 ( 
.A(n_7985),
.Y(n_9690)
);

NAND2xp5_ASAP7_75t_L g9691 ( 
.A(n_8741),
.B(n_7049),
.Y(n_9691)
);

NAND2xp5_ASAP7_75t_L g9692 ( 
.A(n_8753),
.B(n_7076),
.Y(n_9692)
);

INVx2_ASAP7_75t_SL g9693 ( 
.A(n_8153),
.Y(n_9693)
);

OA21x2_ASAP7_75t_L g9694 ( 
.A1(n_8064),
.A2(n_7016),
.B(n_6990),
.Y(n_9694)
);

INVx5_ASAP7_75t_L g9695 ( 
.A(n_7894),
.Y(n_9695)
);

INVx1_ASAP7_75t_L g9696 ( 
.A(n_8828),
.Y(n_9696)
);

AOI22xp33_ASAP7_75t_L g9697 ( 
.A1(n_8014),
.A2(n_7479),
.B1(n_7552),
.B2(n_6930),
.Y(n_9697)
);

AND2x2_ASAP7_75t_L g9698 ( 
.A(n_8309),
.B(n_7414),
.Y(n_9698)
);

INVx1_ASAP7_75t_L g9699 ( 
.A(n_8828),
.Y(n_9699)
);

HB1xp67_ASAP7_75t_L g9700 ( 
.A(n_8321),
.Y(n_9700)
);

OA21x2_ASAP7_75t_L g9701 ( 
.A1(n_8700),
.A2(n_7775),
.B(n_8063),
.Y(n_9701)
);

NAND2xp5_ASAP7_75t_L g9702 ( 
.A(n_8753),
.B(n_8797),
.Y(n_9702)
);

INVx6_ASAP7_75t_L g9703 ( 
.A(n_7867),
.Y(n_9703)
);

INVx2_ASAP7_75t_L g9704 ( 
.A(n_8693),
.Y(n_9704)
);

AND2x2_ASAP7_75t_L g9705 ( 
.A(n_8325),
.B(n_7414),
.Y(n_9705)
);

NAND2x1p5_ASAP7_75t_L g9706 ( 
.A(n_8319),
.B(n_6575),
.Y(n_9706)
);

INVx2_ASAP7_75t_L g9707 ( 
.A(n_8317),
.Y(n_9707)
);

AND2x2_ASAP7_75t_L g9708 ( 
.A(n_8325),
.B(n_7138),
.Y(n_9708)
);

INVx1_ASAP7_75t_L g9709 ( 
.A(n_8835),
.Y(n_9709)
);

INVx1_ASAP7_75t_L g9710 ( 
.A(n_8835),
.Y(n_9710)
);

OAI22xp33_ASAP7_75t_L g9711 ( 
.A1(n_7964),
.A2(n_7374),
.B1(n_7361),
.B2(n_7578),
.Y(n_9711)
);

BUFx3_ASAP7_75t_L g9712 ( 
.A(n_8153),
.Y(n_9712)
);

INVx1_ASAP7_75t_L g9713 ( 
.A(n_8843),
.Y(n_9713)
);

AND2x4_ASAP7_75t_L g9714 ( 
.A(n_8517),
.B(n_7346),
.Y(n_9714)
);

INVx1_ASAP7_75t_L g9715 ( 
.A(n_8843),
.Y(n_9715)
);

HB1xp67_ASAP7_75t_L g9716 ( 
.A(n_8321),
.Y(n_9716)
);

AOI22xp33_ASAP7_75t_L g9717 ( 
.A1(n_7938),
.A2(n_7552),
.B1(n_7187),
.B2(n_6576),
.Y(n_9717)
);

AOI21x1_ASAP7_75t_L g9718 ( 
.A1(n_7696),
.A2(n_7466),
.B(n_7462),
.Y(n_9718)
);

AOI22xp33_ASAP7_75t_L g9719 ( 
.A1(n_8181),
.A2(n_7552),
.B1(n_7187),
.B2(n_6576),
.Y(n_9719)
);

INVx1_ASAP7_75t_L g9720 ( 
.A(n_8844),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_8844),
.Y(n_9721)
);

INVx2_ASAP7_75t_L g9722 ( 
.A(n_8317),
.Y(n_9722)
);

INVx1_ASAP7_75t_L g9723 ( 
.A(n_8854),
.Y(n_9723)
);

OAI21x1_ASAP7_75t_L g9724 ( 
.A1(n_8655),
.A2(n_6735),
.B(n_6723),
.Y(n_9724)
);

AO21x1_ASAP7_75t_L g9725 ( 
.A1(n_8370),
.A2(n_7076),
.B(n_7335),
.Y(n_9725)
);

AOI22xp33_ASAP7_75t_SL g9726 ( 
.A1(n_8120),
.A2(n_7346),
.B1(n_7551),
.B2(n_7496),
.Y(n_9726)
);

HB1xp67_ASAP7_75t_L g9727 ( 
.A(n_8321),
.Y(n_9727)
);

AOI22xp33_ASAP7_75t_L g9728 ( 
.A1(n_7641),
.A2(n_7552),
.B1(n_6576),
.B2(n_6570),
.Y(n_9728)
);

AOI21x1_ASAP7_75t_L g9729 ( 
.A1(n_7696),
.A2(n_7466),
.B(n_7462),
.Y(n_9729)
);

BUFx2_ASAP7_75t_SL g9730 ( 
.A(n_7640),
.Y(n_9730)
);

INVx1_ASAP7_75t_L g9731 ( 
.A(n_8854),
.Y(n_9731)
);

OAI21x1_ASAP7_75t_L g9732 ( 
.A1(n_8655),
.A2(n_6735),
.B(n_6723),
.Y(n_9732)
);

AOI22xp33_ASAP7_75t_L g9733 ( 
.A1(n_7778),
.A2(n_7952),
.B1(n_8551),
.B2(n_8346),
.Y(n_9733)
);

INVx3_ASAP7_75t_L g9734 ( 
.A(n_7894),
.Y(n_9734)
);

BUFx6f_ASAP7_75t_L g9735 ( 
.A(n_8165),
.Y(n_9735)
);

AO21x1_ASAP7_75t_L g9736 ( 
.A1(n_8370),
.A2(n_7396),
.B(n_7335),
.Y(n_9736)
);

BUFx8_ASAP7_75t_L g9737 ( 
.A(n_8892),
.Y(n_9737)
);

AOI21x1_ASAP7_75t_L g9738 ( 
.A1(n_7702),
.A2(n_7481),
.B(n_7478),
.Y(n_9738)
);

AND2x2_ASAP7_75t_L g9739 ( 
.A(n_8325),
.B(n_7138),
.Y(n_9739)
);

OAI22xp5_ASAP7_75t_L g9740 ( 
.A1(n_8166),
.A2(n_7345),
.B1(n_7234),
.B2(n_7361),
.Y(n_9740)
);

CKINVDCx11_ASAP7_75t_R g9741 ( 
.A(n_8685),
.Y(n_9741)
);

INVx8_ASAP7_75t_L g9742 ( 
.A(n_8901),
.Y(n_9742)
);

AOI22xp33_ASAP7_75t_SL g9743 ( 
.A1(n_8120),
.A2(n_7346),
.B1(n_7551),
.B2(n_7496),
.Y(n_9743)
);

BUFx3_ASAP7_75t_L g9744 ( 
.A(n_8165),
.Y(n_9744)
);

INVx1_ASAP7_75t_L g9745 ( 
.A(n_8860),
.Y(n_9745)
);

INVx1_ASAP7_75t_L g9746 ( 
.A(n_8860),
.Y(n_9746)
);

BUFx3_ASAP7_75t_L g9747 ( 
.A(n_8165),
.Y(n_9747)
);

OAI21x1_ASAP7_75t_L g9748 ( 
.A1(n_8655),
.A2(n_6769),
.B(n_6735),
.Y(n_9748)
);

INVx1_ASAP7_75t_L g9749 ( 
.A(n_8906),
.Y(n_9749)
);

AND2x4_ASAP7_75t_L g9750 ( 
.A(n_8517),
.B(n_7496),
.Y(n_9750)
);

INVx1_ASAP7_75t_L g9751 ( 
.A(n_8906),
.Y(n_9751)
);

AND2x4_ASAP7_75t_L g9752 ( 
.A(n_8457),
.B(n_7496),
.Y(n_9752)
);

INVx1_ASAP7_75t_L g9753 ( 
.A(n_8927),
.Y(n_9753)
);

INVx1_ASAP7_75t_L g9754 ( 
.A(n_8927),
.Y(n_9754)
);

INVx3_ASAP7_75t_L g9755 ( 
.A(n_7894),
.Y(n_9755)
);

BUFx6f_ASAP7_75t_L g9756 ( 
.A(n_8165),
.Y(n_9756)
);

INVx1_ASAP7_75t_L g9757 ( 
.A(n_8930),
.Y(n_9757)
);

OAI21x1_ASAP7_75t_SL g9758 ( 
.A1(n_8600),
.A2(n_7426),
.B(n_7420),
.Y(n_9758)
);

OAI21x1_ASAP7_75t_L g9759 ( 
.A1(n_8858),
.A2(n_8700),
.B(n_7611),
.Y(n_9759)
);

AOI22xp33_ASAP7_75t_L g9760 ( 
.A1(n_7952),
.A2(n_8551),
.B1(n_8346),
.B2(n_8003),
.Y(n_9760)
);

INVx3_ASAP7_75t_L g9761 ( 
.A(n_7894),
.Y(n_9761)
);

INVx1_ASAP7_75t_L g9762 ( 
.A(n_8930),
.Y(n_9762)
);

INVx1_ASAP7_75t_L g9763 ( 
.A(n_8935),
.Y(n_9763)
);

CKINVDCx16_ASAP7_75t_R g9764 ( 
.A(n_8554),
.Y(n_9764)
);

INVx2_ASAP7_75t_L g9765 ( 
.A(n_8317),
.Y(n_9765)
);

INVx2_ASAP7_75t_L g9766 ( 
.A(n_8317),
.Y(n_9766)
);

INVx3_ASAP7_75t_L g9767 ( 
.A(n_7894),
.Y(n_9767)
);

OAI21x1_ASAP7_75t_L g9768 ( 
.A1(n_8858),
.A2(n_8700),
.B(n_7611),
.Y(n_9768)
);

AOI22xp33_ASAP7_75t_L g9769 ( 
.A1(n_8003),
.A2(n_8122),
.B1(n_8219),
.B2(n_8756),
.Y(n_9769)
);

INVx2_ASAP7_75t_L g9770 ( 
.A(n_8317),
.Y(n_9770)
);

INVx2_ASAP7_75t_L g9771 ( 
.A(n_8317),
.Y(n_9771)
);

BUFx2_ASAP7_75t_L g9772 ( 
.A(n_8872),
.Y(n_9772)
);

INVx1_ASAP7_75t_L g9773 ( 
.A(n_8935),
.Y(n_9773)
);

AND2x2_ASAP7_75t_L g9774 ( 
.A(n_8390),
.B(n_7138),
.Y(n_9774)
);

HB1xp67_ASAP7_75t_L g9775 ( 
.A(n_8369),
.Y(n_9775)
);

INVx1_ASAP7_75t_L g9776 ( 
.A(n_8936),
.Y(n_9776)
);

OAI21x1_ASAP7_75t_L g9777 ( 
.A1(n_8858),
.A2(n_6769),
.B(n_6735),
.Y(n_9777)
);

HB1xp67_ASAP7_75t_L g9778 ( 
.A(n_8369),
.Y(n_9778)
);

INVx2_ASAP7_75t_L g9779 ( 
.A(n_8349),
.Y(n_9779)
);

INVx1_ASAP7_75t_SL g9780 ( 
.A(n_7985),
.Y(n_9780)
);

INVx1_ASAP7_75t_L g9781 ( 
.A(n_8936),
.Y(n_9781)
);

INVx3_ASAP7_75t_L g9782 ( 
.A(n_8020),
.Y(n_9782)
);

AND2x4_ASAP7_75t_L g9783 ( 
.A(n_8457),
.B(n_7496),
.Y(n_9783)
);

INVx2_ASAP7_75t_L g9784 ( 
.A(n_8349),
.Y(n_9784)
);

INVx2_ASAP7_75t_L g9785 ( 
.A(n_8349),
.Y(n_9785)
);

INVx4_ASAP7_75t_L g9786 ( 
.A(n_8042),
.Y(n_9786)
);

OAI21x1_ASAP7_75t_L g9787 ( 
.A1(n_7611),
.A2(n_6769),
.B(n_6735),
.Y(n_9787)
);

INVx2_ASAP7_75t_L g9788 ( 
.A(n_8349),
.Y(n_9788)
);

NAND2xp5_ASAP7_75t_L g9789 ( 
.A(n_8797),
.B(n_6770),
.Y(n_9789)
);

AND2x2_ASAP7_75t_L g9790 ( 
.A(n_8390),
.B(n_7138),
.Y(n_9790)
);

INVxp67_ASAP7_75t_L g9791 ( 
.A(n_7999),
.Y(n_9791)
);

OAI21x1_ASAP7_75t_L g9792 ( 
.A1(n_7692),
.A2(n_6769),
.B(n_6735),
.Y(n_9792)
);

AOI22xp5_ASAP7_75t_L g9793 ( 
.A1(n_7623),
.A2(n_7468),
.B1(n_6656),
.B2(n_7499),
.Y(n_9793)
);

BUFx3_ASAP7_75t_L g9794 ( 
.A(n_8195),
.Y(n_9794)
);

INVx2_ASAP7_75t_L g9795 ( 
.A(n_8349),
.Y(n_9795)
);

AND2x2_ASAP7_75t_L g9796 ( 
.A(n_8390),
.B(n_8410),
.Y(n_9796)
);

NAND2xp5_ASAP7_75t_L g9797 ( 
.A(n_8832),
.B(n_8840),
.Y(n_9797)
);

INVx2_ASAP7_75t_L g9798 ( 
.A(n_8349),
.Y(n_9798)
);

NAND2xp5_ASAP7_75t_L g9799 ( 
.A(n_8832),
.B(n_6770),
.Y(n_9799)
);

AOI22xp33_ASAP7_75t_L g9800 ( 
.A1(n_8122),
.A2(n_7552),
.B1(n_6576),
.B2(n_6570),
.Y(n_9800)
);

INVx1_ASAP7_75t_L g9801 ( 
.A(n_8945),
.Y(n_9801)
);

AOI21x1_ASAP7_75t_L g9802 ( 
.A1(n_7702),
.A2(n_7481),
.B(n_7478),
.Y(n_9802)
);

CKINVDCx5p33_ASAP7_75t_R g9803 ( 
.A(n_8279),
.Y(n_9803)
);

AOI22xp33_ASAP7_75t_SL g9804 ( 
.A1(n_7779),
.A2(n_7570),
.B1(n_7551),
.B2(n_7552),
.Y(n_9804)
);

NAND2xp5_ASAP7_75t_L g9805 ( 
.A(n_8840),
.B(n_8905),
.Y(n_9805)
);

INVx1_ASAP7_75t_L g9806 ( 
.A(n_8945),
.Y(n_9806)
);

INVx2_ASAP7_75t_L g9807 ( 
.A(n_8350),
.Y(n_9807)
);

AND2x2_ASAP7_75t_L g9808 ( 
.A(n_8410),
.B(n_7138),
.Y(n_9808)
);

INVx1_ASAP7_75t_L g9809 ( 
.A(n_8949),
.Y(n_9809)
);

INVx6_ASAP7_75t_L g9810 ( 
.A(n_7867),
.Y(n_9810)
);

INVx2_ASAP7_75t_L g9811 ( 
.A(n_8350),
.Y(n_9811)
);

BUFx2_ASAP7_75t_L g9812 ( 
.A(n_8159),
.Y(n_9812)
);

INVx1_ASAP7_75t_L g9813 ( 
.A(n_8949),
.Y(n_9813)
);

INVx2_ASAP7_75t_L g9814 ( 
.A(n_8350),
.Y(n_9814)
);

BUFx3_ASAP7_75t_L g9815 ( 
.A(n_8195),
.Y(n_9815)
);

INVx2_ASAP7_75t_L g9816 ( 
.A(n_8350),
.Y(n_9816)
);

OAI21x1_ASAP7_75t_L g9817 ( 
.A1(n_7692),
.A2(n_6774),
.B(n_6769),
.Y(n_9817)
);

INVx2_ASAP7_75t_L g9818 ( 
.A(n_8350),
.Y(n_9818)
);

AOI22xp33_ASAP7_75t_L g9819 ( 
.A1(n_8219),
.A2(n_8758),
.B1(n_8756),
.B2(n_8610),
.Y(n_9819)
);

INVx2_ASAP7_75t_L g9820 ( 
.A(n_8350),
.Y(n_9820)
);

INVx2_ASAP7_75t_L g9821 ( 
.A(n_7670),
.Y(n_9821)
);

INVx1_ASAP7_75t_L g9822 ( 
.A(n_8230),
.Y(n_9822)
);

AOI21x1_ASAP7_75t_L g9823 ( 
.A1(n_7728),
.A2(n_7481),
.B(n_7478),
.Y(n_9823)
);

AND2x2_ASAP7_75t_L g9824 ( 
.A(n_8410),
.B(n_7138),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_8230),
.Y(n_9825)
);

AOI22xp33_ASAP7_75t_L g9826 ( 
.A1(n_8758),
.A2(n_6576),
.B1(n_6570),
.B2(n_7499),
.Y(n_9826)
);

INVx2_ASAP7_75t_L g9827 ( 
.A(n_7670),
.Y(n_9827)
);

AOI22xp33_ASAP7_75t_L g9828 ( 
.A1(n_8610),
.A2(n_6576),
.B1(n_6570),
.B2(n_7468),
.Y(n_9828)
);

AOI22xp33_ASAP7_75t_SL g9829 ( 
.A1(n_7790),
.A2(n_7570),
.B1(n_7551),
.B2(n_7461),
.Y(n_9829)
);

INVx2_ASAP7_75t_L g9830 ( 
.A(n_7670),
.Y(n_9830)
);

AOI22xp33_ASAP7_75t_L g9831 ( 
.A1(n_8617),
.A2(n_6576),
.B1(n_6570),
.B2(n_7551),
.Y(n_9831)
);

INVx2_ASAP7_75t_L g9832 ( 
.A(n_7670),
.Y(n_9832)
);

INVx1_ASAP7_75t_L g9833 ( 
.A(n_8244),
.Y(n_9833)
);

AOI22xp5_ASAP7_75t_L g9834 ( 
.A1(n_7623),
.A2(n_7374),
.B1(n_7361),
.B2(n_7351),
.Y(n_9834)
);

OAI21xp33_ASAP7_75t_L g9835 ( 
.A1(n_8039),
.A2(n_6868),
.B(n_6838),
.Y(n_9835)
);

BUFx2_ASAP7_75t_R g9836 ( 
.A(n_7651),
.Y(n_9836)
);

BUFx3_ASAP7_75t_L g9837 ( 
.A(n_8195),
.Y(n_9837)
);

HB1xp67_ASAP7_75t_L g9838 ( 
.A(n_8415),
.Y(n_9838)
);

AND2x4_ASAP7_75t_L g9839 ( 
.A(n_8457),
.B(n_7551),
.Y(n_9839)
);

BUFx3_ASAP7_75t_L g9840 ( 
.A(n_8195),
.Y(n_9840)
);

INVx2_ASAP7_75t_L g9841 ( 
.A(n_7679),
.Y(n_9841)
);

INVx1_ASAP7_75t_L g9842 ( 
.A(n_8244),
.Y(n_9842)
);

INVx2_ASAP7_75t_L g9843 ( 
.A(n_7679),
.Y(n_9843)
);

INVx2_ASAP7_75t_L g9844 ( 
.A(n_7679),
.Y(n_9844)
);

OAI22xp33_ASAP7_75t_L g9845 ( 
.A1(n_7964),
.A2(n_7578),
.B1(n_7603),
.B2(n_6919),
.Y(n_9845)
);

INVx2_ASAP7_75t_L g9846 ( 
.A(n_7679),
.Y(n_9846)
);

INVx2_ASAP7_75t_L g9847 ( 
.A(n_7682),
.Y(n_9847)
);

AOI22xp33_ASAP7_75t_SL g9848 ( 
.A1(n_8136),
.A2(n_7461),
.B1(n_7517),
.B2(n_7484),
.Y(n_9848)
);

INVx1_ASAP7_75t_L g9849 ( 
.A(n_8266),
.Y(n_9849)
);

OAI21x1_ASAP7_75t_L g9850 ( 
.A1(n_7692),
.A2(n_6774),
.B(n_6769),
.Y(n_9850)
);

INVx2_ASAP7_75t_L g9851 ( 
.A(n_7682),
.Y(n_9851)
);

OAI21x1_ASAP7_75t_L g9852 ( 
.A1(n_8877),
.A2(n_6785),
.B(n_6774),
.Y(n_9852)
);

AND2x4_ASAP7_75t_L g9853 ( 
.A(n_8457),
.B(n_7570),
.Y(n_9853)
);

INVx2_ASAP7_75t_L g9854 ( 
.A(n_7682),
.Y(n_9854)
);

BUFx3_ASAP7_75t_L g9855 ( 
.A(n_8226),
.Y(n_9855)
);

NAND2xp5_ASAP7_75t_L g9856 ( 
.A(n_8905),
.B(n_6793),
.Y(n_9856)
);

INVx2_ASAP7_75t_L g9857 ( 
.A(n_7682),
.Y(n_9857)
);

AO21x1_ASAP7_75t_L g9858 ( 
.A1(n_8049),
.A2(n_8082),
.B(n_7672),
.Y(n_9858)
);

INVx2_ASAP7_75t_L g9859 ( 
.A(n_7722),
.Y(n_9859)
);

OAI21x1_ASAP7_75t_L g9860 ( 
.A1(n_8877),
.A2(n_6785),
.B(n_6774),
.Y(n_9860)
);

INVx1_ASAP7_75t_L g9861 ( 
.A(n_8266),
.Y(n_9861)
);

HB1xp67_ASAP7_75t_L g9862 ( 
.A(n_8513),
.Y(n_9862)
);

NAND2x1p5_ASAP7_75t_L g9863 ( 
.A(n_8319),
.B(n_6575),
.Y(n_9863)
);

INVx1_ASAP7_75t_L g9864 ( 
.A(n_8286),
.Y(n_9864)
);

AND2x2_ASAP7_75t_L g9865 ( 
.A(n_8438),
.B(n_7344),
.Y(n_9865)
);

HB1xp67_ASAP7_75t_L g9866 ( 
.A(n_8513),
.Y(n_9866)
);

INVx2_ASAP7_75t_L g9867 ( 
.A(n_7722),
.Y(n_9867)
);

INVx2_ASAP7_75t_L g9868 ( 
.A(n_7722),
.Y(n_9868)
);

HB1xp67_ASAP7_75t_L g9869 ( 
.A(n_8635),
.Y(n_9869)
);

OA21x2_ASAP7_75t_L g9870 ( 
.A1(n_7775),
.A2(n_7016),
.B(n_6990),
.Y(n_9870)
);

AOI22xp33_ASAP7_75t_L g9871 ( 
.A1(n_8617),
.A2(n_6576),
.B1(n_6570),
.B2(n_7570),
.Y(n_9871)
);

OA21x2_ASAP7_75t_L g9872 ( 
.A1(n_7775),
.A2(n_7016),
.B(n_6990),
.Y(n_9872)
);

AOI22xp5_ASAP7_75t_L g9873 ( 
.A1(n_7718),
.A2(n_7461),
.B1(n_7517),
.B2(n_7484),
.Y(n_9873)
);

INVx1_ASAP7_75t_L g9874 ( 
.A(n_8286),
.Y(n_9874)
);

INVx1_ASAP7_75t_L g9875 ( 
.A(n_8289),
.Y(n_9875)
);

AND2x2_ASAP7_75t_L g9876 ( 
.A(n_8438),
.B(n_7344),
.Y(n_9876)
);

INVx2_ASAP7_75t_L g9877 ( 
.A(n_7722),
.Y(n_9877)
);

INVx2_ASAP7_75t_L g9878 ( 
.A(n_7742),
.Y(n_9878)
);

INVx1_ASAP7_75t_L g9879 ( 
.A(n_8289),
.Y(n_9879)
);

AND2x4_ASAP7_75t_L g9880 ( 
.A(n_8482),
.B(n_7570),
.Y(n_9880)
);

AO21x1_ASAP7_75t_SL g9881 ( 
.A1(n_8463),
.A2(n_7328),
.B(n_7331),
.Y(n_9881)
);

INVx2_ASAP7_75t_L g9882 ( 
.A(n_7742),
.Y(n_9882)
);

AO21x1_ASAP7_75t_L g9883 ( 
.A1(n_8049),
.A2(n_7396),
.B(n_7084),
.Y(n_9883)
);

INVx2_ASAP7_75t_L g9884 ( 
.A(n_7742),
.Y(n_9884)
);

INVx1_ASAP7_75t_L g9885 ( 
.A(n_8294),
.Y(n_9885)
);

BUFx2_ASAP7_75t_L g9886 ( 
.A(n_8159),
.Y(n_9886)
);

OAI22xp5_ASAP7_75t_L g9887 ( 
.A1(n_8166),
.A2(n_7328),
.B1(n_7541),
.B2(n_7540),
.Y(n_9887)
);

BUFx2_ASAP7_75t_SL g9888 ( 
.A(n_7651),
.Y(n_9888)
);

INVx2_ASAP7_75t_L g9889 ( 
.A(n_7742),
.Y(n_9889)
);

HB1xp67_ASAP7_75t_L g9890 ( 
.A(n_8415),
.Y(n_9890)
);

AND2x2_ASAP7_75t_L g9891 ( 
.A(n_8438),
.B(n_8493),
.Y(n_9891)
);

INVx1_ASAP7_75t_L g9892 ( 
.A(n_8294),
.Y(n_9892)
);

OAI21x1_ASAP7_75t_L g9893 ( 
.A1(n_8877),
.A2(n_6785),
.B(n_6774),
.Y(n_9893)
);

INVx1_ASAP7_75t_L g9894 ( 
.A(n_8295),
.Y(n_9894)
);

BUFx6f_ASAP7_75t_L g9895 ( 
.A(n_8226),
.Y(n_9895)
);

NOR2xp33_ASAP7_75t_L g9896 ( 
.A(n_8329),
.B(n_7461),
.Y(n_9896)
);

BUFx6f_ASAP7_75t_L g9897 ( 
.A(n_8226),
.Y(n_9897)
);

INVx2_ASAP7_75t_L g9898 ( 
.A(n_7751),
.Y(n_9898)
);

INVx1_ASAP7_75t_L g9899 ( 
.A(n_8295),
.Y(n_9899)
);

OAI21x1_ASAP7_75t_L g9900 ( 
.A1(n_8885),
.A2(n_6785),
.B(n_6774),
.Y(n_9900)
);

INVx2_ASAP7_75t_L g9901 ( 
.A(n_7751),
.Y(n_9901)
);

INVx1_ASAP7_75t_L g9902 ( 
.A(n_8299),
.Y(n_9902)
);

INVx1_ASAP7_75t_L g9903 ( 
.A(n_8299),
.Y(n_9903)
);

INVx1_ASAP7_75t_L g9904 ( 
.A(n_8302),
.Y(n_9904)
);

INVx2_ASAP7_75t_L g9905 ( 
.A(n_7751),
.Y(n_9905)
);

AND2x2_ASAP7_75t_L g9906 ( 
.A(n_8493),
.B(n_7344),
.Y(n_9906)
);

NAND2xp5_ASAP7_75t_L g9907 ( 
.A(n_8684),
.B(n_6793),
.Y(n_9907)
);

AND2x2_ASAP7_75t_L g9908 ( 
.A(n_8493),
.B(n_7344),
.Y(n_9908)
);

INVx3_ASAP7_75t_L g9909 ( 
.A(n_8020),
.Y(n_9909)
);

CKINVDCx14_ASAP7_75t_R g9910 ( 
.A(n_8213),
.Y(n_9910)
);

INVx1_ASAP7_75t_L g9911 ( 
.A(n_8302),
.Y(n_9911)
);

NAND2xp5_ASAP7_75t_L g9912 ( 
.A(n_8684),
.B(n_6799),
.Y(n_9912)
);

AOI22xp33_ASAP7_75t_L g9913 ( 
.A1(n_8144),
.A2(n_8322),
.B1(n_8298),
.B2(n_8233),
.Y(n_9913)
);

AND2x2_ASAP7_75t_L g9914 ( 
.A(n_8494),
.B(n_7526),
.Y(n_9914)
);

CKINVDCx11_ASAP7_75t_R g9915 ( 
.A(n_7651),
.Y(n_9915)
);

INVx2_ASAP7_75t_L g9916 ( 
.A(n_7751),
.Y(n_9916)
);

INVx1_ASAP7_75t_L g9917 ( 
.A(n_8305),
.Y(n_9917)
);

INVx3_ASAP7_75t_L g9918 ( 
.A(n_8020),
.Y(n_9918)
);

BUFx12f_ASAP7_75t_L g9919 ( 
.A(n_8132),
.Y(n_9919)
);

INVx2_ASAP7_75t_L g9920 ( 
.A(n_7760),
.Y(n_9920)
);

OAI22xp5_ASAP7_75t_L g9921 ( 
.A1(n_7931),
.A2(n_7541),
.B1(n_7540),
.B2(n_7331),
.Y(n_9921)
);

INVx2_ASAP7_75t_L g9922 ( 
.A(n_7760),
.Y(n_9922)
);

BUFx6f_ASAP7_75t_L g9923 ( 
.A(n_8226),
.Y(n_9923)
);

INVx1_ASAP7_75t_L g9924 ( 
.A(n_8305),
.Y(n_9924)
);

INVx2_ASAP7_75t_L g9925 ( 
.A(n_7760),
.Y(n_9925)
);

BUFx3_ASAP7_75t_L g9926 ( 
.A(n_8241),
.Y(n_9926)
);

OAI21x1_ASAP7_75t_L g9927 ( 
.A1(n_8885),
.A2(n_6794),
.B(n_6785),
.Y(n_9927)
);

BUFx6f_ASAP7_75t_L g9928 ( 
.A(n_8241),
.Y(n_9928)
);

INVx2_ASAP7_75t_L g9929 ( 
.A(n_7760),
.Y(n_9929)
);

OA21x2_ASAP7_75t_L g9930 ( 
.A1(n_8063),
.A2(n_7059),
.B(n_7058),
.Y(n_9930)
);

INVx2_ASAP7_75t_L g9931 ( 
.A(n_7805),
.Y(n_9931)
);

CKINVDCx16_ASAP7_75t_R g9932 ( 
.A(n_8554),
.Y(n_9932)
);

OAI22xp5_ASAP7_75t_L g9933 ( 
.A1(n_7931),
.A2(n_7287),
.B1(n_7593),
.B2(n_7578),
.Y(n_9933)
);

OAI22xp33_ASAP7_75t_L g9934 ( 
.A1(n_7713),
.A2(n_7578),
.B1(n_7603),
.B2(n_6919),
.Y(n_9934)
);

BUFx12f_ASAP7_75t_L g9935 ( 
.A(n_8250),
.Y(n_9935)
);

INVx1_ASAP7_75t_L g9936 ( 
.A(n_7915),
.Y(n_9936)
);

INVx2_ASAP7_75t_L g9937 ( 
.A(n_7805),
.Y(n_9937)
);

OAI21xp5_ASAP7_75t_L g9938 ( 
.A1(n_7815),
.A2(n_6876),
.B(n_7287),
.Y(n_9938)
);

INVx4_ASAP7_75t_L g9939 ( 
.A(n_8042),
.Y(n_9939)
);

INVx2_ASAP7_75t_SL g9940 ( 
.A(n_8241),
.Y(n_9940)
);

OA21x2_ASAP7_75t_L g9941 ( 
.A1(n_8063),
.A2(n_7059),
.B(n_7058),
.Y(n_9941)
);

AOI22xp33_ASAP7_75t_SL g9942 ( 
.A1(n_7790),
.A2(n_7570),
.B1(n_7517),
.B2(n_7554),
.Y(n_9942)
);

HB1xp67_ASAP7_75t_L g9943 ( 
.A(n_8635),
.Y(n_9943)
);

INVx1_ASAP7_75t_L g9944 ( 
.A(n_7915),
.Y(n_9944)
);

INVx2_ASAP7_75t_L g9945 ( 
.A(n_7805),
.Y(n_9945)
);

INVx1_ASAP7_75t_L g9946 ( 
.A(n_7917),
.Y(n_9946)
);

AO21x2_ASAP7_75t_L g9947 ( 
.A1(n_8570),
.A2(n_7577),
.B(n_6661),
.Y(n_9947)
);

INVx2_ASAP7_75t_L g9948 ( 
.A(n_7805),
.Y(n_9948)
);

INVx1_ASAP7_75t_SL g9949 ( 
.A(n_8022),
.Y(n_9949)
);

AOI21x1_ASAP7_75t_L g9950 ( 
.A1(n_7728),
.A2(n_7533),
.B(n_7485),
.Y(n_9950)
);

INVx1_ASAP7_75t_L g9951 ( 
.A(n_7917),
.Y(n_9951)
);

BUFx12f_ASAP7_75t_L g9952 ( 
.A(n_8250),
.Y(n_9952)
);

NOR2xp33_ASAP7_75t_L g9953 ( 
.A(n_8329),
.B(n_7484),
.Y(n_9953)
);

INVx2_ASAP7_75t_L g9954 ( 
.A(n_7853),
.Y(n_9954)
);

INVx1_ASAP7_75t_L g9955 ( 
.A(n_7928),
.Y(n_9955)
);

AND2x2_ASAP7_75t_L g9956 ( 
.A(n_8494),
.B(n_7526),
.Y(n_9956)
);

INVx1_ASAP7_75t_L g9957 ( 
.A(n_7928),
.Y(n_9957)
);

OAI21x1_ASAP7_75t_L g9958 ( 
.A1(n_8885),
.A2(n_6794),
.B(n_6785),
.Y(n_9958)
);

INVx1_ASAP7_75t_L g9959 ( 
.A(n_7929),
.Y(n_9959)
);

CKINVDCx5p33_ASAP7_75t_R g9960 ( 
.A(n_8745),
.Y(n_9960)
);

INVx1_ASAP7_75t_L g9961 ( 
.A(n_7929),
.Y(n_9961)
);

AND2x2_ASAP7_75t_L g9962 ( 
.A(n_8494),
.B(n_7526),
.Y(n_9962)
);

AO21x1_ASAP7_75t_SL g9963 ( 
.A1(n_8198),
.A2(n_8799),
.B(n_8755),
.Y(n_9963)
);

INVx2_ASAP7_75t_L g9964 ( 
.A(n_7853),
.Y(n_9964)
);

CKINVDCx11_ASAP7_75t_R g9965 ( 
.A(n_8161),
.Y(n_9965)
);

OAI22xp5_ASAP7_75t_L g9966 ( 
.A1(n_7962),
.A2(n_7287),
.B1(n_7603),
.B2(n_6941),
.Y(n_9966)
);

INVx6_ASAP7_75t_L g9967 ( 
.A(n_7867),
.Y(n_9967)
);

INVx1_ASAP7_75t_L g9968 ( 
.A(n_7934),
.Y(n_9968)
);

INVx2_ASAP7_75t_L g9969 ( 
.A(n_7853),
.Y(n_9969)
);

AND2x4_ASAP7_75t_SL g9970 ( 
.A(n_8042),
.B(n_6690),
.Y(n_9970)
);

CKINVDCx11_ASAP7_75t_R g9971 ( 
.A(n_8161),
.Y(n_9971)
);

OAI21x1_ASAP7_75t_L g9972 ( 
.A1(n_8762),
.A2(n_6839),
.B(n_6794),
.Y(n_9972)
);

NAND2x1p5_ASAP7_75t_L g9973 ( 
.A(n_8319),
.B(n_6575),
.Y(n_9973)
);

INVx1_ASAP7_75t_L g9974 ( 
.A(n_7934),
.Y(n_9974)
);

BUFx3_ASAP7_75t_L g9975 ( 
.A(n_8241),
.Y(n_9975)
);

AO21x2_ASAP7_75t_L g9976 ( 
.A1(n_8570),
.A2(n_7577),
.B(n_6661),
.Y(n_9976)
);

INVx1_ASAP7_75t_L g9977 ( 
.A(n_7935),
.Y(n_9977)
);

AOI22xp33_ASAP7_75t_L g9978 ( 
.A1(n_8144),
.A2(n_6570),
.B1(n_7570),
.B2(n_7086),
.Y(n_9978)
);

INVx2_ASAP7_75t_L g9979 ( 
.A(n_7853),
.Y(n_9979)
);

AOI22xp5_ASAP7_75t_L g9980 ( 
.A1(n_7718),
.A2(n_7517),
.B1(n_7554),
.B2(n_7484),
.Y(n_9980)
);

HB1xp67_ASAP7_75t_L g9981 ( 
.A(n_8640),
.Y(n_9981)
);

INVx2_ASAP7_75t_L g9982 ( 
.A(n_7871),
.Y(n_9982)
);

INVx2_ASAP7_75t_L g9983 ( 
.A(n_7871),
.Y(n_9983)
);

INVx2_ASAP7_75t_L g9984 ( 
.A(n_7871),
.Y(n_9984)
);

INVx2_ASAP7_75t_L g9985 ( 
.A(n_7871),
.Y(n_9985)
);

HB1xp67_ASAP7_75t_L g9986 ( 
.A(n_8640),
.Y(n_9986)
);

BUFx2_ASAP7_75t_L g9987 ( 
.A(n_8159),
.Y(n_9987)
);

INVx1_ASAP7_75t_L g9988 ( 
.A(n_7935),
.Y(n_9988)
);

INVx6_ASAP7_75t_L g9989 ( 
.A(n_7867),
.Y(n_9989)
);

OAI21x1_ASAP7_75t_L g9990 ( 
.A1(n_8762),
.A2(n_6839),
.B(n_6794),
.Y(n_9990)
);

INVx2_ASAP7_75t_L g9991 ( 
.A(n_7877),
.Y(n_9991)
);

BUFx2_ASAP7_75t_L g9992 ( 
.A(n_8159),
.Y(n_9992)
);

INVx3_ASAP7_75t_SL g9993 ( 
.A(n_8712),
.Y(n_9993)
);

INVx2_ASAP7_75t_L g9994 ( 
.A(n_7877),
.Y(n_9994)
);

INVx1_ASAP7_75t_L g9995 ( 
.A(n_7957),
.Y(n_9995)
);

NAND2x1p5_ASAP7_75t_L g9996 ( 
.A(n_8319),
.B(n_6575),
.Y(n_9996)
);

INVx3_ASAP7_75t_L g9997 ( 
.A(n_8020),
.Y(n_9997)
);

INVx1_ASAP7_75t_L g9998 ( 
.A(n_7957),
.Y(n_9998)
);

NAND2xp5_ASAP7_75t_L g9999 ( 
.A(n_8744),
.B(n_6799),
.Y(n_9999)
);

CKINVDCx6p67_ASAP7_75t_R g10000 ( 
.A(n_7788),
.Y(n_10000)
);

BUFx3_ASAP7_75t_L g10001 ( 
.A(n_8292),
.Y(n_10001)
);

OAI21x1_ASAP7_75t_L g10002 ( 
.A1(n_8762),
.A2(n_6839),
.B(n_6794),
.Y(n_10002)
);

NAND2xp5_ASAP7_75t_L g10003 ( 
.A(n_8744),
.B(n_6807),
.Y(n_10003)
);

BUFx3_ASAP7_75t_L g10004 ( 
.A(n_8292),
.Y(n_10004)
);

INVx3_ASAP7_75t_L g10005 ( 
.A(n_8020),
.Y(n_10005)
);

INVx1_ASAP7_75t_L g10006 ( 
.A(n_7965),
.Y(n_10006)
);

INVx1_ASAP7_75t_L g10007 ( 
.A(n_7965),
.Y(n_10007)
);

AND2x4_ASAP7_75t_L g10008 ( 
.A(n_8482),
.B(n_7570),
.Y(n_10008)
);

INVx1_ASAP7_75t_L g10009 ( 
.A(n_7976),
.Y(n_10009)
);

INVx1_ASAP7_75t_L g10010 ( 
.A(n_7976),
.Y(n_10010)
);

INVx2_ASAP7_75t_L g10011 ( 
.A(n_7877),
.Y(n_10011)
);

INVx1_ASAP7_75t_L g10012 ( 
.A(n_7992),
.Y(n_10012)
);

INVx1_ASAP7_75t_SL g10013 ( 
.A(n_8022),
.Y(n_10013)
);

OAI21xp5_ASAP7_75t_L g10014 ( 
.A1(n_7815),
.A2(n_6876),
.B(n_7237),
.Y(n_10014)
);

INVx2_ASAP7_75t_SL g10015 ( 
.A(n_8292),
.Y(n_10015)
);

INVx1_ASAP7_75t_SL g10016 ( 
.A(n_8102),
.Y(n_10016)
);

AO21x2_ASAP7_75t_L g10017 ( 
.A1(n_8570),
.A2(n_6661),
.B(n_7263),
.Y(n_10017)
);

BUFx2_ASAP7_75t_L g10018 ( 
.A(n_8159),
.Y(n_10018)
);

OAI22xp33_ASAP7_75t_L g10019 ( 
.A1(n_7713),
.A2(n_6919),
.B1(n_7255),
.B2(n_6690),
.Y(n_10019)
);

AOI21x1_ASAP7_75t_L g10020 ( 
.A1(n_8479),
.A2(n_7533),
.B(n_7485),
.Y(n_10020)
);

INVx1_ASAP7_75t_L g10021 ( 
.A(n_7992),
.Y(n_10021)
);

OAI21x1_ASAP7_75t_L g10022 ( 
.A1(n_7810),
.A2(n_6839),
.B(n_6794),
.Y(n_10022)
);

BUFx3_ASAP7_75t_L g10023 ( 
.A(n_8292),
.Y(n_10023)
);

OAI22xp5_ASAP7_75t_L g10024 ( 
.A1(n_7962),
.A2(n_6941),
.B1(n_6952),
.B2(n_6912),
.Y(n_10024)
);

AOI22xp33_ASAP7_75t_L g10025 ( 
.A1(n_8144),
.A2(n_6570),
.B1(n_7570),
.B2(n_7086),
.Y(n_10025)
);

OAI21x1_ASAP7_75t_L g10026 ( 
.A1(n_7810),
.A2(n_6843),
.B(n_6839),
.Y(n_10026)
);

INVx1_ASAP7_75t_L g10027 ( 
.A(n_7996),
.Y(n_10027)
);

AOI22xp33_ASAP7_75t_L g10028 ( 
.A1(n_8322),
.A2(n_7570),
.B1(n_7069),
.B2(n_7094),
.Y(n_10028)
);

BUFx2_ASAP7_75t_L g10029 ( 
.A(n_8159),
.Y(n_10029)
);

INVx1_ASAP7_75t_L g10030 ( 
.A(n_7996),
.Y(n_10030)
);

INVx1_ASAP7_75t_L g10031 ( 
.A(n_7997),
.Y(n_10031)
);

AOI22xp33_ASAP7_75t_SL g10032 ( 
.A1(n_8136),
.A2(n_7554),
.B1(n_6941),
.B2(n_6952),
.Y(n_10032)
);

INVxp67_ASAP7_75t_SL g10033 ( 
.A(n_8839),
.Y(n_10033)
);

BUFx2_ASAP7_75t_R g10034 ( 
.A(n_8161),
.Y(n_10034)
);

INVx2_ASAP7_75t_L g10035 ( 
.A(n_7877),
.Y(n_10035)
);

CKINVDCx11_ASAP7_75t_R g10036 ( 
.A(n_8542),
.Y(n_10036)
);

INVx2_ASAP7_75t_L g10037 ( 
.A(n_7885),
.Y(n_10037)
);

INVx1_ASAP7_75t_L g10038 ( 
.A(n_7997),
.Y(n_10038)
);

INVx2_ASAP7_75t_L g10039 ( 
.A(n_7885),
.Y(n_10039)
);

CKINVDCx5p33_ASAP7_75t_R g10040 ( 
.A(n_8745),
.Y(n_10040)
);

INVx2_ASAP7_75t_L g10041 ( 
.A(n_7885),
.Y(n_10041)
);

AOI22xp33_ASAP7_75t_L g10042 ( 
.A1(n_8298),
.A2(n_7069),
.B1(n_7094),
.B2(n_7086),
.Y(n_10042)
);

INVx1_ASAP7_75t_L g10043 ( 
.A(n_8001),
.Y(n_10043)
);

OR2x6_ASAP7_75t_L g10044 ( 
.A(n_7609),
.B(n_7077),
.Y(n_10044)
);

INVx2_ASAP7_75t_L g10045 ( 
.A(n_7885),
.Y(n_10045)
);

INVx1_ASAP7_75t_L g10046 ( 
.A(n_8001),
.Y(n_10046)
);

INVx2_ASAP7_75t_L g10047 ( 
.A(n_7897),
.Y(n_10047)
);

INVx2_ASAP7_75t_L g10048 ( 
.A(n_7897),
.Y(n_10048)
);

INVx2_ASAP7_75t_L g10049 ( 
.A(n_7897),
.Y(n_10049)
);

AOI22xp33_ASAP7_75t_SL g10050 ( 
.A1(n_8082),
.A2(n_7554),
.B1(n_6941),
.B2(n_6952),
.Y(n_10050)
);

AOI22xp33_ASAP7_75t_L g10051 ( 
.A1(n_8233),
.A2(n_7069),
.B1(n_7094),
.B2(n_7086),
.Y(n_10051)
);

INVx1_ASAP7_75t_L g10052 ( 
.A(n_8008),
.Y(n_10052)
);

INVx1_ASAP7_75t_L g10053 ( 
.A(n_8008),
.Y(n_10053)
);

INVx2_ASAP7_75t_L g10054 ( 
.A(n_7897),
.Y(n_10054)
);

CKINVDCx14_ASAP7_75t_R g10055 ( 
.A(n_8213),
.Y(n_10055)
);

AO21x2_ASAP7_75t_L g10056 ( 
.A1(n_7738),
.A2(n_7263),
.B(n_7288),
.Y(n_10056)
);

INVx1_ASAP7_75t_L g10057 ( 
.A(n_8025),
.Y(n_10057)
);

BUFx8_ASAP7_75t_L g10058 ( 
.A(n_8892),
.Y(n_10058)
);

INVx1_ASAP7_75t_L g10059 ( 
.A(n_8025),
.Y(n_10059)
);

INVx1_ASAP7_75t_L g10060 ( 
.A(n_8028),
.Y(n_10060)
);

BUFx2_ASAP7_75t_L g10061 ( 
.A(n_8159),
.Y(n_10061)
);

INVx1_ASAP7_75t_L g10062 ( 
.A(n_8028),
.Y(n_10062)
);

INVx1_ASAP7_75t_L g10063 ( 
.A(n_8034),
.Y(n_10063)
);

BUFx2_ASAP7_75t_L g10064 ( 
.A(n_8159),
.Y(n_10064)
);

BUFx6f_ASAP7_75t_L g10065 ( 
.A(n_8320),
.Y(n_10065)
);

OAI22xp33_ASAP7_75t_L g10066 ( 
.A1(n_8018),
.A2(n_8078),
.B1(n_7862),
.B2(n_8364),
.Y(n_10066)
);

AND2x4_ASAP7_75t_L g10067 ( 
.A(n_8482),
.B(n_7069),
.Y(n_10067)
);

AO21x1_ASAP7_75t_L g10068 ( 
.A1(n_7672),
.A2(n_7084),
.B(n_7080),
.Y(n_10068)
);

INVx1_ASAP7_75t_L g10069 ( 
.A(n_8034),
.Y(n_10069)
);

BUFx8_ASAP7_75t_SL g10070 ( 
.A(n_8712),
.Y(n_10070)
);

INVx2_ASAP7_75t_L g10071 ( 
.A(n_7904),
.Y(n_10071)
);

OAI22xp5_ASAP7_75t_L g10072 ( 
.A1(n_8164),
.A2(n_6952),
.B1(n_6961),
.B2(n_6912),
.Y(n_10072)
);

BUFx2_ASAP7_75t_L g10073 ( 
.A(n_8631),
.Y(n_10073)
);

AOI22xp33_ASAP7_75t_L g10074 ( 
.A1(n_7876),
.A2(n_7094),
.B1(n_7122),
.B2(n_7119),
.Y(n_10074)
);

INVx6_ASAP7_75t_L g10075 ( 
.A(n_7867),
.Y(n_10075)
);

HB1xp67_ASAP7_75t_L g10076 ( 
.A(n_8643),
.Y(n_10076)
);

OA21x2_ASAP7_75t_L g10077 ( 
.A1(n_8477),
.A2(n_7059),
.B(n_7058),
.Y(n_10077)
);

BUFx3_ASAP7_75t_L g10078 ( 
.A(n_8320),
.Y(n_10078)
);

INVx2_ASAP7_75t_SL g10079 ( 
.A(n_8320),
.Y(n_10079)
);

AOI22xp33_ASAP7_75t_L g10080 ( 
.A1(n_7876),
.A2(n_7119),
.B1(n_7165),
.B2(n_7122),
.Y(n_10080)
);

INVx2_ASAP7_75t_L g10081 ( 
.A(n_7904),
.Y(n_10081)
);

INVx1_ASAP7_75t_L g10082 ( 
.A(n_8040),
.Y(n_10082)
);

INVx1_ASAP7_75t_L g10083 ( 
.A(n_8040),
.Y(n_10083)
);

INVx3_ASAP7_75t_L g10084 ( 
.A(n_8020),
.Y(n_10084)
);

INVx2_ASAP7_75t_L g10085 ( 
.A(n_7904),
.Y(n_10085)
);

NAND2x1p5_ASAP7_75t_L g10086 ( 
.A(n_8319),
.B(n_6651),
.Y(n_10086)
);

NAND2xp5_ASAP7_75t_L g10087 ( 
.A(n_8807),
.B(n_8907),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_7904),
.Y(n_10088)
);

INVx3_ASAP7_75t_L g10089 ( 
.A(n_8020),
.Y(n_10089)
);

INVx1_ASAP7_75t_L g10090 ( 
.A(n_8045),
.Y(n_10090)
);

INVx1_ASAP7_75t_L g10091 ( 
.A(n_8045),
.Y(n_10091)
);

INVx1_ASAP7_75t_L g10092 ( 
.A(n_8048),
.Y(n_10092)
);

INVx1_ASAP7_75t_L g10093 ( 
.A(n_8048),
.Y(n_10093)
);

INVx1_ASAP7_75t_L g10094 ( 
.A(n_8061),
.Y(n_10094)
);

AOI22xp33_ASAP7_75t_L g10095 ( 
.A1(n_7876),
.A2(n_7119),
.B1(n_7165),
.B2(n_7122),
.Y(n_10095)
);

INVx2_ASAP7_75t_L g10096 ( 
.A(n_7913),
.Y(n_10096)
);

OAI21x1_ASAP7_75t_L g10097 ( 
.A1(n_7810),
.A2(n_8096),
.B(n_7948),
.Y(n_10097)
);

CKINVDCx20_ASAP7_75t_R g10098 ( 
.A(n_8481),
.Y(n_10098)
);

INVx1_ASAP7_75t_L g10099 ( 
.A(n_8061),
.Y(n_10099)
);

INVx1_ASAP7_75t_L g10100 ( 
.A(n_8067),
.Y(n_10100)
);

OAI22xp5_ASAP7_75t_L g10101 ( 
.A1(n_8164),
.A2(n_6961),
.B1(n_6979),
.B2(n_6912),
.Y(n_10101)
);

INVx2_ASAP7_75t_L g10102 ( 
.A(n_7913),
.Y(n_10102)
);

OAI22xp33_ASAP7_75t_L g10103 ( 
.A1(n_8018),
.A2(n_6919),
.B1(n_7255),
.B2(n_6690),
.Y(n_10103)
);

INVx1_ASAP7_75t_L g10104 ( 
.A(n_8067),
.Y(n_10104)
);

INVx2_ASAP7_75t_L g10105 ( 
.A(n_7913),
.Y(n_10105)
);

INVx2_ASAP7_75t_L g10106 ( 
.A(n_7913),
.Y(n_10106)
);

INVx2_ASAP7_75t_L g10107 ( 
.A(n_8749),
.Y(n_10107)
);

INVx1_ASAP7_75t_L g10108 ( 
.A(n_8071),
.Y(n_10108)
);

INVx1_ASAP7_75t_L g10109 ( 
.A(n_8071),
.Y(n_10109)
);

HB1xp67_ASAP7_75t_L g10110 ( 
.A(n_8650),
.Y(n_10110)
);

INVx2_ASAP7_75t_SL g10111 ( 
.A(n_8320),
.Y(n_10111)
);

INVx2_ASAP7_75t_L g10112 ( 
.A(n_8749),
.Y(n_10112)
);

INVx8_ASAP7_75t_L g10113 ( 
.A(n_8901),
.Y(n_10113)
);

BUFx8_ASAP7_75t_L g10114 ( 
.A(n_8892),
.Y(n_10114)
);

INVx1_ASAP7_75t_L g10115 ( 
.A(n_8085),
.Y(n_10115)
);

INVx1_ASAP7_75t_L g10116 ( 
.A(n_8085),
.Y(n_10116)
);

INVx1_ASAP7_75t_L g10117 ( 
.A(n_8092),
.Y(n_10117)
);

HB1xp67_ASAP7_75t_L g10118 ( 
.A(n_8643),
.Y(n_10118)
);

INVx2_ASAP7_75t_L g10119 ( 
.A(n_8749),
.Y(n_10119)
);

AOI22xp33_ASAP7_75t_L g10120 ( 
.A1(n_7876),
.A2(n_8270),
.B1(n_8273),
.B2(n_8594),
.Y(n_10120)
);

AOI21xp5_ASAP7_75t_L g10121 ( 
.A1(n_7834),
.A2(n_7288),
.B(n_7340),
.Y(n_10121)
);

AND2x2_ASAP7_75t_L g10122 ( 
.A(n_8605),
.B(n_7602),
.Y(n_10122)
);

BUFx2_ASAP7_75t_SL g10123 ( 
.A(n_8042),
.Y(n_10123)
);

INVx2_ASAP7_75t_L g10124 ( 
.A(n_8749),
.Y(n_10124)
);

NOR2xp33_ASAP7_75t_SL g10125 ( 
.A(n_8670),
.B(n_7486),
.Y(n_10125)
);

AOI21x1_ASAP7_75t_L g10126 ( 
.A1(n_8479),
.A2(n_7533),
.B(n_7485),
.Y(n_10126)
);

AOI22xp33_ASAP7_75t_L g10127 ( 
.A1(n_7876),
.A2(n_7119),
.B1(n_7146),
.B2(n_7122),
.Y(n_10127)
);

BUFx10_ASAP7_75t_L g10128 ( 
.A(n_8257),
.Y(n_10128)
);

INVx1_ASAP7_75t_L g10129 ( 
.A(n_8092),
.Y(n_10129)
);

INVx2_ASAP7_75t_L g10130 ( 
.A(n_8749),
.Y(n_10130)
);

INVx2_ASAP7_75t_L g10131 ( 
.A(n_8749),
.Y(n_10131)
);

INVx1_ASAP7_75t_SL g10132 ( 
.A(n_8102),
.Y(n_10132)
);

INVx1_ASAP7_75t_L g10133 ( 
.A(n_8097),
.Y(n_10133)
);

INVx1_ASAP7_75t_L g10134 ( 
.A(n_8097),
.Y(n_10134)
);

INVx2_ASAP7_75t_L g10135 ( 
.A(n_8406),
.Y(n_10135)
);

INVx1_ASAP7_75t_L g10136 ( 
.A(n_8101),
.Y(n_10136)
);

INVx1_ASAP7_75t_L g10137 ( 
.A(n_8101),
.Y(n_10137)
);

INVx3_ASAP7_75t_L g10138 ( 
.A(n_8020),
.Y(n_10138)
);

AND2x2_ASAP7_75t_L g10139 ( 
.A(n_8605),
.B(n_7602),
.Y(n_10139)
);

INVx1_ASAP7_75t_L g10140 ( 
.A(n_8106),
.Y(n_10140)
);

INVx4_ASAP7_75t_L g10141 ( 
.A(n_8042),
.Y(n_10141)
);

OAI22xp5_ASAP7_75t_SL g10142 ( 
.A1(n_8505),
.A2(n_7433),
.B1(n_7465),
.B2(n_7366),
.Y(n_10142)
);

INVx1_ASAP7_75t_L g10143 ( 
.A(n_8106),
.Y(n_10143)
);

INVxp33_ASAP7_75t_L g10144 ( 
.A(n_8182),
.Y(n_10144)
);

INVx1_ASAP7_75t_L g10145 ( 
.A(n_8107),
.Y(n_10145)
);

AOI22xp5_ASAP7_75t_L g10146 ( 
.A1(n_7685),
.A2(n_7340),
.B1(n_7467),
.B2(n_7465),
.Y(n_10146)
);

AOI22xp5_ASAP7_75t_L g10147 ( 
.A1(n_7685),
.A2(n_7340),
.B1(n_7521),
.B2(n_7467),
.Y(n_10147)
);

INVx1_ASAP7_75t_L g10148 ( 
.A(n_8107),
.Y(n_10148)
);

AOI22xp33_ASAP7_75t_L g10149 ( 
.A1(n_8270),
.A2(n_7146),
.B1(n_7280),
.B2(n_7165),
.Y(n_10149)
);

INVx2_ASAP7_75t_L g10150 ( 
.A(n_8406),
.Y(n_10150)
);

INVx3_ASAP7_75t_L g10151 ( 
.A(n_8168),
.Y(n_10151)
);

INVx1_ASAP7_75t_L g10152 ( 
.A(n_8110),
.Y(n_10152)
);

INVx1_ASAP7_75t_L g10153 ( 
.A(n_8110),
.Y(n_10153)
);

INVx1_ASAP7_75t_L g10154 ( 
.A(n_8112),
.Y(n_10154)
);

INVx2_ASAP7_75t_L g10155 ( 
.A(n_8406),
.Y(n_10155)
);

INVx2_ASAP7_75t_L g10156 ( 
.A(n_8422),
.Y(n_10156)
);

HB1xp67_ASAP7_75t_L g10157 ( 
.A(n_8650),
.Y(n_10157)
);

INVx1_ASAP7_75t_L g10158 ( 
.A(n_8112),
.Y(n_10158)
);

INVx2_ASAP7_75t_SL g10159 ( 
.A(n_8374),
.Y(n_10159)
);

HB1xp67_ASAP7_75t_L g10160 ( 
.A(n_8658),
.Y(n_10160)
);

BUFx4f_ASAP7_75t_L g10161 ( 
.A(n_8851),
.Y(n_10161)
);

INVx4_ASAP7_75t_SL g10162 ( 
.A(n_8542),
.Y(n_10162)
);

HB1xp67_ASAP7_75t_L g10163 ( 
.A(n_8658),
.Y(n_10163)
);

BUFx6f_ASAP7_75t_L g10164 ( 
.A(n_8374),
.Y(n_10164)
);

BUFx3_ASAP7_75t_L g10165 ( 
.A(n_8374),
.Y(n_10165)
);

INVx6_ASAP7_75t_L g10166 ( 
.A(n_8052),
.Y(n_10166)
);

AOI22xp33_ASAP7_75t_L g10167 ( 
.A1(n_8594),
.A2(n_7146),
.B1(n_7280),
.B2(n_7165),
.Y(n_10167)
);

NAND2xp5_ASAP7_75t_L g10168 ( 
.A(n_8807),
.B(n_6807),
.Y(n_10168)
);

OA21x2_ASAP7_75t_L g10169 ( 
.A1(n_8477),
.A2(n_7081),
.B(n_7062),
.Y(n_10169)
);

INVx5_ASAP7_75t_L g10170 ( 
.A(n_8168),
.Y(n_10170)
);

INVx2_ASAP7_75t_L g10171 ( 
.A(n_8422),
.Y(n_10171)
);

OAI22xp5_ASAP7_75t_L g10172 ( 
.A1(n_7719),
.A2(n_6961),
.B1(n_6979),
.B2(n_6912),
.Y(n_10172)
);

INVx2_ASAP7_75t_L g10173 ( 
.A(n_8422),
.Y(n_10173)
);

OAI22xp5_ASAP7_75t_L g10174 ( 
.A1(n_7719),
.A2(n_6979),
.B1(n_6986),
.B2(n_6961),
.Y(n_10174)
);

HB1xp67_ASAP7_75t_L g10175 ( 
.A(n_8724),
.Y(n_10175)
);

BUFx6f_ASAP7_75t_L g10176 ( 
.A(n_8374),
.Y(n_10176)
);

OAI22xp5_ASAP7_75t_L g10177 ( 
.A1(n_8134),
.A2(n_6986),
.B1(n_6998),
.B2(n_6979),
.Y(n_10177)
);

OAI21x1_ASAP7_75t_L g10178 ( 
.A1(n_8096),
.A2(n_6843),
.B(n_6839),
.Y(n_10178)
);

INVx2_ASAP7_75t_L g10179 ( 
.A(n_8428),
.Y(n_10179)
);

INVx8_ASAP7_75t_L g10180 ( 
.A(n_8901),
.Y(n_10180)
);

NAND2x1p5_ASAP7_75t_L g10181 ( 
.A(n_8319),
.B(n_6651),
.Y(n_10181)
);

INVx2_ASAP7_75t_L g10182 ( 
.A(n_8428),
.Y(n_10182)
);

CKINVDCx11_ASAP7_75t_R g10183 ( 
.A(n_8542),
.Y(n_10183)
);

AOI22xp33_ASAP7_75t_L g10184 ( 
.A1(n_8596),
.A2(n_7146),
.B1(n_7280),
.B2(n_6792),
.Y(n_10184)
);

HB1xp67_ASAP7_75t_L g10185 ( 
.A(n_8707),
.Y(n_10185)
);

AOI21x1_ASAP7_75t_L g10186 ( 
.A1(n_8479),
.A2(n_7560),
.B(n_7539),
.Y(n_10186)
);

INVx2_ASAP7_75t_L g10187 ( 
.A(n_8428),
.Y(n_10187)
);

INVx1_ASAP7_75t_SL g10188 ( 
.A(n_8306),
.Y(n_10188)
);

INVx1_ASAP7_75t_L g10189 ( 
.A(n_8114),
.Y(n_10189)
);

INVx1_ASAP7_75t_SL g10190 ( 
.A(n_8306),
.Y(n_10190)
);

AO21x1_ASAP7_75t_SL g10191 ( 
.A1(n_8198),
.A2(n_8799),
.B(n_8755),
.Y(n_10191)
);

OAI21x1_ASAP7_75t_L g10192 ( 
.A1(n_7947),
.A2(n_6859),
.B(n_6843),
.Y(n_10192)
);

INVx1_ASAP7_75t_SL g10193 ( 
.A(n_8351),
.Y(n_10193)
);

BUFx3_ASAP7_75t_L g10194 ( 
.A(n_8448),
.Y(n_10194)
);

INVx1_ASAP7_75t_L g10195 ( 
.A(n_8114),
.Y(n_10195)
);

BUFx4f_ASAP7_75t_L g10196 ( 
.A(n_8851),
.Y(n_10196)
);

AOI22xp33_ASAP7_75t_L g10197 ( 
.A1(n_8596),
.A2(n_7280),
.B1(n_6792),
.B2(n_6459),
.Y(n_10197)
);

INVx2_ASAP7_75t_L g10198 ( 
.A(n_8431),
.Y(n_10198)
);

OAI21x1_ASAP7_75t_SL g10199 ( 
.A1(n_8600),
.A2(n_7443),
.B(n_7428),
.Y(n_10199)
);

HB1xp67_ASAP7_75t_L g10200 ( 
.A(n_8707),
.Y(n_10200)
);

AND2x2_ASAP7_75t_L g10201 ( 
.A(n_8605),
.B(n_7602),
.Y(n_10201)
);

AND2x2_ASAP7_75t_L g10202 ( 
.A(n_8713),
.B(n_7602),
.Y(n_10202)
);

BUFx8_ASAP7_75t_SL g10203 ( 
.A(n_8739),
.Y(n_10203)
);

NAND2x1p5_ASAP7_75t_L g10204 ( 
.A(n_8319),
.B(n_6651),
.Y(n_10204)
);

INVx3_ASAP7_75t_L g10205 ( 
.A(n_8168),
.Y(n_10205)
);

BUFx8_ASAP7_75t_L g10206 ( 
.A(n_8892),
.Y(n_10206)
);

INVx2_ASAP7_75t_L g10207 ( 
.A(n_8431),
.Y(n_10207)
);

INVx2_ASAP7_75t_L g10208 ( 
.A(n_8431),
.Y(n_10208)
);

INVx2_ASAP7_75t_SL g10209 ( 
.A(n_8448),
.Y(n_10209)
);

INVx1_ASAP7_75t_L g10210 ( 
.A(n_8119),
.Y(n_10210)
);

INVx1_ASAP7_75t_L g10211 ( 
.A(n_8119),
.Y(n_10211)
);

INVx2_ASAP7_75t_L g10212 ( 
.A(n_8435),
.Y(n_10212)
);

AND2x4_ASAP7_75t_L g10213 ( 
.A(n_8482),
.B(n_7397),
.Y(n_10213)
);

INVx1_ASAP7_75t_L g10214 ( 
.A(n_8121),
.Y(n_10214)
);

AOI22xp33_ASAP7_75t_L g10215 ( 
.A1(n_8669),
.A2(n_6792),
.B1(n_6459),
.B2(n_6477),
.Y(n_10215)
);

INVx1_ASAP7_75t_L g10216 ( 
.A(n_8121),
.Y(n_10216)
);

INVx3_ASAP7_75t_L g10217 ( 
.A(n_8168),
.Y(n_10217)
);

INVx1_ASAP7_75t_L g10218 ( 
.A(n_8124),
.Y(n_10218)
);

HB1xp67_ASAP7_75t_L g10219 ( 
.A(n_8724),
.Y(n_10219)
);

INVx1_ASAP7_75t_L g10220 ( 
.A(n_8124),
.Y(n_10220)
);

AOI22xp33_ASAP7_75t_L g10221 ( 
.A1(n_8669),
.A2(n_6792),
.B1(n_6459),
.B2(n_6477),
.Y(n_10221)
);

OAI21x1_ASAP7_75t_L g10222 ( 
.A1(n_7947),
.A2(n_6859),
.B(n_6843),
.Y(n_10222)
);

HB1xp67_ASAP7_75t_L g10223 ( 
.A(n_8731),
.Y(n_10223)
);

AOI22xp5_ASAP7_75t_L g10224 ( 
.A1(n_8134),
.A2(n_7748),
.B1(n_7688),
.B2(n_7733),
.Y(n_10224)
);

AO21x1_ASAP7_75t_L g10225 ( 
.A1(n_8133),
.A2(n_7080),
.B(n_6831),
.Y(n_10225)
);

OA21x2_ASAP7_75t_L g10226 ( 
.A1(n_8477),
.A2(n_7081),
.B(n_7062),
.Y(n_10226)
);

INVx2_ASAP7_75t_L g10227 ( 
.A(n_8435),
.Y(n_10227)
);

INVx1_ASAP7_75t_L g10228 ( 
.A(n_8126),
.Y(n_10228)
);

INVx1_ASAP7_75t_L g10229 ( 
.A(n_8126),
.Y(n_10229)
);

INVx1_ASAP7_75t_L g10230 ( 
.A(n_8142),
.Y(n_10230)
);

AND2x2_ASAP7_75t_L g10231 ( 
.A(n_8713),
.B(n_7602),
.Y(n_10231)
);

OAI21x1_ASAP7_75t_L g10232 ( 
.A1(n_7947),
.A2(n_6859),
.B(n_6843),
.Y(n_10232)
);

AOI22xp33_ASAP7_75t_SL g10233 ( 
.A1(n_8773),
.A2(n_6998),
.B1(n_7052),
.B2(n_6986),
.Y(n_10233)
);

OA21x2_ASAP7_75t_L g10234 ( 
.A1(n_8478),
.A2(n_7081),
.B(n_7062),
.Y(n_10234)
);

OAI21x1_ASAP7_75t_L g10235 ( 
.A1(n_7948),
.A2(n_6859),
.B(n_6843),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_8142),
.Y(n_10236)
);

BUFx6f_ASAP7_75t_L g10237 ( 
.A(n_8448),
.Y(n_10237)
);

AND2x2_ASAP7_75t_L g10238 ( 
.A(n_8713),
.B(n_7602),
.Y(n_10238)
);

OAI21xp5_ASAP7_75t_L g10239 ( 
.A1(n_7821),
.A2(n_7237),
.B(n_6831),
.Y(n_10239)
);

INVx1_ASAP7_75t_L g10240 ( 
.A(n_8145),
.Y(n_10240)
);

AOI22xp33_ASAP7_75t_SL g10241 ( 
.A1(n_8773),
.A2(n_7724),
.B1(n_8078),
.B2(n_7739),
.Y(n_10241)
);

NOR2x1_ASAP7_75t_L g10242 ( 
.A(n_8516),
.B(n_7384),
.Y(n_10242)
);

INVx1_ASAP7_75t_L g10243 ( 
.A(n_8145),
.Y(n_10243)
);

CKINVDCx5p33_ASAP7_75t_R g10244 ( 
.A(n_8257),
.Y(n_10244)
);

INVx1_ASAP7_75t_L g10245 ( 
.A(n_8167),
.Y(n_10245)
);

AOI22xp33_ASAP7_75t_L g10246 ( 
.A1(n_7733),
.A2(n_8163),
.B1(n_8773),
.B2(n_8130),
.Y(n_10246)
);

OR2x2_ASAP7_75t_L g10247 ( 
.A(n_7797),
.B(n_7215),
.Y(n_10247)
);

NAND2x1p5_ASAP7_75t_L g10248 ( 
.A(n_8641),
.B(n_6651),
.Y(n_10248)
);

INVx2_ASAP7_75t_L g10249 ( 
.A(n_8435),
.Y(n_10249)
);

NAND2xp5_ASAP7_75t_L g10250 ( 
.A(n_8907),
.B(n_8607),
.Y(n_10250)
);

BUFx4f_ASAP7_75t_L g10251 ( 
.A(n_8851),
.Y(n_10251)
);

OAI21x1_ASAP7_75t_L g10252 ( 
.A1(n_7948),
.A2(n_6885),
.B(n_6859),
.Y(n_10252)
);

AO21x1_ASAP7_75t_L g10253 ( 
.A1(n_8133),
.A2(n_6826),
.B(n_6911),
.Y(n_10253)
);

OA21x2_ASAP7_75t_L g10254 ( 
.A1(n_8478),
.A2(n_7087),
.B(n_7085),
.Y(n_10254)
);

INVx1_ASAP7_75t_L g10255 ( 
.A(n_8167),
.Y(n_10255)
);

AO21x2_ASAP7_75t_L g10256 ( 
.A1(n_7738),
.A2(n_7263),
.B(n_6860),
.Y(n_10256)
);

AOI22xp5_ASAP7_75t_L g10257 ( 
.A1(n_7688),
.A2(n_7521),
.B1(n_7564),
.B2(n_7542),
.Y(n_10257)
);

INVx1_ASAP7_75t_L g10258 ( 
.A(n_8172),
.Y(n_10258)
);

INVx1_ASAP7_75t_L g10259 ( 
.A(n_8172),
.Y(n_10259)
);

INVx1_ASAP7_75t_L g10260 ( 
.A(n_8173),
.Y(n_10260)
);

INVx2_ASAP7_75t_L g10261 ( 
.A(n_8437),
.Y(n_10261)
);

INVx1_ASAP7_75t_L g10262 ( 
.A(n_8173),
.Y(n_10262)
);

INVx1_ASAP7_75t_L g10263 ( 
.A(n_8176),
.Y(n_10263)
);

BUFx8_ASAP7_75t_SL g10264 ( 
.A(n_8739),
.Y(n_10264)
);

INVx1_ASAP7_75t_L g10265 ( 
.A(n_8176),
.Y(n_10265)
);

NAND2x1p5_ASAP7_75t_L g10266 ( 
.A(n_8641),
.B(n_6651),
.Y(n_10266)
);

CKINVDCx20_ASAP7_75t_R g10267 ( 
.A(n_8481),
.Y(n_10267)
);

INVx2_ASAP7_75t_L g10268 ( 
.A(n_8437),
.Y(n_10268)
);

INVx1_ASAP7_75t_L g10269 ( 
.A(n_8178),
.Y(n_10269)
);

INVx1_ASAP7_75t_L g10270 ( 
.A(n_8178),
.Y(n_10270)
);

OA21x2_ASAP7_75t_L g10271 ( 
.A1(n_8478),
.A2(n_7087),
.B(n_7085),
.Y(n_10271)
);

INVx2_ASAP7_75t_L g10272 ( 
.A(n_8437),
.Y(n_10272)
);

OAI22xp33_ASAP7_75t_L g10273 ( 
.A1(n_7862),
.A2(n_7314),
.B1(n_7255),
.B2(n_6894),
.Y(n_10273)
);

INVx1_ASAP7_75t_L g10274 ( 
.A(n_8188),
.Y(n_10274)
);

OAI21x1_ASAP7_75t_L g10275 ( 
.A1(n_8577),
.A2(n_6885),
.B(n_6859),
.Y(n_10275)
);

HB1xp67_ASAP7_75t_L g10276 ( 
.A(n_8731),
.Y(n_10276)
);

OA21x2_ASAP7_75t_L g10277 ( 
.A1(n_8348),
.A2(n_7087),
.B(n_7085),
.Y(n_10277)
);

HB1xp67_ASAP7_75t_L g10278 ( 
.A(n_8785),
.Y(n_10278)
);

INVx2_ASAP7_75t_L g10279 ( 
.A(n_8446),
.Y(n_10279)
);

INVx2_ASAP7_75t_L g10280 ( 
.A(n_8446),
.Y(n_10280)
);

OR2x2_ASAP7_75t_L g10281 ( 
.A(n_7797),
.B(n_7253),
.Y(n_10281)
);

INVx2_ASAP7_75t_L g10282 ( 
.A(n_8446),
.Y(n_10282)
);

INVx2_ASAP7_75t_L g10283 ( 
.A(n_8456),
.Y(n_10283)
);

AND2x2_ASAP7_75t_L g10284 ( 
.A(n_8729),
.B(n_7526),
.Y(n_10284)
);

INVx2_ASAP7_75t_L g10285 ( 
.A(n_8456),
.Y(n_10285)
);

AO21x1_ASAP7_75t_SL g10286 ( 
.A1(n_8722),
.A2(n_6988),
.B(n_6982),
.Y(n_10286)
);

INVx1_ASAP7_75t_L g10287 ( 
.A(n_8188),
.Y(n_10287)
);

INVx3_ASAP7_75t_L g10288 ( 
.A(n_8168),
.Y(n_10288)
);

CKINVDCx6p67_ASAP7_75t_R g10289 ( 
.A(n_8542),
.Y(n_10289)
);

INVx2_ASAP7_75t_L g10290 ( 
.A(n_8456),
.Y(n_10290)
);

AND2x2_ASAP7_75t_L g10291 ( 
.A(n_8729),
.B(n_7526),
.Y(n_10291)
);

INVx2_ASAP7_75t_L g10292 ( 
.A(n_9821),
.Y(n_10292)
);

OAI21xp5_ASAP7_75t_L g10293 ( 
.A1(n_9321),
.A2(n_7821),
.B(n_8039),
.Y(n_10293)
);

HB1xp67_ASAP7_75t_L g10294 ( 
.A(n_9614),
.Y(n_10294)
);

INVx1_ASAP7_75t_L g10295 ( 
.A(n_8956),
.Y(n_10295)
);

INVx2_ASAP7_75t_L g10296 ( 
.A(n_9821),
.Y(n_10296)
);

INVx1_ASAP7_75t_L g10297 ( 
.A(n_8956),
.Y(n_10297)
);

INVx3_ASAP7_75t_L g10298 ( 
.A(n_9695),
.Y(n_10298)
);

AOI22xp33_ASAP7_75t_SL g10299 ( 
.A1(n_9495),
.A2(n_7724),
.B1(n_7739),
.B2(n_7738),
.Y(n_10299)
);

HB1xp67_ASAP7_75t_L g10300 ( 
.A(n_9614),
.Y(n_10300)
);

INVx1_ASAP7_75t_L g10301 ( 
.A(n_8958),
.Y(n_10301)
);

INVx5_ASAP7_75t_L g10302 ( 
.A(n_9109),
.Y(n_10302)
);

AND2x2_ASAP7_75t_L g10303 ( 
.A(n_8966),
.B(n_9572),
.Y(n_10303)
);

INVx2_ASAP7_75t_L g10304 ( 
.A(n_9821),
.Y(n_10304)
);

NAND2xp5_ASAP7_75t_L g10305 ( 
.A(n_10224),
.B(n_8083),
.Y(n_10305)
);

INVx2_ASAP7_75t_L g10306 ( 
.A(n_9827),
.Y(n_10306)
);

BUFx3_ASAP7_75t_L g10307 ( 
.A(n_9320),
.Y(n_10307)
);

OAI21x1_ASAP7_75t_L g10308 ( 
.A1(n_10242),
.A2(n_8584),
.B(n_8561),
.Y(n_10308)
);

AOI22xp33_ASAP7_75t_L g10309 ( 
.A1(n_9009),
.A2(n_8047),
.B1(n_8130),
.B2(n_7771),
.Y(n_10309)
);

INVx1_ASAP7_75t_L g10310 ( 
.A(n_8958),
.Y(n_10310)
);

NAND2xp5_ASAP7_75t_L g10311 ( 
.A(n_10224),
.B(n_8083),
.Y(n_10311)
);

INVx1_ASAP7_75t_L g10312 ( 
.A(n_8968),
.Y(n_10312)
);

INVx1_ASAP7_75t_L g10313 ( 
.A(n_8968),
.Y(n_10313)
);

INVx1_ASAP7_75t_L g10314 ( 
.A(n_8970),
.Y(n_10314)
);

AND2x2_ASAP7_75t_L g10315 ( 
.A(n_8966),
.B(n_7662),
.Y(n_10315)
);

INVx1_ASAP7_75t_L g10316 ( 
.A(n_8970),
.Y(n_10316)
);

BUFx2_ASAP7_75t_L g10317 ( 
.A(n_9109),
.Y(n_10317)
);

INVx2_ASAP7_75t_L g10318 ( 
.A(n_9827),
.Y(n_10318)
);

OAI21x1_ASAP7_75t_L g10319 ( 
.A1(n_10242),
.A2(n_8584),
.B(n_8561),
.Y(n_10319)
);

HB1xp67_ASAP7_75t_L g10320 ( 
.A(n_8972),
.Y(n_10320)
);

INVxp67_ASAP7_75t_L g10321 ( 
.A(n_9028),
.Y(n_10321)
);

INVx1_ASAP7_75t_L g10322 ( 
.A(n_8971),
.Y(n_10322)
);

NAND2xp5_ASAP7_75t_L g10323 ( 
.A(n_9321),
.B(n_8128),
.Y(n_10323)
);

AO21x1_ASAP7_75t_SL g10324 ( 
.A1(n_9399),
.A2(n_8695),
.B(n_8688),
.Y(n_10324)
);

AND2x2_ASAP7_75t_L g10325 ( 
.A(n_9572),
.B(n_7662),
.Y(n_10325)
);

INVx2_ASAP7_75t_L g10326 ( 
.A(n_9827),
.Y(n_10326)
);

INVx2_ASAP7_75t_SL g10327 ( 
.A(n_9196),
.Y(n_10327)
);

INVx3_ASAP7_75t_L g10328 ( 
.A(n_9695),
.Y(n_10328)
);

INVx1_ASAP7_75t_L g10329 ( 
.A(n_8971),
.Y(n_10329)
);

INVx2_ASAP7_75t_L g10330 ( 
.A(n_9830),
.Y(n_10330)
);

INVx1_ASAP7_75t_L g10331 ( 
.A(n_8976),
.Y(n_10331)
);

INVx1_ASAP7_75t_L g10332 ( 
.A(n_8976),
.Y(n_10332)
);

AND2x2_ASAP7_75t_L g10333 ( 
.A(n_9592),
.B(n_7662),
.Y(n_10333)
);

INVx3_ASAP7_75t_L g10334 ( 
.A(n_9695),
.Y(n_10334)
);

OAI21x1_ASAP7_75t_L g10335 ( 
.A1(n_9182),
.A2(n_8584),
.B(n_8561),
.Y(n_10335)
);

INVx1_ASAP7_75t_L g10336 ( 
.A(n_8978),
.Y(n_10336)
);

INVx1_ASAP7_75t_L g10337 ( 
.A(n_8978),
.Y(n_10337)
);

INVx1_ASAP7_75t_SL g10338 ( 
.A(n_9028),
.Y(n_10338)
);

INVx1_ASAP7_75t_L g10339 ( 
.A(n_8983),
.Y(n_10339)
);

OAI21x1_ASAP7_75t_L g10340 ( 
.A1(n_9182),
.A2(n_8784),
.B(n_8779),
.Y(n_10340)
);

INVx1_ASAP7_75t_L g10341 ( 
.A(n_8983),
.Y(n_10341)
);

INVx2_ASAP7_75t_L g10342 ( 
.A(n_9830),
.Y(n_10342)
);

AND2x2_ASAP7_75t_L g10343 ( 
.A(n_9592),
.B(n_9663),
.Y(n_10343)
);

INVx1_ASAP7_75t_L g10344 ( 
.A(n_8984),
.Y(n_10344)
);

INVx1_ASAP7_75t_L g10345 ( 
.A(n_8984),
.Y(n_10345)
);

OA21x2_ASAP7_75t_L g10346 ( 
.A1(n_9858),
.A2(n_8348),
.B(n_8503),
.Y(n_10346)
);

INVx1_ASAP7_75t_L g10347 ( 
.A(n_8985),
.Y(n_10347)
);

CKINVDCx5p33_ASAP7_75t_R g10348 ( 
.A(n_9035),
.Y(n_10348)
);

AND2x2_ASAP7_75t_L g10349 ( 
.A(n_9663),
.B(n_7666),
.Y(n_10349)
);

BUFx2_ASAP7_75t_L g10350 ( 
.A(n_9109),
.Y(n_10350)
);

BUFx6f_ASAP7_75t_L g10351 ( 
.A(n_9243),
.Y(n_10351)
);

AND2x4_ASAP7_75t_L g10352 ( 
.A(n_9127),
.B(n_7794),
.Y(n_10352)
);

INVx1_ASAP7_75t_L g10353 ( 
.A(n_8985),
.Y(n_10353)
);

INVx1_ASAP7_75t_L g10354 ( 
.A(n_8992),
.Y(n_10354)
);

CKINVDCx6p67_ASAP7_75t_R g10355 ( 
.A(n_9320),
.Y(n_10355)
);

INVx2_ASAP7_75t_SL g10356 ( 
.A(n_9196),
.Y(n_10356)
);

NAND2x1p5_ASAP7_75t_L g10357 ( 
.A(n_9695),
.B(n_8641),
.Y(n_10357)
);

INVx1_ASAP7_75t_L g10358 ( 
.A(n_8992),
.Y(n_10358)
);

NAND2xp5_ASAP7_75t_L g10359 ( 
.A(n_9181),
.B(n_8128),
.Y(n_10359)
);

BUFx6f_ASAP7_75t_L g10360 ( 
.A(n_9243),
.Y(n_10360)
);

INVx1_ASAP7_75t_L g10361 ( 
.A(n_8995),
.Y(n_10361)
);

BUFx2_ASAP7_75t_L g10362 ( 
.A(n_9243),
.Y(n_10362)
);

OAI21xp5_ASAP7_75t_L g10363 ( 
.A1(n_9495),
.A2(n_7749),
.B(n_8234),
.Y(n_10363)
);

OR2x6_ASAP7_75t_L g10364 ( 
.A(n_10123),
.B(n_8901),
.Y(n_10364)
);

OAI21xp5_ASAP7_75t_L g10365 ( 
.A1(n_9094),
.A2(n_7749),
.B(n_8234),
.Y(n_10365)
);

INVx1_ASAP7_75t_L g10366 ( 
.A(n_8995),
.Y(n_10366)
);

AND2x2_ASAP7_75t_L g10367 ( 
.A(n_9772),
.B(n_7666),
.Y(n_10367)
);

HB1xp67_ASAP7_75t_L g10368 ( 
.A(n_8991),
.Y(n_10368)
);

INVx2_ASAP7_75t_L g10369 ( 
.A(n_9830),
.Y(n_10369)
);

BUFx2_ASAP7_75t_L g10370 ( 
.A(n_9273),
.Y(n_10370)
);

AND2x4_ASAP7_75t_L g10371 ( 
.A(n_9127),
.B(n_7794),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_8999),
.Y(n_10372)
);

INVx1_ASAP7_75t_L g10373 ( 
.A(n_8999),
.Y(n_10373)
);

INVx2_ASAP7_75t_L g10374 ( 
.A(n_9832),
.Y(n_10374)
);

HB1xp67_ASAP7_75t_L g10375 ( 
.A(n_9014),
.Y(n_10375)
);

OR2x6_ASAP7_75t_L g10376 ( 
.A(n_10123),
.B(n_8271),
.Y(n_10376)
);

INVx2_ASAP7_75t_L g10377 ( 
.A(n_9832),
.Y(n_10377)
);

OR2x2_ASAP7_75t_L g10378 ( 
.A(n_8955),
.B(n_7839),
.Y(n_10378)
);

INVx1_ASAP7_75t_L g10379 ( 
.A(n_9000),
.Y(n_10379)
);

BUFx2_ASAP7_75t_L g10380 ( 
.A(n_9273),
.Y(n_10380)
);

AO21x2_ASAP7_75t_L g10381 ( 
.A1(n_9634),
.A2(n_7771),
.B(n_7739),
.Y(n_10381)
);

CKINVDCx11_ASAP7_75t_R g10382 ( 
.A(n_9320),
.Y(n_10382)
);

INVx1_ASAP7_75t_L g10383 ( 
.A(n_9000),
.Y(n_10383)
);

INVx1_ASAP7_75t_L g10384 ( 
.A(n_9001),
.Y(n_10384)
);

INVx2_ASAP7_75t_L g10385 ( 
.A(n_9832),
.Y(n_10385)
);

AO21x2_ASAP7_75t_L g10386 ( 
.A1(n_10068),
.A2(n_7771),
.B(n_7628),
.Y(n_10386)
);

INVx1_ASAP7_75t_L g10387 ( 
.A(n_9001),
.Y(n_10387)
);

BUFx3_ASAP7_75t_L g10388 ( 
.A(n_9404),
.Y(n_10388)
);

INVx1_ASAP7_75t_L g10389 ( 
.A(n_9002),
.Y(n_10389)
);

INVx1_ASAP7_75t_L g10390 ( 
.A(n_9002),
.Y(n_10390)
);

INVx2_ASAP7_75t_L g10391 ( 
.A(n_9841),
.Y(n_10391)
);

AOI21x1_ASAP7_75t_L g10392 ( 
.A1(n_9410),
.A2(n_8742),
.B(n_8737),
.Y(n_10392)
);

INVx2_ASAP7_75t_L g10393 ( 
.A(n_9841),
.Y(n_10393)
);

BUFx6f_ASAP7_75t_L g10394 ( 
.A(n_9273),
.Y(n_10394)
);

BUFx2_ASAP7_75t_L g10395 ( 
.A(n_9475),
.Y(n_10395)
);

OAI21xp5_ASAP7_75t_L g10396 ( 
.A1(n_9668),
.A2(n_8044),
.B(n_7675),
.Y(n_10396)
);

AOI22xp5_ASAP7_75t_L g10397 ( 
.A1(n_9858),
.A2(n_8282),
.B1(n_8277),
.B2(n_8275),
.Y(n_10397)
);

INVx3_ASAP7_75t_L g10398 ( 
.A(n_9695),
.Y(n_10398)
);

AND2x4_ASAP7_75t_L g10399 ( 
.A(n_9365),
.B(n_7794),
.Y(n_10399)
);

INVx2_ASAP7_75t_L g10400 ( 
.A(n_9841),
.Y(n_10400)
);

OAI21x1_ASAP7_75t_L g10401 ( 
.A1(n_9182),
.A2(n_8784),
.B(n_8779),
.Y(n_10401)
);

HB1xp67_ASAP7_75t_L g10402 ( 
.A(n_9024),
.Y(n_10402)
);

BUFx2_ASAP7_75t_L g10403 ( 
.A(n_9475),
.Y(n_10403)
);

INVx1_ASAP7_75t_SL g10404 ( 
.A(n_9103),
.Y(n_10404)
);

INVx2_ASAP7_75t_L g10405 ( 
.A(n_9843),
.Y(n_10405)
);

AND2x4_ASAP7_75t_L g10406 ( 
.A(n_9365),
.B(n_7794),
.Y(n_10406)
);

AND2x4_ASAP7_75t_SL g10407 ( 
.A(n_9467),
.B(n_8271),
.Y(n_10407)
);

INVx1_ASAP7_75t_L g10408 ( 
.A(n_9012),
.Y(n_10408)
);

INVx1_ASAP7_75t_L g10409 ( 
.A(n_9012),
.Y(n_10409)
);

INVx3_ASAP7_75t_L g10410 ( 
.A(n_9695),
.Y(n_10410)
);

INVx2_ASAP7_75t_L g10411 ( 
.A(n_9843),
.Y(n_10411)
);

INVx2_ASAP7_75t_L g10412 ( 
.A(n_9843),
.Y(n_10412)
);

INVx1_ASAP7_75t_L g10413 ( 
.A(n_9017),
.Y(n_10413)
);

INVxp33_ASAP7_75t_SL g10414 ( 
.A(n_10125),
.Y(n_10414)
);

AND2x2_ASAP7_75t_L g10415 ( 
.A(n_9772),
.B(n_7666),
.Y(n_10415)
);

INVx1_ASAP7_75t_L g10416 ( 
.A(n_9017),
.Y(n_10416)
);

NAND2xp5_ASAP7_75t_L g10417 ( 
.A(n_9202),
.B(n_9436),
.Y(n_10417)
);

INVx1_ASAP7_75t_L g10418 ( 
.A(n_9020),
.Y(n_10418)
);

AOI21xp5_ASAP7_75t_L g10419 ( 
.A1(n_9224),
.A2(n_7879),
.B(n_8275),
.Y(n_10419)
);

HB1xp67_ASAP7_75t_L g10420 ( 
.A(n_9039),
.Y(n_10420)
);

INVx2_ASAP7_75t_L g10421 ( 
.A(n_9844),
.Y(n_10421)
);

AOI21x1_ASAP7_75t_L g10422 ( 
.A1(n_9410),
.A2(n_9652),
.B(n_10068),
.Y(n_10422)
);

INVx2_ASAP7_75t_L g10423 ( 
.A(n_9844),
.Y(n_10423)
);

INVx1_ASAP7_75t_L g10424 ( 
.A(n_9020),
.Y(n_10424)
);

INVx1_ASAP7_75t_SL g10425 ( 
.A(n_9103),
.Y(n_10425)
);

BUFx10_ASAP7_75t_L g10426 ( 
.A(n_8954),
.Y(n_10426)
);

BUFx6f_ASAP7_75t_L g10427 ( 
.A(n_8954),
.Y(n_10427)
);

BUFx2_ASAP7_75t_SL g10428 ( 
.A(n_10098),
.Y(n_10428)
);

HB1xp67_ASAP7_75t_L g10429 ( 
.A(n_9050),
.Y(n_10429)
);

AND2x2_ASAP7_75t_L g10430 ( 
.A(n_8960),
.B(n_9007),
.Y(n_10430)
);

INVx2_ASAP7_75t_SL g10431 ( 
.A(n_9196),
.Y(n_10431)
);

INVx2_ASAP7_75t_SL g10432 ( 
.A(n_9196),
.Y(n_10432)
);

INVx2_ASAP7_75t_L g10433 ( 
.A(n_9844),
.Y(n_10433)
);

OR2x2_ASAP7_75t_L g10434 ( 
.A(n_8955),
.B(n_7839),
.Y(n_10434)
);

HB1xp67_ASAP7_75t_L g10435 ( 
.A(n_9110),
.Y(n_10435)
);

AND2x2_ASAP7_75t_L g10436 ( 
.A(n_8960),
.B(n_7706),
.Y(n_10436)
);

AND2x2_ASAP7_75t_L g10437 ( 
.A(n_9007),
.B(n_7706),
.Y(n_10437)
);

INVx1_ASAP7_75t_L g10438 ( 
.A(n_9022),
.Y(n_10438)
);

INVx1_ASAP7_75t_L g10439 ( 
.A(n_9022),
.Y(n_10439)
);

INVx2_ASAP7_75t_L g10440 ( 
.A(n_9846),
.Y(n_10440)
);

AOI22xp33_ASAP7_75t_L g10441 ( 
.A1(n_9009),
.A2(n_8047),
.B1(n_8220),
.B2(n_7748),
.Y(n_10441)
);

INVx1_ASAP7_75t_L g10442 ( 
.A(n_9025),
.Y(n_10442)
);

INVx2_ASAP7_75t_L g10443 ( 
.A(n_9846),
.Y(n_10443)
);

OAI21x1_ASAP7_75t_SL g10444 ( 
.A1(n_10225),
.A2(n_7756),
.B(n_8271),
.Y(n_10444)
);

INVx1_ASAP7_75t_L g10445 ( 
.A(n_9025),
.Y(n_10445)
);

INVx3_ASAP7_75t_L g10446 ( 
.A(n_9695),
.Y(n_10446)
);

BUFx2_ASAP7_75t_L g10447 ( 
.A(n_9475),
.Y(n_10447)
);

INVxp67_ASAP7_75t_L g10448 ( 
.A(n_9105),
.Y(n_10448)
);

INVx2_ASAP7_75t_L g10449 ( 
.A(n_9846),
.Y(n_10449)
);

INVx1_ASAP7_75t_L g10450 ( 
.A(n_9027),
.Y(n_10450)
);

AND2x2_ASAP7_75t_L g10451 ( 
.A(n_9038),
.B(n_7706),
.Y(n_10451)
);

HB1xp67_ASAP7_75t_L g10452 ( 
.A(n_9118),
.Y(n_10452)
);

HB1xp67_ASAP7_75t_L g10453 ( 
.A(n_9131),
.Y(n_10453)
);

INVx1_ASAP7_75t_L g10454 ( 
.A(n_9027),
.Y(n_10454)
);

INVx1_ASAP7_75t_L g10455 ( 
.A(n_9031),
.Y(n_10455)
);

INVx1_ASAP7_75t_L g10456 ( 
.A(n_9031),
.Y(n_10456)
);

INVx1_ASAP7_75t_L g10457 ( 
.A(n_9036),
.Y(n_10457)
);

NOR2x1_ASAP7_75t_R g10458 ( 
.A(n_9404),
.B(n_8271),
.Y(n_10458)
);

INVx1_ASAP7_75t_L g10459 ( 
.A(n_9036),
.Y(n_10459)
);

OAI21x1_ASAP7_75t_L g10460 ( 
.A1(n_9777),
.A2(n_8784),
.B(n_8779),
.Y(n_10460)
);

INVx2_ASAP7_75t_L g10461 ( 
.A(n_9847),
.Y(n_10461)
);

HB1xp67_ASAP7_75t_L g10462 ( 
.A(n_9147),
.Y(n_10462)
);

NOR2x1_ASAP7_75t_SL g10463 ( 
.A(n_9070),
.B(n_7746),
.Y(n_10463)
);

HB1xp67_ASAP7_75t_L g10464 ( 
.A(n_9164),
.Y(n_10464)
);

INVx1_ASAP7_75t_L g10465 ( 
.A(n_9041),
.Y(n_10465)
);

INVx1_ASAP7_75t_L g10466 ( 
.A(n_9041),
.Y(n_10466)
);

INVx1_ASAP7_75t_L g10467 ( 
.A(n_9043),
.Y(n_10467)
);

AOI211xp5_ASAP7_75t_L g10468 ( 
.A1(n_9286),
.A2(n_7607),
.B(n_8220),
.C(n_7879),
.Y(n_10468)
);

AND2x2_ASAP7_75t_L g10469 ( 
.A(n_9038),
.B(n_7734),
.Y(n_10469)
);

INVx1_ASAP7_75t_L g10470 ( 
.A(n_9043),
.Y(n_10470)
);

INVx1_ASAP7_75t_L g10471 ( 
.A(n_9045),
.Y(n_10471)
);

INVx1_ASAP7_75t_L g10472 ( 
.A(n_9045),
.Y(n_10472)
);

INVx1_ASAP7_75t_L g10473 ( 
.A(n_9048),
.Y(n_10473)
);

NOR2xp33_ASAP7_75t_L g10474 ( 
.A(n_9489),
.B(n_8505),
.Y(n_10474)
);

AOI22xp33_ASAP7_75t_L g10475 ( 
.A1(n_9560),
.A2(n_7809),
.B1(n_8163),
.B2(n_7750),
.Y(n_10475)
);

INVx1_ASAP7_75t_L g10476 ( 
.A(n_9048),
.Y(n_10476)
);

BUFx2_ASAP7_75t_L g10477 ( 
.A(n_9475),
.Y(n_10477)
);

AOI21x1_ASAP7_75t_L g10478 ( 
.A1(n_9652),
.A2(n_9593),
.B(n_9494),
.Y(n_10478)
);

INVx2_ASAP7_75t_L g10479 ( 
.A(n_9847),
.Y(n_10479)
);

INVx1_ASAP7_75t_L g10480 ( 
.A(n_9052),
.Y(n_10480)
);

BUFx12f_ASAP7_75t_L g10481 ( 
.A(n_9404),
.Y(n_10481)
);

INVx1_ASAP7_75t_L g10482 ( 
.A(n_9052),
.Y(n_10482)
);

AND2x4_ASAP7_75t_L g10483 ( 
.A(n_9469),
.B(n_7794),
.Y(n_10483)
);

INVx1_ASAP7_75t_L g10484 ( 
.A(n_9056),
.Y(n_10484)
);

AO22x1_ASAP7_75t_L g10485 ( 
.A1(n_9032),
.A2(n_8867),
.B1(n_8448),
.B2(n_8379),
.Y(n_10485)
);

INVx1_ASAP7_75t_L g10486 ( 
.A(n_9056),
.Y(n_10486)
);

AND2x4_ASAP7_75t_L g10487 ( 
.A(n_9469),
.B(n_8490),
.Y(n_10487)
);

BUFx2_ASAP7_75t_L g10488 ( 
.A(n_9737),
.Y(n_10488)
);

INVx1_ASAP7_75t_L g10489 ( 
.A(n_9057),
.Y(n_10489)
);

INVxp67_ASAP7_75t_L g10490 ( 
.A(n_9105),
.Y(n_10490)
);

INVx2_ASAP7_75t_L g10491 ( 
.A(n_9847),
.Y(n_10491)
);

INVx2_ASAP7_75t_L g10492 ( 
.A(n_9851),
.Y(n_10492)
);

INVx2_ASAP7_75t_L g10493 ( 
.A(n_9851),
.Y(n_10493)
);

INVx1_ASAP7_75t_L g10494 ( 
.A(n_9057),
.Y(n_10494)
);

INVx1_ASAP7_75t_L g10495 ( 
.A(n_9058),
.Y(n_10495)
);

INVx1_ASAP7_75t_L g10496 ( 
.A(n_9058),
.Y(n_10496)
);

INVx1_ASAP7_75t_L g10497 ( 
.A(n_9061),
.Y(n_10497)
);

INVx1_ASAP7_75t_L g10498 ( 
.A(n_9061),
.Y(n_10498)
);

AOI22xp33_ASAP7_75t_SL g10499 ( 
.A1(n_9394),
.A2(n_7724),
.B1(n_7842),
.B2(n_7829),
.Y(n_10499)
);

INVx2_ASAP7_75t_L g10500 ( 
.A(n_9851),
.Y(n_10500)
);

HB1xp67_ASAP7_75t_L g10501 ( 
.A(n_9166),
.Y(n_10501)
);

INVx1_ASAP7_75t_L g10502 ( 
.A(n_9069),
.Y(n_10502)
);

OR2x2_ASAP7_75t_L g10503 ( 
.A(n_9667),
.B(n_7684),
.Y(n_10503)
);

INVx2_ASAP7_75t_L g10504 ( 
.A(n_9854),
.Y(n_10504)
);

OA21x2_ASAP7_75t_L g10505 ( 
.A1(n_10225),
.A2(n_8348),
.B(n_8503),
.Y(n_10505)
);

INVx2_ASAP7_75t_L g10506 ( 
.A(n_9854),
.Y(n_10506)
);

NAND2x1p5_ASAP7_75t_L g10507 ( 
.A(n_10170),
.B(n_8641),
.Y(n_10507)
);

INVx2_ASAP7_75t_L g10508 ( 
.A(n_9854),
.Y(n_10508)
);

INVx1_ASAP7_75t_L g10509 ( 
.A(n_9069),
.Y(n_10509)
);

INVx1_ASAP7_75t_L g10510 ( 
.A(n_9075),
.Y(n_10510)
);

AND2x6_ASAP7_75t_L g10511 ( 
.A(n_8954),
.B(n_8357),
.Y(n_10511)
);

INVx1_ASAP7_75t_L g10512 ( 
.A(n_9075),
.Y(n_10512)
);

INVx1_ASAP7_75t_L g10513 ( 
.A(n_9080),
.Y(n_10513)
);

BUFx2_ASAP7_75t_L g10514 ( 
.A(n_9737),
.Y(n_10514)
);

INVx2_ASAP7_75t_L g10515 ( 
.A(n_9857),
.Y(n_10515)
);

INVx2_ASAP7_75t_L g10516 ( 
.A(n_9857),
.Y(n_10516)
);

INVx1_ASAP7_75t_L g10517 ( 
.A(n_9080),
.Y(n_10517)
);

INVx1_ASAP7_75t_L g10518 ( 
.A(n_9082),
.Y(n_10518)
);

NAND2xp5_ASAP7_75t_L g10519 ( 
.A(n_9453),
.B(n_8772),
.Y(n_10519)
);

CKINVDCx5p33_ASAP7_75t_R g10520 ( 
.A(n_10070),
.Y(n_10520)
);

INVx1_ASAP7_75t_L g10521 ( 
.A(n_9082),
.Y(n_10521)
);

AOI21x1_ASAP7_75t_L g10522 ( 
.A1(n_9494),
.A2(n_9643),
.B(n_9593),
.Y(n_10522)
);

AO21x2_ASAP7_75t_L g10523 ( 
.A1(n_9883),
.A2(n_7628),
.B(n_8752),
.Y(n_10523)
);

INVx2_ASAP7_75t_SL g10524 ( 
.A(n_9497),
.Y(n_10524)
);

CKINVDCx6p67_ASAP7_75t_R g10525 ( 
.A(n_9599),
.Y(n_10525)
);

AOI22xp5_ASAP7_75t_L g10526 ( 
.A1(n_9394),
.A2(n_8282),
.B1(n_8277),
.B2(n_8364),
.Y(n_10526)
);

INVx1_ASAP7_75t_L g10527 ( 
.A(n_9083),
.Y(n_10527)
);

BUFx2_ASAP7_75t_L g10528 ( 
.A(n_9737),
.Y(n_10528)
);

NAND2xp33_ASAP7_75t_R g10529 ( 
.A(n_9070),
.B(n_8281),
.Y(n_10529)
);

HB1xp67_ASAP7_75t_L g10530 ( 
.A(n_9172),
.Y(n_10530)
);

BUFx3_ASAP7_75t_L g10531 ( 
.A(n_9599),
.Y(n_10531)
);

INVx2_ASAP7_75t_L g10532 ( 
.A(n_9857),
.Y(n_10532)
);

OAI22xp5_ASAP7_75t_L g10533 ( 
.A1(n_9769),
.A2(n_8324),
.B1(n_8314),
.B2(n_7675),
.Y(n_10533)
);

INVx1_ASAP7_75t_L g10534 ( 
.A(n_9083),
.Y(n_10534)
);

BUFx6f_ASAP7_75t_L g10535 ( 
.A(n_8954),
.Y(n_10535)
);

BUFx3_ASAP7_75t_L g10536 ( 
.A(n_9599),
.Y(n_10536)
);

INVx1_ASAP7_75t_SL g10537 ( 
.A(n_9191),
.Y(n_10537)
);

INVx1_ASAP7_75t_SL g10538 ( 
.A(n_9191),
.Y(n_10538)
);

AO22x1_ASAP7_75t_L g10539 ( 
.A1(n_9032),
.A2(n_8867),
.B1(n_8379),
.B2(n_8452),
.Y(n_10539)
);

AND2x2_ASAP7_75t_L g10540 ( 
.A(n_9148),
.B(n_7734),
.Y(n_10540)
);

AND2x2_ASAP7_75t_L g10541 ( 
.A(n_9148),
.B(n_7734),
.Y(n_10541)
);

INVx1_ASAP7_75t_L g10542 ( 
.A(n_9088),
.Y(n_10542)
);

BUFx3_ASAP7_75t_L g10543 ( 
.A(n_9609),
.Y(n_10543)
);

INVx3_ASAP7_75t_L g10544 ( 
.A(n_10170),
.Y(n_10544)
);

OAI21x1_ASAP7_75t_L g10545 ( 
.A1(n_9777),
.A2(n_8804),
.B(n_8803),
.Y(n_10545)
);

INVx1_ASAP7_75t_L g10546 ( 
.A(n_9088),
.Y(n_10546)
);

HB1xp67_ASAP7_75t_L g10547 ( 
.A(n_9198),
.Y(n_10547)
);

BUFx6f_ASAP7_75t_L g10548 ( 
.A(n_8954),
.Y(n_10548)
);

HB1xp67_ASAP7_75t_L g10549 ( 
.A(n_9260),
.Y(n_10549)
);

HB1xp67_ASAP7_75t_L g10550 ( 
.A(n_9281),
.Y(n_10550)
);

BUFx3_ASAP7_75t_L g10551 ( 
.A(n_9609),
.Y(n_10551)
);

AND2x2_ASAP7_75t_L g10552 ( 
.A(n_9159),
.B(n_7711),
.Y(n_10552)
);

INVx1_ASAP7_75t_L g10553 ( 
.A(n_9091),
.Y(n_10553)
);

AOI22xp33_ASAP7_75t_SL g10554 ( 
.A1(n_9242),
.A2(n_7724),
.B1(n_7842),
.B2(n_7829),
.Y(n_10554)
);

HB1xp67_ASAP7_75t_L g10555 ( 
.A(n_9293),
.Y(n_10555)
);

HB1xp67_ASAP7_75t_L g10556 ( 
.A(n_9327),
.Y(n_10556)
);

INVx2_ASAP7_75t_L g10557 ( 
.A(n_9859),
.Y(n_10557)
);

BUFx2_ASAP7_75t_L g10558 ( 
.A(n_9737),
.Y(n_10558)
);

INVx1_ASAP7_75t_L g10559 ( 
.A(n_9091),
.Y(n_10559)
);

BUFx6f_ASAP7_75t_L g10560 ( 
.A(n_8954),
.Y(n_10560)
);

BUFx3_ASAP7_75t_L g10561 ( 
.A(n_9609),
.Y(n_10561)
);

INVx1_ASAP7_75t_L g10562 ( 
.A(n_9092),
.Y(n_10562)
);

INVx2_ASAP7_75t_L g10563 ( 
.A(n_9859),
.Y(n_10563)
);

OAI21x1_ASAP7_75t_L g10564 ( 
.A1(n_9777),
.A2(n_8804),
.B(n_8803),
.Y(n_10564)
);

AND2x2_ASAP7_75t_L g10565 ( 
.A(n_9159),
.B(n_7711),
.Y(n_10565)
);

BUFx3_ASAP7_75t_L g10566 ( 
.A(n_9919),
.Y(n_10566)
);

AO31x2_ASAP7_75t_L g10567 ( 
.A1(n_10253),
.A2(n_7628),
.A3(n_8663),
.B(n_7802),
.Y(n_10567)
);

INVx2_ASAP7_75t_L g10568 ( 
.A(n_9859),
.Y(n_10568)
);

INVx1_ASAP7_75t_L g10569 ( 
.A(n_9092),
.Y(n_10569)
);

OAI21x1_ASAP7_75t_L g10570 ( 
.A1(n_9634),
.A2(n_8804),
.B(n_8803),
.Y(n_10570)
);

BUFx6f_ASAP7_75t_L g10571 ( 
.A(n_9013),
.Y(n_10571)
);

BUFx3_ASAP7_75t_L g10572 ( 
.A(n_9919),
.Y(n_10572)
);

BUFx3_ASAP7_75t_L g10573 ( 
.A(n_9919),
.Y(n_10573)
);

INVx1_ASAP7_75t_L g10574 ( 
.A(n_9095),
.Y(n_10574)
);

BUFx6f_ASAP7_75t_L g10575 ( 
.A(n_9013),
.Y(n_10575)
);

AOI21x1_ASAP7_75t_L g10576 ( 
.A1(n_9643),
.A2(n_8742),
.B(n_8737),
.Y(n_10576)
);

AND2x2_ASAP7_75t_L g10577 ( 
.A(n_9161),
.B(n_7711),
.Y(n_10577)
);

AOI21x1_ASAP7_75t_L g10578 ( 
.A1(n_9718),
.A2(n_8742),
.B(n_8737),
.Y(n_10578)
);

INVx2_ASAP7_75t_L g10579 ( 
.A(n_9867),
.Y(n_10579)
);

HB1xp67_ASAP7_75t_L g10580 ( 
.A(n_10087),
.Y(n_10580)
);

NAND2xp5_ASAP7_75t_L g10581 ( 
.A(n_9583),
.B(n_8772),
.Y(n_10581)
);

INVx1_ASAP7_75t_L g10582 ( 
.A(n_9095),
.Y(n_10582)
);

HB1xp67_ASAP7_75t_L g10583 ( 
.A(n_10087),
.Y(n_10583)
);

INVx1_ASAP7_75t_L g10584 ( 
.A(n_9099),
.Y(n_10584)
);

AND2x2_ASAP7_75t_L g10585 ( 
.A(n_9161),
.B(n_7711),
.Y(n_10585)
);

INVx1_ASAP7_75t_L g10586 ( 
.A(n_9099),
.Y(n_10586)
);

OR2x2_ASAP7_75t_L g10587 ( 
.A(n_9667),
.B(n_10247),
.Y(n_10587)
);

INVx2_ASAP7_75t_L g10588 ( 
.A(n_9867),
.Y(n_10588)
);

AND2x2_ASAP7_75t_L g10589 ( 
.A(n_9184),
.B(n_7711),
.Y(n_10589)
);

INVx1_ASAP7_75t_L g10590 ( 
.A(n_9101),
.Y(n_10590)
);

INVx2_ASAP7_75t_L g10591 ( 
.A(n_9867),
.Y(n_10591)
);

INVx1_ASAP7_75t_L g10592 ( 
.A(n_9101),
.Y(n_10592)
);

OR2x6_ASAP7_75t_L g10593 ( 
.A(n_9070),
.B(n_8271),
.Y(n_10593)
);

INVx1_ASAP7_75t_L g10594 ( 
.A(n_9102),
.Y(n_10594)
);

OAI21x1_ASAP7_75t_L g10595 ( 
.A1(n_9758),
.A2(n_8810),
.B(n_8503),
.Y(n_10595)
);

INVx2_ASAP7_75t_L g10596 ( 
.A(n_9868),
.Y(n_10596)
);

INVx1_ASAP7_75t_L g10597 ( 
.A(n_9102),
.Y(n_10597)
);

INVx1_ASAP7_75t_L g10598 ( 
.A(n_9107),
.Y(n_10598)
);

OA21x2_ASAP7_75t_L g10599 ( 
.A1(n_9119),
.A2(n_8447),
.B(n_8442),
.Y(n_10599)
);

INVx2_ASAP7_75t_L g10600 ( 
.A(n_9868),
.Y(n_10600)
);

HB1xp67_ASAP7_75t_L g10601 ( 
.A(n_9344),
.Y(n_10601)
);

BUFx3_ASAP7_75t_L g10602 ( 
.A(n_9935),
.Y(n_10602)
);

OR2x2_ASAP7_75t_L g10603 ( 
.A(n_10247),
.B(n_7684),
.Y(n_10603)
);

INVx1_ASAP7_75t_L g10604 ( 
.A(n_9107),
.Y(n_10604)
);

INVx3_ASAP7_75t_L g10605 ( 
.A(n_10170),
.Y(n_10605)
);

INVx1_ASAP7_75t_L g10606 ( 
.A(n_9108),
.Y(n_10606)
);

INVx1_ASAP7_75t_L g10607 ( 
.A(n_9108),
.Y(n_10607)
);

HB1xp67_ASAP7_75t_L g10608 ( 
.A(n_9354),
.Y(n_10608)
);

OAI21x1_ASAP7_75t_L g10609 ( 
.A1(n_9758),
.A2(n_8810),
.B(n_8522),
.Y(n_10609)
);

BUFx2_ASAP7_75t_L g10610 ( 
.A(n_10058),
.Y(n_10610)
);

AO21x2_ASAP7_75t_L g10611 ( 
.A1(n_9883),
.A2(n_8752),
.B(n_7605),
.Y(n_10611)
);

INVx1_ASAP7_75t_L g10612 ( 
.A(n_9116),
.Y(n_10612)
);

OAI21xp5_ASAP7_75t_L g10613 ( 
.A1(n_8988),
.A2(n_8044),
.B(n_7862),
.Y(n_10613)
);

INVx1_ASAP7_75t_L g10614 ( 
.A(n_9116),
.Y(n_10614)
);

INVx2_ASAP7_75t_L g10615 ( 
.A(n_9868),
.Y(n_10615)
);

OAI21x1_ASAP7_75t_L g10616 ( 
.A1(n_10199),
.A2(n_8810),
.B(n_8522),
.Y(n_10616)
);

HB1xp67_ASAP7_75t_L g10617 ( 
.A(n_9389),
.Y(n_10617)
);

INVx1_ASAP7_75t_L g10618 ( 
.A(n_9117),
.Y(n_10618)
);

OAI21x1_ASAP7_75t_L g10619 ( 
.A1(n_10199),
.A2(n_8522),
.B(n_8447),
.Y(n_10619)
);

AND2x4_ASAP7_75t_L g10620 ( 
.A(n_10213),
.B(n_8490),
.Y(n_10620)
);

INVx1_ASAP7_75t_L g10621 ( 
.A(n_9117),
.Y(n_10621)
);

AO31x2_ASAP7_75t_L g10622 ( 
.A1(n_10253),
.A2(n_8663),
.A3(n_7802),
.B(n_8476),
.Y(n_10622)
);

OR2x6_ASAP7_75t_L g10623 ( 
.A(n_9070),
.B(n_8379),
.Y(n_10623)
);

INVx1_ASAP7_75t_L g10624 ( 
.A(n_9125),
.Y(n_10624)
);

INVx2_ASAP7_75t_L g10625 ( 
.A(n_9877),
.Y(n_10625)
);

BUFx2_ASAP7_75t_L g10626 ( 
.A(n_10058),
.Y(n_10626)
);

BUFx2_ASAP7_75t_L g10627 ( 
.A(n_10058),
.Y(n_10627)
);

AOI22xp33_ASAP7_75t_SL g10628 ( 
.A1(n_9242),
.A2(n_7724),
.B1(n_7842),
.B2(n_7829),
.Y(n_10628)
);

INVx1_ASAP7_75t_L g10629 ( 
.A(n_9125),
.Y(n_10629)
);

HB1xp67_ASAP7_75t_L g10630 ( 
.A(n_9400),
.Y(n_10630)
);

BUFx2_ASAP7_75t_L g10631 ( 
.A(n_10058),
.Y(n_10631)
);

INVx2_ASAP7_75t_SL g10632 ( 
.A(n_9497),
.Y(n_10632)
);

BUFx3_ASAP7_75t_L g10633 ( 
.A(n_9935),
.Y(n_10633)
);

AO21x2_ASAP7_75t_L g10634 ( 
.A1(n_9319),
.A2(n_9353),
.B(n_10273),
.Y(n_10634)
);

INVx2_ASAP7_75t_L g10635 ( 
.A(n_9877),
.Y(n_10635)
);

NAND2x1_ASAP7_75t_L g10636 ( 
.A(n_9557),
.B(n_7605),
.Y(n_10636)
);

HB1xp67_ASAP7_75t_L g10637 ( 
.A(n_9460),
.Y(n_10637)
);

NAND2xp5_ASAP7_75t_L g10638 ( 
.A(n_9583),
.B(n_8776),
.Y(n_10638)
);

INVx3_ASAP7_75t_L g10639 ( 
.A(n_10170),
.Y(n_10639)
);

INVx2_ASAP7_75t_L g10640 ( 
.A(n_9877),
.Y(n_10640)
);

INVx1_ASAP7_75t_L g10641 ( 
.A(n_9137),
.Y(n_10641)
);

INVx2_ASAP7_75t_L g10642 ( 
.A(n_9878),
.Y(n_10642)
);

INVx2_ASAP7_75t_L g10643 ( 
.A(n_9878),
.Y(n_10643)
);

AND2x2_ASAP7_75t_L g10644 ( 
.A(n_9184),
.B(n_7744),
.Y(n_10644)
);

BUFx6f_ASAP7_75t_L g10645 ( 
.A(n_9013),
.Y(n_10645)
);

NAND3xp33_ASAP7_75t_L g10646 ( 
.A(n_10246),
.B(n_7809),
.C(n_7970),
.Y(n_10646)
);

OA21x2_ASAP7_75t_L g10647 ( 
.A1(n_9119),
.A2(n_8447),
.B(n_8442),
.Y(n_10647)
);

NAND2xp5_ASAP7_75t_SL g10648 ( 
.A(n_9326),
.B(n_7756),
.Y(n_10648)
);

INVx2_ASAP7_75t_L g10649 ( 
.A(n_9878),
.Y(n_10649)
);

INVx4_ASAP7_75t_SL g10650 ( 
.A(n_8959),
.Y(n_10650)
);

INVx2_ASAP7_75t_L g10651 ( 
.A(n_9882),
.Y(n_10651)
);

INVx1_ASAP7_75t_L g10652 ( 
.A(n_9137),
.Y(n_10652)
);

OA21x2_ASAP7_75t_L g10653 ( 
.A1(n_9119),
.A2(n_8442),
.B(n_8342),
.Y(n_10653)
);

INVx2_ASAP7_75t_L g10654 ( 
.A(n_9882),
.Y(n_10654)
);

INVx1_ASAP7_75t_L g10655 ( 
.A(n_9138),
.Y(n_10655)
);

INVx1_ASAP7_75t_L g10656 ( 
.A(n_9138),
.Y(n_10656)
);

INVx1_ASAP7_75t_L g10657 ( 
.A(n_9141),
.Y(n_10657)
);

AND2x4_ASAP7_75t_L g10658 ( 
.A(n_10213),
.B(n_8490),
.Y(n_10658)
);

OR2x6_ASAP7_75t_L g10659 ( 
.A(n_9070),
.B(n_8379),
.Y(n_10659)
);

BUFx6f_ASAP7_75t_L g10660 ( 
.A(n_9013),
.Y(n_10660)
);

INVx1_ASAP7_75t_L g10661 ( 
.A(n_9141),
.Y(n_10661)
);

INVx2_ASAP7_75t_L g10662 ( 
.A(n_9882),
.Y(n_10662)
);

OR2x2_ASAP7_75t_L g10663 ( 
.A(n_10281),
.B(n_8904),
.Y(n_10663)
);

INVx2_ASAP7_75t_SL g10664 ( 
.A(n_9497),
.Y(n_10664)
);

INVx1_ASAP7_75t_L g10665 ( 
.A(n_9149),
.Y(n_10665)
);

INVx1_ASAP7_75t_L g10666 ( 
.A(n_9149),
.Y(n_10666)
);

INVx2_ASAP7_75t_L g10667 ( 
.A(n_9884),
.Y(n_10667)
);

OA21x2_ASAP7_75t_L g10668 ( 
.A1(n_9759),
.A2(n_8342),
.B(n_8848),
.Y(n_10668)
);

INVx1_ASAP7_75t_L g10669 ( 
.A(n_9157),
.Y(n_10669)
);

AND2x4_ASAP7_75t_L g10670 ( 
.A(n_10213),
.B(n_8490),
.Y(n_10670)
);

INVx1_ASAP7_75t_L g10671 ( 
.A(n_9157),
.Y(n_10671)
);

OAI21x1_ASAP7_75t_L g10672 ( 
.A1(n_9852),
.A2(n_8894),
.B(n_8814),
.Y(n_10672)
);

INVx1_ASAP7_75t_L g10673 ( 
.A(n_9160),
.Y(n_10673)
);

OR2x6_ASAP7_75t_L g10674 ( 
.A(n_9065),
.B(n_8379),
.Y(n_10674)
);

AND2x2_ASAP7_75t_L g10675 ( 
.A(n_9351),
.B(n_9466),
.Y(n_10675)
);

HB1xp67_ASAP7_75t_L g10676 ( 
.A(n_9482),
.Y(n_10676)
);

INVxp33_ASAP7_75t_L g10677 ( 
.A(n_9485),
.Y(n_10677)
);

INVx2_ASAP7_75t_L g10678 ( 
.A(n_9884),
.Y(n_10678)
);

INVx1_ASAP7_75t_L g10679 ( 
.A(n_9160),
.Y(n_10679)
);

HB1xp67_ASAP7_75t_L g10680 ( 
.A(n_9484),
.Y(n_10680)
);

INVx3_ASAP7_75t_L g10681 ( 
.A(n_10170),
.Y(n_10681)
);

INVx2_ASAP7_75t_L g10682 ( 
.A(n_9884),
.Y(n_10682)
);

INVxp67_ASAP7_75t_L g10683 ( 
.A(n_9567),
.Y(n_10683)
);

NAND2x1p5_ASAP7_75t_L g10684 ( 
.A(n_10170),
.B(n_8641),
.Y(n_10684)
);

BUFx3_ASAP7_75t_L g10685 ( 
.A(n_9935),
.Y(n_10685)
);

AOI22xp33_ASAP7_75t_L g10686 ( 
.A1(n_9059),
.A2(n_7750),
.B1(n_8197),
.B2(n_7832),
.Y(n_10686)
);

INVx1_ASAP7_75t_L g10687 ( 
.A(n_9162),
.Y(n_10687)
);

AOI22xp33_ASAP7_75t_SL g10688 ( 
.A1(n_10174),
.A2(n_7724),
.B1(n_7842),
.B2(n_7750),
.Y(n_10688)
);

INVx1_ASAP7_75t_L g10689 ( 
.A(n_9162),
.Y(n_10689)
);

INVx1_ASAP7_75t_L g10690 ( 
.A(n_9169),
.Y(n_10690)
);

INVx1_ASAP7_75t_L g10691 ( 
.A(n_9169),
.Y(n_10691)
);

AOI22xp33_ASAP7_75t_L g10692 ( 
.A1(n_9059),
.A2(n_7750),
.B1(n_8197),
.B2(n_7832),
.Y(n_10692)
);

NAND2xp5_ASAP7_75t_L g10693 ( 
.A(n_9648),
.B(n_8776),
.Y(n_10693)
);

OR2x6_ASAP7_75t_L g10694 ( 
.A(n_9065),
.B(n_8452),
.Y(n_10694)
);

INVx2_ASAP7_75t_L g10695 ( 
.A(n_9889),
.Y(n_10695)
);

OR2x2_ASAP7_75t_L g10696 ( 
.A(n_10281),
.B(n_8904),
.Y(n_10696)
);

INVx2_ASAP7_75t_L g10697 ( 
.A(n_9889),
.Y(n_10697)
);

INVx2_ASAP7_75t_L g10698 ( 
.A(n_9889),
.Y(n_10698)
);

NAND2xp5_ASAP7_75t_L g10699 ( 
.A(n_9648),
.B(n_8884),
.Y(n_10699)
);

INVx1_ASAP7_75t_L g10700 ( 
.A(n_9171),
.Y(n_10700)
);

INVx2_ASAP7_75t_L g10701 ( 
.A(n_9898),
.Y(n_10701)
);

INVx1_ASAP7_75t_L g10702 ( 
.A(n_9171),
.Y(n_10702)
);

INVx1_ASAP7_75t_L g10703 ( 
.A(n_9173),
.Y(n_10703)
);

INVx2_ASAP7_75t_L g10704 ( 
.A(n_9898),
.Y(n_10704)
);

INVx1_ASAP7_75t_L g10705 ( 
.A(n_9173),
.Y(n_10705)
);

AOI221xp5_ASAP7_75t_SL g10706 ( 
.A1(n_10172),
.A2(n_8476),
.B1(n_8272),
.B2(n_8265),
.C(n_8516),
.Y(n_10706)
);

OAI21x1_ASAP7_75t_L g10707 ( 
.A1(n_9852),
.A2(n_8894),
.B(n_8814),
.Y(n_10707)
);

NOR2x1_ASAP7_75t_L g10708 ( 
.A(n_9289),
.B(n_8452),
.Y(n_10708)
);

BUFx2_ASAP7_75t_L g10709 ( 
.A(n_10114),
.Y(n_10709)
);

INVx1_ASAP7_75t_L g10710 ( 
.A(n_9175),
.Y(n_10710)
);

INVx1_ASAP7_75t_L g10711 ( 
.A(n_9175),
.Y(n_10711)
);

BUFx2_ASAP7_75t_L g10712 ( 
.A(n_10114),
.Y(n_10712)
);

INVx2_ASAP7_75t_L g10713 ( 
.A(n_9898),
.Y(n_10713)
);

AND2x2_ASAP7_75t_L g10714 ( 
.A(n_9351),
.B(n_7744),
.Y(n_10714)
);

INVx3_ASAP7_75t_L g10715 ( 
.A(n_10170),
.Y(n_10715)
);

OR2x6_ASAP7_75t_L g10716 ( 
.A(n_9065),
.B(n_8452),
.Y(n_10716)
);

INVx1_ASAP7_75t_L g10717 ( 
.A(n_9177),
.Y(n_10717)
);

AO21x1_ASAP7_75t_SL g10718 ( 
.A1(n_9399),
.A2(n_8695),
.B(n_8688),
.Y(n_10718)
);

OAI21xp5_ASAP7_75t_L g10719 ( 
.A1(n_8988),
.A2(n_8243),
.B(n_8924),
.Y(n_10719)
);

INVx1_ASAP7_75t_L g10720 ( 
.A(n_9177),
.Y(n_10720)
);

OR2x2_ASAP7_75t_L g10721 ( 
.A(n_9702),
.B(n_8904),
.Y(n_10721)
);

INVx1_ASAP7_75t_L g10722 ( 
.A(n_9178),
.Y(n_10722)
);

INVx2_ASAP7_75t_L g10723 ( 
.A(n_9901),
.Y(n_10723)
);

INVx2_ASAP7_75t_L g10724 ( 
.A(n_9901),
.Y(n_10724)
);

NOR2xp33_ASAP7_75t_L g10725 ( 
.A(n_9489),
.B(n_7960),
.Y(n_10725)
);

INVx2_ASAP7_75t_L g10726 ( 
.A(n_9901),
.Y(n_10726)
);

OAI21x1_ASAP7_75t_L g10727 ( 
.A1(n_9852),
.A2(n_9893),
.B(n_9860),
.Y(n_10727)
);

OR2x6_ASAP7_75t_L g10728 ( 
.A(n_9065),
.B(n_9150),
.Y(n_10728)
);

INVx2_ASAP7_75t_L g10729 ( 
.A(n_9905),
.Y(n_10729)
);

INVx2_ASAP7_75t_L g10730 ( 
.A(n_9905),
.Y(n_10730)
);

INVx2_ASAP7_75t_L g10731 ( 
.A(n_9905),
.Y(n_10731)
);

INVx2_ASAP7_75t_L g10732 ( 
.A(n_9916),
.Y(n_10732)
);

INVx1_ASAP7_75t_L g10733 ( 
.A(n_9178),
.Y(n_10733)
);

INVx1_ASAP7_75t_L g10734 ( 
.A(n_9186),
.Y(n_10734)
);

INVx1_ASAP7_75t_L g10735 ( 
.A(n_9186),
.Y(n_10735)
);

INVx2_ASAP7_75t_L g10736 ( 
.A(n_9916),
.Y(n_10736)
);

AOI22xp33_ASAP7_75t_L g10737 ( 
.A1(n_9913),
.A2(n_7750),
.B1(n_7832),
.B2(n_7649),
.Y(n_10737)
);

INVx1_ASAP7_75t_L g10738 ( 
.A(n_9188),
.Y(n_10738)
);

BUFx2_ASAP7_75t_L g10739 ( 
.A(n_10114),
.Y(n_10739)
);

NOR2x1_ASAP7_75t_R g10740 ( 
.A(n_9627),
.B(n_8452),
.Y(n_10740)
);

CKINVDCx5p33_ASAP7_75t_R g10741 ( 
.A(n_10203),
.Y(n_10741)
);

INVx2_ASAP7_75t_SL g10742 ( 
.A(n_9497),
.Y(n_10742)
);

INVx2_ASAP7_75t_L g10743 ( 
.A(n_9916),
.Y(n_10743)
);

BUFx3_ASAP7_75t_L g10744 ( 
.A(n_9952),
.Y(n_10744)
);

HB1xp67_ASAP7_75t_L g10745 ( 
.A(n_9504),
.Y(n_10745)
);

INVx2_ASAP7_75t_L g10746 ( 
.A(n_9920),
.Y(n_10746)
);

INVx2_ASAP7_75t_SL g10747 ( 
.A(n_9624),
.Y(n_10747)
);

INVx1_ASAP7_75t_L g10748 ( 
.A(n_9188),
.Y(n_10748)
);

NOR2xp33_ASAP7_75t_L g10749 ( 
.A(n_9764),
.B(n_7960),
.Y(n_10749)
);

HB1xp67_ASAP7_75t_L g10750 ( 
.A(n_9775),
.Y(n_10750)
);

INVx1_ASAP7_75t_L g10751 ( 
.A(n_9189),
.Y(n_10751)
);

NOR2xp33_ASAP7_75t_L g10752 ( 
.A(n_9764),
.B(n_8823),
.Y(n_10752)
);

INVx2_ASAP7_75t_L g10753 ( 
.A(n_9920),
.Y(n_10753)
);

INVx2_ASAP7_75t_L g10754 ( 
.A(n_9920),
.Y(n_10754)
);

OAI21x1_ASAP7_75t_L g10755 ( 
.A1(n_9860),
.A2(n_8894),
.B(n_8814),
.Y(n_10755)
);

INVx1_ASAP7_75t_L g10756 ( 
.A(n_9189),
.Y(n_10756)
);

OAI22xp33_ASAP7_75t_L g10757 ( 
.A1(n_10146),
.A2(n_10147),
.B1(n_9055),
.B2(n_10172),
.Y(n_10757)
);

INVx1_ASAP7_75t_L g10758 ( 
.A(n_9190),
.Y(n_10758)
);

INVx1_ASAP7_75t_L g10759 ( 
.A(n_9190),
.Y(n_10759)
);

OAI21x1_ASAP7_75t_L g10760 ( 
.A1(n_9860),
.A2(n_9900),
.B(n_9893),
.Y(n_10760)
);

INVx1_ASAP7_75t_L g10761 ( 
.A(n_9195),
.Y(n_10761)
);

INVx2_ASAP7_75t_L g10762 ( 
.A(n_9922),
.Y(n_10762)
);

INVx2_ASAP7_75t_L g10763 ( 
.A(n_9922),
.Y(n_10763)
);

INVx2_ASAP7_75t_L g10764 ( 
.A(n_9922),
.Y(n_10764)
);

HB1xp67_ASAP7_75t_L g10765 ( 
.A(n_9778),
.Y(n_10765)
);

INVx3_ASAP7_75t_L g10766 ( 
.A(n_9706),
.Y(n_10766)
);

AND2x2_ASAP7_75t_L g10767 ( 
.A(n_9466),
.B(n_7744),
.Y(n_10767)
);

BUFx3_ASAP7_75t_L g10768 ( 
.A(n_9952),
.Y(n_10768)
);

HB1xp67_ASAP7_75t_L g10769 ( 
.A(n_9838),
.Y(n_10769)
);

INVx1_ASAP7_75t_L g10770 ( 
.A(n_9195),
.Y(n_10770)
);

INVx1_ASAP7_75t_L g10771 ( 
.A(n_9197),
.Y(n_10771)
);

INVx3_ASAP7_75t_L g10772 ( 
.A(n_9706),
.Y(n_10772)
);

INVx2_ASAP7_75t_L g10773 ( 
.A(n_9925),
.Y(n_10773)
);

INVx1_ASAP7_75t_L g10774 ( 
.A(n_9197),
.Y(n_10774)
);

OAI21x1_ASAP7_75t_L g10775 ( 
.A1(n_9893),
.A2(n_8819),
.B(n_8812),
.Y(n_10775)
);

BUFx3_ASAP7_75t_L g10776 ( 
.A(n_9952),
.Y(n_10776)
);

INVx2_ASAP7_75t_SL g10777 ( 
.A(n_9624),
.Y(n_10777)
);

AND2x2_ASAP7_75t_L g10778 ( 
.A(n_9470),
.B(n_7744),
.Y(n_10778)
);

INVx1_ASAP7_75t_L g10779 ( 
.A(n_9205),
.Y(n_10779)
);

INVx2_ASAP7_75t_L g10780 ( 
.A(n_9925),
.Y(n_10780)
);

HB1xp67_ASAP7_75t_L g10781 ( 
.A(n_9862),
.Y(n_10781)
);

INVx2_ASAP7_75t_L g10782 ( 
.A(n_9925),
.Y(n_10782)
);

INVx1_ASAP7_75t_L g10783 ( 
.A(n_9205),
.Y(n_10783)
);

BUFx3_ASAP7_75t_L g10784 ( 
.A(n_10114),
.Y(n_10784)
);

INVx2_ASAP7_75t_SL g10785 ( 
.A(n_9624),
.Y(n_10785)
);

INVx1_ASAP7_75t_L g10786 ( 
.A(n_9207),
.Y(n_10786)
);

OAI21x1_ASAP7_75t_L g10787 ( 
.A1(n_9900),
.A2(n_8819),
.B(n_8812),
.Y(n_10787)
);

INVx2_ASAP7_75t_L g10788 ( 
.A(n_9929),
.Y(n_10788)
);

AND2x2_ASAP7_75t_L g10789 ( 
.A(n_9470),
.B(n_7744),
.Y(n_10789)
);

AND2x2_ASAP7_75t_L g10790 ( 
.A(n_9496),
.B(n_8768),
.Y(n_10790)
);

INVx1_ASAP7_75t_L g10791 ( 
.A(n_9207),
.Y(n_10791)
);

INVx1_ASAP7_75t_L g10792 ( 
.A(n_9208),
.Y(n_10792)
);

AND2x2_ASAP7_75t_L g10793 ( 
.A(n_9496),
.B(n_9498),
.Y(n_10793)
);

AOI22xp33_ASAP7_75t_L g10794 ( 
.A1(n_9345),
.A2(n_7832),
.B1(n_7649),
.B2(n_7737),
.Y(n_10794)
);

OAI21xp5_ASAP7_75t_L g10795 ( 
.A1(n_10174),
.A2(n_8243),
.B(n_8924),
.Y(n_10795)
);

AOI22xp33_ASAP7_75t_SL g10796 ( 
.A1(n_9380),
.A2(n_9464),
.B1(n_10055),
.B2(n_9910),
.Y(n_10796)
);

INVx1_ASAP7_75t_L g10797 ( 
.A(n_9208),
.Y(n_10797)
);

INVx1_ASAP7_75t_L g10798 ( 
.A(n_9209),
.Y(n_10798)
);

INVx1_ASAP7_75t_L g10799 ( 
.A(n_9209),
.Y(n_10799)
);

INVx1_ASAP7_75t_L g10800 ( 
.A(n_9211),
.Y(n_10800)
);

AND2x2_ASAP7_75t_L g10801 ( 
.A(n_9498),
.B(n_8768),
.Y(n_10801)
);

INVx2_ASAP7_75t_SL g10802 ( 
.A(n_9624),
.Y(n_10802)
);

NAND2xp5_ASAP7_75t_L g10803 ( 
.A(n_9304),
.B(n_8884),
.Y(n_10803)
);

INVx2_ASAP7_75t_L g10804 ( 
.A(n_9929),
.Y(n_10804)
);

INVx2_ASAP7_75t_SL g10805 ( 
.A(n_10128),
.Y(n_10805)
);

AND2x2_ASAP7_75t_L g10806 ( 
.A(n_10213),
.B(n_9291),
.Y(n_10806)
);

HB1xp67_ASAP7_75t_L g10807 ( 
.A(n_9866),
.Y(n_10807)
);

NAND2xp5_ASAP7_75t_L g10808 ( 
.A(n_9304),
.B(n_8005),
.Y(n_10808)
);

INVx1_ASAP7_75t_L g10809 ( 
.A(n_9211),
.Y(n_10809)
);

AO21x2_ASAP7_75t_L g10810 ( 
.A1(n_9319),
.A2(n_7605),
.B(n_8663),
.Y(n_10810)
);

INVx2_ASAP7_75t_L g10811 ( 
.A(n_9929),
.Y(n_10811)
);

OAI21x1_ASAP7_75t_L g10812 ( 
.A1(n_9900),
.A2(n_8819),
.B(n_8812),
.Y(n_10812)
);

NAND2xp5_ASAP7_75t_L g10813 ( 
.A(n_9123),
.B(n_8005),
.Y(n_10813)
);

INVx2_ASAP7_75t_L g10814 ( 
.A(n_9931),
.Y(n_10814)
);

INVx1_ASAP7_75t_L g10815 ( 
.A(n_9215),
.Y(n_10815)
);

BUFx2_ASAP7_75t_L g10816 ( 
.A(n_10206),
.Y(n_10816)
);

INVx1_ASAP7_75t_L g10817 ( 
.A(n_9215),
.Y(n_10817)
);

INVx1_ASAP7_75t_L g10818 ( 
.A(n_9217),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_9217),
.Y(n_10819)
);

INVx1_ASAP7_75t_L g10820 ( 
.A(n_9219),
.Y(n_10820)
);

AND2x2_ASAP7_75t_L g10821 ( 
.A(n_9291),
.B(n_8768),
.Y(n_10821)
);

INVx2_ASAP7_75t_L g10822 ( 
.A(n_9931),
.Y(n_10822)
);

INVx3_ASAP7_75t_L g10823 ( 
.A(n_9706),
.Y(n_10823)
);

HB1xp67_ASAP7_75t_L g10824 ( 
.A(n_9869),
.Y(n_10824)
);

HB1xp67_ASAP7_75t_L g10825 ( 
.A(n_9890),
.Y(n_10825)
);

INVx1_ASAP7_75t_L g10826 ( 
.A(n_9219),
.Y(n_10826)
);

INVx1_ASAP7_75t_L g10827 ( 
.A(n_9220),
.Y(n_10827)
);

OAI21xp5_ASAP7_75t_L g10828 ( 
.A1(n_9326),
.A2(n_8743),
.B(n_8706),
.Y(n_10828)
);

NAND2xp33_ASAP7_75t_SL g10829 ( 
.A(n_9277),
.B(n_8281),
.Y(n_10829)
);

INVx1_ASAP7_75t_L g10830 ( 
.A(n_9220),
.Y(n_10830)
);

CKINVDCx20_ASAP7_75t_R g10831 ( 
.A(n_9174),
.Y(n_10831)
);

INVx1_ASAP7_75t_L g10832 ( 
.A(n_9222),
.Y(n_10832)
);

INVx2_ASAP7_75t_L g10833 ( 
.A(n_9931),
.Y(n_10833)
);

INVx4_ASAP7_75t_L g10834 ( 
.A(n_9013),
.Y(n_10834)
);

INVx4_ASAP7_75t_L g10835 ( 
.A(n_9013),
.Y(n_10835)
);

AND2x2_ASAP7_75t_L g10836 ( 
.A(n_9298),
.B(n_8863),
.Y(n_10836)
);

INVx2_ASAP7_75t_L g10837 ( 
.A(n_9937),
.Y(n_10837)
);

INVx2_ASAP7_75t_SL g10838 ( 
.A(n_10128),
.Y(n_10838)
);

HB1xp67_ASAP7_75t_L g10839 ( 
.A(n_9943),
.Y(n_10839)
);

AOI22xp5_ASAP7_75t_L g10840 ( 
.A1(n_9380),
.A2(n_8909),
.B1(n_7819),
.B2(n_7607),
.Y(n_10840)
);

OAI21x1_ASAP7_75t_L g10841 ( 
.A1(n_9927),
.A2(n_8829),
.B(n_8826),
.Y(n_10841)
);

INVx3_ASAP7_75t_L g10842 ( 
.A(n_9863),
.Y(n_10842)
);

INVx2_ASAP7_75t_L g10843 ( 
.A(n_9937),
.Y(n_10843)
);

INVx3_ASAP7_75t_L g10844 ( 
.A(n_9863),
.Y(n_10844)
);

INVx1_ASAP7_75t_L g10845 ( 
.A(n_9222),
.Y(n_10845)
);

NAND2xp5_ASAP7_75t_L g10846 ( 
.A(n_9123),
.B(n_8024),
.Y(n_10846)
);

AOI22xp33_ASAP7_75t_L g10847 ( 
.A1(n_9345),
.A2(n_7832),
.B1(n_7737),
.B2(n_8221),
.Y(n_10847)
);

INVx2_ASAP7_75t_L g10848 ( 
.A(n_9937),
.Y(n_10848)
);

INVx1_ASAP7_75t_L g10849 ( 
.A(n_9230),
.Y(n_10849)
);

BUFx3_ASAP7_75t_L g10850 ( 
.A(n_10206),
.Y(n_10850)
);

INVx1_ASAP7_75t_L g10851 ( 
.A(n_9230),
.Y(n_10851)
);

AO21x1_ASAP7_75t_SL g10852 ( 
.A1(n_9282),
.A2(n_8678),
.B(n_8465),
.Y(n_10852)
);

OAI21x1_ASAP7_75t_L g10853 ( 
.A1(n_9927),
.A2(n_8829),
.B(n_8826),
.Y(n_10853)
);

INVx1_ASAP7_75t_L g10854 ( 
.A(n_9231),
.Y(n_10854)
);

OAI21x1_ASAP7_75t_L g10855 ( 
.A1(n_9927),
.A2(n_8829),
.B(n_8826),
.Y(n_10855)
);

INVx1_ASAP7_75t_L g10856 ( 
.A(n_9231),
.Y(n_10856)
);

OAI21x1_ASAP7_75t_L g10857 ( 
.A1(n_9958),
.A2(n_8845),
.B(n_8841),
.Y(n_10857)
);

AND2x2_ASAP7_75t_L g10858 ( 
.A(n_9298),
.B(n_8863),
.Y(n_10858)
);

CKINVDCx20_ASAP7_75t_R g10859 ( 
.A(n_9185),
.Y(n_10859)
);

OAI22xp5_ASAP7_75t_L g10860 ( 
.A1(n_9760),
.A2(n_9112),
.B1(n_9733),
.B2(n_9932),
.Y(n_10860)
);

AND2x4_ASAP7_75t_L g10861 ( 
.A(n_9416),
.B(n_8556),
.Y(n_10861)
);

INVx2_ASAP7_75t_L g10862 ( 
.A(n_9945),
.Y(n_10862)
);

OR2x2_ASAP7_75t_L g10863 ( 
.A(n_9702),
.B(n_9797),
.Y(n_10863)
);

INVx2_ASAP7_75t_L g10864 ( 
.A(n_9945),
.Y(n_10864)
);

OAI21x1_ASAP7_75t_L g10865 ( 
.A1(n_9958),
.A2(n_8845),
.B(n_8841),
.Y(n_10865)
);

NAND2xp5_ASAP7_75t_L g10866 ( 
.A(n_9140),
.B(n_9605),
.Y(n_10866)
);

OAI21x1_ASAP7_75t_L g10867 ( 
.A1(n_9958),
.A2(n_8845),
.B(n_8841),
.Y(n_10867)
);

INVx2_ASAP7_75t_L g10868 ( 
.A(n_9945),
.Y(n_10868)
);

INVx1_ASAP7_75t_L g10869 ( 
.A(n_9235),
.Y(n_10869)
);

HB1xp67_ASAP7_75t_L g10870 ( 
.A(n_9981),
.Y(n_10870)
);

INVx1_ASAP7_75t_SL g10871 ( 
.A(n_9567),
.Y(n_10871)
);

HB1xp67_ASAP7_75t_L g10872 ( 
.A(n_9986),
.Y(n_10872)
);

INVx3_ASAP7_75t_L g10873 ( 
.A(n_9863),
.Y(n_10873)
);

INVx2_ASAP7_75t_L g10874 ( 
.A(n_9948),
.Y(n_10874)
);

BUFx12f_ASAP7_75t_L g10875 ( 
.A(n_9651),
.Y(n_10875)
);

HB1xp67_ASAP7_75t_L g10876 ( 
.A(n_10076),
.Y(n_10876)
);

INVx1_ASAP7_75t_L g10877 ( 
.A(n_9235),
.Y(n_10877)
);

NAND2xp5_ASAP7_75t_L g10878 ( 
.A(n_9140),
.B(n_8024),
.Y(n_10878)
);

INVx1_ASAP7_75t_L g10879 ( 
.A(n_9250),
.Y(n_10879)
);

INVx2_ASAP7_75t_SL g10880 ( 
.A(n_10128),
.Y(n_10880)
);

OAI21xp5_ASAP7_75t_L g10881 ( 
.A1(n_9873),
.A2(n_9980),
.B(n_9938),
.Y(n_10881)
);

INVx2_ASAP7_75t_L g10882 ( 
.A(n_9948),
.Y(n_10882)
);

INVx1_ASAP7_75t_L g10883 ( 
.A(n_9250),
.Y(n_10883)
);

INVx1_ASAP7_75t_SL g10884 ( 
.A(n_9836),
.Y(n_10884)
);

BUFx4f_ASAP7_75t_L g10885 ( 
.A(n_9026),
.Y(n_10885)
);

INVx1_ASAP7_75t_L g10886 ( 
.A(n_9251),
.Y(n_10886)
);

INVx1_ASAP7_75t_L g10887 ( 
.A(n_9251),
.Y(n_10887)
);

AOI22xp33_ASAP7_75t_L g10888 ( 
.A1(n_9049),
.A2(n_7737),
.B1(n_8221),
.B2(n_7700),
.Y(n_10888)
);

NAND3x1_ASAP7_75t_L g10889 ( 
.A(n_9873),
.B(n_8670),
.C(n_8395),
.Y(n_10889)
);

INVx1_ASAP7_75t_L g10890 ( 
.A(n_9936),
.Y(n_10890)
);

OR2x2_ASAP7_75t_L g10891 ( 
.A(n_9797),
.B(n_8576),
.Y(n_10891)
);

INVx1_ASAP7_75t_L g10892 ( 
.A(n_9936),
.Y(n_10892)
);

AO21x1_ASAP7_75t_SL g10893 ( 
.A1(n_9283),
.A2(n_8678),
.B(n_8465),
.Y(n_10893)
);

INVx2_ASAP7_75t_L g10894 ( 
.A(n_9948),
.Y(n_10894)
);

INVx1_ASAP7_75t_L g10895 ( 
.A(n_9944),
.Y(n_10895)
);

INVx1_ASAP7_75t_L g10896 ( 
.A(n_9944),
.Y(n_10896)
);

INVx1_ASAP7_75t_L g10897 ( 
.A(n_9946),
.Y(n_10897)
);

AND2x2_ASAP7_75t_L g10898 ( 
.A(n_9891),
.B(n_8863),
.Y(n_10898)
);

BUFx3_ASAP7_75t_L g10899 ( 
.A(n_10206),
.Y(n_10899)
);

HB1xp67_ASAP7_75t_L g10900 ( 
.A(n_10110),
.Y(n_10900)
);

AND2x2_ASAP7_75t_L g10901 ( 
.A(n_9891),
.B(n_8875),
.Y(n_10901)
);

INVxp67_ASAP7_75t_L g10902 ( 
.A(n_8979),
.Y(n_10902)
);

AND2x2_ASAP7_75t_L g10903 ( 
.A(n_10067),
.B(n_8875),
.Y(n_10903)
);

INVxp33_ASAP7_75t_L g10904 ( 
.A(n_9485),
.Y(n_10904)
);

HB1xp67_ASAP7_75t_L g10905 ( 
.A(n_10118),
.Y(n_10905)
);

OAI21x1_ASAP7_75t_L g10906 ( 
.A1(n_9346),
.A2(n_8870),
.B(n_8869),
.Y(n_10906)
);

OAI21x1_ASAP7_75t_L g10907 ( 
.A1(n_9346),
.A2(n_8870),
.B(n_8869),
.Y(n_10907)
);

INVx1_ASAP7_75t_L g10908 ( 
.A(n_9946),
.Y(n_10908)
);

INVx1_ASAP7_75t_L g10909 ( 
.A(n_9951),
.Y(n_10909)
);

INVx1_ASAP7_75t_L g10910 ( 
.A(n_9951),
.Y(n_10910)
);

HB1xp67_ASAP7_75t_L g10911 ( 
.A(n_10157),
.Y(n_10911)
);

AND2x2_ASAP7_75t_L g10912 ( 
.A(n_10067),
.B(n_8875),
.Y(n_10912)
);

INVx1_ASAP7_75t_L g10913 ( 
.A(n_9955),
.Y(n_10913)
);

AO21x2_ASAP7_75t_L g10914 ( 
.A1(n_9736),
.A2(n_8752),
.B(n_7874),
.Y(n_10914)
);

INVx2_ASAP7_75t_L g10915 ( 
.A(n_9954),
.Y(n_10915)
);

AND2x4_ASAP7_75t_L g10916 ( 
.A(n_9416),
.B(n_8556),
.Y(n_10916)
);

HB1xp67_ASAP7_75t_L g10917 ( 
.A(n_10160),
.Y(n_10917)
);

INVx1_ASAP7_75t_L g10918 ( 
.A(n_9955),
.Y(n_10918)
);

INVx1_ASAP7_75t_L g10919 ( 
.A(n_9957),
.Y(n_10919)
);

INVx2_ASAP7_75t_L g10920 ( 
.A(n_9954),
.Y(n_10920)
);

BUFx3_ASAP7_75t_L g10921 ( 
.A(n_10206),
.Y(n_10921)
);

INVx1_ASAP7_75t_L g10922 ( 
.A(n_9957),
.Y(n_10922)
);

INVx1_ASAP7_75t_L g10923 ( 
.A(n_9959),
.Y(n_10923)
);

INVx2_ASAP7_75t_L g10924 ( 
.A(n_9954),
.Y(n_10924)
);

NAND2xp5_ASAP7_75t_L g10925 ( 
.A(n_9791),
.B(n_8084),
.Y(n_10925)
);

OAI21x1_ASAP7_75t_SL g10926 ( 
.A1(n_9306),
.A2(n_7802),
.B(n_8371),
.Y(n_10926)
);

OAI21x1_ASAP7_75t_L g10927 ( 
.A1(n_9346),
.A2(n_8870),
.B(n_8869),
.Y(n_10927)
);

INVx2_ASAP7_75t_L g10928 ( 
.A(n_9964),
.Y(n_10928)
);

INVx1_ASAP7_75t_L g10929 ( 
.A(n_9959),
.Y(n_10929)
);

INVx2_ASAP7_75t_L g10930 ( 
.A(n_9964),
.Y(n_10930)
);

AOI22xp5_ASAP7_75t_L g10931 ( 
.A1(n_10066),
.A2(n_8909),
.B1(n_7819),
.B2(n_8492),
.Y(n_10931)
);

INVx1_ASAP7_75t_L g10932 ( 
.A(n_9961),
.Y(n_10932)
);

INVx1_ASAP7_75t_L g10933 ( 
.A(n_9961),
.Y(n_10933)
);

INVx1_ASAP7_75t_L g10934 ( 
.A(n_9968),
.Y(n_10934)
);

AND2x2_ASAP7_75t_L g10935 ( 
.A(n_10067),
.B(n_8939),
.Y(n_10935)
);

INVx2_ASAP7_75t_L g10936 ( 
.A(n_9964),
.Y(n_10936)
);

CKINVDCx12_ASAP7_75t_R g10937 ( 
.A(n_9464),
.Y(n_10937)
);

INVx2_ASAP7_75t_L g10938 ( 
.A(n_9969),
.Y(n_10938)
);

AND2x4_ASAP7_75t_L g10939 ( 
.A(n_9416),
.B(n_8556),
.Y(n_10939)
);

INVx1_ASAP7_75t_L g10940 ( 
.A(n_9968),
.Y(n_10940)
);

INVx1_ASAP7_75t_L g10941 ( 
.A(n_9974),
.Y(n_10941)
);

AOI22xp33_ASAP7_75t_L g10942 ( 
.A1(n_9049),
.A2(n_7737),
.B1(n_7700),
.B2(n_8311),
.Y(n_10942)
);

INVx1_ASAP7_75t_L g10943 ( 
.A(n_9974),
.Y(n_10943)
);

INVx2_ASAP7_75t_L g10944 ( 
.A(n_9969),
.Y(n_10944)
);

BUFx2_ASAP7_75t_L g10945 ( 
.A(n_9467),
.Y(n_10945)
);

BUFx3_ASAP7_75t_L g10946 ( 
.A(n_10128),
.Y(n_10946)
);

BUFx3_ASAP7_75t_L g10947 ( 
.A(n_9097),
.Y(n_10947)
);

AND2x2_ASAP7_75t_L g10948 ( 
.A(n_10067),
.B(n_8939),
.Y(n_10948)
);

INVx1_ASAP7_75t_L g10949 ( 
.A(n_9977),
.Y(n_10949)
);

HB1xp67_ASAP7_75t_L g10950 ( 
.A(n_10163),
.Y(n_10950)
);

BUFx2_ASAP7_75t_L g10951 ( 
.A(n_9467),
.Y(n_10951)
);

INVx2_ASAP7_75t_L g10952 ( 
.A(n_9969),
.Y(n_10952)
);

INVx2_ASAP7_75t_L g10953 ( 
.A(n_9979),
.Y(n_10953)
);

INVx1_ASAP7_75t_L g10954 ( 
.A(n_9977),
.Y(n_10954)
);

BUFx4f_ASAP7_75t_SL g10955 ( 
.A(n_9026),
.Y(n_10955)
);

OAI21x1_ASAP7_75t_L g10956 ( 
.A1(n_9388),
.A2(n_8880),
.B(n_8871),
.Y(n_10956)
);

INVx2_ASAP7_75t_L g10957 ( 
.A(n_9979),
.Y(n_10957)
);

INVx2_ASAP7_75t_L g10958 ( 
.A(n_9979),
.Y(n_10958)
);

INVx2_ASAP7_75t_L g10959 ( 
.A(n_9982),
.Y(n_10959)
);

AND2x4_ASAP7_75t_L g10960 ( 
.A(n_9416),
.B(n_8556),
.Y(n_10960)
);

INVx2_ASAP7_75t_L g10961 ( 
.A(n_9982),
.Y(n_10961)
);

BUFx3_ASAP7_75t_L g10962 ( 
.A(n_9097),
.Y(n_10962)
);

BUFx2_ASAP7_75t_L g10963 ( 
.A(n_9618),
.Y(n_10963)
);

INVx1_ASAP7_75t_L g10964 ( 
.A(n_9988),
.Y(n_10964)
);

BUFx4f_ASAP7_75t_SL g10965 ( 
.A(n_9026),
.Y(n_10965)
);

INVx1_ASAP7_75t_L g10966 ( 
.A(n_9988),
.Y(n_10966)
);

NAND2xp5_ASAP7_75t_L g10967 ( 
.A(n_9034),
.B(n_8084),
.Y(n_10967)
);

AND2x2_ASAP7_75t_L g10968 ( 
.A(n_9796),
.B(n_8939),
.Y(n_10968)
);

INVx3_ASAP7_75t_L g10969 ( 
.A(n_9973),
.Y(n_10969)
);

INVx1_ASAP7_75t_L g10970 ( 
.A(n_9995),
.Y(n_10970)
);

INVx2_ASAP7_75t_L g10971 ( 
.A(n_9982),
.Y(n_10971)
);

OA21x2_ASAP7_75t_L g10972 ( 
.A1(n_9759),
.A2(n_8342),
.B(n_8848),
.Y(n_10972)
);

OAI21x1_ASAP7_75t_L g10973 ( 
.A1(n_9388),
.A2(n_8880),
.B(n_8871),
.Y(n_10973)
);

INVxp67_ASAP7_75t_L g10974 ( 
.A(n_8979),
.Y(n_10974)
);

INVx1_ASAP7_75t_L g10975 ( 
.A(n_9995),
.Y(n_10975)
);

INVx1_ASAP7_75t_L g10976 ( 
.A(n_9998),
.Y(n_10976)
);

INVx3_ASAP7_75t_L g10977 ( 
.A(n_9973),
.Y(n_10977)
);

INVx3_ASAP7_75t_L g10978 ( 
.A(n_9973),
.Y(n_10978)
);

NOR2xp33_ASAP7_75t_L g10979 ( 
.A(n_9932),
.B(n_8823),
.Y(n_10979)
);

INVx1_ASAP7_75t_L g10980 ( 
.A(n_9998),
.Y(n_10980)
);

INVx2_ASAP7_75t_L g10981 ( 
.A(n_9983),
.Y(n_10981)
);

INVx2_ASAP7_75t_L g10982 ( 
.A(n_9983),
.Y(n_10982)
);

OAI211xp5_ASAP7_75t_L g10983 ( 
.A1(n_9938),
.A2(n_8310),
.B(n_7970),
.C(n_7981),
.Y(n_10983)
);

OAI21x1_ASAP7_75t_L g10984 ( 
.A1(n_9388),
.A2(n_9431),
.B(n_9718),
.Y(n_10984)
);

INVx2_ASAP7_75t_L g10985 ( 
.A(n_9983),
.Y(n_10985)
);

INVx2_ASAP7_75t_L g10986 ( 
.A(n_9984),
.Y(n_10986)
);

INVx1_ASAP7_75t_L g10987 ( 
.A(n_10006),
.Y(n_10987)
);

INVx1_ASAP7_75t_L g10988 ( 
.A(n_10006),
.Y(n_10988)
);

AND2x2_ASAP7_75t_L g10989 ( 
.A(n_9796),
.B(n_7777),
.Y(n_10989)
);

OR2x6_ASAP7_75t_L g10990 ( 
.A(n_9065),
.B(n_7926),
.Y(n_10990)
);

INVx1_ASAP7_75t_L g10991 ( 
.A(n_10007),
.Y(n_10991)
);

O2A1O1Ixp5_ASAP7_75t_L g10992 ( 
.A1(n_9725),
.A2(n_8699),
.B(n_8815),
.C(n_8383),
.Y(n_10992)
);

INVx1_ASAP7_75t_L g10993 ( 
.A(n_10007),
.Y(n_10993)
);

INVx1_ASAP7_75t_L g10994 ( 
.A(n_10009),
.Y(n_10994)
);

OAI21xp5_ASAP7_75t_L g10995 ( 
.A1(n_9980),
.A2(n_8743),
.B(n_8706),
.Y(n_10995)
);

INVx1_ASAP7_75t_L g10996 ( 
.A(n_10009),
.Y(n_10996)
);

OAI22xp5_ASAP7_75t_L g10997 ( 
.A1(n_9133),
.A2(n_8324),
.B1(n_8314),
.B2(n_8205),
.Y(n_10997)
);

INVx2_ASAP7_75t_L g10998 ( 
.A(n_9984),
.Y(n_10998)
);

CKINVDCx5p33_ASAP7_75t_R g10999 ( 
.A(n_10264),
.Y(n_10999)
);

INVx1_ASAP7_75t_SL g11000 ( 
.A(n_9836),
.Y(n_11000)
);

HB1xp67_ASAP7_75t_L g11001 ( 
.A(n_10175),
.Y(n_11001)
);

INVx1_ASAP7_75t_L g11002 ( 
.A(n_10010),
.Y(n_11002)
);

OAI21x1_ASAP7_75t_L g11003 ( 
.A1(n_9431),
.A2(n_9738),
.B(n_9729),
.Y(n_11003)
);

INVx2_ASAP7_75t_L g11004 ( 
.A(n_9984),
.Y(n_11004)
);

OAI21x1_ASAP7_75t_L g11005 ( 
.A1(n_9431),
.A2(n_9738),
.B(n_9729),
.Y(n_11005)
);

AOI21xp5_ASAP7_75t_L g11006 ( 
.A1(n_9412),
.A2(n_8624),
.B(n_8533),
.Y(n_11006)
);

INVx2_ASAP7_75t_L g11007 ( 
.A(n_9985),
.Y(n_11007)
);

AND2x2_ASAP7_75t_L g11008 ( 
.A(n_9055),
.B(n_7777),
.Y(n_11008)
);

BUFx6f_ASAP7_75t_L g11009 ( 
.A(n_9026),
.Y(n_11009)
);

HB1xp67_ASAP7_75t_L g11010 ( 
.A(n_10185),
.Y(n_11010)
);

AO21x2_ASAP7_75t_L g11011 ( 
.A1(n_9736),
.A2(n_7874),
.B(n_8108),
.Y(n_11011)
);

INVx2_ASAP7_75t_L g11012 ( 
.A(n_9985),
.Y(n_11012)
);

OAI21xp5_ASAP7_75t_L g11013 ( 
.A1(n_9819),
.A2(n_7981),
.B(n_8265),
.Y(n_11013)
);

INVx1_ASAP7_75t_L g11014 ( 
.A(n_10010),
.Y(n_11014)
);

BUFx2_ASAP7_75t_SL g11015 ( 
.A(n_10267),
.Y(n_11015)
);

INVx2_ASAP7_75t_L g11016 ( 
.A(n_9985),
.Y(n_11016)
);

INVx4_ASAP7_75t_L g11017 ( 
.A(n_9026),
.Y(n_11017)
);

INVx2_ASAP7_75t_L g11018 ( 
.A(n_9991),
.Y(n_11018)
);

BUFx2_ASAP7_75t_L g11019 ( 
.A(n_9618),
.Y(n_11019)
);

NAND2xp5_ASAP7_75t_L g11020 ( 
.A(n_9034),
.B(n_8177),
.Y(n_11020)
);

AND2x4_ASAP7_75t_L g11021 ( 
.A(n_9416),
.B(n_8579),
.Y(n_11021)
);

NAND2xp33_ASAP7_75t_R g11022 ( 
.A(n_9656),
.B(n_8514),
.Y(n_11022)
);

INVx1_ASAP7_75t_L g11023 ( 
.A(n_10012),
.Y(n_11023)
);

INVx1_ASAP7_75t_L g11024 ( 
.A(n_10012),
.Y(n_11024)
);

AND2x2_ASAP7_75t_L g11025 ( 
.A(n_9914),
.B(n_7777),
.Y(n_11025)
);

AND2x2_ASAP7_75t_L g11026 ( 
.A(n_9914),
.B(n_7777),
.Y(n_11026)
);

OR2x6_ASAP7_75t_L g11027 ( 
.A(n_9150),
.B(n_7926),
.Y(n_11027)
);

OAI21x1_ASAP7_75t_L g11028 ( 
.A1(n_9802),
.A2(n_8880),
.B(n_8871),
.Y(n_11028)
);

INVx1_ASAP7_75t_L g11029 ( 
.A(n_10021),
.Y(n_11029)
);

INVx1_ASAP7_75t_L g11030 ( 
.A(n_10021),
.Y(n_11030)
);

INVx1_ASAP7_75t_L g11031 ( 
.A(n_10027),
.Y(n_11031)
);

INVx2_ASAP7_75t_L g11032 ( 
.A(n_9991),
.Y(n_11032)
);

INVx1_ASAP7_75t_L g11033 ( 
.A(n_10027),
.Y(n_11033)
);

INVx1_ASAP7_75t_L g11034 ( 
.A(n_10030),
.Y(n_11034)
);

INVx2_ASAP7_75t_L g11035 ( 
.A(n_9991),
.Y(n_11035)
);

INVx1_ASAP7_75t_L g11036 ( 
.A(n_10030),
.Y(n_11036)
);

BUFx3_ASAP7_75t_L g11037 ( 
.A(n_9097),
.Y(n_11037)
);

OAI21x1_ASAP7_75t_L g11038 ( 
.A1(n_9802),
.A2(n_8926),
.B(n_8881),
.Y(n_11038)
);

INVx2_ASAP7_75t_L g11039 ( 
.A(n_9994),
.Y(n_11039)
);

INVx1_ASAP7_75t_L g11040 ( 
.A(n_10031),
.Y(n_11040)
);

BUFx6f_ASAP7_75t_L g11041 ( 
.A(n_9026),
.Y(n_11041)
);

INVx1_ASAP7_75t_L g11042 ( 
.A(n_10031),
.Y(n_11042)
);

OAI21x1_ASAP7_75t_L g11043 ( 
.A1(n_9823),
.A2(n_9950),
.B(n_9549),
.Y(n_11043)
);

INVx1_ASAP7_75t_L g11044 ( 
.A(n_10038),
.Y(n_11044)
);

INVx2_ASAP7_75t_L g11045 ( 
.A(n_9994),
.Y(n_11045)
);

INVx2_ASAP7_75t_L g11046 ( 
.A(n_9994),
.Y(n_11046)
);

INVx2_ASAP7_75t_L g11047 ( 
.A(n_10011),
.Y(n_11047)
);

INVx1_ASAP7_75t_L g11048 ( 
.A(n_10038),
.Y(n_11048)
);

AND2x2_ASAP7_75t_L g11049 ( 
.A(n_9956),
.B(n_7777),
.Y(n_11049)
);

HB1xp67_ASAP7_75t_SL g11050 ( 
.A(n_9661),
.Y(n_11050)
);

INVx2_ASAP7_75t_L g11051 ( 
.A(n_10011),
.Y(n_11051)
);

INVx1_ASAP7_75t_L g11052 ( 
.A(n_10043),
.Y(n_11052)
);

AOI22xp33_ASAP7_75t_SL g11053 ( 
.A1(n_9638),
.A2(n_7842),
.B1(n_7843),
.B2(n_8108),
.Y(n_11053)
);

OA21x2_ASAP7_75t_L g11054 ( 
.A1(n_9759),
.A2(n_8848),
.B(n_8676),
.Y(n_11054)
);

INVx2_ASAP7_75t_L g11055 ( 
.A(n_10011),
.Y(n_11055)
);

BUFx2_ASAP7_75t_L g11056 ( 
.A(n_9618),
.Y(n_11056)
);

OR2x2_ASAP7_75t_L g11057 ( 
.A(n_9805),
.B(n_8576),
.Y(n_11057)
);

INVx1_ASAP7_75t_L g11058 ( 
.A(n_10043),
.Y(n_11058)
);

INVx1_ASAP7_75t_L g11059 ( 
.A(n_10046),
.Y(n_11059)
);

HB1xp67_ASAP7_75t_SL g11060 ( 
.A(n_9661),
.Y(n_11060)
);

INVx1_ASAP7_75t_L g11061 ( 
.A(n_10046),
.Y(n_11061)
);

INVx1_ASAP7_75t_L g11062 ( 
.A(n_10052),
.Y(n_11062)
);

INVx2_ASAP7_75t_L g11063 ( 
.A(n_10035),
.Y(n_11063)
);

INVx2_ASAP7_75t_L g11064 ( 
.A(n_10035),
.Y(n_11064)
);

INVx2_ASAP7_75t_L g11065 ( 
.A(n_10035),
.Y(n_11065)
);

AO31x2_ASAP7_75t_L g11066 ( 
.A1(n_9725),
.A2(n_7669),
.A3(n_7608),
.B(n_8837),
.Y(n_11066)
);

INVx2_ASAP7_75t_L g11067 ( 
.A(n_10037),
.Y(n_11067)
);

INVx3_ASAP7_75t_L g11068 ( 
.A(n_9996),
.Y(n_11068)
);

AOI22xp33_ASAP7_75t_L g11069 ( 
.A1(n_9412),
.A2(n_7737),
.B1(n_7700),
.B2(n_8311),
.Y(n_11069)
);

NAND2xp5_ASAP7_75t_L g11070 ( 
.A(n_9060),
.B(n_8177),
.Y(n_11070)
);

AND2x2_ASAP7_75t_L g11071 ( 
.A(n_9956),
.B(n_7787),
.Y(n_11071)
);

AND2x2_ASAP7_75t_L g11072 ( 
.A(n_9962),
.B(n_7787),
.Y(n_11072)
);

BUFx2_ASAP7_75t_SL g11073 ( 
.A(n_9066),
.Y(n_11073)
);

INVx1_ASAP7_75t_L g11074 ( 
.A(n_10052),
.Y(n_11074)
);

NAND2xp5_ASAP7_75t_SL g11075 ( 
.A(n_9848),
.B(n_8719),
.Y(n_11075)
);

NAND2xp5_ASAP7_75t_L g11076 ( 
.A(n_9060),
.B(n_8264),
.Y(n_11076)
);

BUFx2_ASAP7_75t_L g11077 ( 
.A(n_10000),
.Y(n_11077)
);

INVx2_ASAP7_75t_L g11078 ( 
.A(n_10037),
.Y(n_11078)
);

AND2x2_ASAP7_75t_L g11079 ( 
.A(n_9962),
.B(n_7787),
.Y(n_11079)
);

INVx2_ASAP7_75t_L g11080 ( 
.A(n_10037),
.Y(n_11080)
);

AND2x2_ASAP7_75t_L g11081 ( 
.A(n_10122),
.B(n_7787),
.Y(n_11081)
);

NAND2x1_ASAP7_75t_L g11082 ( 
.A(n_9557),
.B(n_8790),
.Y(n_11082)
);

BUFx2_ASAP7_75t_L g11083 ( 
.A(n_10000),
.Y(n_11083)
);

AO21x2_ASAP7_75t_L g11084 ( 
.A1(n_9319),
.A2(n_7874),
.B(n_8108),
.Y(n_11084)
);

AO21x2_ASAP7_75t_L g11085 ( 
.A1(n_9319),
.A2(n_8050),
.B(n_8068),
.Y(n_11085)
);

INVx1_ASAP7_75t_L g11086 ( 
.A(n_10053),
.Y(n_11086)
);

OA21x2_ASAP7_75t_L g11087 ( 
.A1(n_9768),
.A2(n_8676),
.B(n_8675),
.Y(n_11087)
);

BUFx2_ASAP7_75t_L g11088 ( 
.A(n_10000),
.Y(n_11088)
);

INVx2_ASAP7_75t_L g11089 ( 
.A(n_10039),
.Y(n_11089)
);

INVx1_ASAP7_75t_L g11090 ( 
.A(n_10053),
.Y(n_11090)
);

OAI21x1_ASAP7_75t_L g11091 ( 
.A1(n_9823),
.A2(n_8926),
.B(n_8881),
.Y(n_11091)
);

INVx1_ASAP7_75t_L g11092 ( 
.A(n_10057),
.Y(n_11092)
);

OAI21x1_ASAP7_75t_L g11093 ( 
.A1(n_9950),
.A2(n_8926),
.B(n_8881),
.Y(n_11093)
);

AO21x2_ASAP7_75t_L g11094 ( 
.A1(n_9621),
.A2(n_8815),
.B(n_8344),
.Y(n_11094)
);

AND2x2_ASAP7_75t_L g11095 ( 
.A(n_10122),
.B(n_7787),
.Y(n_11095)
);

INVx1_ASAP7_75t_L g11096 ( 
.A(n_10057),
.Y(n_11096)
);

INVx2_ASAP7_75t_L g11097 ( 
.A(n_10039),
.Y(n_11097)
);

AND2x2_ASAP7_75t_L g11098 ( 
.A(n_10139),
.B(n_7789),
.Y(n_11098)
);

INVx3_ASAP7_75t_L g11099 ( 
.A(n_9996),
.Y(n_11099)
);

INVx2_ASAP7_75t_L g11100 ( 
.A(n_10039),
.Y(n_11100)
);

INVx1_ASAP7_75t_L g11101 ( 
.A(n_10059),
.Y(n_11101)
);

INVx1_ASAP7_75t_L g11102 ( 
.A(n_10059),
.Y(n_11102)
);

INVx1_ASAP7_75t_L g11103 ( 
.A(n_10060),
.Y(n_11103)
);

AND2x2_ASAP7_75t_L g11104 ( 
.A(n_10139),
.B(n_10201),
.Y(n_11104)
);

AND2x2_ASAP7_75t_L g11105 ( 
.A(n_10201),
.B(n_7789),
.Y(n_11105)
);

INVx2_ASAP7_75t_L g11106 ( 
.A(n_10041),
.Y(n_11106)
);

NAND2xp5_ASAP7_75t_L g11107 ( 
.A(n_9165),
.B(n_9433),
.Y(n_11107)
);

INVx2_ASAP7_75t_L g11108 ( 
.A(n_10041),
.Y(n_11108)
);

AND2x2_ASAP7_75t_L g11109 ( 
.A(n_10202),
.B(n_7789),
.Y(n_11109)
);

INVx2_ASAP7_75t_L g11110 ( 
.A(n_10041),
.Y(n_11110)
);

OR2x2_ASAP7_75t_L g11111 ( 
.A(n_9805),
.B(n_8800),
.Y(n_11111)
);

AO21x2_ASAP7_75t_L g11112 ( 
.A1(n_9621),
.A2(n_8344),
.B(n_8486),
.Y(n_11112)
);

INVx1_ASAP7_75t_L g11113 ( 
.A(n_10060),
.Y(n_11113)
);

INVx1_ASAP7_75t_L g11114 ( 
.A(n_10062),
.Y(n_11114)
);

INVx1_ASAP7_75t_L g11115 ( 
.A(n_10062),
.Y(n_11115)
);

INVx3_ASAP7_75t_L g11116 ( 
.A(n_9996),
.Y(n_11116)
);

INVx2_ASAP7_75t_L g11117 ( 
.A(n_10045),
.Y(n_11117)
);

OAI21x1_ASAP7_75t_L g11118 ( 
.A1(n_9385),
.A2(n_8258),
.B(n_8237),
.Y(n_11118)
);

BUFx6f_ASAP7_75t_L g11119 ( 
.A(n_9033),
.Y(n_11119)
);

AOI22xp33_ASAP7_75t_L g11120 ( 
.A1(n_9412),
.A2(n_7700),
.B1(n_8532),
.B2(n_7792),
.Y(n_11120)
);

INVx2_ASAP7_75t_L g11121 ( 
.A(n_10045),
.Y(n_11121)
);

AO21x2_ASAP7_75t_L g11122 ( 
.A1(n_9418),
.A2(n_8486),
.B(n_8395),
.Y(n_11122)
);

INVx1_ASAP7_75t_L g11123 ( 
.A(n_10063),
.Y(n_11123)
);

INVx2_ASAP7_75t_L g11124 ( 
.A(n_10045),
.Y(n_11124)
);

INVx1_ASAP7_75t_L g11125 ( 
.A(n_10063),
.Y(n_11125)
);

HB1xp67_ASAP7_75t_L g11126 ( 
.A(n_10200),
.Y(n_11126)
);

INVx1_ASAP7_75t_L g11127 ( 
.A(n_10069),
.Y(n_11127)
);

INVx1_ASAP7_75t_L g11128 ( 
.A(n_10069),
.Y(n_11128)
);

INVx2_ASAP7_75t_L g11129 ( 
.A(n_10047),
.Y(n_11129)
);

BUFx4f_ASAP7_75t_L g11130 ( 
.A(n_9033),
.Y(n_11130)
);

INVx1_ASAP7_75t_L g11131 ( 
.A(n_10082),
.Y(n_11131)
);

INVx1_ASAP7_75t_L g11132 ( 
.A(n_10082),
.Y(n_11132)
);

INVx1_ASAP7_75t_L g11133 ( 
.A(n_10083),
.Y(n_11133)
);

OAI21x1_ASAP7_75t_L g11134 ( 
.A1(n_9385),
.A2(n_8258),
.B(n_8237),
.Y(n_11134)
);

CKINVDCx5p33_ASAP7_75t_R g11135 ( 
.A(n_9295),
.Y(n_11135)
);

INVx2_ASAP7_75t_L g11136 ( 
.A(n_10047),
.Y(n_11136)
);

AND2x2_ASAP7_75t_L g11137 ( 
.A(n_10202),
.B(n_7789),
.Y(n_11137)
);

INVx1_ASAP7_75t_L g11138 ( 
.A(n_10083),
.Y(n_11138)
);

INVx1_ASAP7_75t_L g11139 ( 
.A(n_10090),
.Y(n_11139)
);

INVx1_ASAP7_75t_L g11140 ( 
.A(n_10090),
.Y(n_11140)
);

AOI221x1_ASAP7_75t_L g11141 ( 
.A1(n_9021),
.A2(n_8310),
.B1(n_8859),
.B2(n_8368),
.C(n_8842),
.Y(n_11141)
);

OA21x2_ASAP7_75t_L g11142 ( 
.A1(n_9768),
.A2(n_8676),
.B(n_8675),
.Y(n_11142)
);

BUFx3_ASAP7_75t_L g11143 ( 
.A(n_9097),
.Y(n_11143)
);

INVx2_ASAP7_75t_L g11144 ( 
.A(n_10047),
.Y(n_11144)
);

AND2x2_ASAP7_75t_L g11145 ( 
.A(n_10231),
.B(n_7789),
.Y(n_11145)
);

INVx1_ASAP7_75t_L g11146 ( 
.A(n_10091),
.Y(n_11146)
);

INVxp67_ASAP7_75t_SL g11147 ( 
.A(n_9306),
.Y(n_11147)
);

INVx2_ASAP7_75t_L g11148 ( 
.A(n_10048),
.Y(n_11148)
);

OAI21x1_ASAP7_75t_SL g11149 ( 
.A1(n_9347),
.A2(n_8738),
.B(n_8371),
.Y(n_11149)
);

INVx1_ASAP7_75t_L g11150 ( 
.A(n_10091),
.Y(n_11150)
);

INVx1_ASAP7_75t_L g11151 ( 
.A(n_10092),
.Y(n_11151)
);

BUFx3_ASAP7_75t_L g11152 ( 
.A(n_9134),
.Y(n_11152)
);

OAI22xp5_ASAP7_75t_L g11153 ( 
.A1(n_8963),
.A2(n_8205),
.B1(n_8361),
.B2(n_8680),
.Y(n_11153)
);

INVx2_ASAP7_75t_L g11154 ( 
.A(n_10048),
.Y(n_11154)
);

INVx2_ASAP7_75t_L g11155 ( 
.A(n_10048),
.Y(n_11155)
);

INVx1_ASAP7_75t_L g11156 ( 
.A(n_10092),
.Y(n_11156)
);

AO21x2_ASAP7_75t_L g11157 ( 
.A1(n_9418),
.A2(n_9552),
.B(n_9486),
.Y(n_11157)
);

INVx2_ASAP7_75t_L g11158 ( 
.A(n_10049),
.Y(n_11158)
);

INVx1_ASAP7_75t_L g11159 ( 
.A(n_10093),
.Y(n_11159)
);

HB1xp67_ASAP7_75t_L g11160 ( 
.A(n_10219),
.Y(n_11160)
);

INVx2_ASAP7_75t_L g11161 ( 
.A(n_10049),
.Y(n_11161)
);

OAI21xp5_ASAP7_75t_L g11162 ( 
.A1(n_9412),
.A2(n_8272),
.B(n_7834),
.Y(n_11162)
);

INVx1_ASAP7_75t_L g11163 ( 
.A(n_10093),
.Y(n_11163)
);

AND2x2_ASAP7_75t_L g11164 ( 
.A(n_10231),
.B(n_7840),
.Y(n_11164)
);

AND2x2_ASAP7_75t_L g11165 ( 
.A(n_10238),
.B(n_7840),
.Y(n_11165)
);

INVx2_ASAP7_75t_L g11166 ( 
.A(n_10049),
.Y(n_11166)
);

BUFx2_ASAP7_75t_L g11167 ( 
.A(n_10289),
.Y(n_11167)
);

INVx2_ASAP7_75t_L g11168 ( 
.A(n_10054),
.Y(n_11168)
);

OAI21x1_ASAP7_75t_L g11169 ( 
.A1(n_9385),
.A2(n_8258),
.B(n_8237),
.Y(n_11169)
);

INVx1_ASAP7_75t_L g11170 ( 
.A(n_10094),
.Y(n_11170)
);

BUFx3_ASAP7_75t_L g11171 ( 
.A(n_9134),
.Y(n_11171)
);

INVx2_ASAP7_75t_L g11172 ( 
.A(n_10054),
.Y(n_11172)
);

OAI21x1_ASAP7_75t_L g11173 ( 
.A1(n_9549),
.A2(n_8262),
.B(n_8260),
.Y(n_11173)
);

AND2x2_ASAP7_75t_L g11174 ( 
.A(n_10238),
.B(n_7840),
.Y(n_11174)
);

INVx2_ASAP7_75t_L g11175 ( 
.A(n_10054),
.Y(n_11175)
);

INVx1_ASAP7_75t_L g11176 ( 
.A(n_10094),
.Y(n_11176)
);

INVx1_ASAP7_75t_L g11177 ( 
.A(n_10099),
.Y(n_11177)
);

INVx1_ASAP7_75t_L g11178 ( 
.A(n_10099),
.Y(n_11178)
);

AOI22xp33_ASAP7_75t_L g11179 ( 
.A1(n_9412),
.A2(n_7700),
.B1(n_8532),
.B2(n_7792),
.Y(n_11179)
);

BUFx6f_ASAP7_75t_L g11180 ( 
.A(n_9033),
.Y(n_11180)
);

INVx2_ASAP7_75t_L g11181 ( 
.A(n_10071),
.Y(n_11181)
);

BUFx12f_ASAP7_75t_L g11182 ( 
.A(n_9676),
.Y(n_11182)
);

INVx4_ASAP7_75t_L g11183 ( 
.A(n_9033),
.Y(n_11183)
);

INVx1_ASAP7_75t_L g11184 ( 
.A(n_10100),
.Y(n_11184)
);

INVx2_ASAP7_75t_L g11185 ( 
.A(n_10071),
.Y(n_11185)
);

OR2x2_ASAP7_75t_L g11186 ( 
.A(n_9789),
.B(n_8800),
.Y(n_11186)
);

AND2x2_ASAP7_75t_L g11187 ( 
.A(n_10284),
.B(n_7840),
.Y(n_11187)
);

INVx2_ASAP7_75t_L g11188 ( 
.A(n_10071),
.Y(n_11188)
);

INVx1_ASAP7_75t_L g11189 ( 
.A(n_10100),
.Y(n_11189)
);

INVx1_ASAP7_75t_L g11190 ( 
.A(n_10104),
.Y(n_11190)
);

OAI21x1_ASAP7_75t_L g11191 ( 
.A1(n_9549),
.A2(n_8262),
.B(n_8260),
.Y(n_11191)
);

INVx1_ASAP7_75t_L g11192 ( 
.A(n_10104),
.Y(n_11192)
);

INVx2_ASAP7_75t_L g11193 ( 
.A(n_10081),
.Y(n_11193)
);

AO21x2_ASAP7_75t_L g11194 ( 
.A1(n_9353),
.A2(n_9180),
.B(n_9347),
.Y(n_11194)
);

INVx1_ASAP7_75t_L g11195 ( 
.A(n_10108),
.Y(n_11195)
);

BUFx6f_ASAP7_75t_L g11196 ( 
.A(n_9033),
.Y(n_11196)
);

BUFx2_ASAP7_75t_L g11197 ( 
.A(n_10289),
.Y(n_11197)
);

INVx2_ASAP7_75t_L g11198 ( 
.A(n_10081),
.Y(n_11198)
);

INVx1_ASAP7_75t_L g11199 ( 
.A(n_10108),
.Y(n_11199)
);

INVx2_ASAP7_75t_L g11200 ( 
.A(n_10081),
.Y(n_11200)
);

NAND2x1_ASAP7_75t_L g11201 ( 
.A(n_9703),
.B(n_9810),
.Y(n_11201)
);

INVx1_ASAP7_75t_L g11202 ( 
.A(n_10109),
.Y(n_11202)
);

INVx1_ASAP7_75t_L g11203 ( 
.A(n_10109),
.Y(n_11203)
);

INVxp67_ASAP7_75t_L g11204 ( 
.A(n_10034),
.Y(n_11204)
);

INVx3_ASAP7_75t_L g11205 ( 
.A(n_10086),
.Y(n_11205)
);

INVx2_ASAP7_75t_L g11206 ( 
.A(n_10085),
.Y(n_11206)
);

NAND2x1p5_ASAP7_75t_L g11207 ( 
.A(n_9690),
.B(n_8641),
.Y(n_11207)
);

AND2x2_ASAP7_75t_L g11208 ( 
.A(n_10284),
.B(n_7840),
.Y(n_11208)
);

INVx2_ASAP7_75t_L g11209 ( 
.A(n_10085),
.Y(n_11209)
);

HB1xp67_ASAP7_75t_L g11210 ( 
.A(n_10223),
.Y(n_11210)
);

INVx2_ASAP7_75t_L g11211 ( 
.A(n_10085),
.Y(n_11211)
);

INVxp33_ASAP7_75t_SL g11212 ( 
.A(n_10125),
.Y(n_11212)
);

AOI22xp33_ASAP7_75t_L g11213 ( 
.A1(n_9129),
.A2(n_7792),
.B1(n_7895),
.B2(n_8524),
.Y(n_11213)
);

INVx2_ASAP7_75t_SL g11214 ( 
.A(n_9150),
.Y(n_11214)
);

INVx1_ASAP7_75t_L g11215 ( 
.A(n_10115),
.Y(n_11215)
);

NAND2xp5_ASAP7_75t_L g11216 ( 
.A(n_9165),
.B(n_8264),
.Y(n_11216)
);

INVx2_ASAP7_75t_L g11217 ( 
.A(n_10088),
.Y(n_11217)
);

INVx1_ASAP7_75t_L g11218 ( 
.A(n_10115),
.Y(n_11218)
);

AO21x1_ASAP7_75t_SL g11219 ( 
.A1(n_9324),
.A2(n_8722),
.B(n_8361),
.Y(n_11219)
);

INVx1_ASAP7_75t_L g11220 ( 
.A(n_10116),
.Y(n_11220)
);

NOR2xp33_ASAP7_75t_L g11221 ( 
.A(n_9066),
.B(n_8514),
.Y(n_11221)
);

INVx2_ASAP7_75t_L g11222 ( 
.A(n_10088),
.Y(n_11222)
);

BUFx2_ASAP7_75t_L g11223 ( 
.A(n_10289),
.Y(n_11223)
);

INVx1_ASAP7_75t_L g11224 ( 
.A(n_10116),
.Y(n_11224)
);

OR2x2_ASAP7_75t_L g11225 ( 
.A(n_9789),
.B(n_8800),
.Y(n_11225)
);

INVx3_ASAP7_75t_L g11226 ( 
.A(n_10086),
.Y(n_11226)
);

CKINVDCx5p33_ASAP7_75t_R g11227 ( 
.A(n_9295),
.Y(n_11227)
);

INVx1_ASAP7_75t_L g11228 ( 
.A(n_10117),
.Y(n_11228)
);

AOI21xp33_ASAP7_75t_L g11229 ( 
.A1(n_9845),
.A2(n_10033),
.B(n_9611),
.Y(n_11229)
);

INVx3_ASAP7_75t_L g11230 ( 
.A(n_10086),
.Y(n_11230)
);

INVx2_ASAP7_75t_L g11231 ( 
.A(n_10088),
.Y(n_11231)
);

INVx1_ASAP7_75t_L g11232 ( 
.A(n_10117),
.Y(n_11232)
);

HB1xp67_ASAP7_75t_L g11233 ( 
.A(n_10276),
.Y(n_11233)
);

INVx1_ASAP7_75t_L g11234 ( 
.A(n_10129),
.Y(n_11234)
);

CKINVDCx8_ASAP7_75t_R g11235 ( 
.A(n_9021),
.Y(n_11235)
);

BUFx3_ASAP7_75t_L g11236 ( 
.A(n_9134),
.Y(n_11236)
);

OR2x2_ASAP7_75t_L g11237 ( 
.A(n_9799),
.B(n_8817),
.Y(n_11237)
);

INVx2_ASAP7_75t_SL g11238 ( 
.A(n_9150),
.Y(n_11238)
);

OAI21x1_ASAP7_75t_L g11239 ( 
.A1(n_9972),
.A2(n_8262),
.B(n_8260),
.Y(n_11239)
);

HB1xp67_ASAP7_75t_L g11240 ( 
.A(n_10278),
.Y(n_11240)
);

INVx1_ASAP7_75t_L g11241 ( 
.A(n_10129),
.Y(n_11241)
);

OAI21x1_ASAP7_75t_L g11242 ( 
.A1(n_9972),
.A2(n_8267),
.B(n_7786),
.Y(n_11242)
);

AOI22xp33_ASAP7_75t_SL g11243 ( 
.A1(n_9638),
.A2(n_7842),
.B1(n_7843),
.B2(n_7841),
.Y(n_11243)
);

INVx2_ASAP7_75t_L g11244 ( 
.A(n_10096),
.Y(n_11244)
);

INVx2_ASAP7_75t_SL g11245 ( 
.A(n_9150),
.Y(n_11245)
);

OAI21x1_ASAP7_75t_L g11246 ( 
.A1(n_9972),
.A2(n_8267),
.B(n_7786),
.Y(n_11246)
);

INVx2_ASAP7_75t_L g11247 ( 
.A(n_10096),
.Y(n_11247)
);

HB1xp67_ASAP7_75t_SL g11248 ( 
.A(n_10034),
.Y(n_11248)
);

AO21x2_ASAP7_75t_L g11249 ( 
.A1(n_9353),
.A2(n_9180),
.B(n_9486),
.Y(n_11249)
);

INVx2_ASAP7_75t_L g11250 ( 
.A(n_10096),
.Y(n_11250)
);

INVx1_ASAP7_75t_SL g11251 ( 
.A(n_9741),
.Y(n_11251)
);

BUFx12f_ASAP7_75t_L g11252 ( 
.A(n_10036),
.Y(n_11252)
);

INVx1_ASAP7_75t_L g11253 ( 
.A(n_10133),
.Y(n_11253)
);

HB1xp67_ASAP7_75t_L g11254 ( 
.A(n_9690),
.Y(n_11254)
);

INVx1_ASAP7_75t_L g11255 ( 
.A(n_10133),
.Y(n_11255)
);

AOI21x1_ASAP7_75t_L g11256 ( 
.A1(n_9074),
.A2(n_8383),
.B(n_8338),
.Y(n_11256)
);

AND2x2_ASAP7_75t_L g11257 ( 
.A(n_10291),
.B(n_7860),
.Y(n_11257)
);

INVx2_ASAP7_75t_L g11258 ( 
.A(n_10102),
.Y(n_11258)
);

AND2x2_ASAP7_75t_L g11259 ( 
.A(n_10291),
.B(n_7860),
.Y(n_11259)
);

OAI21x1_ASAP7_75t_L g11260 ( 
.A1(n_9990),
.A2(n_8267),
.B(n_7786),
.Y(n_11260)
);

BUFx2_ASAP7_75t_L g11261 ( 
.A(n_9200),
.Y(n_11261)
);

INVx1_ASAP7_75t_L g11262 ( 
.A(n_10134),
.Y(n_11262)
);

INVx1_ASAP7_75t_L g11263 ( 
.A(n_10134),
.Y(n_11263)
);

INVx2_ASAP7_75t_L g11264 ( 
.A(n_10102),
.Y(n_11264)
);

INVx1_ASAP7_75t_L g11265 ( 
.A(n_10136),
.Y(n_11265)
);

OR2x6_ASAP7_75t_L g11266 ( 
.A(n_9210),
.B(n_7746),
.Y(n_11266)
);

INVx1_ASAP7_75t_L g11267 ( 
.A(n_10136),
.Y(n_11267)
);

BUFx2_ASAP7_75t_L g11268 ( 
.A(n_9200),
.Y(n_11268)
);

INVx1_ASAP7_75t_L g11269 ( 
.A(n_10137),
.Y(n_11269)
);

HB1xp67_ASAP7_75t_L g11270 ( 
.A(n_9780),
.Y(n_11270)
);

HB1xp67_ASAP7_75t_L g11271 ( 
.A(n_9780),
.Y(n_11271)
);

OR2x2_ASAP7_75t_L g11272 ( 
.A(n_9799),
.B(n_8817),
.Y(n_11272)
);

INVx1_ASAP7_75t_L g11273 ( 
.A(n_10137),
.Y(n_11273)
);

AND2x2_ASAP7_75t_L g11274 ( 
.A(n_10286),
.B(n_7860),
.Y(n_11274)
);

BUFx2_ASAP7_75t_L g11275 ( 
.A(n_9200),
.Y(n_11275)
);

INVx1_ASAP7_75t_L g11276 ( 
.A(n_10140),
.Y(n_11276)
);

INVx2_ASAP7_75t_L g11277 ( 
.A(n_10102),
.Y(n_11277)
);

INVx2_ASAP7_75t_L g11278 ( 
.A(n_10105),
.Y(n_11278)
);

INVx2_ASAP7_75t_SL g11279 ( 
.A(n_9571),
.Y(n_11279)
);

INVx2_ASAP7_75t_L g11280 ( 
.A(n_10105),
.Y(n_11280)
);

O2A1O1Ixp5_ASAP7_75t_L g11281 ( 
.A1(n_10014),
.A2(n_8699),
.B(n_8459),
.C(n_8338),
.Y(n_11281)
);

INVx2_ASAP7_75t_L g11282 ( 
.A(n_10105),
.Y(n_11282)
);

NAND2xp5_ASAP7_75t_L g11283 ( 
.A(n_9433),
.B(n_8882),
.Y(n_11283)
);

INVx1_ASAP7_75t_L g11284 ( 
.A(n_10140),
.Y(n_11284)
);

INVx2_ASAP7_75t_L g11285 ( 
.A(n_10106),
.Y(n_11285)
);

INVx2_ASAP7_75t_L g11286 ( 
.A(n_10106),
.Y(n_11286)
);

INVx2_ASAP7_75t_L g11287 ( 
.A(n_10106),
.Y(n_11287)
);

AO21x2_ASAP7_75t_L g11288 ( 
.A1(n_9552),
.A2(n_8076),
.B(n_8790),
.Y(n_11288)
);

AND2x2_ASAP7_75t_L g11289 ( 
.A(n_10286),
.B(n_7860),
.Y(n_11289)
);

INVx3_ASAP7_75t_L g11290 ( 
.A(n_10181),
.Y(n_11290)
);

INVx4_ASAP7_75t_L g11291 ( 
.A(n_9033),
.Y(n_11291)
);

OAI21x1_ASAP7_75t_SL g11292 ( 
.A1(n_9537),
.A2(n_9272),
.B(n_9074),
.Y(n_11292)
);

INVx3_ASAP7_75t_L g11293 ( 
.A(n_10181),
.Y(n_11293)
);

AND2x2_ASAP7_75t_L g11294 ( 
.A(n_9114),
.B(n_7860),
.Y(n_11294)
);

INVx2_ASAP7_75t_L g11295 ( 
.A(n_9865),
.Y(n_11295)
);

INVx1_ASAP7_75t_L g11296 ( 
.A(n_10143),
.Y(n_11296)
);

HB1xp67_ASAP7_75t_L g11297 ( 
.A(n_9949),
.Y(n_11297)
);

BUFx4f_ASAP7_75t_L g11298 ( 
.A(n_9086),
.Y(n_11298)
);

OAI21x1_ASAP7_75t_L g11299 ( 
.A1(n_9990),
.A2(n_8664),
.B(n_8293),
.Y(n_11299)
);

INVx2_ASAP7_75t_L g11300 ( 
.A(n_9865),
.Y(n_11300)
);

HB1xp67_ASAP7_75t_L g11301 ( 
.A(n_9949),
.Y(n_11301)
);

AND2x4_ASAP7_75t_L g11302 ( 
.A(n_10162),
.B(n_8579),
.Y(n_11302)
);

OAI22xp33_ASAP7_75t_L g11303 ( 
.A1(n_10146),
.A2(n_7668),
.B1(n_7754),
.B2(n_8943),
.Y(n_11303)
);

NAND2xp5_ASAP7_75t_L g11304 ( 
.A(n_9566),
.B(n_8882),
.Y(n_11304)
);

AOI21x1_ASAP7_75t_L g11305 ( 
.A1(n_9272),
.A2(n_8459),
.B(n_8887),
.Y(n_11305)
);

INVx1_ASAP7_75t_L g11306 ( 
.A(n_10143),
.Y(n_11306)
);

INVx1_ASAP7_75t_L g11307 ( 
.A(n_10145),
.Y(n_11307)
);

INVx2_ASAP7_75t_L g11308 ( 
.A(n_9876),
.Y(n_11308)
);

AND2x2_ASAP7_75t_L g11309 ( 
.A(n_9114),
.B(n_7898),
.Y(n_11309)
);

INVx2_ASAP7_75t_L g11310 ( 
.A(n_9876),
.Y(n_11310)
);

O2A1O1Ixp33_ASAP7_75t_SL g11311 ( 
.A1(n_9442),
.A2(n_8747),
.B(n_8455),
.C(n_8585),
.Y(n_11311)
);

INVx1_ASAP7_75t_L g11312 ( 
.A(n_10145),
.Y(n_11312)
);

INVx1_ASAP7_75t_L g11313 ( 
.A(n_10148),
.Y(n_11313)
);

NAND2xp5_ASAP7_75t_L g11314 ( 
.A(n_9566),
.B(n_7664),
.Y(n_11314)
);

OR2x2_ASAP7_75t_L g11315 ( 
.A(n_9856),
.B(n_8817),
.Y(n_11315)
);

INVx1_ASAP7_75t_L g11316 ( 
.A(n_10148),
.Y(n_11316)
);

INVx2_ASAP7_75t_L g11317 ( 
.A(n_9906),
.Y(n_11317)
);

AND2x4_ASAP7_75t_L g11318 ( 
.A(n_10162),
.B(n_8579),
.Y(n_11318)
);

INVxp67_ASAP7_75t_L g11319 ( 
.A(n_9210),
.Y(n_11319)
);

INVx2_ASAP7_75t_L g11320 ( 
.A(n_9906),
.Y(n_11320)
);

INVx1_ASAP7_75t_L g11321 ( 
.A(n_10152),
.Y(n_11321)
);

AND2x2_ASAP7_75t_L g11322 ( 
.A(n_9151),
.B(n_7898),
.Y(n_11322)
);

AOI21x1_ASAP7_75t_L g11323 ( 
.A1(n_10020),
.A2(n_8887),
.B(n_8004),
.Y(n_11323)
);

AND2x4_ASAP7_75t_L g11324 ( 
.A(n_10162),
.B(n_8579),
.Y(n_11324)
);

INVx4_ASAP7_75t_L g11325 ( 
.A(n_9086),
.Y(n_11325)
);

AOI22xp33_ASAP7_75t_L g11326 ( 
.A1(n_9129),
.A2(n_7895),
.B1(n_8524),
.B2(n_7754),
.Y(n_11326)
);

INVx1_ASAP7_75t_L g11327 ( 
.A(n_10152),
.Y(n_11327)
);

INVx1_ASAP7_75t_L g11328 ( 
.A(n_10153),
.Y(n_11328)
);

HB1xp67_ASAP7_75t_L g11329 ( 
.A(n_10013),
.Y(n_11329)
);

INVx1_ASAP7_75t_L g11330 ( 
.A(n_10153),
.Y(n_11330)
);

INVx3_ASAP7_75t_L g11331 ( 
.A(n_10181),
.Y(n_11331)
);

AOI21xp5_ASAP7_75t_L g11332 ( 
.A1(n_9225),
.A2(n_8624),
.B(n_8533),
.Y(n_11332)
);

INVx1_ASAP7_75t_L g11333 ( 
.A(n_10154),
.Y(n_11333)
);

INVx1_ASAP7_75t_L g11334 ( 
.A(n_10154),
.Y(n_11334)
);

OR2x6_ASAP7_75t_L g11335 ( 
.A(n_9730),
.B(n_7770),
.Y(n_11335)
);

INVx3_ASAP7_75t_L g11336 ( 
.A(n_10204),
.Y(n_11336)
);

INVx2_ASAP7_75t_L g11337 ( 
.A(n_9908),
.Y(n_11337)
);

AND2x2_ASAP7_75t_L g11338 ( 
.A(n_9151),
.B(n_7898),
.Y(n_11338)
);

INVx2_ASAP7_75t_L g11339 ( 
.A(n_9908),
.Y(n_11339)
);

INVx2_ASAP7_75t_L g11340 ( 
.A(n_9616),
.Y(n_11340)
);

OR2x2_ASAP7_75t_L g11341 ( 
.A(n_9856),
.B(n_8818),
.Y(n_11341)
);

INVx1_ASAP7_75t_L g11342 ( 
.A(n_10158),
.Y(n_11342)
);

INVx2_ASAP7_75t_L g11343 ( 
.A(n_9616),
.Y(n_11343)
);

AOI222xp33_ASAP7_75t_L g11344 ( 
.A1(n_9835),
.A2(n_9225),
.B1(n_10250),
.B2(n_9492),
.C1(n_9563),
.C2(n_9046),
.Y(n_11344)
);

INVx1_ASAP7_75t_L g11345 ( 
.A(n_10158),
.Y(n_11345)
);

INVx1_ASAP7_75t_L g11346 ( 
.A(n_10189),
.Y(n_11346)
);

INVx2_ASAP7_75t_SL g11347 ( 
.A(n_9571),
.Y(n_11347)
);

INVx1_ASAP7_75t_L g11348 ( 
.A(n_10189),
.Y(n_11348)
);

AND2x2_ASAP7_75t_L g11349 ( 
.A(n_9204),
.B(n_7898),
.Y(n_11349)
);

INVx1_ASAP7_75t_L g11350 ( 
.A(n_10195),
.Y(n_11350)
);

HB1xp67_ASAP7_75t_L g11351 ( 
.A(n_10016),
.Y(n_11351)
);

INVx1_ASAP7_75t_L g11352 ( 
.A(n_10195),
.Y(n_11352)
);

INVx1_ASAP7_75t_L g11353 ( 
.A(n_10210),
.Y(n_11353)
);

INVx1_ASAP7_75t_L g11354 ( 
.A(n_10210),
.Y(n_11354)
);

HB1xp67_ASAP7_75t_L g11355 ( 
.A(n_10016),
.Y(n_11355)
);

INVx2_ASAP7_75t_L g11356 ( 
.A(n_9617),
.Y(n_11356)
);

BUFx2_ASAP7_75t_SL g11357 ( 
.A(n_9134),
.Y(n_11357)
);

OAI21x1_ASAP7_75t_L g11358 ( 
.A1(n_9990),
.A2(n_8664),
.B(n_8293),
.Y(n_11358)
);

AND2x2_ASAP7_75t_L g11359 ( 
.A(n_9204),
.B(n_7898),
.Y(n_11359)
);

BUFx2_ASAP7_75t_SL g11360 ( 
.A(n_8965),
.Y(n_11360)
);

INVx2_ASAP7_75t_SL g11361 ( 
.A(n_9664),
.Y(n_11361)
);

BUFx6f_ASAP7_75t_L g11362 ( 
.A(n_9086),
.Y(n_11362)
);

INVx3_ASAP7_75t_L g11363 ( 
.A(n_10204),
.Y(n_11363)
);

INVx1_ASAP7_75t_L g11364 ( 
.A(n_10211),
.Y(n_11364)
);

BUFx2_ASAP7_75t_SL g11365 ( 
.A(n_9167),
.Y(n_11365)
);

INVx1_ASAP7_75t_L g11366 ( 
.A(n_10211),
.Y(n_11366)
);

INVxp67_ASAP7_75t_SL g11367 ( 
.A(n_8986),
.Y(n_11367)
);

BUFx2_ASAP7_75t_L g11368 ( 
.A(n_9223),
.Y(n_11368)
);

NAND2xp5_ASAP7_75t_L g11369 ( 
.A(n_9569),
.B(n_7664),
.Y(n_11369)
);

INVx5_ASAP7_75t_L g11370 ( 
.A(n_9086),
.Y(n_11370)
);

INVx1_ASAP7_75t_L g11371 ( 
.A(n_10214),
.Y(n_11371)
);

INVx1_ASAP7_75t_L g11372 ( 
.A(n_10214),
.Y(n_11372)
);

OAI21x1_ASAP7_75t_L g11373 ( 
.A1(n_10002),
.A2(n_8664),
.B(n_8293),
.Y(n_11373)
);

AO21x2_ASAP7_75t_L g11374 ( 
.A1(n_9353),
.A2(n_9145),
.B(n_9037),
.Y(n_11374)
);

INVx2_ASAP7_75t_L g11375 ( 
.A(n_9617),
.Y(n_11375)
);

INVx2_ASAP7_75t_L g11376 ( 
.A(n_9698),
.Y(n_11376)
);

INVx2_ASAP7_75t_L g11377 ( 
.A(n_9698),
.Y(n_11377)
);

INVx3_ASAP7_75t_L g11378 ( 
.A(n_10204),
.Y(n_11378)
);

INVx1_ASAP7_75t_L g11379 ( 
.A(n_10216),
.Y(n_11379)
);

INVx2_ASAP7_75t_L g11380 ( 
.A(n_9705),
.Y(n_11380)
);

OAI21xp5_ASAP7_75t_L g11381 ( 
.A1(n_10147),
.A2(n_7668),
.B(n_7884),
.Y(n_11381)
);

INVx1_ASAP7_75t_SL g11382 ( 
.A(n_9915),
.Y(n_11382)
);

INVxp67_ASAP7_75t_L g11383 ( 
.A(n_9730),
.Y(n_11383)
);

INVx1_ASAP7_75t_L g11384 ( 
.A(n_10216),
.Y(n_11384)
);

INVx1_ASAP7_75t_L g11385 ( 
.A(n_10218),
.Y(n_11385)
);

INVx1_ASAP7_75t_L g11386 ( 
.A(n_10218),
.Y(n_11386)
);

HB1xp67_ASAP7_75t_L g11387 ( 
.A(n_10013),
.Y(n_11387)
);

INVx1_ASAP7_75t_L g11388 ( 
.A(n_10220),
.Y(n_11388)
);

INVx1_ASAP7_75t_L g11389 ( 
.A(n_10220),
.Y(n_11389)
);

INVx1_ASAP7_75t_L g11390 ( 
.A(n_10228),
.Y(n_11390)
);

AOI21x1_ASAP7_75t_L g11391 ( 
.A1(n_10020),
.A2(n_8887),
.B(n_8004),
.Y(n_11391)
);

HB1xp67_ASAP7_75t_L g11392 ( 
.A(n_10132),
.Y(n_11392)
);

AND2x2_ASAP7_75t_L g11393 ( 
.A(n_9216),
.B(n_9228),
.Y(n_11393)
);

INVx2_ASAP7_75t_L g11394 ( 
.A(n_9705),
.Y(n_11394)
);

INVx2_ASAP7_75t_L g11395 ( 
.A(n_9812),
.Y(n_11395)
);

BUFx2_ASAP7_75t_L g11396 ( 
.A(n_9223),
.Y(n_11396)
);

OAI21x1_ASAP7_75t_L g11397 ( 
.A1(n_10002),
.A2(n_9218),
.B(n_9768),
.Y(n_11397)
);

AND2x4_ASAP7_75t_L g11398 ( 
.A(n_10162),
.B(n_8791),
.Y(n_11398)
);

CKINVDCx5p33_ASAP7_75t_R g11399 ( 
.A(n_9649),
.Y(n_11399)
);

BUFx3_ASAP7_75t_L g11400 ( 
.A(n_9993),
.Y(n_11400)
);

INVx2_ASAP7_75t_L g11401 ( 
.A(n_9812),
.Y(n_11401)
);

INVx2_ASAP7_75t_L g11402 ( 
.A(n_9886),
.Y(n_11402)
);

INVx1_ASAP7_75t_L g11403 ( 
.A(n_10228),
.Y(n_11403)
);

INVx1_ASAP7_75t_L g11404 ( 
.A(n_10229),
.Y(n_11404)
);

INVx2_ASAP7_75t_L g11405 ( 
.A(n_9886),
.Y(n_11405)
);

INVx2_ASAP7_75t_L g11406 ( 
.A(n_9987),
.Y(n_11406)
);

OR2x2_ASAP7_75t_L g11407 ( 
.A(n_9657),
.B(n_8818),
.Y(n_11407)
);

AND2x2_ASAP7_75t_L g11408 ( 
.A(n_9216),
.B(n_9228),
.Y(n_11408)
);

INVx1_ASAP7_75t_L g11409 ( 
.A(n_10229),
.Y(n_11409)
);

INVx1_ASAP7_75t_L g11410 ( 
.A(n_10230),
.Y(n_11410)
);

OAI21x1_ASAP7_75t_L g11411 ( 
.A1(n_10002),
.A2(n_8280),
.B(n_8080),
.Y(n_11411)
);

INVx1_ASAP7_75t_L g11412 ( 
.A(n_10230),
.Y(n_11412)
);

INVx1_ASAP7_75t_L g11413 ( 
.A(n_10236),
.Y(n_11413)
);

AND2x4_ASAP7_75t_L g11414 ( 
.A(n_10162),
.B(n_8791),
.Y(n_11414)
);

INVx2_ASAP7_75t_L g11415 ( 
.A(n_9987),
.Y(n_11415)
);

HB1xp67_ASAP7_75t_L g11416 ( 
.A(n_10132),
.Y(n_11416)
);

INVx1_ASAP7_75t_L g11417 ( 
.A(n_10236),
.Y(n_11417)
);

INVx1_ASAP7_75t_L g11418 ( 
.A(n_10240),
.Y(n_11418)
);

HB1xp67_ASAP7_75t_L g11419 ( 
.A(n_10188),
.Y(n_11419)
);

INVx2_ASAP7_75t_L g11420 ( 
.A(n_9992),
.Y(n_11420)
);

AND2x2_ASAP7_75t_L g11421 ( 
.A(n_9301),
.B(n_7916),
.Y(n_11421)
);

NAND2xp5_ASAP7_75t_L g11422 ( 
.A(n_9569),
.B(n_7689),
.Y(n_11422)
);

BUFx2_ASAP7_75t_L g11423 ( 
.A(n_9223),
.Y(n_11423)
);

INVx2_ASAP7_75t_L g11424 ( 
.A(n_9992),
.Y(n_11424)
);

INVx2_ASAP7_75t_L g11425 ( 
.A(n_10018),
.Y(n_11425)
);

INVx2_ASAP7_75t_L g11426 ( 
.A(n_10018),
.Y(n_11426)
);

OR2x2_ASAP7_75t_L g11427 ( 
.A(n_9657),
.B(n_8818),
.Y(n_11427)
);

OR2x2_ASAP7_75t_L g11428 ( 
.A(n_9691),
.B(n_8868),
.Y(n_11428)
);

INVx2_ASAP7_75t_L g11429 ( 
.A(n_10029),
.Y(n_11429)
);

INVx1_ASAP7_75t_L g11430 ( 
.A(n_10240),
.Y(n_11430)
);

BUFx2_ASAP7_75t_L g11431 ( 
.A(n_8998),
.Y(n_11431)
);

INVx2_ASAP7_75t_L g11432 ( 
.A(n_10029),
.Y(n_11432)
);

BUFx3_ASAP7_75t_L g11433 ( 
.A(n_9993),
.Y(n_11433)
);

NAND2xp5_ASAP7_75t_L g11434 ( 
.A(n_10250),
.B(n_7689),
.Y(n_11434)
);

OAI22xp33_ASAP7_75t_L g11435 ( 
.A1(n_9003),
.A2(n_8943),
.B1(n_8473),
.B2(n_8660),
.Y(n_11435)
);

INVx1_ASAP7_75t_L g11436 ( 
.A(n_10243),
.Y(n_11436)
);

BUFx3_ASAP7_75t_L g11437 ( 
.A(n_9993),
.Y(n_11437)
);

CKINVDCx20_ASAP7_75t_R g11438 ( 
.A(n_9288),
.Y(n_11438)
);

BUFx2_ASAP7_75t_L g11439 ( 
.A(n_8998),
.Y(n_11439)
);

INVx2_ASAP7_75t_L g11440 ( 
.A(n_10061),
.Y(n_11440)
);

INVx2_ASAP7_75t_L g11441 ( 
.A(n_10061),
.Y(n_11441)
);

AOI21xp5_ASAP7_75t_L g11442 ( 
.A1(n_10293),
.A2(n_9193),
.B(n_9835),
.Y(n_11442)
);

INVx1_ASAP7_75t_L g11443 ( 
.A(n_10890),
.Y(n_11443)
);

AOI22xp33_ASAP7_75t_L g11444 ( 
.A1(n_10363),
.A2(n_9963),
.B1(n_10191),
.B2(n_9564),
.Y(n_11444)
);

AND2x2_ASAP7_75t_L g11445 ( 
.A(n_10806),
.B(n_9289),
.Y(n_11445)
);

AND2x2_ASAP7_75t_L g11446 ( 
.A(n_10806),
.B(n_9289),
.Y(n_11446)
);

NOR2xp33_ASAP7_75t_SL g11447 ( 
.A(n_10414),
.B(n_8182),
.Y(n_11447)
);

HB1xp67_ASAP7_75t_L g11448 ( 
.A(n_10294),
.Y(n_11448)
);

AOI22xp33_ASAP7_75t_L g11449 ( 
.A1(n_10365),
.A2(n_9963),
.B1(n_10191),
.B2(n_9564),
.Y(n_11449)
);

HB1xp67_ASAP7_75t_L g11450 ( 
.A(n_10300),
.Y(n_11450)
);

INVx5_ASAP7_75t_L g11451 ( 
.A(n_10481),
.Y(n_11451)
);

AND2x2_ASAP7_75t_L g11452 ( 
.A(n_11008),
.B(n_9316),
.Y(n_11452)
);

OAI21xp5_ASAP7_75t_L g11453 ( 
.A1(n_10889),
.A2(n_10014),
.B(n_10241),
.Y(n_11453)
);

NAND3xp33_ASAP7_75t_L g11454 ( 
.A(n_10309),
.B(n_10239),
.C(n_9563),
.Y(n_11454)
);

AND2x2_ASAP7_75t_L g11455 ( 
.A(n_11008),
.B(n_9316),
.Y(n_11455)
);

BUFx6f_ASAP7_75t_SL g11456 ( 
.A(n_10307),
.Y(n_11456)
);

BUFx10_ASAP7_75t_L g11457 ( 
.A(n_11399),
.Y(n_11457)
);

INVx3_ASAP7_75t_L g11458 ( 
.A(n_11252),
.Y(n_11458)
);

NAND2xp5_ASAP7_75t_L g11459 ( 
.A(n_10441),
.B(n_9290),
.Y(n_11459)
);

BUFx4f_ASAP7_75t_L g11460 ( 
.A(n_10481),
.Y(n_11460)
);

OAI211xp5_ASAP7_75t_L g11461 ( 
.A1(n_10309),
.A2(n_10257),
.B(n_9793),
.C(n_10239),
.Y(n_11461)
);

AOI211xp5_ASAP7_75t_L g11462 ( 
.A1(n_11229),
.A2(n_9933),
.B(n_9711),
.C(n_9455),
.Y(n_11462)
);

OAI22xp33_ASAP7_75t_L g11463 ( 
.A1(n_10397),
.A2(n_9455),
.B1(n_9003),
.B2(n_8975),
.Y(n_11463)
);

AOI22xp33_ASAP7_75t_L g11464 ( 
.A1(n_10942),
.A2(n_9008),
.B1(n_9042),
.B2(n_9597),
.Y(n_11464)
);

INVx1_ASAP7_75t_L g11465 ( 
.A(n_10892),
.Y(n_11465)
);

INVx1_ASAP7_75t_L g11466 ( 
.A(n_10895),
.Y(n_11466)
);

O2A1O1Ixp33_ASAP7_75t_L g11467 ( 
.A1(n_10533),
.A2(n_9316),
.B(n_9933),
.C(n_9212),
.Y(n_11467)
);

AOI22xp33_ASAP7_75t_SL g11468 ( 
.A1(n_10997),
.A2(n_9492),
.B1(n_9740),
.B2(n_9132),
.Y(n_11468)
);

AOI22xp33_ASAP7_75t_L g11469 ( 
.A1(n_10942),
.A2(n_9678),
.B1(n_9597),
.B2(n_9073),
.Y(n_11469)
);

NAND2xp5_ASAP7_75t_SL g11470 ( 
.A(n_10468),
.B(n_9510),
.Y(n_11470)
);

AOI22xp33_ASAP7_75t_L g11471 ( 
.A1(n_10888),
.A2(n_11013),
.B1(n_10613),
.B2(n_10396),
.Y(n_11471)
);

OAI211xp5_ASAP7_75t_L g11472 ( 
.A1(n_10796),
.A2(n_10257),
.B(n_9793),
.C(n_9158),
.Y(n_11472)
);

OAI21xp33_ASAP7_75t_SL g11473 ( 
.A1(n_11344),
.A2(n_9187),
.B(n_9143),
.Y(n_11473)
);

HB1xp67_ASAP7_75t_L g11474 ( 
.A(n_11254),
.Y(n_11474)
);

OAI22xp33_ASAP7_75t_L g11475 ( 
.A1(n_10526),
.A2(n_8975),
.B1(n_8989),
.B2(n_9500),
.Y(n_11475)
);

OAI211xp5_ASAP7_75t_L g11476 ( 
.A1(n_10299),
.A2(n_9500),
.B(n_10032),
.C(n_9848),
.Y(n_11476)
);

NAND4xp25_ASAP7_75t_SL g11477 ( 
.A(n_10419),
.B(n_8969),
.C(n_8719),
.D(n_9371),
.Y(n_11477)
);

AND2x2_ASAP7_75t_L g11478 ( 
.A(n_10474),
.B(n_9277),
.Y(n_11478)
);

INVx1_ASAP7_75t_L g11479 ( 
.A(n_10896),
.Y(n_11479)
);

HB1xp67_ASAP7_75t_L g11480 ( 
.A(n_11270),
.Y(n_11480)
);

AOI221xp5_ASAP7_75t_L g11481 ( 
.A1(n_10847),
.A2(n_9578),
.B1(n_9179),
.B2(n_9201),
.C(n_9966),
.Y(n_11481)
);

AOI22xp33_ASAP7_75t_L g11482 ( 
.A1(n_10888),
.A2(n_9678),
.B1(n_9597),
.B2(n_9544),
.Y(n_11482)
);

OAI221xp5_ASAP7_75t_L g11483 ( 
.A1(n_10881),
.A2(n_9463),
.B1(n_9371),
.B2(n_9443),
.C(n_9386),
.Y(n_11483)
);

NAND2xp33_ASAP7_75t_R g11484 ( 
.A(n_10414),
.B(n_9803),
.Y(n_11484)
);

AOI22xp33_ASAP7_75t_L g11485 ( 
.A1(n_10646),
.A2(n_9678),
.B1(n_9597),
.B2(n_9544),
.Y(n_11485)
);

AOI22xp33_ASAP7_75t_L g11486 ( 
.A1(n_10648),
.A2(n_9678),
.B1(n_9597),
.B2(n_9544),
.Y(n_11486)
);

AOI21xp33_ASAP7_75t_L g11487 ( 
.A1(n_10386),
.A2(n_9678),
.B(n_9544),
.Y(n_11487)
);

AOI21x1_ASAP7_75t_L g11488 ( 
.A1(n_10422),
.A2(n_9372),
.B(n_10126),
.Y(n_11488)
);

NAND2xp5_ASAP7_75t_L g11489 ( 
.A(n_10441),
.B(n_9290),
.Y(n_11489)
);

AOI22xp33_ASAP7_75t_L g11490 ( 
.A1(n_10648),
.A2(n_9544),
.B1(n_9740),
.B2(n_9881),
.Y(n_11490)
);

INVx1_ASAP7_75t_L g11491 ( 
.A(n_10897),
.Y(n_11491)
);

BUFx2_ASAP7_75t_L g11492 ( 
.A(n_11252),
.Y(n_11492)
);

AOI22xp33_ASAP7_75t_SL g11493 ( 
.A1(n_10860),
.A2(n_9132),
.B1(n_9067),
.B2(n_9212),
.Y(n_11493)
);

AOI22xp33_ASAP7_75t_L g11494 ( 
.A1(n_10475),
.A2(n_10852),
.B1(n_10893),
.B2(n_11219),
.Y(n_11494)
);

OAI22xp5_ASAP7_75t_L g11495 ( 
.A1(n_10889),
.A2(n_9341),
.B1(n_9294),
.B2(n_8989),
.Y(n_11495)
);

AOI221xp5_ASAP7_75t_L g11496 ( 
.A1(n_10847),
.A2(n_9179),
.B1(n_9966),
.B2(n_9912),
.C(n_9907),
.Y(n_11496)
);

OR2x2_ASAP7_75t_L g11497 ( 
.A(n_10866),
.B(n_9691),
.Y(n_11497)
);

BUFx8_ASAP7_75t_SL g11498 ( 
.A(n_11135),
.Y(n_11498)
);

INVx2_ASAP7_75t_L g11499 ( 
.A(n_11400),
.Y(n_11499)
);

AOI221xp5_ASAP7_75t_L g11500 ( 
.A1(n_10475),
.A2(n_9912),
.B1(n_9907),
.B2(n_8981),
.C(n_10121),
.Y(n_11500)
);

OAI22xp5_ASAP7_75t_L g11501 ( 
.A1(n_11248),
.A2(n_9341),
.B1(n_9111),
.B2(n_10050),
.Y(n_11501)
);

OAI22xp5_ASAP7_75t_L g11502 ( 
.A1(n_10840),
.A2(n_10050),
.B1(n_9602),
.B2(n_9292),
.Y(n_11502)
);

CKINVDCx6p67_ASAP7_75t_R g11503 ( 
.A(n_10382),
.Y(n_11503)
);

AOI22xp33_ASAP7_75t_L g11504 ( 
.A1(n_10757),
.A2(n_9881),
.B1(n_9261),
.B2(n_9271),
.Y(n_11504)
);

A2O1A1Ixp33_ASAP7_75t_L g11505 ( 
.A1(n_10992),
.A2(n_10983),
.B(n_11281),
.C(n_10323),
.Y(n_11505)
);

AOI22xp5_ASAP7_75t_L g11506 ( 
.A1(n_10937),
.A2(n_9888),
.B1(n_9081),
.B2(n_9067),
.Y(n_11506)
);

OAI22xp5_ASAP7_75t_L g11507 ( 
.A1(n_10686),
.A2(n_9602),
.B1(n_9307),
.B2(n_9834),
.Y(n_11507)
);

AOI22xp33_ASAP7_75t_L g11508 ( 
.A1(n_10686),
.A2(n_9261),
.B1(n_10120),
.B2(n_9090),
.Y(n_11508)
);

AOI22xp33_ASAP7_75t_L g11509 ( 
.A1(n_10692),
.A2(n_11326),
.B1(n_10499),
.B2(n_11075),
.Y(n_11509)
);

AND2x2_ASAP7_75t_L g11510 ( 
.A(n_10474),
.B(n_9277),
.Y(n_11510)
);

AOI222xp33_ASAP7_75t_L g11511 ( 
.A1(n_10305),
.A2(n_10024),
.B1(n_9921),
.B2(n_9887),
.C1(n_9302),
.C2(n_9193),
.Y(n_11511)
);

AOI21xp5_ASAP7_75t_L g11512 ( 
.A1(n_11311),
.A2(n_11075),
.B(n_11212),
.Y(n_11512)
);

INVx1_ASAP7_75t_L g11513 ( 
.A(n_10908),
.Y(n_11513)
);

BUFx2_ASAP7_75t_L g11514 ( 
.A(n_10875),
.Y(n_11514)
);

OAI22xp33_ASAP7_75t_L g11515 ( 
.A1(n_10931),
.A2(n_9834),
.B1(n_9238),
.B2(n_9249),
.Y(n_11515)
);

AO21x2_ASAP7_75t_L g11516 ( 
.A1(n_11147),
.A2(n_9255),
.B(n_10107),
.Y(n_11516)
);

OAI22xp33_ASAP7_75t_L g11517 ( 
.A1(n_11141),
.A2(n_10795),
.B1(n_10828),
.B2(n_11283),
.Y(n_11517)
);

AOI221xp5_ASAP7_75t_SL g11518 ( 
.A1(n_11303),
.A2(n_9076),
.B1(n_9384),
.B2(n_10121),
.C(n_9408),
.Y(n_11518)
);

AND2x2_ASAP7_75t_L g11519 ( 
.A(n_10749),
.B(n_8998),
.Y(n_11519)
);

OR2x2_ASAP7_75t_L g11520 ( 
.A(n_10417),
.B(n_9692),
.Y(n_11520)
);

AND2x2_ASAP7_75t_L g11521 ( 
.A(n_10749),
.B(n_8998),
.Y(n_11521)
);

INVx1_ASAP7_75t_L g11522 ( 
.A(n_10909),
.Y(n_11522)
);

BUFx6f_ASAP7_75t_L g11523 ( 
.A(n_10382),
.Y(n_11523)
);

NAND2xp5_ASAP7_75t_SL g11524 ( 
.A(n_11212),
.B(n_9510),
.Y(n_11524)
);

AOI221xp5_ASAP7_75t_L g11525 ( 
.A1(n_10794),
.A2(n_10064),
.B1(n_10073),
.B2(n_9214),
.C(n_9268),
.Y(n_11525)
);

AOI221xp5_ASAP7_75t_L g11526 ( 
.A1(n_10794),
.A2(n_10073),
.B1(n_10064),
.B2(n_9213),
.C(n_9248),
.Y(n_11526)
);

AOI222xp33_ASAP7_75t_L g11527 ( 
.A1(n_10311),
.A2(n_10024),
.B1(n_9921),
.B2(n_9887),
.C1(n_9332),
.C2(n_9358),
.Y(n_11527)
);

INVx1_ASAP7_75t_L g11528 ( 
.A(n_10910),
.Y(n_11528)
);

HB1xp67_ASAP7_75t_L g11529 ( 
.A(n_11271),
.Y(n_11529)
);

OAI22xp5_ASAP7_75t_L g11530 ( 
.A1(n_10692),
.A2(n_9087),
.B1(n_10032),
.B2(n_9122),
.Y(n_11530)
);

AOI221xp5_ASAP7_75t_L g11531 ( 
.A1(n_10737),
.A2(n_9248),
.B1(n_9384),
.B2(n_10101),
.C(n_10072),
.Y(n_11531)
);

AOI22xp5_ASAP7_75t_L g11532 ( 
.A1(n_10937),
.A2(n_9888),
.B1(n_9081),
.B2(n_9942),
.Y(n_11532)
);

AND2x2_ASAP7_75t_L g11533 ( 
.A(n_10725),
.B(n_9325),
.Y(n_11533)
);

AND2x4_ASAP7_75t_L g11534 ( 
.A(n_10708),
.B(n_10327),
.Y(n_11534)
);

INVx1_ASAP7_75t_L g11535 ( 
.A(n_10913),
.Y(n_11535)
);

AOI22xp33_ASAP7_75t_SL g11536 ( 
.A1(n_10386),
.A2(n_9332),
.B1(n_9358),
.B2(n_7843),
.Y(n_11536)
);

OR2x2_ASAP7_75t_L g11537 ( 
.A(n_10359),
.B(n_9692),
.Y(n_11537)
);

AOI22xp33_ASAP7_75t_L g11538 ( 
.A1(n_11326),
.A2(n_9090),
.B1(n_8969),
.B2(n_9239),
.Y(n_11538)
);

AOI221xp5_ASAP7_75t_L g11539 ( 
.A1(n_10737),
.A2(n_10101),
.B1(n_10072),
.B2(n_10177),
.C(n_9541),
.Y(n_11539)
);

INVx2_ASAP7_75t_L g11540 ( 
.A(n_11400),
.Y(n_11540)
);

AND2x2_ASAP7_75t_L g11541 ( 
.A(n_10725),
.B(n_9325),
.Y(n_11541)
);

AOI22xp33_ASAP7_75t_L g11542 ( 
.A1(n_11069),
.A2(n_9239),
.B1(n_9697),
.B2(n_10233),
.Y(n_11542)
);

AND2x2_ASAP7_75t_L g11543 ( 
.A(n_10821),
.B(n_9325),
.Y(n_11543)
);

BUFx2_ASAP7_75t_L g11544 ( 
.A(n_10875),
.Y(n_11544)
);

OAI21x1_ASAP7_75t_L g11545 ( 
.A1(n_11043),
.A2(n_8990),
.B(n_8986),
.Y(n_11545)
);

HB1xp67_ASAP7_75t_L g11546 ( 
.A(n_11297),
.Y(n_11546)
);

INVx1_ASAP7_75t_L g11547 ( 
.A(n_10918),
.Y(n_11547)
);

AOI21xp33_ASAP7_75t_SL g11548 ( 
.A1(n_10321),
.A2(n_10490),
.B(n_10448),
.Y(n_11548)
);

INVx2_ASAP7_75t_L g11549 ( 
.A(n_11433),
.Y(n_11549)
);

HB1xp67_ASAP7_75t_L g11550 ( 
.A(n_11301),
.Y(n_11550)
);

OAI21xp5_ASAP7_75t_L g11551 ( 
.A1(n_11069),
.A2(n_9804),
.B(n_10177),
.Y(n_11551)
);

AOI22xp33_ASAP7_75t_L g11552 ( 
.A1(n_11162),
.A2(n_9625),
.B1(n_9717),
.B2(n_9829),
.Y(n_11552)
);

AOI22xp33_ASAP7_75t_L g11553 ( 
.A1(n_11073),
.A2(n_8959),
.B1(n_9206),
.B2(n_9044),
.Y(n_11553)
);

AOI22xp33_ASAP7_75t_L g11554 ( 
.A1(n_11153),
.A2(n_8959),
.B1(n_9206),
.B2(n_9044),
.Y(n_11554)
);

AOI22xp33_ASAP7_75t_L g11555 ( 
.A1(n_11213),
.A2(n_8959),
.B1(n_9206),
.B2(n_9044),
.Y(n_11555)
);

INVx1_ASAP7_75t_L g11556 ( 
.A(n_10919),
.Y(n_11556)
);

INVx1_ASAP7_75t_L g11557 ( 
.A(n_10922),
.Y(n_11557)
);

OAI211xp5_ASAP7_75t_L g11558 ( 
.A1(n_11213),
.A2(n_9471),
.B(n_9639),
.C(n_9511),
.Y(n_11558)
);

AOI222xp33_ASAP7_75t_L g11559 ( 
.A1(n_10808),
.A2(n_9305),
.B1(n_9328),
.B2(n_9249),
.C1(n_9238),
.C2(n_8948),
.Y(n_11559)
);

AOI22xp33_ASAP7_75t_SL g11560 ( 
.A1(n_10343),
.A2(n_7843),
.B1(n_9328),
.B2(n_9305),
.Y(n_11560)
);

AOI221xp5_ASAP7_75t_SL g11561 ( 
.A1(n_11435),
.A2(n_9934),
.B1(n_8473),
.B2(n_7669),
.C(n_7608),
.Y(n_11561)
);

OAI221xp5_ASAP7_75t_L g11562 ( 
.A1(n_10719),
.A2(n_9743),
.B1(n_9726),
.B2(n_9359),
.C(n_9680),
.Y(n_11562)
);

NAND2xp5_ASAP7_75t_L g11563 ( 
.A(n_11434),
.B(n_10581),
.Y(n_11563)
);

OAI21xp5_ASAP7_75t_L g11564 ( 
.A1(n_11120),
.A2(n_9545),
.B(n_10144),
.Y(n_11564)
);

OAI211xp5_ASAP7_75t_L g11565 ( 
.A1(n_11120),
.A2(n_11179),
.B(n_11243),
.C(n_10688),
.Y(n_11565)
);

AOI22xp33_ASAP7_75t_L g11566 ( 
.A1(n_10324),
.A2(n_8959),
.B1(n_9206),
.B2(n_9044),
.Y(n_11566)
);

INVx1_ASAP7_75t_L g11567 ( 
.A(n_10923),
.Y(n_11567)
);

OAI22x1_ASAP7_75t_L g11568 ( 
.A1(n_10343),
.A2(n_9537),
.B1(n_9068),
.B2(n_9115),
.Y(n_11568)
);

AND2x2_ASAP7_75t_SL g11569 ( 
.A(n_10752),
.B(n_9510),
.Y(n_11569)
);

AOI22xp33_ASAP7_75t_L g11570 ( 
.A1(n_10718),
.A2(n_9044),
.B1(n_9275),
.B2(n_9206),
.Y(n_11570)
);

OAI22xp5_ASAP7_75t_L g11571 ( 
.A1(n_11235),
.A2(n_9279),
.B1(n_9331),
.B2(n_9493),
.Y(n_11571)
);

OAI22xp33_ASAP7_75t_L g11572 ( 
.A1(n_11304),
.A2(n_8660),
.B1(n_8534),
.B2(n_9387),
.Y(n_11572)
);

INVx1_ASAP7_75t_SL g11573 ( 
.A(n_11050),
.Y(n_11573)
);

AOI22xp33_ASAP7_75t_L g11574 ( 
.A1(n_11053),
.A2(n_9275),
.B1(n_9826),
.B2(n_9828),
.Y(n_11574)
);

OAI21xp5_ASAP7_75t_L g11575 ( 
.A1(n_11179),
.A2(n_9377),
.B(n_9654),
.Y(n_11575)
);

AOI22xp33_ASAP7_75t_L g11576 ( 
.A1(n_10554),
.A2(n_9275),
.B1(n_9379),
.B2(n_9831),
.Y(n_11576)
);

AOI22xp33_ASAP7_75t_L g11577 ( 
.A1(n_10628),
.A2(n_9275),
.B1(n_9379),
.B2(n_9871),
.Y(n_11577)
);

AOI221xp5_ASAP7_75t_L g11578 ( 
.A1(n_11311),
.A2(n_7669),
.B1(n_7608),
.B2(n_8878),
.C(n_8674),
.Y(n_11578)
);

AOI221xp5_ASAP7_75t_L g11579 ( 
.A1(n_10967),
.A2(n_8674),
.B1(n_8878),
.B2(n_8466),
.C(n_8948),
.Y(n_11579)
);

INVx1_ASAP7_75t_L g11580 ( 
.A(n_10929),
.Y(n_11580)
);

AOI21xp5_ASAP7_75t_L g11581 ( 
.A1(n_10829),
.A2(n_10458),
.B(n_11020),
.Y(n_11581)
);

AOI22xp33_ASAP7_75t_L g11582 ( 
.A1(n_11070),
.A2(n_9275),
.B1(n_9379),
.B2(n_9053),
.Y(n_11582)
);

OAI22xp5_ASAP7_75t_L g11583 ( 
.A1(n_11235),
.A2(n_9374),
.B1(n_9383),
.B2(n_9538),
.Y(n_11583)
);

AOI21xp5_ASAP7_75t_L g11584 ( 
.A1(n_10829),
.A2(n_9510),
.B(n_10161),
.Y(n_11584)
);

INVx1_ASAP7_75t_L g11585 ( 
.A(n_10932),
.Y(n_11585)
);

NAND2xp5_ASAP7_75t_L g11586 ( 
.A(n_10638),
.B(n_9029),
.Y(n_11586)
);

OAI22xp5_ASAP7_75t_L g11587 ( 
.A1(n_11060),
.A2(n_9551),
.B1(n_9662),
.B2(n_9603),
.Y(n_11587)
);

AOI22xp5_ASAP7_75t_L g11588 ( 
.A1(n_10529),
.A2(n_9536),
.B1(n_9501),
.B2(n_9513),
.Y(n_11588)
);

AOI22xp33_ASAP7_75t_L g11589 ( 
.A1(n_11381),
.A2(n_9379),
.B1(n_9053),
.B2(n_9054),
.Y(n_11589)
);

AOI22xp33_ASAP7_75t_L g11590 ( 
.A1(n_10523),
.A2(n_9379),
.B1(n_9053),
.B2(n_9054),
.Y(n_11590)
);

OAI22xp5_ASAP7_75t_L g11591 ( 
.A1(n_10683),
.A2(n_9642),
.B1(n_9637),
.B2(n_9588),
.Y(n_11591)
);

AOI22xp33_ASAP7_75t_L g11592 ( 
.A1(n_10523),
.A2(n_9053),
.B1(n_9054),
.B2(n_9800),
.Y(n_11592)
);

OAI22xp33_ASAP7_75t_L g11593 ( 
.A1(n_10529),
.A2(n_10699),
.B1(n_10693),
.B2(n_10995),
.Y(n_11593)
);

AOI22xp33_ASAP7_75t_L g11594 ( 
.A1(n_10813),
.A2(n_9054),
.B1(n_9093),
.B2(n_9086),
.Y(n_11594)
);

OAI22xp33_ASAP7_75t_L g11595 ( 
.A1(n_11266),
.A2(n_8534),
.B1(n_9501),
.B2(n_9387),
.Y(n_11595)
);

INVx3_ASAP7_75t_L g11596 ( 
.A(n_10357),
.Y(n_11596)
);

INVx2_ASAP7_75t_L g11597 ( 
.A(n_11433),
.Y(n_11597)
);

AOI22xp5_ASAP7_75t_L g11598 ( 
.A1(n_10706),
.A2(n_9501),
.B1(n_9513),
.B2(n_9387),
.Y(n_11598)
);

INVx1_ASAP7_75t_L g11599 ( 
.A(n_10933),
.Y(n_11599)
);

INVx3_ASAP7_75t_L g11600 ( 
.A(n_10357),
.Y(n_11600)
);

INVx1_ASAP7_75t_L g11601 ( 
.A(n_10934),
.Y(n_11601)
);

AOI22xp33_ASAP7_75t_L g11602 ( 
.A1(n_10846),
.A2(n_9086),
.B1(n_9152),
.B2(n_9093),
.Y(n_11602)
);

AOI222xp33_ASAP7_75t_L g11603 ( 
.A1(n_10925),
.A2(n_8303),
.B1(n_8312),
.B2(n_10142),
.C1(n_8886),
.C2(n_8842),
.Y(n_11603)
);

AOI21xp5_ASAP7_75t_L g11604 ( 
.A1(n_10878),
.A2(n_10196),
.B(n_10161),
.Y(n_11604)
);

INVx1_ASAP7_75t_L g11605 ( 
.A(n_10940),
.Y(n_11605)
);

AOI22xp33_ASAP7_75t_L g11606 ( 
.A1(n_10677),
.A2(n_9093),
.B1(n_9152),
.B2(n_9719),
.Y(n_11606)
);

AOI222xp33_ASAP7_75t_L g11607 ( 
.A1(n_11204),
.A2(n_8303),
.B1(n_8312),
.B2(n_10142),
.C1(n_8899),
.C2(n_8886),
.Y(n_11607)
);

AND2x4_ASAP7_75t_L g11608 ( 
.A(n_10327),
.B(n_9233),
.Y(n_11608)
);

AOI22xp33_ASAP7_75t_L g11609 ( 
.A1(n_10677),
.A2(n_10904),
.B1(n_10317),
.B2(n_10362),
.Y(n_11609)
);

NOR2xp33_ASAP7_75t_L g11610 ( 
.A(n_10355),
.B(n_10525),
.Y(n_11610)
);

INVx3_ASAP7_75t_L g11611 ( 
.A(n_10507),
.Y(n_11611)
);

INVx2_ASAP7_75t_L g11612 ( 
.A(n_11437),
.Y(n_11612)
);

OAI21x1_ASAP7_75t_L g11613 ( 
.A1(n_11043),
.A2(n_8990),
.B(n_8986),
.Y(n_11613)
);

OAI22xp33_ASAP7_75t_L g11614 ( 
.A1(n_11266),
.A2(n_9501),
.B1(n_9513),
.B2(n_9387),
.Y(n_11614)
);

NAND2xp33_ASAP7_75t_R g11615 ( 
.A(n_11399),
.B(n_8525),
.Y(n_11615)
);

INVx1_ASAP7_75t_L g11616 ( 
.A(n_10941),
.Y(n_11616)
);

AOI22xp33_ASAP7_75t_L g11617 ( 
.A1(n_10904),
.A2(n_9093),
.B1(n_9152),
.B2(n_9554),
.Y(n_11617)
);

INVx1_ASAP7_75t_L g11618 ( 
.A(n_10943),
.Y(n_11618)
);

AND2x2_ASAP7_75t_L g11619 ( 
.A(n_10821),
.B(n_9378),
.Y(n_11619)
);

AND2x4_ASAP7_75t_L g11620 ( 
.A(n_10356),
.B(n_9233),
.Y(n_11620)
);

BUFx3_ASAP7_75t_L g11621 ( 
.A(n_10831),
.Y(n_11621)
);

INVx2_ASAP7_75t_L g11622 ( 
.A(n_11437),
.Y(n_11622)
);

OAI21xp33_ASAP7_75t_L g11623 ( 
.A1(n_10325),
.A2(n_9689),
.B(n_9683),
.Y(n_11623)
);

INVx2_ASAP7_75t_L g11624 ( 
.A(n_10427),
.Y(n_11624)
);

INVx1_ASAP7_75t_L g11625 ( 
.A(n_10949),
.Y(n_11625)
);

AOI21xp5_ASAP7_75t_L g11626 ( 
.A1(n_10740),
.A2(n_10196),
.B(n_10161),
.Y(n_11626)
);

OAI221xp5_ASAP7_75t_L g11627 ( 
.A1(n_10902),
.A2(n_8990),
.B1(n_10028),
.B2(n_9728),
.C(n_9442),
.Y(n_11627)
);

HB1xp67_ASAP7_75t_L g11628 ( 
.A(n_11329),
.Y(n_11628)
);

INVx4_ASAP7_75t_L g11629 ( 
.A(n_10355),
.Y(n_11629)
);

NAND2xp5_ASAP7_75t_L g11630 ( 
.A(n_10580),
.B(n_9029),
.Y(n_11630)
);

OAI21x1_ASAP7_75t_L g11631 ( 
.A1(n_10478),
.A2(n_10578),
.B(n_10576),
.Y(n_11631)
);

OAI221xp5_ASAP7_75t_L g11632 ( 
.A1(n_10974),
.A2(n_10051),
.B1(n_10149),
.B2(n_9269),
.C(n_10042),
.Y(n_11632)
);

AND2x2_ASAP7_75t_L g11633 ( 
.A(n_10836),
.B(n_9378),
.Y(n_11633)
);

AND2x4_ASAP7_75t_L g11634 ( 
.A(n_10356),
.B(n_9233),
.Y(n_11634)
);

OAI22xp5_ASAP7_75t_L g11635 ( 
.A1(n_10338),
.A2(n_8918),
.B1(n_8639),
.B2(n_8883),
.Y(n_11635)
);

AOI22xp33_ASAP7_75t_SL g11636 ( 
.A1(n_11157),
.A2(n_7843),
.B1(n_7619),
.B2(n_7686),
.Y(n_11636)
);

OR2x2_ASAP7_75t_L g11637 ( 
.A(n_10587),
.B(n_9999),
.Y(n_11637)
);

HB1xp67_ASAP7_75t_L g11638 ( 
.A(n_11351),
.Y(n_11638)
);

INVx2_ASAP7_75t_L g11639 ( 
.A(n_10427),
.Y(n_11639)
);

CKINVDCx20_ASAP7_75t_R g11640 ( 
.A(n_10831),
.Y(n_11640)
);

BUFx12f_ASAP7_75t_L g11641 ( 
.A(n_10348),
.Y(n_11641)
);

INVx1_ASAP7_75t_L g11642 ( 
.A(n_10954),
.Y(n_11642)
);

AOI221xp5_ASAP7_75t_L g11643 ( 
.A1(n_10583),
.A2(n_8466),
.B1(n_9037),
.B2(n_9247),
.C(n_9145),
.Y(n_11643)
);

OAI22xp5_ASAP7_75t_L g11644 ( 
.A1(n_10404),
.A2(n_8918),
.B1(n_8639),
.B2(n_8883),
.Y(n_11644)
);

AOI221xp5_ASAP7_75t_L g11645 ( 
.A1(n_11157),
.A2(n_9145),
.B1(n_9247),
.B2(n_9037),
.C(n_8788),
.Y(n_11645)
);

HB1xp67_ASAP7_75t_L g11646 ( 
.A(n_11355),
.Y(n_11646)
);

OAI211xp5_ASAP7_75t_L g11647 ( 
.A1(n_11305),
.A2(n_9965),
.B(n_9971),
.C(n_8274),
.Y(n_11647)
);

OR2x6_ASAP7_75t_L g11648 ( 
.A(n_11357),
.B(n_9093),
.Y(n_11648)
);

AOI22xp33_ASAP7_75t_L g11649 ( 
.A1(n_10350),
.A2(n_9093),
.B1(n_9152),
.B2(n_9554),
.Y(n_11649)
);

NAND3xp33_ASAP7_75t_L g11650 ( 
.A(n_10539),
.B(n_10485),
.C(n_11319),
.Y(n_11650)
);

OR2x2_ASAP7_75t_L g11651 ( 
.A(n_10587),
.B(n_9999),
.Y(n_11651)
);

AOI21xp33_ASAP7_75t_L g11652 ( 
.A1(n_10914),
.A2(n_10019),
.B(n_8982),
.Y(n_11652)
);

AOI22xp33_ASAP7_75t_L g11653 ( 
.A1(n_10370),
.A2(n_9152),
.B1(n_9596),
.B2(n_9554),
.Y(n_11653)
);

AND2x2_ASAP7_75t_L g11654 ( 
.A(n_10836),
.B(n_10858),
.Y(n_11654)
);

AOI22xp33_ASAP7_75t_L g11655 ( 
.A1(n_10380),
.A2(n_9152),
.B1(n_9596),
.B2(n_9554),
.Y(n_11655)
);

INVx3_ASAP7_75t_L g11656 ( 
.A(n_10507),
.Y(n_11656)
);

INVx1_ASAP7_75t_L g11657 ( 
.A(n_10964),
.Y(n_11657)
);

OAI22xp5_ASAP7_75t_L g11658 ( 
.A1(n_10425),
.A2(n_9532),
.B1(n_9524),
.B2(n_9629),
.Y(n_11658)
);

NAND3xp33_ASAP7_75t_L g11659 ( 
.A(n_11383),
.B(n_7686),
.C(n_7619),
.Y(n_11659)
);

INVxp67_ASAP7_75t_SL g11660 ( 
.A(n_10303),
.Y(n_11660)
);

INVx3_ASAP7_75t_L g11661 ( 
.A(n_10684),
.Y(n_11661)
);

INVx1_ASAP7_75t_L g11662 ( 
.A(n_10966),
.Y(n_11662)
);

AND2x2_ASAP7_75t_L g11663 ( 
.A(n_10858),
.B(n_9378),
.Y(n_11663)
);

OAI211xp5_ASAP7_75t_L g11664 ( 
.A1(n_11332),
.A2(n_8274),
.B(n_7686),
.C(n_7619),
.Y(n_11664)
);

OAI22xp5_ASAP7_75t_L g11665 ( 
.A1(n_10537),
.A2(n_8760),
.B1(n_8775),
.B2(n_8769),
.Y(n_11665)
);

AND2x2_ASAP7_75t_L g11666 ( 
.A(n_10315),
.B(n_10352),
.Y(n_11666)
);

OAI221xp5_ASAP7_75t_L g11667 ( 
.A1(n_10945),
.A2(n_9953),
.B1(n_9896),
.B2(n_9487),
.C(n_9529),
.Y(n_11667)
);

INVx5_ASAP7_75t_L g11668 ( 
.A(n_10351),
.Y(n_11668)
);

OAI211xp5_ASAP7_75t_L g11669 ( 
.A1(n_10392),
.A2(n_7686),
.B(n_7619),
.C(n_10183),
.Y(n_11669)
);

AOI22xp33_ASAP7_75t_L g11670 ( 
.A1(n_10914),
.A2(n_10403),
.B1(n_10447),
.B2(n_10395),
.Y(n_11670)
);

AOI22xp5_ASAP7_75t_L g11671 ( 
.A1(n_10538),
.A2(n_9501),
.B1(n_9513),
.B2(n_9387),
.Y(n_11671)
);

AOI221xp5_ASAP7_75t_L g11672 ( 
.A1(n_10444),
.A2(n_10325),
.B1(n_10333),
.B2(n_10926),
.C(n_11122),
.Y(n_11672)
);

XOR2xp5_ASAP7_75t_L g11673 ( 
.A(n_10859),
.B(n_9030),
.Y(n_11673)
);

OR2x6_ASAP7_75t_L g11674 ( 
.A(n_10728),
.B(n_9446),
.Y(n_11674)
);

AOI22xp33_ASAP7_75t_L g11675 ( 
.A1(n_10477),
.A2(n_9596),
.B1(n_9786),
.B2(n_9671),
.Y(n_11675)
);

OAI22xp33_ASAP7_75t_L g11676 ( 
.A1(n_11266),
.A2(n_9501),
.B1(n_9513),
.B2(n_9387),
.Y(n_11676)
);

AOI22xp33_ASAP7_75t_L g11677 ( 
.A1(n_10488),
.A2(n_9596),
.B1(n_9786),
.B2(n_9671),
.Y(n_11677)
);

AOI22xp33_ASAP7_75t_L g11678 ( 
.A1(n_10514),
.A2(n_10558),
.B1(n_10610),
.B2(n_10528),
.Y(n_11678)
);

OAI22xp5_ASAP7_75t_L g11679 ( 
.A1(n_10871),
.A2(n_8760),
.B1(n_8775),
.B2(n_8769),
.Y(n_11679)
);

OR2x2_ASAP7_75t_L g11680 ( 
.A(n_10519),
.B(n_10003),
.Y(n_11680)
);

AOI22xp5_ASAP7_75t_L g11681 ( 
.A1(n_10884),
.A2(n_9517),
.B1(n_9565),
.B2(n_9513),
.Y(n_11681)
);

OAI21xp5_ASAP7_75t_L g11682 ( 
.A1(n_11006),
.A2(n_10196),
.B(n_10161),
.Y(n_11682)
);

OAI22xp5_ASAP7_75t_L g11683 ( 
.A1(n_11000),
.A2(n_8680),
.B1(n_10025),
.B2(n_9978),
.Y(n_11683)
);

OR2x2_ASAP7_75t_L g11684 ( 
.A(n_10378),
.B(n_10003),
.Y(n_11684)
);

INVx1_ASAP7_75t_L g11685 ( 
.A(n_10970),
.Y(n_11685)
);

AOI22xp33_ASAP7_75t_L g11686 ( 
.A1(n_10626),
.A2(n_9671),
.B1(n_9939),
.B2(n_9786),
.Y(n_11686)
);

BUFx6f_ASAP7_75t_L g11687 ( 
.A(n_10307),
.Y(n_11687)
);

OAI22xp5_ASAP7_75t_L g11688 ( 
.A1(n_11266),
.A2(n_9403),
.B1(n_9401),
.B2(n_10167),
.Y(n_11688)
);

AND2x2_ASAP7_75t_L g11689 ( 
.A(n_10315),
.B(n_9458),
.Y(n_11689)
);

INVxp33_ASAP7_75t_L g11690 ( 
.A(n_11221),
.Y(n_11690)
);

HB1xp67_ASAP7_75t_L g11691 ( 
.A(n_11387),
.Y(n_11691)
);

AOI22xp5_ASAP7_75t_L g11692 ( 
.A1(n_11221),
.A2(n_9565),
.B1(n_9570),
.B2(n_9517),
.Y(n_11692)
);

AOI22xp33_ASAP7_75t_SL g11693 ( 
.A1(n_10333),
.A2(n_11122),
.B1(n_10367),
.B2(n_10415),
.Y(n_11693)
);

OR2x6_ASAP7_75t_L g11694 ( 
.A(n_10728),
.B(n_9446),
.Y(n_11694)
);

AOI22xp33_ASAP7_75t_SL g11695 ( 
.A1(n_10349),
.A2(n_7843),
.B1(n_7619),
.B2(n_7686),
.Y(n_11695)
);

INVx1_ASAP7_75t_L g11696 ( 
.A(n_10975),
.Y(n_11696)
);

AOI22xp33_ASAP7_75t_SL g11697 ( 
.A1(n_10349),
.A2(n_7619),
.B1(n_7686),
.B2(n_7683),
.Y(n_11697)
);

HB1xp67_ASAP7_75t_L g11698 ( 
.A(n_11392),
.Y(n_11698)
);

OAI22xp33_ASAP7_75t_L g11699 ( 
.A1(n_11335),
.A2(n_9565),
.B1(n_9570),
.B2(n_9517),
.Y(n_11699)
);

INVx1_ASAP7_75t_L g11700 ( 
.A(n_10976),
.Y(n_11700)
);

NOR2x1_ASAP7_75t_SL g11701 ( 
.A(n_11335),
.B(n_10044),
.Y(n_11701)
);

INVx2_ASAP7_75t_L g11702 ( 
.A(n_10427),
.Y(n_11702)
);

BUFx2_ASAP7_75t_L g11703 ( 
.A(n_11182),
.Y(n_11703)
);

INVx6_ASAP7_75t_L g11704 ( 
.A(n_10302),
.Y(n_11704)
);

BUFx3_ASAP7_75t_L g11705 ( 
.A(n_10859),
.Y(n_11705)
);

INVx1_ASAP7_75t_L g11706 ( 
.A(n_10980),
.Y(n_11706)
);

INVx2_ASAP7_75t_L g11707 ( 
.A(n_10427),
.Y(n_11707)
);

OAI211xp5_ASAP7_75t_SL g11708 ( 
.A1(n_11251),
.A2(n_9104),
.B(n_10080),
.C(n_10074),
.Y(n_11708)
);

CKINVDCx5p33_ASAP7_75t_R g11709 ( 
.A(n_11022),
.Y(n_11709)
);

NAND2xp5_ASAP7_75t_L g11710 ( 
.A(n_10803),
.B(n_9068),
.Y(n_11710)
);

AOI22xp33_ASAP7_75t_L g11711 ( 
.A1(n_10627),
.A2(n_9786),
.B1(n_9939),
.B2(n_9671),
.Y(n_11711)
);

AOI22xp5_ASAP7_75t_L g11712 ( 
.A1(n_10951),
.A2(n_9565),
.B1(n_9570),
.B2(n_9517),
.Y(n_11712)
);

AND2x4_ASAP7_75t_L g11713 ( 
.A(n_10431),
.B(n_9233),
.Y(n_11713)
);

INVx2_ASAP7_75t_SL g11714 ( 
.A(n_10388),
.Y(n_11714)
);

OAI22xp5_ASAP7_75t_L g11715 ( 
.A1(n_11335),
.A2(n_9636),
.B1(n_10251),
.B2(n_10196),
.Y(n_11715)
);

NAND3xp33_ASAP7_75t_L g11716 ( 
.A(n_10346),
.B(n_10141),
.C(n_9939),
.Y(n_11716)
);

OAI22xp5_ASAP7_75t_L g11717 ( 
.A1(n_11335),
.A2(n_10251),
.B1(n_9576),
.B2(n_10184),
.Y(n_11717)
);

AOI221xp5_ASAP7_75t_L g11718 ( 
.A1(n_10367),
.A2(n_9145),
.B1(n_9247),
.B2(n_9037),
.C(n_8788),
.Y(n_11718)
);

OAI22xp33_ASAP7_75t_L g11719 ( 
.A1(n_10990),
.A2(n_9565),
.B1(n_9570),
.B2(n_9517),
.Y(n_11719)
);

BUFx6f_ASAP7_75t_L g11720 ( 
.A(n_10388),
.Y(n_11720)
);

INVx2_ASAP7_75t_L g11721 ( 
.A(n_10535),
.Y(n_11721)
);

INVx11_ASAP7_75t_L g11722 ( 
.A(n_11182),
.Y(n_11722)
);

AOI22xp33_ASAP7_75t_SL g11723 ( 
.A1(n_10415),
.A2(n_7654),
.B1(n_7683),
.B2(n_9255),
.Y(n_11723)
);

AND2x2_ASAP7_75t_L g11724 ( 
.A(n_10352),
.B(n_9458),
.Y(n_11724)
);

OAI221xp5_ASAP7_75t_L g11725 ( 
.A1(n_10963),
.A2(n_9490),
.B1(n_9529),
.B2(n_9487),
.C(n_9446),
.Y(n_11725)
);

INVxp67_ASAP7_75t_L g11726 ( 
.A(n_11261),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_10987),
.Y(n_11727)
);

INVx1_ASAP7_75t_L g11728 ( 
.A(n_10988),
.Y(n_11728)
);

NOR2xp67_ASAP7_75t_L g11729 ( 
.A(n_10302),
.B(n_9446),
.Y(n_11729)
);

OAI22xp5_ASAP7_75t_L g11730 ( 
.A1(n_10752),
.A2(n_10251),
.B1(n_9481),
.B2(n_9507),
.Y(n_11730)
);

AOI22xp33_ASAP7_75t_L g11731 ( 
.A1(n_10631),
.A2(n_10712),
.B1(n_10739),
.B2(n_10709),
.Y(n_11731)
);

CKINVDCx5p33_ASAP7_75t_R g11732 ( 
.A(n_11022),
.Y(n_11732)
);

AOI21xp5_ASAP7_75t_L g11733 ( 
.A1(n_10885),
.A2(n_10251),
.B(n_8761),
.Y(n_11733)
);

INVx2_ASAP7_75t_SL g11734 ( 
.A(n_10531),
.Y(n_11734)
);

OAI211xp5_ASAP7_75t_L g11735 ( 
.A1(n_10303),
.A2(n_8228),
.B(n_7804),
.C(n_8913),
.Y(n_11735)
);

OAI22xp33_ASAP7_75t_L g11736 ( 
.A1(n_10990),
.A2(n_9565),
.B1(n_9570),
.B2(n_9517),
.Y(n_11736)
);

BUFx3_ASAP7_75t_L g11737 ( 
.A(n_10531),
.Y(n_11737)
);

AOI22xp33_ASAP7_75t_L g11738 ( 
.A1(n_10816),
.A2(n_10141),
.B1(n_9939),
.B2(n_9586),
.Y(n_11738)
);

OAI22xp33_ASAP7_75t_L g11739 ( 
.A1(n_10990),
.A2(n_9586),
.B1(n_9604),
.B2(n_9570),
.Y(n_11739)
);

AOI21xp33_ASAP7_75t_L g11740 ( 
.A1(n_10990),
.A2(n_8967),
.B(n_10141),
.Y(n_11740)
);

CKINVDCx6p67_ASAP7_75t_R g11741 ( 
.A(n_10525),
.Y(n_11741)
);

NAND2x1_ASAP7_75t_L g11742 ( 
.A(n_11149),
.B(n_11292),
.Y(n_11742)
);

OAI21xp5_ASAP7_75t_L g11743 ( 
.A1(n_11027),
.A2(n_7884),
.B(n_9372),
.Y(n_11743)
);

BUFx2_ASAP7_75t_L g11744 ( 
.A(n_10536),
.Y(n_11744)
);

OR2x2_ASAP7_75t_L g11745 ( 
.A(n_10378),
.B(n_10168),
.Y(n_11745)
);

AOI21xp5_ASAP7_75t_L g11746 ( 
.A1(n_10885),
.A2(n_8761),
.B(n_8533),
.Y(n_11746)
);

OAI221xp5_ASAP7_75t_SL g11747 ( 
.A1(n_11027),
.A2(n_10127),
.B1(n_10095),
.B2(n_8612),
.C(n_8834),
.Y(n_11747)
);

OA21x2_ASAP7_75t_L g11748 ( 
.A1(n_11003),
.A2(n_11005),
.B(n_10319),
.Y(n_11748)
);

INVx2_ASAP7_75t_L g11749 ( 
.A(n_10535),
.Y(n_11749)
);

AOI22xp33_ASAP7_75t_L g11750 ( 
.A1(n_11027),
.A2(n_10141),
.B1(n_9604),
.B2(n_9632),
.Y(n_11750)
);

OAI22xp33_ASAP7_75t_L g11751 ( 
.A1(n_11027),
.A2(n_10623),
.B1(n_10659),
.B2(n_10593),
.Y(n_11751)
);

AND2x2_ASAP7_75t_L g11752 ( 
.A(n_10352),
.B(n_9458),
.Y(n_11752)
);

AOI221xp5_ASAP7_75t_L g11753 ( 
.A1(n_11249),
.A2(n_9247),
.B1(n_8816),
.B2(n_8899),
.C(n_8839),
.Y(n_11753)
);

AOI21xp5_ASAP7_75t_L g11754 ( 
.A1(n_10885),
.A2(n_8533),
.B(n_8941),
.Y(n_11754)
);

BUFx3_ASAP7_75t_L g11755 ( 
.A(n_10536),
.Y(n_11755)
);

INVx2_ASAP7_75t_L g11756 ( 
.A(n_10535),
.Y(n_11756)
);

AOI22xp33_ASAP7_75t_L g11757 ( 
.A1(n_10784),
.A2(n_9604),
.B1(n_9632),
.B2(n_9586),
.Y(n_11757)
);

INVx1_ASAP7_75t_L g11758 ( 
.A(n_10991),
.Y(n_11758)
);

AND2x2_ASAP7_75t_L g11759 ( 
.A(n_10371),
.B(n_9481),
.Y(n_11759)
);

A2O1A1Ixp33_ASAP7_75t_L g11760 ( 
.A1(n_11130),
.A2(n_8891),
.B(n_8613),
.C(n_8811),
.Y(n_11760)
);

OAI22xp5_ASAP7_75t_L g11761 ( 
.A1(n_10979),
.A2(n_9507),
.B1(n_9543),
.B2(n_9481),
.Y(n_11761)
);

OAI22xp5_ASAP7_75t_L g11762 ( 
.A1(n_10979),
.A2(n_9543),
.B1(n_9507),
.B2(n_8856),
.Y(n_11762)
);

OAI221xp5_ASAP7_75t_L g11763 ( 
.A1(n_11019),
.A2(n_9529),
.B1(n_9490),
.B2(n_9487),
.C(n_10044),
.Y(n_11763)
);

HB1xp67_ASAP7_75t_L g11764 ( 
.A(n_11416),
.Y(n_11764)
);

NOR3xp33_ASAP7_75t_L g11765 ( 
.A(n_11431),
.B(n_9490),
.C(n_9487),
.Y(n_11765)
);

AOI22xp33_ASAP7_75t_L g11766 ( 
.A1(n_10784),
.A2(n_9604),
.B1(n_9632),
.B2(n_9586),
.Y(n_11766)
);

BUFx3_ASAP7_75t_L g11767 ( 
.A(n_10543),
.Y(n_11767)
);

INVx2_ASAP7_75t_L g11768 ( 
.A(n_10535),
.Y(n_11768)
);

OAI22xp5_ASAP7_75t_L g11769 ( 
.A1(n_11314),
.A2(n_9543),
.B1(n_8856),
.B2(n_8834),
.Y(n_11769)
);

AND2x2_ASAP7_75t_L g11770 ( 
.A(n_10371),
.B(n_9548),
.Y(n_11770)
);

AOI222xp33_ASAP7_75t_L g11771 ( 
.A1(n_11369),
.A2(n_11422),
.B1(n_11107),
.B2(n_10561),
.C1(n_10543),
.C2(n_10551),
.Y(n_11771)
);

OR2x2_ASAP7_75t_SL g11772 ( 
.A(n_10346),
.B(n_9586),
.Y(n_11772)
);

AOI22xp33_ASAP7_75t_L g11773 ( 
.A1(n_10850),
.A2(n_9604),
.B1(n_9632),
.B2(n_9586),
.Y(n_11773)
);

AOI22xp33_ASAP7_75t_L g11774 ( 
.A1(n_10850),
.A2(n_9632),
.B1(n_9735),
.B2(n_9604),
.Y(n_11774)
);

AOI22xp33_ASAP7_75t_L g11775 ( 
.A1(n_10899),
.A2(n_9735),
.B1(n_9756),
.B2(n_9632),
.Y(n_11775)
);

AOI211xp5_ASAP7_75t_L g11776 ( 
.A1(n_11056),
.A2(n_10103),
.B(n_8228),
.C(n_8434),
.Y(n_11776)
);

INVx1_ASAP7_75t_L g11777 ( 
.A(n_10993),
.Y(n_11777)
);

NAND4xp25_ASAP7_75t_L g11778 ( 
.A(n_11268),
.B(n_8612),
.C(n_8891),
.D(n_8531),
.Y(n_11778)
);

INVx2_ASAP7_75t_SL g11779 ( 
.A(n_10551),
.Y(n_11779)
);

INVx1_ASAP7_75t_L g11780 ( 
.A(n_10994),
.Y(n_11780)
);

OAI22xp33_ASAP7_75t_L g11781 ( 
.A1(n_10593),
.A2(n_9756),
.B1(n_9895),
.B2(n_9735),
.Y(n_11781)
);

A2O1A1Ixp33_ASAP7_75t_L g11782 ( 
.A1(n_11130),
.A2(n_11298),
.B(n_10561),
.C(n_10302),
.Y(n_11782)
);

AOI22xp33_ASAP7_75t_L g11783 ( 
.A1(n_10899),
.A2(n_9756),
.B1(n_9895),
.B2(n_9735),
.Y(n_11783)
);

AND2x2_ASAP7_75t_L g11784 ( 
.A(n_10371),
.B(n_9548),
.Y(n_11784)
);

AND2x4_ASAP7_75t_L g11785 ( 
.A(n_10431),
.B(n_9233),
.Y(n_11785)
);

AOI22xp33_ASAP7_75t_L g11786 ( 
.A1(n_10921),
.A2(n_9756),
.B1(n_9895),
.B2(n_9735),
.Y(n_11786)
);

INVx2_ASAP7_75t_L g11787 ( 
.A(n_10548),
.Y(n_11787)
);

AND2x2_ASAP7_75t_L g11788 ( 
.A(n_10399),
.B(n_9548),
.Y(n_11788)
);

AOI22xp33_ASAP7_75t_L g11789 ( 
.A1(n_10921),
.A2(n_9756),
.B1(n_9895),
.B2(n_9735),
.Y(n_11789)
);

NOR2x1p5_ASAP7_75t_L g11790 ( 
.A(n_11135),
.B(n_11227),
.Y(n_11790)
);

AOI22xp33_ASAP7_75t_L g11791 ( 
.A1(n_11011),
.A2(n_9895),
.B1(n_9897),
.B2(n_9756),
.Y(n_11791)
);

AOI21xp5_ASAP7_75t_L g11792 ( 
.A1(n_11130),
.A2(n_8533),
.B(n_8941),
.Y(n_11792)
);

AOI222xp33_ASAP7_75t_L g11793 ( 
.A1(n_11216),
.A2(n_8816),
.B1(n_8366),
.B2(n_8540),
.C1(n_8256),
.C2(n_9681),
.Y(n_11793)
);

INVx3_ASAP7_75t_L g11794 ( 
.A(n_10684),
.Y(n_11794)
);

OAI211xp5_ASAP7_75t_L g11795 ( 
.A1(n_10346),
.A2(n_7804),
.B(n_8913),
.C(n_8545),
.Y(n_11795)
);

AOI22xp33_ASAP7_75t_SL g11796 ( 
.A1(n_11249),
.A2(n_7654),
.B1(n_7683),
.B2(n_8909),
.Y(n_11796)
);

AND2x2_ASAP7_75t_L g11797 ( 
.A(n_10399),
.B(n_9606),
.Y(n_11797)
);

BUFx12f_ASAP7_75t_L g11798 ( 
.A(n_10348),
.Y(n_11798)
);

AND2x2_ASAP7_75t_L g11799 ( 
.A(n_10399),
.B(n_9606),
.Y(n_11799)
);

INVx1_ASAP7_75t_L g11800 ( 
.A(n_10996),
.Y(n_11800)
);

INVx2_ASAP7_75t_SL g11801 ( 
.A(n_10520),
.Y(n_11801)
);

INVx1_ASAP7_75t_L g11802 ( 
.A(n_11002),
.Y(n_11802)
);

OAI221xp5_ASAP7_75t_L g11803 ( 
.A1(n_11077),
.A2(n_11167),
.B1(n_11197),
.B2(n_11088),
.C(n_11083),
.Y(n_11803)
);

AOI22xp33_ASAP7_75t_L g11804 ( 
.A1(n_11011),
.A2(n_9897),
.B1(n_9923),
.B2(n_9895),
.Y(n_11804)
);

BUFx3_ASAP7_75t_L g11805 ( 
.A(n_11438),
.Y(n_11805)
);

INVx2_ASAP7_75t_SL g11806 ( 
.A(n_10520),
.Y(n_11806)
);

AOI22xp33_ASAP7_75t_L g11807 ( 
.A1(n_11223),
.A2(n_9923),
.B1(n_9928),
.B2(n_9897),
.Y(n_11807)
);

INVx4_ASAP7_75t_L g11808 ( 
.A(n_10302),
.Y(n_11808)
);

INVx1_ASAP7_75t_L g11809 ( 
.A(n_11014),
.Y(n_11809)
);

AOI221x1_ASAP7_75t_L g11810 ( 
.A1(n_10834),
.A2(n_9928),
.B1(n_10065),
.B2(n_9923),
.C(n_9897),
.Y(n_11810)
);

OAI221xp5_ASAP7_75t_L g11811 ( 
.A1(n_11439),
.A2(n_9529),
.B1(n_9490),
.B2(n_10044),
.C(n_9078),
.Y(n_11811)
);

AND2x4_ASAP7_75t_L g11812 ( 
.A(n_10432),
.B(n_9257),
.Y(n_11812)
);

AOI21x1_ASAP7_75t_L g11813 ( 
.A1(n_11275),
.A2(n_10186),
.B(n_10126),
.Y(n_11813)
);

OAI221xp5_ASAP7_75t_L g11814 ( 
.A1(n_10593),
.A2(n_10044),
.B1(n_9078),
.B2(n_9120),
.C(n_9064),
.Y(n_11814)
);

OA21x2_ASAP7_75t_L g11815 ( 
.A1(n_11003),
.A2(n_9170),
.B(n_10107),
.Y(n_11815)
);

NAND2xp5_ASAP7_75t_L g11816 ( 
.A(n_11076),
.B(n_9115),
.Y(n_11816)
);

AOI22xp33_ASAP7_75t_SL g11817 ( 
.A1(n_11249),
.A2(n_7654),
.B1(n_7683),
.B2(n_8909),
.Y(n_11817)
);

A2O1A1Ixp33_ASAP7_75t_L g11818 ( 
.A1(n_11298),
.A2(n_8613),
.B(n_8811),
.C(n_8019),
.Y(n_11818)
);

OAI221xp5_ASAP7_75t_L g11819 ( 
.A1(n_10593),
.A2(n_10044),
.B1(n_9078),
.B2(n_9120),
.C(n_9064),
.Y(n_11819)
);

AOI332xp33_ASAP7_75t_L g11820 ( 
.A1(n_11429),
.A2(n_10124),
.A3(n_10112),
.B1(n_10131),
.B2(n_10130),
.B3(n_10119),
.C1(n_10107),
.C2(n_10243),
.Y(n_11820)
);

OR2x2_ASAP7_75t_L g11821 ( 
.A(n_10434),
.B(n_11419),
.Y(n_11821)
);

AOI221xp5_ASAP7_75t_L g11822 ( 
.A1(n_11194),
.A2(n_8607),
.B1(n_8538),
.B2(n_8552),
.C(n_7695),
.Y(n_11822)
);

OAI22xp5_ASAP7_75t_L g11823 ( 
.A1(n_10432),
.A2(n_10197),
.B1(n_7671),
.B2(n_7772),
.Y(n_11823)
);

INVx3_ASAP7_75t_L g11824 ( 
.A(n_11207),
.Y(n_11824)
);

AND2x4_ASAP7_75t_L g11825 ( 
.A(n_10524),
.B(n_9257),
.Y(n_11825)
);

AND2x2_ASAP7_75t_L g11826 ( 
.A(n_10406),
.B(n_9606),
.Y(n_11826)
);

OAI21xp33_ASAP7_75t_L g11827 ( 
.A1(n_10434),
.A2(n_8531),
.B(n_8373),
.Y(n_11827)
);

NAND3xp33_ASAP7_75t_SL g11828 ( 
.A(n_11368),
.B(n_8525),
.C(n_9106),
.Y(n_11828)
);

AOI211xp5_ASAP7_75t_L g11829 ( 
.A1(n_10430),
.A2(n_8434),
.B(n_8426),
.C(n_7989),
.Y(n_11829)
);

AOI22xp33_ASAP7_75t_L g11830 ( 
.A1(n_10351),
.A2(n_9923),
.B1(n_9928),
.B2(n_9897),
.Y(n_11830)
);

NAND2xp5_ASAP7_75t_L g11831 ( 
.A(n_11396),
.B(n_9156),
.Y(n_11831)
);

INVx4_ASAP7_75t_L g11832 ( 
.A(n_10302),
.Y(n_11832)
);

OAI22xp5_ASAP7_75t_L g11833 ( 
.A1(n_10524),
.A2(n_7671),
.B1(n_7772),
.B2(n_7609),
.Y(n_11833)
);

OAI211xp5_ASAP7_75t_SL g11834 ( 
.A1(n_11382),
.A2(n_10168),
.B(n_9241),
.C(n_9390),
.Y(n_11834)
);

CKINVDCx5p33_ASAP7_75t_R g11835 ( 
.A(n_10741),
.Y(n_11835)
);

OAI22xp5_ASAP7_75t_L g11836 ( 
.A1(n_10632),
.A2(n_7671),
.B1(n_7772),
.B2(n_7609),
.Y(n_11836)
);

AND2x2_ASAP7_75t_L g11837 ( 
.A(n_10406),
.B(n_9646),
.Y(n_11837)
);

AOI22xp33_ASAP7_75t_L g11838 ( 
.A1(n_10351),
.A2(n_9923),
.B1(n_9928),
.B2(n_9897),
.Y(n_11838)
);

OAI22xp5_ASAP7_75t_L g11839 ( 
.A1(n_10632),
.A2(n_10742),
.B1(n_10747),
.B2(n_10664),
.Y(n_11839)
);

INVx2_ASAP7_75t_L g11840 ( 
.A(n_10548),
.Y(n_11840)
);

OAI21x1_ASAP7_75t_L g11841 ( 
.A1(n_10522),
.A2(n_10186),
.B(n_9491),
.Y(n_11841)
);

AOI22xp33_ASAP7_75t_L g11842 ( 
.A1(n_10351),
.A2(n_10394),
.B1(n_10360),
.B2(n_10623),
.Y(n_11842)
);

AOI22xp33_ASAP7_75t_SL g11843 ( 
.A1(n_11194),
.A2(n_7654),
.B1(n_7683),
.B2(n_7770),
.Y(n_11843)
);

INVx2_ASAP7_75t_L g11844 ( 
.A(n_10548),
.Y(n_11844)
);

OAI211xp5_ASAP7_75t_L g11845 ( 
.A1(n_11423),
.A2(n_7804),
.B(n_8545),
.C(n_8540),
.Y(n_11845)
);

INVx2_ASAP7_75t_L g11846 ( 
.A(n_10548),
.Y(n_11846)
);

AOI221xp5_ASAP7_75t_L g11847 ( 
.A1(n_11194),
.A2(n_8538),
.B1(n_8552),
.B2(n_7695),
.C(n_10256),
.Y(n_11847)
);

NAND2xp5_ASAP7_75t_L g11848 ( 
.A(n_10664),
.B(n_9156),
.Y(n_11848)
);

INVx5_ASAP7_75t_L g11849 ( 
.A(n_10360),
.Y(n_11849)
);

INVx4_ASAP7_75t_L g11850 ( 
.A(n_10360),
.Y(n_11850)
);

BUFx4f_ASAP7_75t_SL g11851 ( 
.A(n_11438),
.Y(n_11851)
);

AOI22xp33_ASAP7_75t_SL g11852 ( 
.A1(n_10463),
.A2(n_7654),
.B1(n_7828),
.B2(n_7770),
.Y(n_11852)
);

AOI22xp33_ASAP7_75t_L g11853 ( 
.A1(n_10360),
.A2(n_9928),
.B1(n_10065),
.B2(n_9923),
.Y(n_11853)
);

OAI221xp5_ASAP7_75t_L g11854 ( 
.A1(n_10623),
.A2(n_10659),
.B1(n_11298),
.B2(n_10747),
.C(n_10777),
.Y(n_11854)
);

AOI22xp33_ASAP7_75t_L g11855 ( 
.A1(n_10394),
.A2(n_10065),
.B1(n_10164),
.B2(n_9928),
.Y(n_11855)
);

OAI22xp33_ASAP7_75t_L g11856 ( 
.A1(n_10623),
.A2(n_10164),
.B1(n_10176),
.B2(n_10065),
.Y(n_11856)
);

INVx2_ASAP7_75t_L g11857 ( 
.A(n_10560),
.Y(n_11857)
);

AOI22xp33_ASAP7_75t_SL g11858 ( 
.A1(n_10611),
.A2(n_8013),
.B1(n_7828),
.B2(n_7841),
.Y(n_11858)
);

AOI22xp33_ASAP7_75t_SL g11859 ( 
.A1(n_10611),
.A2(n_10381),
.B1(n_10634),
.B2(n_11084),
.Y(n_11859)
);

OAI21xp5_ASAP7_75t_L g11860 ( 
.A1(n_10319),
.A2(n_8546),
.B(n_8398),
.Y(n_11860)
);

BUFx6f_ASAP7_75t_L g11861 ( 
.A(n_10394),
.Y(n_11861)
);

OAI22xp33_ASAP7_75t_L g11862 ( 
.A1(n_10659),
.A2(n_10164),
.B1(n_10176),
.B2(n_10065),
.Y(n_11862)
);

INVx2_ASAP7_75t_L g11863 ( 
.A(n_10560),
.Y(n_11863)
);

INVx2_ASAP7_75t_L g11864 ( 
.A(n_10560),
.Y(n_11864)
);

OAI21x1_ASAP7_75t_SL g11865 ( 
.A1(n_10742),
.A2(n_9390),
.B(n_9241),
.Y(n_11865)
);

AOI221xp5_ASAP7_75t_SL g11866 ( 
.A1(n_10436),
.A2(n_8824),
.B1(n_8859),
.B2(n_8838),
.C(n_8781),
.Y(n_11866)
);

AOI221xp5_ASAP7_75t_L g11867 ( 
.A1(n_10381),
.A2(n_10256),
.B1(n_8824),
.B2(n_8366),
.C(n_8462),
.Y(n_11867)
);

INVx1_ASAP7_75t_L g11868 ( 
.A(n_11023),
.Y(n_11868)
);

CKINVDCx20_ASAP7_75t_R g11869 ( 
.A(n_10741),
.Y(n_11869)
);

OAI221xp5_ASAP7_75t_L g11870 ( 
.A1(n_10659),
.A2(n_9120),
.B1(n_9064),
.B2(n_9712),
.C(n_9646),
.Y(n_11870)
);

INVx2_ASAP7_75t_L g11871 ( 
.A(n_10560),
.Y(n_11871)
);

AND2x2_ASAP7_75t_L g11872 ( 
.A(n_10406),
.B(n_9646),
.Y(n_11872)
);

OAI22xp5_ASAP7_75t_L g11873 ( 
.A1(n_10777),
.A2(n_7671),
.B1(n_7772),
.B2(n_7609),
.Y(n_11873)
);

OR2x6_ASAP7_75t_L g11874 ( 
.A(n_10728),
.B(n_8911),
.Y(n_11874)
);

INVx1_ASAP7_75t_L g11875 ( 
.A(n_11024),
.Y(n_11875)
);

AND2x2_ASAP7_75t_L g11876 ( 
.A(n_10483),
.B(n_9712),
.Y(n_11876)
);

AOI21xp5_ASAP7_75t_L g11877 ( 
.A1(n_10728),
.A2(n_8426),
.B(n_8155),
.Y(n_11877)
);

AND2x2_ASAP7_75t_L g11878 ( 
.A(n_10483),
.B(n_9712),
.Y(n_11878)
);

BUFx4f_ASAP7_75t_SL g11879 ( 
.A(n_10566),
.Y(n_11879)
);

INVx2_ASAP7_75t_L g11880 ( 
.A(n_10571),
.Y(n_11880)
);

INVx1_ASAP7_75t_L g11881 ( 
.A(n_11029),
.Y(n_11881)
);

INVxp67_ASAP7_75t_L g11882 ( 
.A(n_10320),
.Y(n_11882)
);

BUFx6f_ASAP7_75t_L g11883 ( 
.A(n_10394),
.Y(n_11883)
);

OAI22xp5_ASAP7_75t_L g11884 ( 
.A1(n_10785),
.A2(n_9226),
.B1(n_10221),
.B2(n_10215),
.Y(n_11884)
);

OA21x2_ASAP7_75t_L g11885 ( 
.A1(n_11005),
.A2(n_9170),
.B(n_10112),
.Y(n_11885)
);

AOI21xp33_ASAP7_75t_L g11886 ( 
.A1(n_11084),
.A2(n_9515),
.B(n_9509),
.Y(n_11886)
);

CKINVDCx11_ASAP7_75t_R g11887 ( 
.A(n_10566),
.Y(n_11887)
);

OAI211xp5_ASAP7_75t_L g11888 ( 
.A1(n_11391),
.A2(n_7804),
.B(n_8897),
.C(n_8256),
.Y(n_11888)
);

INVx1_ASAP7_75t_L g11889 ( 
.A(n_11030),
.Y(n_11889)
);

CKINVDCx5p33_ASAP7_75t_R g11890 ( 
.A(n_10999),
.Y(n_11890)
);

AOI22xp33_ASAP7_75t_L g11891 ( 
.A1(n_10572),
.A2(n_10065),
.B1(n_10176),
.B2(n_10164),
.Y(n_11891)
);

AOI221xp5_ASAP7_75t_L g11892 ( 
.A1(n_10381),
.A2(n_10256),
.B1(n_8462),
.B2(n_7841),
.C(n_8468),
.Y(n_11892)
);

INVx1_ASAP7_75t_L g11893 ( 
.A(n_11031),
.Y(n_11893)
);

AND2x2_ASAP7_75t_L g11894 ( 
.A(n_10483),
.B(n_9744),
.Y(n_11894)
);

AND2x2_ASAP7_75t_L g11895 ( 
.A(n_10487),
.B(n_9744),
.Y(n_11895)
);

OR2x2_ASAP7_75t_L g11896 ( 
.A(n_10863),
.B(n_7895),
.Y(n_11896)
);

INVx1_ASAP7_75t_L g11897 ( 
.A(n_11033),
.Y(n_11897)
);

OAI22xp5_ASAP7_75t_L g11898 ( 
.A1(n_10785),
.A2(n_8657),
.B1(n_8430),
.B2(n_9744),
.Y(n_11898)
);

OAI31xp33_ASAP7_75t_L g11899 ( 
.A1(n_10407),
.A2(n_9794),
.A3(n_9815),
.B(n_9747),
.Y(n_11899)
);

AOI221xp5_ASAP7_75t_L g11900 ( 
.A1(n_10634),
.A2(n_11084),
.B1(n_10402),
.B2(n_10420),
.C(n_10375),
.Y(n_11900)
);

BUFx2_ASAP7_75t_L g11901 ( 
.A(n_10947),
.Y(n_11901)
);

OAI211xp5_ASAP7_75t_L g11902 ( 
.A1(n_11323),
.A2(n_7804),
.B(n_8897),
.C(n_8081),
.Y(n_11902)
);

OAI22xp5_ASAP7_75t_L g11903 ( 
.A1(n_10802),
.A2(n_8657),
.B1(n_8430),
.B2(n_9747),
.Y(n_11903)
);

HB1xp67_ASAP7_75t_L g11904 ( 
.A(n_10750),
.Y(n_11904)
);

OAI22xp5_ASAP7_75t_L g11905 ( 
.A1(n_10802),
.A2(n_9794),
.B1(n_9815),
.B2(n_9747),
.Y(n_11905)
);

NOR2xp33_ASAP7_75t_L g11906 ( 
.A(n_11227),
.B(n_9664),
.Y(n_11906)
);

AOI21xp5_ASAP7_75t_L g11907 ( 
.A1(n_10634),
.A2(n_8155),
.B(n_9264),
.Y(n_11907)
);

OAI21x1_ASAP7_75t_L g11908 ( 
.A1(n_11207),
.A2(n_9491),
.B(n_10248),
.Y(n_11908)
);

OAI22xp33_ASAP7_75t_L g11909 ( 
.A1(n_10955),
.A2(n_10176),
.B1(n_10237),
.B2(n_10164),
.Y(n_11909)
);

AOI222xp33_ASAP7_75t_L g11910 ( 
.A1(n_10955),
.A2(n_8373),
.B1(n_8339),
.B2(n_8439),
.C1(n_8468),
.C2(n_8648),
.Y(n_11910)
);

INVx1_ASAP7_75t_L g11911 ( 
.A(n_11034),
.Y(n_11911)
);

NAND2xp5_ASAP7_75t_L g11912 ( 
.A(n_10805),
.B(n_10838),
.Y(n_11912)
);

AO221x2_ASAP7_75t_L g11913 ( 
.A1(n_11441),
.A2(n_8859),
.B1(n_8474),
.B2(n_8801),
.C(n_8853),
.Y(n_11913)
);

AOI22xp33_ASAP7_75t_SL g11914 ( 
.A1(n_11112),
.A2(n_8013),
.B1(n_7828),
.B2(n_7852),
.Y(n_11914)
);

OR2x2_ASAP7_75t_L g11915 ( 
.A(n_10863),
.B(n_7895),
.Y(n_11915)
);

AOI22xp33_ASAP7_75t_SL g11916 ( 
.A1(n_11112),
.A2(n_8013),
.B1(n_7852),
.B2(n_8394),
.Y(n_11916)
);

INVx6_ASAP7_75t_SL g11917 ( 
.A(n_10674),
.Y(n_11917)
);

OAI221xp5_ASAP7_75t_SL g11918 ( 
.A1(n_10674),
.A2(n_7989),
.B1(n_7914),
.B2(n_8015),
.C(n_8698),
.Y(n_11918)
);

OAI22xp33_ASAP7_75t_L g11919 ( 
.A1(n_10965),
.A2(n_10176),
.B1(n_10237),
.B2(n_10164),
.Y(n_11919)
);

NAND2xp5_ASAP7_75t_L g11920 ( 
.A(n_10805),
.B(n_9509),
.Y(n_11920)
);

INVx1_ASAP7_75t_L g11921 ( 
.A(n_11036),
.Y(n_11921)
);

AOI22xp33_ASAP7_75t_L g11922 ( 
.A1(n_10572),
.A2(n_10237),
.B1(n_10176),
.B2(n_9794),
.Y(n_11922)
);

NAND2xp5_ASAP7_75t_L g11923 ( 
.A(n_10838),
.B(n_10880),
.Y(n_11923)
);

AOI22xp33_ASAP7_75t_L g11924 ( 
.A1(n_10573),
.A2(n_10237),
.B1(n_9815),
.B2(n_9840),
.Y(n_11924)
);

OR2x2_ASAP7_75t_L g11925 ( 
.A(n_10503),
.B(n_7895),
.Y(n_11925)
);

AND2x4_ASAP7_75t_SL g11926 ( 
.A(n_10426),
.B(n_9315),
.Y(n_11926)
);

INVx2_ASAP7_75t_L g11927 ( 
.A(n_10571),
.Y(n_11927)
);

INVx2_ASAP7_75t_L g11928 ( 
.A(n_10571),
.Y(n_11928)
);

AND2x2_ASAP7_75t_L g11929 ( 
.A(n_10487),
.B(n_9837),
.Y(n_11929)
);

A2O1A1Ixp33_ASAP7_75t_L g11930 ( 
.A1(n_10407),
.A2(n_8019),
.B(n_8507),
.C(n_8475),
.Y(n_11930)
);

OAI21xp5_ASAP7_75t_L g11931 ( 
.A1(n_10308),
.A2(n_8546),
.B(n_8398),
.Y(n_11931)
);

NAND2xp5_ASAP7_75t_L g11932 ( 
.A(n_10880),
.B(n_9515),
.Y(n_11932)
);

AOI22xp33_ASAP7_75t_L g11933 ( 
.A1(n_10573),
.A2(n_10237),
.B1(n_9840),
.B2(n_9855),
.Y(n_11933)
);

INVx2_ASAP7_75t_L g11934 ( 
.A(n_10571),
.Y(n_11934)
);

OAI22xp33_ASAP7_75t_SL g11935 ( 
.A1(n_10376),
.A2(n_9491),
.B1(n_9810),
.B2(n_9703),
.Y(n_11935)
);

AOI221xp5_ASAP7_75t_L g11936 ( 
.A1(n_10368),
.A2(n_10256),
.B1(n_8801),
.B2(n_7620),
.C(n_7637),
.Y(n_11936)
);

OAI22xp5_ASAP7_75t_L g11937 ( 
.A1(n_10946),
.A2(n_10965),
.B1(n_10962),
.B2(n_10947),
.Y(n_11937)
);

AO21x2_ASAP7_75t_L g11938 ( 
.A1(n_11374),
.A2(n_10119),
.B(n_10112),
.Y(n_11938)
);

OAI21xp5_ASAP7_75t_L g11939 ( 
.A1(n_10308),
.A2(n_8546),
.B(n_8398),
.Y(n_11939)
);

OAI22xp33_ASAP7_75t_L g11940 ( 
.A1(n_10364),
.A2(n_10237),
.B1(n_9840),
.B2(n_9855),
.Y(n_11940)
);

OAI22xp5_ASAP7_75t_L g11941 ( 
.A1(n_10946),
.A2(n_9855),
.B1(n_9926),
.B2(n_9837),
.Y(n_11941)
);

AOI22xp33_ASAP7_75t_L g11942 ( 
.A1(n_10602),
.A2(n_9926),
.B1(n_9975),
.B2(n_9837),
.Y(n_11942)
);

OAI21xp5_ASAP7_75t_SL g11943 ( 
.A1(n_11279),
.A2(n_8507),
.B(n_8475),
.Y(n_11943)
);

AND2x2_ASAP7_75t_L g11944 ( 
.A(n_10487),
.B(n_9926),
.Y(n_11944)
);

NOR2xp33_ASAP7_75t_L g11945 ( 
.A(n_10999),
.B(n_9267),
.Y(n_11945)
);

OAI222xp33_ASAP7_75t_L g11946 ( 
.A1(n_10674),
.A2(n_8852),
.B1(n_8648),
.B2(n_8394),
.C1(n_9562),
.C2(n_9558),
.Y(n_11946)
);

INVx1_ASAP7_75t_L g11947 ( 
.A(n_11040),
.Y(n_11947)
);

NAND2xp5_ASAP7_75t_L g11948 ( 
.A(n_10429),
.B(n_9558),
.Y(n_11948)
);

AOI21xp5_ASAP7_75t_L g11949 ( 
.A1(n_10674),
.A2(n_9473),
.B(n_9428),
.Y(n_11949)
);

INVx3_ASAP7_75t_L g11950 ( 
.A(n_10426),
.Y(n_11950)
);

AOI221xp5_ASAP7_75t_L g11951 ( 
.A1(n_10435),
.A2(n_7620),
.B1(n_7637),
.B2(n_7629),
.C(n_7618),
.Y(n_11951)
);

AND2x4_ASAP7_75t_L g11952 ( 
.A(n_10962),
.B(n_9257),
.Y(n_11952)
);

AOI22xp33_ASAP7_75t_L g11953 ( 
.A1(n_10602),
.A2(n_10001),
.B1(n_10004),
.B2(n_9975),
.Y(n_11953)
);

OAI211xp5_ASAP7_75t_SL g11954 ( 
.A1(n_11214),
.A2(n_9693),
.B(n_9940),
.C(n_9562),
.Y(n_11954)
);

AND2x4_ASAP7_75t_L g11955 ( 
.A(n_11037),
.B(n_9257),
.Y(n_11955)
);

OAI221xp5_ASAP7_75t_L g11956 ( 
.A1(n_10694),
.A2(n_10004),
.B1(n_10023),
.B2(n_10001),
.C(n_9975),
.Y(n_11956)
);

OAI22xp5_ASAP7_75t_L g11957 ( 
.A1(n_11037),
.A2(n_10004),
.B1(n_10023),
.B2(n_10001),
.Y(n_11957)
);

OAI22xp5_ASAP7_75t_L g11958 ( 
.A1(n_11143),
.A2(n_10078),
.B1(n_10165),
.B2(n_10023),
.Y(n_11958)
);

AOI22xp33_ASAP7_75t_L g11959 ( 
.A1(n_10633),
.A2(n_10744),
.B1(n_10768),
.B2(n_10685),
.Y(n_11959)
);

HB1xp67_ASAP7_75t_L g11960 ( 
.A(n_10765),
.Y(n_11960)
);

OAI22xp5_ASAP7_75t_L g11961 ( 
.A1(n_11143),
.A2(n_10165),
.B1(n_10194),
.B2(n_10078),
.Y(n_11961)
);

INVx1_ASAP7_75t_L g11962 ( 
.A(n_11042),
.Y(n_11962)
);

INVx1_ASAP7_75t_L g11963 ( 
.A(n_11044),
.Y(n_11963)
);

BUFx2_ASAP7_75t_L g11964 ( 
.A(n_11152),
.Y(n_11964)
);

CKINVDCx5p33_ASAP7_75t_R g11965 ( 
.A(n_10428),
.Y(n_11965)
);

OAI22xp33_ASAP7_75t_L g11966 ( 
.A1(n_10364),
.A2(n_10165),
.B1(n_10194),
.B2(n_10078),
.Y(n_11966)
);

BUFx6f_ASAP7_75t_L g11967 ( 
.A(n_10633),
.Y(n_11967)
);

AOI221xp5_ASAP7_75t_L g11968 ( 
.A1(n_10452),
.A2(n_7620),
.B1(n_7637),
.B2(n_7629),
.C(n_7618),
.Y(n_11968)
);

OAI22xp5_ASAP7_75t_L g11969 ( 
.A1(n_11152),
.A2(n_10194),
.B1(n_8698),
.B2(n_8718),
.Y(n_11969)
);

AND2x2_ASAP7_75t_L g11970 ( 
.A(n_10436),
.B(n_10437),
.Y(n_11970)
);

AOI221xp5_ASAP7_75t_L g11971 ( 
.A1(n_10453),
.A2(n_7620),
.B1(n_7637),
.B2(n_7629),
.C(n_7618),
.Y(n_11971)
);

OAI22xp5_ASAP7_75t_L g11972 ( 
.A1(n_11171),
.A2(n_8718),
.B1(n_8345),
.B2(n_8358),
.Y(n_11972)
);

OR2x2_ASAP7_75t_L g11973 ( 
.A(n_10503),
.B(n_9693),
.Y(n_11973)
);

AND2x2_ASAP7_75t_L g11974 ( 
.A(n_10437),
.B(n_9940),
.Y(n_11974)
);

INVx1_ASAP7_75t_L g11975 ( 
.A(n_11048),
.Y(n_11975)
);

OAI21x1_ASAP7_75t_L g11976 ( 
.A1(n_11256),
.A2(n_10266),
.B(n_10248),
.Y(n_11976)
);

HB1xp67_ASAP7_75t_L g11977 ( 
.A(n_10769),
.Y(n_11977)
);

AOI222xp33_ASAP7_75t_L g11978 ( 
.A1(n_10685),
.A2(n_10768),
.B1(n_10776),
.B2(n_10744),
.C1(n_11236),
.C2(n_11171),
.Y(n_11978)
);

INVx4_ASAP7_75t_L g11979 ( 
.A(n_10776),
.Y(n_11979)
);

AND2x2_ASAP7_75t_L g11980 ( 
.A(n_10451),
.B(n_10469),
.Y(n_11980)
);

OAI221xp5_ASAP7_75t_L g11981 ( 
.A1(n_10694),
.A2(n_10079),
.B1(n_10159),
.B2(n_10111),
.C(n_10015),
.Y(n_11981)
);

INVx3_ASAP7_75t_L g11982 ( 
.A(n_10426),
.Y(n_11982)
);

INVx1_ASAP7_75t_L g11983 ( 
.A(n_11052),
.Y(n_11983)
);

OAI211xp5_ASAP7_75t_L g11984 ( 
.A1(n_10505),
.A2(n_7804),
.B(n_8081),
.C(n_7914),
.Y(n_11984)
);

AND2x2_ASAP7_75t_L g11985 ( 
.A(n_10451),
.B(n_10015),
.Y(n_11985)
);

AOI22xp5_ASAP7_75t_L g11986 ( 
.A1(n_11214),
.A2(n_11238),
.B1(n_11245),
.B2(n_11236),
.Y(n_11986)
);

NAND2xp5_ASAP7_75t_L g11987 ( 
.A(n_10462),
.B(n_10079),
.Y(n_11987)
);

OAI21xp33_ASAP7_75t_L g11988 ( 
.A1(n_10469),
.A2(n_10541),
.B(n_10540),
.Y(n_11988)
);

AOI22xp33_ASAP7_75t_L g11989 ( 
.A1(n_11238),
.A2(n_9783),
.B1(n_9839),
.B2(n_9752),
.Y(n_11989)
);

BUFx4f_ASAP7_75t_SL g11990 ( 
.A(n_11279),
.Y(n_11990)
);

NAND2xp5_ASAP7_75t_L g11991 ( 
.A(n_10464),
.B(n_10111),
.Y(n_11991)
);

INVx2_ASAP7_75t_L g11992 ( 
.A(n_10575),
.Y(n_11992)
);

NAND2xp5_ASAP7_75t_L g11993 ( 
.A(n_10501),
.B(n_10159),
.Y(n_11993)
);

INVx2_ASAP7_75t_L g11994 ( 
.A(n_10575),
.Y(n_11994)
);

AOI22xp5_ASAP7_75t_L g11995 ( 
.A1(n_11245),
.A2(n_11361),
.B1(n_11347),
.B2(n_10835),
.Y(n_11995)
);

OAI22xp5_ASAP7_75t_L g11996 ( 
.A1(n_11370),
.A2(n_8345),
.B1(n_8358),
.B2(n_10209),
.Y(n_11996)
);

AOI22xp33_ASAP7_75t_L g11997 ( 
.A1(n_10575),
.A2(n_9752),
.B1(n_9839),
.B2(n_9783),
.Y(n_11997)
);

AOI22xp33_ASAP7_75t_L g11998 ( 
.A1(n_10575),
.A2(n_9752),
.B1(n_9839),
.B2(n_9783),
.Y(n_11998)
);

AOI21xp33_ASAP7_75t_L g11999 ( 
.A1(n_10834),
.A2(n_10209),
.B(n_7717),
.Y(n_11999)
);

OAI22xp33_ASAP7_75t_L g12000 ( 
.A1(n_10364),
.A2(n_8492),
.B1(n_8852),
.B2(n_8929),
.Y(n_12000)
);

NAND2xp5_ASAP7_75t_L g12001 ( 
.A(n_10530),
.B(n_8770),
.Y(n_12001)
);

NAND2xp5_ASAP7_75t_L g12002 ( 
.A(n_10547),
.B(n_10549),
.Y(n_12002)
);

AOI221xp5_ASAP7_75t_L g12003 ( 
.A1(n_10550),
.A2(n_7629),
.B1(n_7639),
.B2(n_7638),
.C(n_7618),
.Y(n_12003)
);

AOI22xp33_ASAP7_75t_L g12004 ( 
.A1(n_10645),
.A2(n_9752),
.B1(n_9839),
.B2(n_9783),
.Y(n_12004)
);

INVx1_ASAP7_75t_L g12005 ( 
.A(n_11058),
.Y(n_12005)
);

OAI22xp5_ASAP7_75t_L g12006 ( 
.A1(n_11370),
.A2(n_10376),
.B1(n_8820),
.B2(n_10364),
.Y(n_12006)
);

AOI22xp33_ASAP7_75t_L g12007 ( 
.A1(n_10645),
.A2(n_10660),
.B1(n_11041),
.B2(n_11009),
.Y(n_12007)
);

NOR2x1_ASAP7_75t_SL g12008 ( 
.A(n_11288),
.B(n_9301),
.Y(n_12008)
);

INVx1_ASAP7_75t_L g12009 ( 
.A(n_11059),
.Y(n_12009)
);

AOI21xp5_ASAP7_75t_L g12010 ( 
.A1(n_10694),
.A2(n_7486),
.B(n_9364),
.Y(n_12010)
);

OAI22xp5_ASAP7_75t_L g12011 ( 
.A1(n_11370),
.A2(n_8820),
.B1(n_9810),
.B2(n_9703),
.Y(n_12011)
);

INVx1_ASAP7_75t_L g12012 ( 
.A(n_11061),
.Y(n_12012)
);

OAI22xp33_ASAP7_75t_L g12013 ( 
.A1(n_10376),
.A2(n_11201),
.B1(n_10505),
.B2(n_11370),
.Y(n_12013)
);

OAI211xp5_ASAP7_75t_L g12014 ( 
.A1(n_10505),
.A2(n_8015),
.B(n_8601),
.C(n_8529),
.Y(n_12014)
);

HB1xp67_ASAP7_75t_L g12015 ( 
.A(n_10781),
.Y(n_12015)
);

INVx2_ASAP7_75t_L g12016 ( 
.A(n_10645),
.Y(n_12016)
);

OAI22xp5_ASAP7_75t_L g12017 ( 
.A1(n_11370),
.A2(n_9703),
.B1(n_9967),
.B2(n_9810),
.Y(n_12017)
);

INVx2_ASAP7_75t_L g12018 ( 
.A(n_10645),
.Y(n_12018)
);

AOI22xp33_ASAP7_75t_L g12019 ( 
.A1(n_10660),
.A2(n_11041),
.B1(n_11119),
.B2(n_11009),
.Y(n_12019)
);

AOI22xp33_ASAP7_75t_L g12020 ( 
.A1(n_10660),
.A2(n_9880),
.B1(n_10008),
.B2(n_9853),
.Y(n_12020)
);

AND2x2_ASAP7_75t_L g12021 ( 
.A(n_10540),
.B(n_9308),
.Y(n_12021)
);

OAI211xp5_ASAP7_75t_L g12022 ( 
.A1(n_10834),
.A2(n_8601),
.B(n_8529),
.C(n_8527),
.Y(n_12022)
);

INVx2_ASAP7_75t_L g12023 ( 
.A(n_10660),
.Y(n_12023)
);

OAI22xp33_ASAP7_75t_L g12024 ( 
.A1(n_10376),
.A2(n_8934),
.B1(n_8929),
.B2(n_8716),
.Y(n_12024)
);

OAI22xp5_ASAP7_75t_L g12025 ( 
.A1(n_10694),
.A2(n_9703),
.B1(n_9967),
.B2(n_9810),
.Y(n_12025)
);

AOI221xp5_ASAP7_75t_L g12026 ( 
.A1(n_10555),
.A2(n_7639),
.B1(n_7655),
.B2(n_7647),
.C(n_7638),
.Y(n_12026)
);

AND2x2_ASAP7_75t_L g12027 ( 
.A(n_10541),
.B(n_9308),
.Y(n_12027)
);

AOI22xp33_ASAP7_75t_SL g12028 ( 
.A1(n_11274),
.A2(n_7852),
.B1(n_8323),
.B2(n_7864),
.Y(n_12028)
);

OAI22xp5_ASAP7_75t_L g12029 ( 
.A1(n_10716),
.A2(n_9967),
.B1(n_10075),
.B2(n_9989),
.Y(n_12029)
);

BUFx12f_ASAP7_75t_L g12030 ( 
.A(n_11347),
.Y(n_12030)
);

OR2x6_ASAP7_75t_L g12031 ( 
.A(n_10716),
.B(n_8911),
.Y(n_12031)
);

AND2x2_ASAP7_75t_L g12032 ( 
.A(n_10861),
.B(n_9337),
.Y(n_12032)
);

AOI221xp5_ASAP7_75t_L g12033 ( 
.A1(n_10556),
.A2(n_7639),
.B1(n_7655),
.B2(n_7647),
.C(n_7638),
.Y(n_12033)
);

INVx4_ASAP7_75t_L g12034 ( 
.A(n_11009),
.Y(n_12034)
);

CKINVDCx6p67_ASAP7_75t_R g12035 ( 
.A(n_11015),
.Y(n_12035)
);

INVx1_ASAP7_75t_L g12036 ( 
.A(n_11062),
.Y(n_12036)
);

AOI221xp5_ASAP7_75t_L g12037 ( 
.A1(n_10807),
.A2(n_7639),
.B1(n_7655),
.B2(n_7647),
.C(n_7638),
.Y(n_12037)
);

INVx2_ASAP7_75t_SL g12038 ( 
.A(n_11009),
.Y(n_12038)
);

OR2x2_ASAP7_75t_L g12039 ( 
.A(n_10603),
.B(n_8232),
.Y(n_12039)
);

INVx1_ASAP7_75t_L g12040 ( 
.A(n_11074),
.Y(n_12040)
);

AOI22xp33_ASAP7_75t_L g12041 ( 
.A1(n_11041),
.A2(n_9880),
.B1(n_10008),
.B2(n_9853),
.Y(n_12041)
);

AOI21xp33_ASAP7_75t_L g12042 ( 
.A1(n_10835),
.A2(n_7717),
.B(n_8050),
.Y(n_12042)
);

INVx1_ASAP7_75t_L g12043 ( 
.A(n_11086),
.Y(n_12043)
);

AOI22xp33_ASAP7_75t_L g12044 ( 
.A1(n_11041),
.A2(n_9880),
.B1(n_10008),
.B2(n_9853),
.Y(n_12044)
);

INVx4_ASAP7_75t_L g12045 ( 
.A(n_11119),
.Y(n_12045)
);

AOI21xp33_ASAP7_75t_L g12046 ( 
.A1(n_10835),
.A2(n_7717),
.B(n_8050),
.Y(n_12046)
);

NOR2xp33_ASAP7_75t_L g12047 ( 
.A(n_11361),
.B(n_8911),
.Y(n_12047)
);

OAI221xp5_ASAP7_75t_L g12048 ( 
.A1(n_10716),
.A2(n_7653),
.B1(n_8592),
.B2(n_8598),
.C(n_9967),
.Y(n_12048)
);

INVx1_ASAP7_75t_L g12049 ( 
.A(n_11090),
.Y(n_12049)
);

AOI22xp33_ASAP7_75t_SL g12050 ( 
.A1(n_11274),
.A2(n_7852),
.B1(n_8323),
.B2(n_7864),
.Y(n_12050)
);

INVx2_ASAP7_75t_L g12051 ( 
.A(n_11119),
.Y(n_12051)
);

INVx1_ASAP7_75t_L g12052 ( 
.A(n_11092),
.Y(n_12052)
);

INVx2_ASAP7_75t_L g12053 ( 
.A(n_11119),
.Y(n_12053)
);

OAI22xp5_ASAP7_75t_L g12054 ( 
.A1(n_10716),
.A2(n_9967),
.B1(n_10075),
.B2(n_9989),
.Y(n_12054)
);

OAI22xp5_ASAP7_75t_L g12055 ( 
.A1(n_10861),
.A2(n_9989),
.B1(n_10166),
.B2(n_10075),
.Y(n_12055)
);

INVx1_ASAP7_75t_L g12056 ( 
.A(n_11096),
.Y(n_12056)
);

OAI22xp5_ASAP7_75t_L g12057 ( 
.A1(n_10861),
.A2(n_9989),
.B1(n_10166),
.B2(n_10075),
.Y(n_12057)
);

AOI22xp33_ASAP7_75t_L g12058 ( 
.A1(n_11180),
.A2(n_9880),
.B1(n_10008),
.B2(n_9853),
.Y(n_12058)
);

NAND3xp33_ASAP7_75t_L g12059 ( 
.A(n_11017),
.B(n_7852),
.C(n_7941),
.Y(n_12059)
);

AOI22xp33_ASAP7_75t_L g12060 ( 
.A1(n_11180),
.A2(n_11362),
.B1(n_11196),
.B2(n_10511),
.Y(n_12060)
);

INVx1_ASAP7_75t_L g12061 ( 
.A(n_11101),
.Y(n_12061)
);

AND2x2_ASAP7_75t_L g12062 ( 
.A(n_10916),
.B(n_9337),
.Y(n_12062)
);

OAI22xp5_ASAP7_75t_L g12063 ( 
.A1(n_10916),
.A2(n_9989),
.B1(n_10166),
.B2(n_10075),
.Y(n_12063)
);

BUFx2_ASAP7_75t_L g12064 ( 
.A(n_11017),
.Y(n_12064)
);

AOI221xp5_ASAP7_75t_L g12065 ( 
.A1(n_10824),
.A2(n_7647),
.B1(n_7655),
.B2(n_8853),
.C(n_8389),
.Y(n_12065)
);

INVx1_ASAP7_75t_L g12066 ( 
.A(n_11102),
.Y(n_12066)
);

AOI22xp33_ASAP7_75t_L g12067 ( 
.A1(n_11180),
.A2(n_11196),
.B1(n_11362),
.B2(n_10511),
.Y(n_12067)
);

INVx1_ASAP7_75t_L g12068 ( 
.A(n_11103),
.Y(n_12068)
);

CKINVDCx5p33_ASAP7_75t_R g12069 ( 
.A(n_11360),
.Y(n_12069)
);

AND2x2_ASAP7_75t_L g12070 ( 
.A(n_10916),
.B(n_9343),
.Y(n_12070)
);

INVx4_ASAP7_75t_L g12071 ( 
.A(n_11180),
.Y(n_12071)
);

BUFx8_ASAP7_75t_SL g12072 ( 
.A(n_11196),
.Y(n_12072)
);

OAI22xp5_ASAP7_75t_L g12073 ( 
.A1(n_10939),
.A2(n_10166),
.B1(n_8362),
.B2(n_8530),
.Y(n_12073)
);

AOI332xp33_ASAP7_75t_L g12074 ( 
.A1(n_11425),
.A2(n_10131),
.A3(n_10124),
.B1(n_10130),
.B2(n_10119),
.B3(n_10258),
.C1(n_10255),
.C2(n_10245),
.Y(n_12074)
);

AND2x2_ASAP7_75t_L g12075 ( 
.A(n_10939),
.B(n_9343),
.Y(n_12075)
);

AOI21xp5_ASAP7_75t_L g12076 ( 
.A1(n_11094),
.A2(n_10810),
.B(n_11017),
.Y(n_12076)
);

NAND3xp33_ASAP7_75t_L g12077 ( 
.A(n_11183),
.B(n_7852),
.C(n_7941),
.Y(n_12077)
);

AOI22xp5_ASAP7_75t_L g12078 ( 
.A1(n_11183),
.A2(n_8934),
.B1(n_8732),
.B2(n_8716),
.Y(n_12078)
);

INVx2_ASAP7_75t_L g12079 ( 
.A(n_11196),
.Y(n_12079)
);

BUFx4f_ASAP7_75t_SL g12080 ( 
.A(n_11362),
.Y(n_12080)
);

OAI21xp33_ASAP7_75t_L g12081 ( 
.A1(n_10603),
.A2(n_8372),
.B(n_8530),
.Y(n_12081)
);

AND2x2_ASAP7_75t_L g12082 ( 
.A(n_10939),
.B(n_9414),
.Y(n_12082)
);

BUFx2_ASAP7_75t_L g12083 ( 
.A(n_11183),
.Y(n_12083)
);

AOI22xp33_ASAP7_75t_SL g12084 ( 
.A1(n_11289),
.A2(n_7864),
.B1(n_8323),
.B2(n_7941),
.Y(n_12084)
);

NAND3xp33_ASAP7_75t_L g12085 ( 
.A(n_11291),
.B(n_7941),
.C(n_8011),
.Y(n_12085)
);

OAI221xp5_ASAP7_75t_L g12086 ( 
.A1(n_11291),
.A2(n_7653),
.B1(n_8592),
.B2(n_8598),
.C(n_10166),
.Y(n_12086)
);

AOI221xp5_ASAP7_75t_L g12087 ( 
.A1(n_10825),
.A2(n_8389),
.B1(n_8671),
.B2(n_8563),
.C(n_8050),
.Y(n_12087)
);

BUFx4f_ASAP7_75t_SL g12088 ( 
.A(n_11362),
.Y(n_12088)
);

OR2x2_ASAP7_75t_L g12089 ( 
.A(n_10891),
.B(n_8232),
.Y(n_12089)
);

AOI221xp5_ASAP7_75t_SL g12090 ( 
.A1(n_10790),
.A2(n_8838),
.B1(n_8781),
.B2(n_8585),
.C(n_8619),
.Y(n_12090)
);

NAND2xp5_ASAP7_75t_L g12091 ( 
.A(n_10839),
.B(n_8770),
.Y(n_12091)
);

OAI22xp33_ASAP7_75t_L g12092 ( 
.A1(n_10636),
.A2(n_8732),
.B1(n_8199),
.B2(n_8919),
.Y(n_12092)
);

OAI22xp5_ASAP7_75t_L g12093 ( 
.A1(n_10960),
.A2(n_8362),
.B1(n_8372),
.B2(n_8474),
.Y(n_12093)
);

AOI22xp33_ASAP7_75t_L g12094 ( 
.A1(n_10511),
.A2(n_9556),
.B1(n_9679),
.B2(n_9364),
.Y(n_12094)
);

NAND2xp5_ASAP7_75t_SL g12095 ( 
.A(n_10960),
.B(n_9257),
.Y(n_12095)
);

BUFx2_ASAP7_75t_L g12096 ( 
.A(n_11291),
.Y(n_12096)
);

AOI22xp33_ASAP7_75t_L g12097 ( 
.A1(n_10511),
.A2(n_9556),
.B1(n_9679),
.B2(n_9364),
.Y(n_12097)
);

AOI21xp5_ASAP7_75t_L g12098 ( 
.A1(n_11094),
.A2(n_9556),
.B(n_9364),
.Y(n_12098)
);

OAI21xp33_ASAP7_75t_L g12099 ( 
.A1(n_10430),
.A2(n_8339),
.B(n_8203),
.Y(n_12099)
);

AOI22xp33_ASAP7_75t_L g12100 ( 
.A1(n_10511),
.A2(n_9556),
.B1(n_9679),
.B2(n_9364),
.Y(n_12100)
);

INVx1_ASAP7_75t_SL g12101 ( 
.A(n_11365),
.Y(n_12101)
);

NOR2x1_ASAP7_75t_SL g12102 ( 
.A(n_11288),
.B(n_9414),
.Y(n_12102)
);

AOI22xp33_ASAP7_75t_L g12103 ( 
.A1(n_11325),
.A2(n_9679),
.B1(n_9742),
.B2(n_9556),
.Y(n_12103)
);

OAI22xp5_ASAP7_75t_L g12104 ( 
.A1(n_10960),
.A2(n_8919),
.B1(n_9970),
.B2(n_9370),
.Y(n_12104)
);

INVx2_ASAP7_75t_L g12105 ( 
.A(n_10298),
.Y(n_12105)
);

INVx1_ASAP7_75t_L g12106 ( 
.A(n_11113),
.Y(n_12106)
);

AOI22xp33_ASAP7_75t_L g12107 ( 
.A1(n_11325),
.A2(n_9742),
.B1(n_10113),
.B2(n_9679),
.Y(n_12107)
);

AOI22xp33_ASAP7_75t_L g12108 ( 
.A1(n_11325),
.A2(n_10113),
.B1(n_10180),
.B2(n_9742),
.Y(n_12108)
);

OAI22xp5_ASAP7_75t_L g12109 ( 
.A1(n_11021),
.A2(n_9970),
.B1(n_9595),
.B2(n_9623),
.Y(n_12109)
);

OAI211xp5_ASAP7_75t_L g12110 ( 
.A1(n_10675),
.A2(n_8527),
.B(n_8616),
.C(n_8011),
.Y(n_12110)
);

AOI22xp33_ASAP7_75t_L g12111 ( 
.A1(n_11021),
.A2(n_10113),
.B1(n_10180),
.B2(n_9742),
.Y(n_12111)
);

AND2x4_ASAP7_75t_L g12112 ( 
.A(n_10650),
.B(n_9970),
.Y(n_12112)
);

AOI33xp33_ASAP7_75t_L g12113 ( 
.A1(n_10675),
.A2(n_8671),
.A3(n_8563),
.B1(n_10190),
.B2(n_10193),
.B3(n_10188),
.Y(n_12113)
);

HB1xp67_ASAP7_75t_L g12114 ( 
.A(n_10870),
.Y(n_12114)
);

OAI22xp33_ASAP7_75t_L g12115 ( 
.A1(n_10872),
.A2(n_8199),
.B1(n_8946),
.B2(n_8010),
.Y(n_12115)
);

INVx1_ASAP7_75t_L g12116 ( 
.A(n_11114),
.Y(n_12116)
);

AOI221xp5_ASAP7_75t_L g12117 ( 
.A1(n_10876),
.A2(n_8050),
.B1(n_10056),
.B2(n_9947),
.C(n_9976),
.Y(n_12117)
);

AOI22xp33_ASAP7_75t_L g12118 ( 
.A1(n_11021),
.A2(n_10113),
.B1(n_10180),
.B2(n_9742),
.Y(n_12118)
);

OAI22xp5_ASAP7_75t_L g12119 ( 
.A1(n_11302),
.A2(n_9357),
.B1(n_8636),
.B2(n_8751),
.Y(n_12119)
);

OAI211xp5_ASAP7_75t_L g12120 ( 
.A1(n_10793),
.A2(n_8616),
.B(n_8011),
.C(n_7941),
.Y(n_12120)
);

OAI22xp5_ASAP7_75t_L g12121 ( 
.A1(n_11302),
.A2(n_8636),
.B1(n_8751),
.B2(n_8628),
.Y(n_12121)
);

NOR2xp33_ASAP7_75t_L g12122 ( 
.A(n_10650),
.B(n_8911),
.Y(n_12122)
);

AND2x2_ASAP7_75t_L g12123 ( 
.A(n_11302),
.B(n_9452),
.Y(n_12123)
);

AOI22xp33_ASAP7_75t_L g12124 ( 
.A1(n_11318),
.A2(n_10180),
.B1(n_10113),
.B2(n_7717),
.Y(n_12124)
);

OAI22xp5_ASAP7_75t_L g12125 ( 
.A1(n_11318),
.A2(n_8628),
.B1(n_7936),
.B2(n_8143),
.Y(n_12125)
);

NAND3xp33_ASAP7_75t_L g12126 ( 
.A(n_10900),
.B(n_7941),
.C(n_8011),
.Y(n_12126)
);

INVx4_ASAP7_75t_L g12127 ( 
.A(n_10650),
.Y(n_12127)
);

AOI22xp33_ASAP7_75t_L g12128 ( 
.A1(n_11318),
.A2(n_10180),
.B1(n_7717),
.B2(n_8914),
.Y(n_12128)
);

INVx1_ASAP7_75t_L g12129 ( 
.A(n_11115),
.Y(n_12129)
);

AOI22xp33_ASAP7_75t_L g12130 ( 
.A1(n_11324),
.A2(n_8790),
.B1(n_8914),
.B2(n_8849),
.Y(n_12130)
);

AOI22xp33_ASAP7_75t_L g12131 ( 
.A1(n_11324),
.A2(n_8914),
.B1(n_8791),
.B2(n_8849),
.Y(n_12131)
);

OA21x2_ASAP7_75t_L g12132 ( 
.A1(n_10984),
.A2(n_9170),
.B(n_10124),
.Y(n_12132)
);

INVx2_ASAP7_75t_L g12133 ( 
.A(n_10298),
.Y(n_12133)
);

INVx1_ASAP7_75t_L g12134 ( 
.A(n_11123),
.Y(n_12134)
);

BUFx12f_ASAP7_75t_L g12135 ( 
.A(n_11324),
.Y(n_12135)
);

OAI211xp5_ASAP7_75t_SL g12136 ( 
.A1(n_11367),
.A2(n_8283),
.B(n_8327),
.C(n_8276),
.Y(n_12136)
);

OAI22xp5_ASAP7_75t_L g12137 ( 
.A1(n_11398),
.A2(n_7936),
.B1(n_8143),
.B2(n_8010),
.Y(n_12137)
);

OAI21x1_ASAP7_75t_L g12138 ( 
.A1(n_10595),
.A2(n_10266),
.B(n_10248),
.Y(n_12138)
);

INVx1_ASAP7_75t_L g12139 ( 
.A(n_11125),
.Y(n_12139)
);

AOI22xp33_ASAP7_75t_L g12140 ( 
.A1(n_11398),
.A2(n_8791),
.B1(n_8849),
.B2(n_8203),
.Y(n_12140)
);

OAI21x1_ASAP7_75t_L g12141 ( 
.A1(n_10595),
.A2(n_10266),
.B(n_9278),
.Y(n_12141)
);

NAND3xp33_ASAP7_75t_L g12142 ( 
.A(n_10905),
.B(n_8011),
.C(n_8709),
.Y(n_12142)
);

INVx1_ASAP7_75t_L g12143 ( 
.A(n_11127),
.Y(n_12143)
);

INVx1_ASAP7_75t_L g12144 ( 
.A(n_11128),
.Y(n_12144)
);

INVx1_ASAP7_75t_L g12145 ( 
.A(n_11131),
.Y(n_12145)
);

OAI22xp5_ASAP7_75t_L g12146 ( 
.A1(n_11398),
.A2(n_7936),
.B1(n_8143),
.B2(n_8010),
.Y(n_12146)
);

OAI22xp33_ASAP7_75t_L g12147 ( 
.A1(n_10911),
.A2(n_8199),
.B1(n_8946),
.B2(n_8191),
.Y(n_12147)
);

OAI221xp5_ASAP7_75t_L g12148 ( 
.A1(n_11082),
.A2(n_8076),
.B1(n_8191),
.B2(n_8193),
.C(n_8170),
.Y(n_12148)
);

AOI22xp33_ASAP7_75t_L g12149 ( 
.A1(n_11414),
.A2(n_8849),
.B1(n_7969),
.B2(n_8191),
.Y(n_12149)
);

AOI22xp33_ASAP7_75t_L g12150 ( 
.A1(n_11414),
.A2(n_7969),
.B1(n_8193),
.B2(n_8170),
.Y(n_12150)
);

INVx2_ASAP7_75t_L g12151 ( 
.A(n_10298),
.Y(n_12151)
);

INVx2_ASAP7_75t_SL g12152 ( 
.A(n_11414),
.Y(n_12152)
);

INVx2_ASAP7_75t_L g12153 ( 
.A(n_10328),
.Y(n_12153)
);

OR2x6_ASAP7_75t_L g12154 ( 
.A(n_10793),
.B(n_6592),
.Y(n_12154)
);

AOI21xp5_ASAP7_75t_L g12155 ( 
.A1(n_10810),
.A2(n_10244),
.B(n_10040),
.Y(n_12155)
);

AOI22xp33_ASAP7_75t_L g12156 ( 
.A1(n_11289),
.A2(n_7969),
.B1(n_8193),
.B2(n_8170),
.Y(n_12156)
);

AOI221xp5_ASAP7_75t_L g12157 ( 
.A1(n_10917),
.A2(n_10056),
.B1(n_9976),
.B2(n_9947),
.C(n_8352),
.Y(n_12157)
);

AOI22xp33_ASAP7_75t_SL g12158 ( 
.A1(n_10810),
.A2(n_8194),
.B1(n_8206),
.B2(n_8183),
.Y(n_12158)
);

OA21x2_ASAP7_75t_L g12159 ( 
.A1(n_10984),
.A2(n_10131),
.B(n_10130),
.Y(n_12159)
);

OAI22xp5_ASAP7_75t_L g12160 ( 
.A1(n_10620),
.A2(n_10670),
.B1(n_10658),
.B2(n_8245),
.Y(n_12160)
);

INVx1_ASAP7_75t_L g12161 ( 
.A(n_11132),
.Y(n_12161)
);

INVx2_ASAP7_75t_L g12162 ( 
.A(n_10328),
.Y(n_12162)
);

AO21x2_ASAP7_75t_L g12163 ( 
.A1(n_11374),
.A2(n_9722),
.B(n_9707),
.Y(n_12163)
);

NAND2xp5_ASAP7_75t_L g12164 ( 
.A(n_10950),
.B(n_8662),
.Y(n_12164)
);

OAI22xp5_ASAP7_75t_L g12165 ( 
.A1(n_10620),
.A2(n_8245),
.B1(n_8354),
.B2(n_8242),
.Y(n_12165)
);

NAND2xp5_ASAP7_75t_L g12166 ( 
.A(n_11001),
.B(n_8662),
.Y(n_12166)
);

NAND2x1_ASAP7_75t_L g12167 ( 
.A(n_10328),
.B(n_10334),
.Y(n_12167)
);

NAND2xp5_ASAP7_75t_L g12168 ( 
.A(n_11010),
.B(n_8705),
.Y(n_12168)
);

BUFx2_ASAP7_75t_L g12169 ( 
.A(n_11126),
.Y(n_12169)
);

AOI22xp33_ASAP7_75t_L g12170 ( 
.A1(n_10620),
.A2(n_7969),
.B1(n_8245),
.B2(n_8242),
.Y(n_12170)
);

INVx1_ASAP7_75t_SL g12171 ( 
.A(n_10790),
.Y(n_12171)
);

AND2x4_ASAP7_75t_L g12172 ( 
.A(n_10658),
.B(n_9011),
.Y(n_12172)
);

AO221x2_ASAP7_75t_L g12173 ( 
.A1(n_11424),
.A2(n_8368),
.B1(n_9722),
.B2(n_9765),
.C(n_9707),
.Y(n_12173)
);

OAI222xp33_ASAP7_75t_L g12174 ( 
.A1(n_10663),
.A2(n_8621),
.B1(n_8619),
.B2(n_9015),
.C1(n_9079),
.C2(n_8973),
.Y(n_12174)
);

AOI22xp33_ASAP7_75t_L g12175 ( 
.A1(n_10670),
.A2(n_7969),
.B1(n_8354),
.B2(n_8242),
.Y(n_12175)
);

NOR2xp33_ASAP7_75t_L g12176 ( 
.A(n_10891),
.B(n_7381),
.Y(n_12176)
);

INVx2_ASAP7_75t_L g12177 ( 
.A(n_10334),
.Y(n_12177)
);

AOI22xp33_ASAP7_75t_L g12178 ( 
.A1(n_10670),
.A2(n_7969),
.B1(n_8461),
.B2(n_8354),
.Y(n_12178)
);

AOI21x1_ASAP7_75t_L g12179 ( 
.A1(n_10801),
.A2(n_9519),
.B(n_9516),
.Y(n_12179)
);

INVx1_ASAP7_75t_L g12180 ( 
.A(n_11133),
.Y(n_12180)
);

OAI33xp33_ASAP7_75t_L g12181 ( 
.A1(n_11138),
.A2(n_10259),
.A3(n_10255),
.B1(n_10260),
.B2(n_10258),
.B3(n_10245),
.Y(n_12181)
);

OAI221xp5_ASAP7_75t_L g12182 ( 
.A1(n_11160),
.A2(n_8710),
.B1(n_8603),
.B2(n_8461),
.C(n_8378),
.Y(n_12182)
);

INVx1_ASAP7_75t_L g12183 ( 
.A(n_11139),
.Y(n_12183)
);

OR2x2_ASAP7_75t_L g12184 ( 
.A(n_11057),
.B(n_8276),
.Y(n_12184)
);

AO21x2_ASAP7_75t_L g12185 ( 
.A1(n_11374),
.A2(n_9722),
.B(n_9707),
.Y(n_12185)
);

AOI22xp33_ASAP7_75t_L g12186 ( 
.A1(n_10658),
.A2(n_7969),
.B1(n_8603),
.B2(n_8461),
.Y(n_12186)
);

AOI22xp33_ASAP7_75t_L g12187 ( 
.A1(n_10903),
.A2(n_8603),
.B1(n_8710),
.B2(n_8673),
.Y(n_12187)
);

INVx1_ASAP7_75t_L g12188 ( 
.A(n_11140),
.Y(n_12188)
);

OAI22xp5_ASAP7_75t_L g12189 ( 
.A1(n_11210),
.A2(n_8710),
.B1(n_8357),
.B2(n_8051),
.Y(n_12189)
);

NAND4xp25_ASAP7_75t_L g12190 ( 
.A(n_10801),
.B(n_8709),
.C(n_8365),
.D(n_8378),
.Y(n_12190)
);

AOI22xp33_ASAP7_75t_L g12191 ( 
.A1(n_10903),
.A2(n_8673),
.B1(n_8409),
.B2(n_9011),
.Y(n_12191)
);

INVx1_ASAP7_75t_L g12192 ( 
.A(n_11146),
.Y(n_12192)
);

AOI22xp33_ASAP7_75t_L g12193 ( 
.A1(n_10912),
.A2(n_8673),
.B1(n_8409),
.B2(n_9011),
.Y(n_12193)
);

AOI22xp33_ASAP7_75t_L g12194 ( 
.A1(n_10912),
.A2(n_8673),
.B1(n_8409),
.B2(n_10935),
.Y(n_12194)
);

AOI22xp5_ASAP7_75t_SL g12195 ( 
.A1(n_11233),
.A2(n_7564),
.B1(n_7542),
.B2(n_9960),
.Y(n_12195)
);

AND2x4_ASAP7_75t_L g12196 ( 
.A(n_10935),
.B(n_9011),
.Y(n_12196)
);

BUFx2_ASAP7_75t_L g12197 ( 
.A(n_11240),
.Y(n_12197)
);

OAI22xp33_ASAP7_75t_L g12198 ( 
.A1(n_10663),
.A2(n_8621),
.B1(n_8194),
.B2(n_8206),
.Y(n_12198)
);

AOI221xp5_ASAP7_75t_L g12199 ( 
.A1(n_10601),
.A2(n_10056),
.B1(n_9976),
.B2(n_9947),
.C(n_8352),
.Y(n_12199)
);

AOI221xp5_ASAP7_75t_L g12200 ( 
.A1(n_10608),
.A2(n_10056),
.B1(n_9976),
.B2(n_9947),
.C(n_8439),
.Y(n_12200)
);

AOI21xp33_ASAP7_75t_L g12201 ( 
.A1(n_10617),
.A2(n_8157),
.B(n_8192),
.Y(n_12201)
);

BUFx12f_ASAP7_75t_L g12202 ( 
.A(n_10948),
.Y(n_12202)
);

CKINVDCx20_ASAP7_75t_R g12203 ( 
.A(n_11393),
.Y(n_12203)
);

AOI22xp5_ASAP7_75t_L g12204 ( 
.A1(n_10948),
.A2(n_9136),
.B1(n_9199),
.B2(n_9047),
.Y(n_12204)
);

INVx1_ASAP7_75t_L g12205 ( 
.A(n_11150),
.Y(n_12205)
);

OAI22xp5_ASAP7_75t_L g12206 ( 
.A1(n_10630),
.A2(n_8357),
.B1(n_8051),
.B2(n_7761),
.Y(n_12206)
);

INVx1_ASAP7_75t_L g12207 ( 
.A(n_11151),
.Y(n_12207)
);

OAI22xp5_ASAP7_75t_L g12208 ( 
.A1(n_10680),
.A2(n_8357),
.B1(n_8051),
.B2(n_7761),
.Y(n_12208)
);

AOI22xp33_ASAP7_75t_L g12209 ( 
.A1(n_10552),
.A2(n_8673),
.B1(n_8409),
.B2(n_9047),
.Y(n_12209)
);

OAI22xp5_ASAP7_75t_L g12210 ( 
.A1(n_10745),
.A2(n_8357),
.B1(n_8051),
.B2(n_7761),
.Y(n_12210)
);

AOI22xp5_ASAP7_75t_L g12211 ( 
.A1(n_10589),
.A2(n_9136),
.B1(n_9199),
.B2(n_9047),
.Y(n_12211)
);

BUFx3_ASAP7_75t_L g12212 ( 
.A(n_10637),
.Y(n_12212)
);

AOI22xp33_ASAP7_75t_SL g12213 ( 
.A1(n_10968),
.A2(n_8194),
.B1(n_8206),
.B2(n_8183),
.Y(n_12213)
);

AOI22xp33_ASAP7_75t_SL g12214 ( 
.A1(n_10968),
.A2(n_8194),
.B1(n_8206),
.B2(n_8183),
.Y(n_12214)
);

OAI221xp5_ASAP7_75t_L g12215 ( 
.A1(n_10676),
.A2(n_8381),
.B1(n_8391),
.B2(n_8365),
.C(n_8222),
.Y(n_12215)
);

AOI22xp33_ASAP7_75t_SL g12216 ( 
.A1(n_10898),
.A2(n_8194),
.B1(n_8206),
.B2(n_8183),
.Y(n_12216)
);

BUFx2_ASAP7_75t_L g12217 ( 
.A(n_11393),
.Y(n_12217)
);

INVx5_ASAP7_75t_SL g12218 ( 
.A(n_11085),
.Y(n_12218)
);

AND2x2_ASAP7_75t_L g12219 ( 
.A(n_11408),
.B(n_9452),
.Y(n_12219)
);

AOI221xp5_ASAP7_75t_L g12220 ( 
.A1(n_11395),
.A2(n_8368),
.B1(n_8809),
.B2(n_8075),
.C(n_8068),
.Y(n_12220)
);

AOI22xp5_ASAP7_75t_L g12221 ( 
.A1(n_10589),
.A2(n_9136),
.B1(n_9199),
.B2(n_9047),
.Y(n_12221)
);

INVx4_ASAP7_75t_SL g12222 ( 
.A(n_10567),
.Y(n_12222)
);

NAND2xp5_ASAP7_75t_L g12223 ( 
.A(n_11057),
.B(n_8705),
.Y(n_12223)
);

CKINVDCx5p33_ASAP7_75t_R g12224 ( 
.A(n_10334),
.Y(n_12224)
);

AND2x2_ASAP7_75t_L g12225 ( 
.A(n_11408),
.B(n_9499),
.Y(n_12225)
);

AOI22xp33_ASAP7_75t_L g12226 ( 
.A1(n_10552),
.A2(n_8409),
.B1(n_9199),
.B2(n_9136),
.Y(n_12226)
);

AOI22xp33_ASAP7_75t_L g12227 ( 
.A1(n_10565),
.A2(n_9254),
.B1(n_9407),
.B2(n_9227),
.Y(n_12227)
);

INVx3_ASAP7_75t_L g12228 ( 
.A(n_10398),
.Y(n_12228)
);

AO21x2_ASAP7_75t_L g12229 ( 
.A1(n_11085),
.A2(n_9766),
.B(n_9765),
.Y(n_12229)
);

OAI221xp5_ASAP7_75t_L g12230 ( 
.A1(n_10766),
.A2(n_8391),
.B1(n_8381),
.B2(n_8222),
.C(n_8809),
.Y(n_12230)
);

INVx1_ASAP7_75t_L g12231 ( 
.A(n_11156),
.Y(n_12231)
);

HB1xp67_ASAP7_75t_L g12232 ( 
.A(n_11395),
.Y(n_12232)
);

AND2x2_ASAP7_75t_L g12233 ( 
.A(n_11294),
.B(n_9499),
.Y(n_12233)
);

OAI21x1_ASAP7_75t_L g12234 ( 
.A1(n_10335),
.A2(n_10619),
.B(n_10616),
.Y(n_12234)
);

HB1xp67_ASAP7_75t_L g12235 ( 
.A(n_11401),
.Y(n_12235)
);

NOR2xp33_ASAP7_75t_L g12236 ( 
.A(n_11407),
.B(n_8747),
.Y(n_12236)
);

INVx1_ASAP7_75t_L g12237 ( 
.A(n_11159),
.Y(n_12237)
);

INVx2_ASAP7_75t_SL g12238 ( 
.A(n_10398),
.Y(n_12238)
);

AOI22xp33_ASAP7_75t_L g12239 ( 
.A1(n_10565),
.A2(n_9254),
.B1(n_9407),
.B2(n_9227),
.Y(n_12239)
);

AOI21xp5_ASAP7_75t_L g12240 ( 
.A1(n_11085),
.A2(n_8455),
.B(n_8425),
.Y(n_12240)
);

AOI222xp33_ASAP7_75t_L g12241 ( 
.A1(n_11401),
.A2(n_7901),
.B1(n_8333),
.B2(n_7642),
.C1(n_10193),
.C2(n_10190),
.Y(n_12241)
);

INVx1_ASAP7_75t_L g12242 ( 
.A(n_11163),
.Y(n_12242)
);

AOI22xp33_ASAP7_75t_L g12243 ( 
.A1(n_10577),
.A2(n_9254),
.B1(n_9407),
.B2(n_9227),
.Y(n_12243)
);

BUFx2_ASAP7_75t_L g12244 ( 
.A(n_10898),
.Y(n_12244)
);

AOI21xp33_ASAP7_75t_L g12245 ( 
.A1(n_11170),
.A2(n_8157),
.B(n_8192),
.Y(n_12245)
);

INVx1_ASAP7_75t_L g12246 ( 
.A(n_11176),
.Y(n_12246)
);

OAI22xp5_ASAP7_75t_L g12247 ( 
.A1(n_11295),
.A2(n_8357),
.B1(n_8051),
.B2(n_7761),
.Y(n_12247)
);

INVx2_ASAP7_75t_L g12248 ( 
.A(n_10398),
.Y(n_12248)
);

AO21x2_ASAP7_75t_L g12249 ( 
.A1(n_11402),
.A2(n_9766),
.B(n_9765),
.Y(n_12249)
);

AND2x4_ASAP7_75t_L g12250 ( 
.A(n_10989),
.B(n_9227),
.Y(n_12250)
);

INVx1_ASAP7_75t_L g12251 ( 
.A(n_11177),
.Y(n_12251)
);

AOI22xp33_ASAP7_75t_L g12252 ( 
.A1(n_10577),
.A2(n_9407),
.B1(n_9520),
.B2(n_9254),
.Y(n_12252)
);

BUFx12f_ASAP7_75t_L g12253 ( 
.A(n_10585),
.Y(n_12253)
);

A2O1A1Ixp33_ASAP7_75t_L g12254 ( 
.A1(n_10619),
.A2(n_10178),
.B(n_10097),
.C(n_9040),
.Y(n_12254)
);

OAI21x1_ASAP7_75t_SL g12255 ( 
.A1(n_11426),
.A2(n_8738),
.B(n_8371),
.Y(n_12255)
);

AOI22xp33_ASAP7_75t_L g12256 ( 
.A1(n_10585),
.A2(n_9527),
.B1(n_9542),
.B2(n_9520),
.Y(n_12256)
);

AOI221xp5_ASAP7_75t_L g12257 ( 
.A1(n_11402),
.A2(n_8075),
.B1(n_8068),
.B2(n_10017),
.C(n_8123),
.Y(n_12257)
);

AOI22xp33_ASAP7_75t_SL g12258 ( 
.A1(n_10901),
.A2(n_8194),
.B1(n_8206),
.B2(n_8183),
.Y(n_12258)
);

AOI21xp33_ASAP7_75t_SL g12259 ( 
.A1(n_10410),
.A2(n_7281),
.B(n_7259),
.Y(n_12259)
);

AOI221xp5_ASAP7_75t_L g12260 ( 
.A1(n_11405),
.A2(n_8075),
.B1(n_8068),
.B2(n_10017),
.C(n_8123),
.Y(n_12260)
);

OAI222xp33_ASAP7_75t_L g12261 ( 
.A1(n_10696),
.A2(n_9015),
.B1(n_9079),
.B2(n_8973),
.C1(n_9561),
.C2(n_7811),
.Y(n_12261)
);

NAND2xp5_ASAP7_75t_L g12262 ( 
.A(n_11428),
.B(n_8413),
.Y(n_12262)
);

BUFx12f_ASAP7_75t_L g12263 ( 
.A(n_10644),
.Y(n_12263)
);

OR2x2_ASAP7_75t_L g12264 ( 
.A(n_11427),
.B(n_8283),
.Y(n_12264)
);

OAI22xp33_ASAP7_75t_L g12265 ( 
.A1(n_10696),
.A2(n_8210),
.B1(n_8239),
.B2(n_8183),
.Y(n_12265)
);

OR2x2_ASAP7_75t_L g12266 ( 
.A(n_11427),
.B(n_8327),
.Y(n_12266)
);

INVx2_ASAP7_75t_L g12267 ( 
.A(n_10410),
.Y(n_12267)
);

BUFx6f_ASAP7_75t_L g12268 ( 
.A(n_10410),
.Y(n_12268)
);

INVx2_ASAP7_75t_L g12269 ( 
.A(n_10446),
.Y(n_12269)
);

NAND2xp5_ASAP7_75t_L g12270 ( 
.A(n_11407),
.B(n_8413),
.Y(n_12270)
);

INVx1_ASAP7_75t_L g12271 ( 
.A(n_11178),
.Y(n_12271)
);

CKINVDCx8_ASAP7_75t_R g12272 ( 
.A(n_10599),
.Y(n_12272)
);

AOI221xp5_ASAP7_75t_L g12273 ( 
.A1(n_11405),
.A2(n_8075),
.B1(n_8068),
.B2(n_10017),
.C(n_8123),
.Y(n_12273)
);

HB1xp67_ASAP7_75t_L g12274 ( 
.A(n_11406),
.Y(n_12274)
);

BUFx3_ASAP7_75t_L g12275 ( 
.A(n_10644),
.Y(n_12275)
);

AOI21xp5_ASAP7_75t_L g12276 ( 
.A1(n_10609),
.A2(n_8467),
.B(n_8425),
.Y(n_12276)
);

AOI22xp33_ASAP7_75t_L g12277 ( 
.A1(n_10714),
.A2(n_9527),
.B1(n_9542),
.B2(n_9520),
.Y(n_12277)
);

AO31x2_ASAP7_75t_L g12278 ( 
.A1(n_11406),
.A2(n_9770),
.A3(n_9771),
.B(n_9766),
.Y(n_12278)
);

INVx2_ASAP7_75t_L g12279 ( 
.A(n_10446),
.Y(n_12279)
);

OAI22xp5_ASAP7_75t_L g12280 ( 
.A1(n_11295),
.A2(n_8357),
.B1(n_8051),
.B2(n_7761),
.Y(n_12280)
);

INVx1_ASAP7_75t_L g12281 ( 
.A(n_11184),
.Y(n_12281)
);

NOR2xp33_ASAP7_75t_SL g12282 ( 
.A(n_10714),
.B(n_7255),
.Y(n_12282)
);

INVx4_ASAP7_75t_L g12283 ( 
.A(n_10446),
.Y(n_12283)
);

OAI22xp33_ASAP7_75t_L g12284 ( 
.A1(n_11300),
.A2(n_8210),
.B1(n_8239),
.B2(n_7314),
.Y(n_12284)
);

AOI222xp33_ASAP7_75t_L g12285 ( 
.A1(n_11415),
.A2(n_7901),
.B1(n_8333),
.B2(n_7642),
.C1(n_9659),
.C2(n_9523),
.Y(n_12285)
);

OA21x2_ASAP7_75t_L g12286 ( 
.A1(n_11397),
.A2(n_9236),
.B(n_9274),
.Y(n_12286)
);

AOI22xp33_ASAP7_75t_L g12287 ( 
.A1(n_10767),
.A2(n_9527),
.B1(n_9542),
.B2(n_9520),
.Y(n_12287)
);

BUFx3_ASAP7_75t_L g12288 ( 
.A(n_10767),
.Y(n_12288)
);

BUFx3_ASAP7_75t_L g12289 ( 
.A(n_10778),
.Y(n_12289)
);

OAI22xp33_ASAP7_75t_L g12290 ( 
.A1(n_11300),
.A2(n_8210),
.B1(n_8239),
.B2(n_7314),
.Y(n_12290)
);

AOI22xp33_ASAP7_75t_L g12291 ( 
.A1(n_10778),
.A2(n_9542),
.B1(n_9608),
.B2(n_9527),
.Y(n_12291)
);

INVx1_ASAP7_75t_SL g12292 ( 
.A(n_10789),
.Y(n_12292)
);

INVx1_ASAP7_75t_L g12293 ( 
.A(n_11189),
.Y(n_12293)
);

INVx4_ASAP7_75t_L g12294 ( 
.A(n_10544),
.Y(n_12294)
);

AOI21xp33_ASAP7_75t_L g12295 ( 
.A1(n_11190),
.A2(n_8157),
.B(n_8192),
.Y(n_12295)
);

AOI22xp33_ASAP7_75t_SL g12296 ( 
.A1(n_10901),
.A2(n_8239),
.B1(n_8210),
.B2(n_8837),
.Y(n_12296)
);

OR2x2_ASAP7_75t_L g12297 ( 
.A(n_11428),
.B(n_8174),
.Y(n_12297)
);

NOR2xp67_ASAP7_75t_L g12298 ( 
.A(n_10544),
.B(n_9682),
.Y(n_12298)
);

OAI22xp33_ASAP7_75t_L g12299 ( 
.A1(n_11308),
.A2(n_8210),
.B1(n_8239),
.B2(n_7314),
.Y(n_12299)
);

AOI22xp5_ASAP7_75t_L g12300 ( 
.A1(n_10789),
.A2(n_9619),
.B1(n_9714),
.B2(n_9608),
.Y(n_12300)
);

AOI22xp5_ASAP7_75t_L g12301 ( 
.A1(n_11340),
.A2(n_9619),
.B1(n_9714),
.B2(n_9608),
.Y(n_12301)
);

INVx1_ASAP7_75t_L g12302 ( 
.A(n_11192),
.Y(n_12302)
);

AND2x4_ASAP7_75t_L g12303 ( 
.A(n_10989),
.B(n_11294),
.Y(n_12303)
);

OAI22xp5_ASAP7_75t_L g12304 ( 
.A1(n_11308),
.A2(n_8392),
.B1(n_8454),
.B2(n_7761),
.Y(n_12304)
);

INVx3_ASAP7_75t_L g12305 ( 
.A(n_10544),
.Y(n_12305)
);

AOI21xp33_ASAP7_75t_L g12306 ( 
.A1(n_11195),
.A2(n_8157),
.B(n_8192),
.Y(n_12306)
);

AO21x2_ASAP7_75t_L g12307 ( 
.A1(n_11415),
.A2(n_9771),
.B(n_9770),
.Y(n_12307)
);

AOI21x1_ASAP7_75t_L g12308 ( 
.A1(n_11420),
.A2(n_9700),
.B(n_9687),
.Y(n_12308)
);

NAND2xp5_ASAP7_75t_L g12309 ( 
.A(n_11111),
.B(n_9716),
.Y(n_12309)
);

OAI22xp5_ASAP7_75t_L g12310 ( 
.A1(n_11310),
.A2(n_8454),
.B1(n_8649),
.B2(n_8392),
.Y(n_12310)
);

OAI21xp33_ASAP7_75t_L g12311 ( 
.A1(n_11111),
.A2(n_8186),
.B(n_8174),
.Y(n_12311)
);

INVx1_ASAP7_75t_L g12312 ( 
.A(n_11199),
.Y(n_12312)
);

NOR2xp33_ASAP7_75t_L g12313 ( 
.A(n_11186),
.B(n_6592),
.Y(n_12313)
);

AOI22xp33_ASAP7_75t_L g12314 ( 
.A1(n_11340),
.A2(n_9619),
.B1(n_9714),
.B2(n_9608),
.Y(n_12314)
);

BUFx3_ASAP7_75t_L g12315 ( 
.A(n_10605),
.Y(n_12315)
);

AOI33xp33_ASAP7_75t_L g12316 ( 
.A1(n_11441),
.A2(n_8541),
.A3(n_8573),
.B1(n_8590),
.B2(n_8565),
.B3(n_9770),
.Y(n_12316)
);

INVx1_ASAP7_75t_L g12317 ( 
.A(n_11202),
.Y(n_12317)
);

OAI22xp33_ASAP7_75t_L g12318 ( 
.A1(n_11310),
.A2(n_8239),
.B1(n_8210),
.B2(n_8641),
.Y(n_12318)
);

AO222x2_ASAP7_75t_L g12319 ( 
.A1(n_10567),
.A2(n_8333),
.B1(n_7642),
.B2(n_7901),
.C1(n_9714),
.C2(n_9619),
.Y(n_12319)
);

OAI21xp33_ASAP7_75t_L g12320 ( 
.A1(n_11186),
.A2(n_8186),
.B(n_8189),
.Y(n_12320)
);

INVx4_ASAP7_75t_L g12321 ( 
.A(n_10605),
.Y(n_12321)
);

OAI22xp5_ASAP7_75t_L g12322 ( 
.A1(n_11317),
.A2(n_8454),
.B1(n_8649),
.B2(n_8392),
.Y(n_12322)
);

INVxp67_ASAP7_75t_L g12323 ( 
.A(n_11203),
.Y(n_12323)
);

AOI22xp33_ASAP7_75t_L g12324 ( 
.A1(n_11343),
.A2(n_9750),
.B1(n_11375),
.B2(n_11356),
.Y(n_12324)
);

CKINVDCx5p33_ASAP7_75t_R g12325 ( 
.A(n_10605),
.Y(n_12325)
);

AOI21xp33_ASAP7_75t_L g12326 ( 
.A1(n_11215),
.A2(n_11220),
.B(n_11218),
.Y(n_12326)
);

AND2x4_ASAP7_75t_L g12327 ( 
.A(n_11309),
.B(n_9750),
.Y(n_12327)
);

INVx1_ASAP7_75t_L g12328 ( 
.A(n_11224),
.Y(n_12328)
);

OR2x2_ASAP7_75t_L g12329 ( 
.A(n_11225),
.B(n_11237),
.Y(n_12329)
);

INVx1_ASAP7_75t_L g12330 ( 
.A(n_11228),
.Y(n_12330)
);

INVx1_ASAP7_75t_L g12331 ( 
.A(n_11232),
.Y(n_12331)
);

AOI221xp5_ASAP7_75t_L g12332 ( 
.A1(n_11420),
.A2(n_8075),
.B1(n_10017),
.B2(n_8123),
.C(n_8509),
.Y(n_12332)
);

AOI22xp33_ASAP7_75t_L g12333 ( 
.A1(n_11343),
.A2(n_9750),
.B1(n_8392),
.B2(n_8649),
.Y(n_12333)
);

INVx2_ASAP7_75t_L g12334 ( 
.A(n_10639),
.Y(n_12334)
);

OAI22xp33_ASAP7_75t_L g12335 ( 
.A1(n_11317),
.A2(n_8711),
.B1(n_8798),
.B2(n_8641),
.Y(n_12335)
);

NAND2xp33_ASAP7_75t_L g12336 ( 
.A(n_10766),
.B(n_7259),
.Y(n_12336)
);

HB1xp67_ASAP7_75t_L g12337 ( 
.A(n_11424),
.Y(n_12337)
);

AOI21xp5_ASAP7_75t_L g12338 ( 
.A1(n_10609),
.A2(n_8467),
.B(n_9750),
.Y(n_12338)
);

AO21x2_ASAP7_75t_L g12339 ( 
.A1(n_11425),
.A2(n_9779),
.B(n_9771),
.Y(n_12339)
);

OAI21xp5_ASAP7_75t_L g12340 ( 
.A1(n_10335),
.A2(n_10097),
.B(n_9218),
.Y(n_12340)
);

BUFx12f_ASAP7_75t_L g12341 ( 
.A(n_10721),
.Y(n_12341)
);

INVx3_ASAP7_75t_L g12342 ( 
.A(n_10639),
.Y(n_12342)
);

AOI22xp33_ASAP7_75t_L g12343 ( 
.A1(n_11356),
.A2(n_8392),
.B1(n_8649),
.B2(n_8454),
.Y(n_12343)
);

AOI22xp33_ASAP7_75t_L g12344 ( 
.A1(n_11375),
.A2(n_8392),
.B1(n_8649),
.B2(n_8454),
.Y(n_12344)
);

AOI22xp5_ASAP7_75t_L g12345 ( 
.A1(n_11376),
.A2(n_9561),
.B1(n_8359),
.B2(n_7823),
.Y(n_12345)
);

OAI211xp5_ASAP7_75t_L g12346 ( 
.A1(n_11426),
.A2(n_8011),
.B(n_7951),
.C(n_7980),
.Y(n_12346)
);

OR2x2_ASAP7_75t_L g12347 ( 
.A(n_11225),
.B(n_8464),
.Y(n_12347)
);

AOI22xp33_ASAP7_75t_L g12348 ( 
.A1(n_11376),
.A2(n_8454),
.B1(n_8649),
.B2(n_7930),
.Y(n_12348)
);

AO21x2_ASAP7_75t_L g12349 ( 
.A1(n_11429),
.A2(n_9784),
.B(n_9779),
.Y(n_12349)
);

AOI22xp33_ASAP7_75t_L g12350 ( 
.A1(n_11377),
.A2(n_7930),
.B1(n_8157),
.B2(n_8359),
.Y(n_12350)
);

AND2x2_ASAP7_75t_L g12351 ( 
.A(n_11309),
.B(n_9808),
.Y(n_12351)
);

AOI22xp33_ASAP7_75t_L g12352 ( 
.A1(n_11377),
.A2(n_7930),
.B1(n_8359),
.B2(n_8367),
.Y(n_12352)
);

NAND2xp5_ASAP7_75t_L g12353 ( 
.A(n_11237),
.B(n_9727),
.Y(n_12353)
);

AOI22xp33_ASAP7_75t_L g12354 ( 
.A1(n_11380),
.A2(n_7930),
.B1(n_8359),
.B2(n_8367),
.Y(n_12354)
);

OAI22xp5_ASAP7_75t_L g12355 ( 
.A1(n_11320),
.A2(n_8565),
.B1(n_8573),
.B2(n_8541),
.Y(n_12355)
);

CKINVDCx5p33_ASAP7_75t_R g12356 ( 
.A(n_10639),
.Y(n_12356)
);

OAI22xp5_ASAP7_75t_L g12357 ( 
.A1(n_11320),
.A2(n_8590),
.B1(n_8711),
.B2(n_8641),
.Y(n_12357)
);

INVx2_ASAP7_75t_SL g12358 ( 
.A(n_10681),
.Y(n_12358)
);

OAI22xp5_ASAP7_75t_L g12359 ( 
.A1(n_11337),
.A2(n_8798),
.B1(n_8711),
.B2(n_6998),
.Y(n_12359)
);

NAND2x1_ASAP7_75t_L g12360 ( 
.A(n_10681),
.B(n_8961),
.Y(n_12360)
);

INVx3_ASAP7_75t_L g12361 ( 
.A(n_10681),
.Y(n_12361)
);

AOI22xp33_ASAP7_75t_L g12362 ( 
.A1(n_11380),
.A2(n_7930),
.B1(n_8359),
.B2(n_8367),
.Y(n_12362)
);

INVx1_ASAP7_75t_L g12363 ( 
.A(n_11234),
.Y(n_12363)
);

AOI22xp33_ASAP7_75t_L g12364 ( 
.A1(n_11394),
.A2(n_7930),
.B1(n_8367),
.B2(n_7924),
.Y(n_12364)
);

AOI22xp33_ASAP7_75t_L g12365 ( 
.A1(n_11394),
.A2(n_8367),
.B1(n_7924),
.B2(n_7925),
.Y(n_12365)
);

AOI21xp33_ASAP7_75t_L g12366 ( 
.A1(n_11241),
.A2(n_8192),
.B(n_7979),
.Y(n_12366)
);

NAND3xp33_ASAP7_75t_L g12367 ( 
.A(n_11253),
.B(n_9168),
.C(n_9072),
.Y(n_12367)
);

OAI22xp33_ASAP7_75t_L g12368 ( 
.A1(n_11337),
.A2(n_8798),
.B1(n_8711),
.B2(n_6894),
.Y(n_12368)
);

INVx1_ASAP7_75t_L g12369 ( 
.A(n_11255),
.Y(n_12369)
);

OAI22xp5_ASAP7_75t_L g12370 ( 
.A1(n_11339),
.A2(n_8798),
.B1(n_8711),
.B2(n_6998),
.Y(n_12370)
);

A2O1A1Ixp33_ASAP7_75t_L g12371 ( 
.A1(n_10616),
.A2(n_10178),
.B(n_10097),
.C(n_9040),
.Y(n_12371)
);

NAND2x1_ASAP7_75t_L g12372 ( 
.A(n_10715),
.B(n_8961),
.Y(n_12372)
);

AND2x2_ASAP7_75t_L g12373 ( 
.A(n_11322),
.B(n_9808),
.Y(n_12373)
);

INVx1_ASAP7_75t_L g12374 ( 
.A(n_11262),
.Y(n_12374)
);

OAI211xp5_ASAP7_75t_SL g12375 ( 
.A1(n_10715),
.A2(n_8974),
.B(n_8997),
.C(n_8961),
.Y(n_12375)
);

AOI22xp5_ASAP7_75t_L g12376 ( 
.A1(n_11322),
.A2(n_7823),
.B1(n_7800),
.B2(n_8002),
.Y(n_12376)
);

OAI22xp5_ASAP7_75t_L g12377 ( 
.A1(n_11339),
.A2(n_8798),
.B1(n_8711),
.B2(n_7052),
.Y(n_12377)
);

AOI22xp33_ASAP7_75t_L g12378 ( 
.A1(n_11338),
.A2(n_7924),
.B1(n_7925),
.B2(n_7922),
.Y(n_12378)
);

OAI21x1_ASAP7_75t_L g12379 ( 
.A1(n_10570),
.A2(n_9278),
.B(n_9274),
.Y(n_12379)
);

INVx1_ASAP7_75t_L g12380 ( 
.A(n_11263),
.Y(n_12380)
);

OAI22xp33_ASAP7_75t_L g12381 ( 
.A1(n_10721),
.A2(n_8798),
.B1(n_8711),
.B2(n_6894),
.Y(n_12381)
);

OAI22xp5_ASAP7_75t_L g12382 ( 
.A1(n_11338),
.A2(n_8798),
.B1(n_8711),
.B2(n_7052),
.Y(n_12382)
);

HB1xp67_ASAP7_75t_L g12383 ( 
.A(n_11432),
.Y(n_12383)
);

AOI22xp33_ASAP7_75t_L g12384 ( 
.A1(n_11349),
.A2(n_7924),
.B1(n_7925),
.B2(n_7922),
.Y(n_12384)
);

AOI22xp33_ASAP7_75t_L g12385 ( 
.A1(n_11349),
.A2(n_7924),
.B1(n_7925),
.B2(n_7922),
.Y(n_12385)
);

AOI221xp5_ASAP7_75t_L g12386 ( 
.A1(n_11432),
.A2(n_8123),
.B1(n_8509),
.B2(n_8562),
.C(n_8484),
.Y(n_12386)
);

INVx2_ASAP7_75t_L g12387 ( 
.A(n_10715),
.Y(n_12387)
);

NAND2xp5_ASAP7_75t_L g12388 ( 
.A(n_11272),
.B(n_8464),
.Y(n_12388)
);

AOI221xp5_ASAP7_75t_L g12389 ( 
.A1(n_11440),
.A2(n_8567),
.B1(n_8562),
.B2(n_8484),
.C(n_9779),
.Y(n_12389)
);

INVx2_ASAP7_75t_L g12390 ( 
.A(n_11359),
.Y(n_12390)
);

OAI22xp5_ASAP7_75t_L g12391 ( 
.A1(n_11359),
.A2(n_8798),
.B1(n_8711),
.B2(n_7052),
.Y(n_12391)
);

AOI22xp33_ASAP7_75t_SL g12392 ( 
.A1(n_10766),
.A2(n_8837),
.B1(n_9310),
.B2(n_8738),
.Y(n_12392)
);

INVxp67_ASAP7_75t_L g12393 ( 
.A(n_11265),
.Y(n_12393)
);

OAI22xp5_ASAP7_75t_L g12394 ( 
.A1(n_11421),
.A2(n_8798),
.B1(n_7061),
.B2(n_6986),
.Y(n_12394)
);

OAI211xp5_ASAP7_75t_L g12395 ( 
.A1(n_11440),
.A2(n_7968),
.B(n_7980),
.C(n_7951),
.Y(n_12395)
);

OR2x2_ASAP7_75t_L g12396 ( 
.A(n_11272),
.B(n_8470),
.Y(n_12396)
);

INVx1_ASAP7_75t_L g12397 ( 
.A(n_11267),
.Y(n_12397)
);

BUFx6f_ASAP7_75t_L g12398 ( 
.A(n_10772),
.Y(n_12398)
);

AOI22xp33_ASAP7_75t_L g12399 ( 
.A1(n_11421),
.A2(n_7925),
.B1(n_7939),
.B2(n_7922),
.Y(n_12399)
);

AOI21xp33_ASAP7_75t_SL g12400 ( 
.A1(n_10567),
.A2(n_7281),
.B(n_5903),
.Y(n_12400)
);

AND2x2_ASAP7_75t_L g12401 ( 
.A(n_11025),
.B(n_9824),
.Y(n_12401)
);

AND2x4_ASAP7_75t_L g12402 ( 
.A(n_11025),
.B(n_9824),
.Y(n_12402)
);

AOI222xp33_ASAP7_75t_L g12403 ( 
.A1(n_11269),
.A2(n_8567),
.B1(n_7555),
.B2(n_7548),
.C1(n_7294),
.C2(n_7275),
.Y(n_12403)
);

INVx4_ASAP7_75t_L g12404 ( 
.A(n_10772),
.Y(n_12404)
);

BUFx12f_ASAP7_75t_L g12405 ( 
.A(n_11315),
.Y(n_12405)
);

BUFx4f_ASAP7_75t_SL g12406 ( 
.A(n_10772),
.Y(n_12406)
);

AND2x4_ASAP7_75t_L g12407 ( 
.A(n_11026),
.B(n_9708),
.Y(n_12407)
);

INVx2_ASAP7_75t_L g12408 ( 
.A(n_11104),
.Y(n_12408)
);

AOI21xp33_ASAP7_75t_L g12409 ( 
.A1(n_11273),
.A2(n_7979),
.B(n_7963),
.Y(n_12409)
);

INVx2_ASAP7_75t_L g12410 ( 
.A(n_11104),
.Y(n_12410)
);

AOI22xp33_ASAP7_75t_L g12411 ( 
.A1(n_10823),
.A2(n_7939),
.B1(n_7944),
.B2(n_7922),
.Y(n_12411)
);

BUFx4f_ASAP7_75t_SL g12412 ( 
.A(n_10823),
.Y(n_12412)
);

OR2x2_ASAP7_75t_L g12413 ( 
.A(n_12002),
.B(n_11315),
.Y(n_12413)
);

INVx2_ASAP7_75t_L g12414 ( 
.A(n_11621),
.Y(n_12414)
);

INVx1_ASAP7_75t_L g12415 ( 
.A(n_11474),
.Y(n_12415)
);

INVx1_ASAP7_75t_L g12416 ( 
.A(n_12232),
.Y(n_12416)
);

AND2x4_ASAP7_75t_SL g12417 ( 
.A(n_11457),
.B(n_8052),
.Y(n_12417)
);

AND2x2_ASAP7_75t_L g12418 ( 
.A(n_11654),
.B(n_11026),
.Y(n_12418)
);

AND2x2_ASAP7_75t_L g12419 ( 
.A(n_11445),
.B(n_11049),
.Y(n_12419)
);

INVx1_ASAP7_75t_L g12420 ( 
.A(n_12235),
.Y(n_12420)
);

HB1xp67_ASAP7_75t_L g12421 ( 
.A(n_12244),
.Y(n_12421)
);

NAND2xp5_ASAP7_75t_L g12422 ( 
.A(n_11505),
.B(n_11341),
.Y(n_12422)
);

INVx2_ASAP7_75t_L g12423 ( 
.A(n_11705),
.Y(n_12423)
);

NOR2xp33_ASAP7_75t_L g12424 ( 
.A(n_11503),
.B(n_11523),
.Y(n_12424)
);

INVx1_ASAP7_75t_L g12425 ( 
.A(n_12274),
.Y(n_12425)
);

INVx2_ASAP7_75t_L g12426 ( 
.A(n_11687),
.Y(n_12426)
);

INVx2_ASAP7_75t_L g12427 ( 
.A(n_11687),
.Y(n_12427)
);

AND2x2_ASAP7_75t_L g12428 ( 
.A(n_11446),
.B(n_11049),
.Y(n_12428)
);

AND2x2_ASAP7_75t_L g12429 ( 
.A(n_11478),
.B(n_11071),
.Y(n_12429)
);

OR2x2_ASAP7_75t_L g12430 ( 
.A(n_11821),
.B(n_11341),
.Y(n_12430)
);

AND2x2_ASAP7_75t_L g12431 ( 
.A(n_11510),
.B(n_11071),
.Y(n_12431)
);

OR2x2_ASAP7_75t_L g12432 ( 
.A(n_11480),
.B(n_11276),
.Y(n_12432)
);

AND2x4_ASAP7_75t_L g12433 ( 
.A(n_11810),
.B(n_11072),
.Y(n_12433)
);

HB1xp67_ASAP7_75t_L g12434 ( 
.A(n_11529),
.Y(n_12434)
);

AND2x2_ASAP7_75t_L g12435 ( 
.A(n_11452),
.B(n_11072),
.Y(n_12435)
);

INVx1_ASAP7_75t_L g12436 ( 
.A(n_12337),
.Y(n_12436)
);

INVx1_ASAP7_75t_L g12437 ( 
.A(n_12383),
.Y(n_12437)
);

INVx2_ASAP7_75t_SL g12438 ( 
.A(n_11457),
.Y(n_12438)
);

HB1xp67_ASAP7_75t_L g12439 ( 
.A(n_11546),
.Y(n_12439)
);

INVxp67_ASAP7_75t_SL g12440 ( 
.A(n_11484),
.Y(n_12440)
);

INVx1_ASAP7_75t_L g12441 ( 
.A(n_11550),
.Y(n_12441)
);

AND2x4_ASAP7_75t_L g12442 ( 
.A(n_11534),
.B(n_11079),
.Y(n_12442)
);

AND2x2_ASAP7_75t_L g12443 ( 
.A(n_11455),
.B(n_11079),
.Y(n_12443)
);

INVx2_ASAP7_75t_L g12444 ( 
.A(n_11687),
.Y(n_12444)
);

AND2x2_ASAP7_75t_L g12445 ( 
.A(n_11543),
.B(n_11081),
.Y(n_12445)
);

INVx1_ASAP7_75t_L g12446 ( 
.A(n_11628),
.Y(n_12446)
);

INVx2_ASAP7_75t_L g12447 ( 
.A(n_11720),
.Y(n_12447)
);

AND2x2_ASAP7_75t_L g12448 ( 
.A(n_11619),
.B(n_11081),
.Y(n_12448)
);

HB1xp67_ASAP7_75t_L g12449 ( 
.A(n_11638),
.Y(n_12449)
);

OR2x2_ASAP7_75t_L g12450 ( 
.A(n_11646),
.B(n_11284),
.Y(n_12450)
);

INVx1_ASAP7_75t_L g12451 ( 
.A(n_11691),
.Y(n_12451)
);

AND2x2_ASAP7_75t_L g12452 ( 
.A(n_11633),
.B(n_11095),
.Y(n_12452)
);

OR2x2_ASAP7_75t_L g12453 ( 
.A(n_11698),
.B(n_11296),
.Y(n_12453)
);

AND2x2_ASAP7_75t_L g12454 ( 
.A(n_11663),
.B(n_11095),
.Y(n_12454)
);

NAND2xp5_ASAP7_75t_L g12455 ( 
.A(n_11471),
.B(n_11306),
.Y(n_12455)
);

INVx1_ASAP7_75t_L g12456 ( 
.A(n_11764),
.Y(n_12456)
);

AND2x4_ASAP7_75t_SL g12457 ( 
.A(n_12035),
.B(n_11640),
.Y(n_12457)
);

INVx1_ASAP7_75t_L g12458 ( 
.A(n_11448),
.Y(n_12458)
);

INVx2_ASAP7_75t_L g12459 ( 
.A(n_11720),
.Y(n_12459)
);

OAI22xp5_ASAP7_75t_L g12460 ( 
.A1(n_11538),
.A2(n_9310),
.B1(n_7798),
.B2(n_7811),
.Y(n_12460)
);

INVxp67_ASAP7_75t_SL g12461 ( 
.A(n_12298),
.Y(n_12461)
);

AND2x2_ASAP7_75t_L g12462 ( 
.A(n_11533),
.B(n_11098),
.Y(n_12462)
);

OR2x2_ASAP7_75t_L g12463 ( 
.A(n_12169),
.B(n_11307),
.Y(n_12463)
);

AND2x2_ASAP7_75t_L g12464 ( 
.A(n_11541),
.B(n_11098),
.Y(n_12464)
);

INVx2_ASAP7_75t_L g12465 ( 
.A(n_11720),
.Y(n_12465)
);

OR2x6_ASAP7_75t_L g12466 ( 
.A(n_11523),
.B(n_6259),
.Y(n_12466)
);

NAND2xp5_ASAP7_75t_L g12467 ( 
.A(n_11548),
.B(n_11312),
.Y(n_12467)
);

INVx1_ASAP7_75t_L g12468 ( 
.A(n_11450),
.Y(n_12468)
);

INVx1_ASAP7_75t_L g12469 ( 
.A(n_11904),
.Y(n_12469)
);

OR2x2_ASAP7_75t_L g12470 ( 
.A(n_12197),
.B(n_11313),
.Y(n_12470)
);

INVx2_ASAP7_75t_L g12471 ( 
.A(n_11737),
.Y(n_12471)
);

INVx1_ASAP7_75t_L g12472 ( 
.A(n_11960),
.Y(n_12472)
);

INVx1_ASAP7_75t_L g12473 ( 
.A(n_11977),
.Y(n_12473)
);

INVx1_ASAP7_75t_L g12474 ( 
.A(n_12015),
.Y(n_12474)
);

INVx2_ASAP7_75t_L g12475 ( 
.A(n_11755),
.Y(n_12475)
);

HB1xp67_ASAP7_75t_L g12476 ( 
.A(n_12217),
.Y(n_12476)
);

AND2x2_ASAP7_75t_L g12477 ( 
.A(n_11666),
.B(n_11105),
.Y(n_12477)
);

INVx2_ASAP7_75t_L g12478 ( 
.A(n_11767),
.Y(n_12478)
);

HB1xp67_ASAP7_75t_L g12479 ( 
.A(n_11970),
.Y(n_12479)
);

INVx1_ASAP7_75t_L g12480 ( 
.A(n_12114),
.Y(n_12480)
);

AND2x2_ASAP7_75t_L g12481 ( 
.A(n_11980),
.B(n_11105),
.Y(n_12481)
);

NAND2xp5_ASAP7_75t_L g12482 ( 
.A(n_11548),
.B(n_11316),
.Y(n_12482)
);

AND2x2_ASAP7_75t_L g12483 ( 
.A(n_12101),
.B(n_11689),
.Y(n_12483)
);

NOR2x1p5_ASAP7_75t_L g12484 ( 
.A(n_11741),
.B(n_6592),
.Y(n_12484)
);

AND2x2_ASAP7_75t_L g12485 ( 
.A(n_11926),
.B(n_11109),
.Y(n_12485)
);

INVx2_ASAP7_75t_L g12486 ( 
.A(n_12268),
.Y(n_12486)
);

AND2x2_ASAP7_75t_L g12487 ( 
.A(n_11744),
.B(n_11109),
.Y(n_12487)
);

AND2x2_ASAP7_75t_L g12488 ( 
.A(n_11519),
.B(n_11137),
.Y(n_12488)
);

INVx2_ASAP7_75t_SL g12489 ( 
.A(n_11722),
.Y(n_12489)
);

AND2x2_ASAP7_75t_L g12490 ( 
.A(n_11521),
.B(n_11137),
.Y(n_12490)
);

AND2x4_ASAP7_75t_L g12491 ( 
.A(n_11534),
.B(n_12152),
.Y(n_12491)
);

NAND2xp5_ASAP7_75t_L g12492 ( 
.A(n_11463),
.B(n_11321),
.Y(n_12492)
);

INVx2_ASAP7_75t_L g12493 ( 
.A(n_12268),
.Y(n_12493)
);

BUFx3_ASAP7_75t_L g12494 ( 
.A(n_11641),
.Y(n_12494)
);

BUFx3_ASAP7_75t_L g12495 ( 
.A(n_11798),
.Y(n_12495)
);

INVx4_ASAP7_75t_SL g12496 ( 
.A(n_11523),
.Y(n_12496)
);

INVx1_ASAP7_75t_L g12497 ( 
.A(n_11443),
.Y(n_12497)
);

INVx1_ASAP7_75t_L g12498 ( 
.A(n_11465),
.Y(n_12498)
);

INVx1_ASAP7_75t_L g12499 ( 
.A(n_11466),
.Y(n_12499)
);

INVx1_ASAP7_75t_L g12500 ( 
.A(n_11479),
.Y(n_12500)
);

INVx4_ASAP7_75t_L g12501 ( 
.A(n_11451),
.Y(n_12501)
);

INVx1_ASAP7_75t_L g12502 ( 
.A(n_11491),
.Y(n_12502)
);

AND2x2_ASAP7_75t_SL g12503 ( 
.A(n_11569),
.B(n_8291),
.Y(n_12503)
);

INVx2_ASAP7_75t_L g12504 ( 
.A(n_12268),
.Y(n_12504)
);

AND2x4_ASAP7_75t_L g12505 ( 
.A(n_11714),
.B(n_11145),
.Y(n_12505)
);

AND2x2_ASAP7_75t_L g12506 ( 
.A(n_12195),
.B(n_11145),
.Y(n_12506)
);

INVx2_ASAP7_75t_L g12507 ( 
.A(n_11805),
.Y(n_12507)
);

INVx1_ASAP7_75t_L g12508 ( 
.A(n_11513),
.Y(n_12508)
);

OR2x2_ASAP7_75t_L g12509 ( 
.A(n_11680),
.B(n_11327),
.Y(n_12509)
);

NOR2x1p5_ASAP7_75t_L g12510 ( 
.A(n_11458),
.B(n_6592),
.Y(n_12510)
);

OR2x2_ASAP7_75t_L g12511 ( 
.A(n_11520),
.B(n_11328),
.Y(n_12511)
);

AND2x2_ASAP7_75t_L g12512 ( 
.A(n_11724),
.B(n_11164),
.Y(n_12512)
);

INVx1_ASAP7_75t_L g12513 ( 
.A(n_11522),
.Y(n_12513)
);

INVxp67_ASAP7_75t_SL g12514 ( 
.A(n_12008),
.Y(n_12514)
);

INVx1_ASAP7_75t_L g12515 ( 
.A(n_11528),
.Y(n_12515)
);

BUFx2_ASAP7_75t_L g12516 ( 
.A(n_12253),
.Y(n_12516)
);

NOR2x1_ASAP7_75t_L g12517 ( 
.A(n_12127),
.B(n_10823),
.Y(n_12517)
);

INVx1_ASAP7_75t_L g12518 ( 
.A(n_11535),
.Y(n_12518)
);

INVxp33_ASAP7_75t_SL g12519 ( 
.A(n_11673),
.Y(n_12519)
);

INVx1_ASAP7_75t_L g12520 ( 
.A(n_11547),
.Y(n_12520)
);

HB1xp67_ASAP7_75t_L g12521 ( 
.A(n_12212),
.Y(n_12521)
);

INVx2_ASAP7_75t_L g12522 ( 
.A(n_12303),
.Y(n_12522)
);

AND2x2_ASAP7_75t_L g12523 ( 
.A(n_11752),
.B(n_11164),
.Y(n_12523)
);

INVx1_ASAP7_75t_L g12524 ( 
.A(n_11556),
.Y(n_12524)
);

INVxp67_ASAP7_75t_L g12525 ( 
.A(n_12064),
.Y(n_12525)
);

OR2x2_ASAP7_75t_L g12526 ( 
.A(n_12171),
.B(n_11330),
.Y(n_12526)
);

BUFx3_ASAP7_75t_L g12527 ( 
.A(n_11498),
.Y(n_12527)
);

OR2x2_ASAP7_75t_L g12528 ( 
.A(n_11497),
.B(n_11333),
.Y(n_12528)
);

AND2x2_ASAP7_75t_L g12529 ( 
.A(n_11759),
.B(n_11165),
.Y(n_12529)
);

AND2x2_ASAP7_75t_L g12530 ( 
.A(n_12032),
.B(n_11165),
.Y(n_12530)
);

AND2x2_ASAP7_75t_L g12531 ( 
.A(n_12062),
.B(n_11174),
.Y(n_12531)
);

INVx1_ASAP7_75t_L g12532 ( 
.A(n_11557),
.Y(n_12532)
);

INVx1_ASAP7_75t_L g12533 ( 
.A(n_11567),
.Y(n_12533)
);

INVx2_ASAP7_75t_L g12534 ( 
.A(n_12303),
.Y(n_12534)
);

NAND2xp5_ASAP7_75t_L g12535 ( 
.A(n_11517),
.B(n_11334),
.Y(n_12535)
);

INVx1_ASAP7_75t_L g12536 ( 
.A(n_11580),
.Y(n_12536)
);

AND2x4_ASAP7_75t_L g12537 ( 
.A(n_11734),
.B(n_11174),
.Y(n_12537)
);

INVx1_ASAP7_75t_L g12538 ( 
.A(n_11585),
.Y(n_12538)
);

INVx2_ASAP7_75t_L g12539 ( 
.A(n_12283),
.Y(n_12539)
);

AND2x2_ASAP7_75t_L g12540 ( 
.A(n_12070),
.B(n_11187),
.Y(n_12540)
);

INVx1_ASAP7_75t_L g12541 ( 
.A(n_11599),
.Y(n_12541)
);

INVx3_ASAP7_75t_L g12542 ( 
.A(n_12135),
.Y(n_12542)
);

HB1xp67_ASAP7_75t_L g12543 ( 
.A(n_12341),
.Y(n_12543)
);

AND2x2_ASAP7_75t_L g12544 ( 
.A(n_12075),
.B(n_11187),
.Y(n_12544)
);

AND2x2_ASAP7_75t_L g12545 ( 
.A(n_12082),
.B(n_11208),
.Y(n_12545)
);

BUFx2_ASAP7_75t_L g12546 ( 
.A(n_12263),
.Y(n_12546)
);

OR2x2_ASAP7_75t_L g12547 ( 
.A(n_11637),
.B(n_11342),
.Y(n_12547)
);

INVx1_ASAP7_75t_L g12548 ( 
.A(n_11601),
.Y(n_12548)
);

INVx2_ASAP7_75t_L g12549 ( 
.A(n_12283),
.Y(n_12549)
);

BUFx3_ASAP7_75t_L g12550 ( 
.A(n_11869),
.Y(n_12550)
);

INVx2_ASAP7_75t_L g12551 ( 
.A(n_12294),
.Y(n_12551)
);

INVx2_ASAP7_75t_L g12552 ( 
.A(n_12294),
.Y(n_12552)
);

AOI21xp33_ASAP7_75t_SL g12553 ( 
.A1(n_11593),
.A2(n_5175),
.B(n_5165),
.Y(n_12553)
);

INVx1_ASAP7_75t_L g12554 ( 
.A(n_11605),
.Y(n_12554)
);

AND2x2_ASAP7_75t_L g12555 ( 
.A(n_12123),
.B(n_11208),
.Y(n_12555)
);

INVxp67_ASAP7_75t_SL g12556 ( 
.A(n_12102),
.Y(n_12556)
);

BUFx4f_ASAP7_75t_L g12557 ( 
.A(n_11458),
.Y(n_12557)
);

AND2x2_ASAP7_75t_L g12558 ( 
.A(n_11492),
.B(n_11257),
.Y(n_12558)
);

INVx2_ASAP7_75t_L g12559 ( 
.A(n_12321),
.Y(n_12559)
);

HB1xp67_ASAP7_75t_L g12560 ( 
.A(n_12405),
.Y(n_12560)
);

AND2x2_ASAP7_75t_L g12561 ( 
.A(n_11895),
.B(n_11257),
.Y(n_12561)
);

INVx2_ASAP7_75t_L g12562 ( 
.A(n_12321),
.Y(n_12562)
);

INVx2_ASAP7_75t_L g12563 ( 
.A(n_11514),
.Y(n_12563)
);

INVx2_ASAP7_75t_L g12564 ( 
.A(n_11544),
.Y(n_12564)
);

CKINVDCx5p33_ASAP7_75t_R g12565 ( 
.A(n_11615),
.Y(n_12565)
);

AND2x2_ASAP7_75t_L g12566 ( 
.A(n_11929),
.B(n_11259),
.Y(n_12566)
);

INVx2_ASAP7_75t_L g12567 ( 
.A(n_11703),
.Y(n_12567)
);

AND2x2_ASAP7_75t_L g12568 ( 
.A(n_11944),
.B(n_11259),
.Y(n_12568)
);

AND2x2_ASAP7_75t_L g12569 ( 
.A(n_11770),
.B(n_9708),
.Y(n_12569)
);

AND2x2_ASAP7_75t_L g12570 ( 
.A(n_11784),
.B(n_9739),
.Y(n_12570)
);

AND2x2_ASAP7_75t_L g12571 ( 
.A(n_11788),
.B(n_9739),
.Y(n_12571)
);

AND2x2_ASAP7_75t_L g12572 ( 
.A(n_11797),
.B(n_9774),
.Y(n_12572)
);

INVx1_ASAP7_75t_L g12573 ( 
.A(n_11616),
.Y(n_12573)
);

INVx2_ASAP7_75t_L g12574 ( 
.A(n_12228),
.Y(n_12574)
);

INVx2_ASAP7_75t_L g12575 ( 
.A(n_12228),
.Y(n_12575)
);

INVxp67_ASAP7_75t_SL g12576 ( 
.A(n_12167),
.Y(n_12576)
);

INVx1_ASAP7_75t_L g12577 ( 
.A(n_11618),
.Y(n_12577)
);

INVx2_ASAP7_75t_SL g12578 ( 
.A(n_11451),
.Y(n_12578)
);

INVx1_ASAP7_75t_L g12579 ( 
.A(n_11625),
.Y(n_12579)
);

NAND2xp5_ASAP7_75t_L g12580 ( 
.A(n_11726),
.B(n_11345),
.Y(n_12580)
);

AND2x2_ASAP7_75t_L g12581 ( 
.A(n_11799),
.B(n_9774),
.Y(n_12581)
);

INVx1_ASAP7_75t_L g12582 ( 
.A(n_11642),
.Y(n_12582)
);

NAND2xp5_ASAP7_75t_L g12583 ( 
.A(n_11509),
.B(n_11346),
.Y(n_12583)
);

BUFx3_ASAP7_75t_L g12584 ( 
.A(n_11851),
.Y(n_12584)
);

INVx2_ASAP7_75t_L g12585 ( 
.A(n_12305),
.Y(n_12585)
);

AND2x2_ASAP7_75t_L g12586 ( 
.A(n_11826),
.B(n_9790),
.Y(n_12586)
);

INVx1_ASAP7_75t_L g12587 ( 
.A(n_11657),
.Y(n_12587)
);

INVx2_ASAP7_75t_SL g12588 ( 
.A(n_11451),
.Y(n_12588)
);

AND2x2_ASAP7_75t_L g12589 ( 
.A(n_11837),
.B(n_9790),
.Y(n_12589)
);

INVx1_ASAP7_75t_L g12590 ( 
.A(n_11662),
.Y(n_12590)
);

AND2x2_ASAP7_75t_L g12591 ( 
.A(n_11872),
.B(n_10842),
.Y(n_12591)
);

AND2x2_ASAP7_75t_L g12592 ( 
.A(n_11876),
.B(n_10842),
.Y(n_12592)
);

NAND2xp5_ASAP7_75t_L g12593 ( 
.A(n_11512),
.B(n_11348),
.Y(n_12593)
);

BUFx2_ASAP7_75t_L g12594 ( 
.A(n_11917),
.Y(n_12594)
);

INVx2_ASAP7_75t_L g12595 ( 
.A(n_12305),
.Y(n_12595)
);

BUFx4f_ASAP7_75t_SL g12596 ( 
.A(n_12030),
.Y(n_12596)
);

INVx2_ASAP7_75t_L g12597 ( 
.A(n_12342),
.Y(n_12597)
);

AND2x2_ASAP7_75t_L g12598 ( 
.A(n_11878),
.B(n_10842),
.Y(n_12598)
);

CKINVDCx10_ASAP7_75t_R g12599 ( 
.A(n_11456),
.Y(n_12599)
);

INVx2_ASAP7_75t_L g12600 ( 
.A(n_12342),
.Y(n_12600)
);

NAND2xp5_ASAP7_75t_L g12601 ( 
.A(n_11468),
.B(n_11350),
.Y(n_12601)
);

NAND2xp5_ASAP7_75t_L g12602 ( 
.A(n_11475),
.B(n_11352),
.Y(n_12602)
);

AND2x2_ASAP7_75t_L g12603 ( 
.A(n_11894),
.B(n_10844),
.Y(n_12603)
);

AND2x2_ASAP7_75t_L g12604 ( 
.A(n_11974),
.B(n_10844),
.Y(n_12604)
);

AND2x4_ASAP7_75t_L g12605 ( 
.A(n_11779),
.B(n_10844),
.Y(n_12605)
);

BUFx6f_ASAP7_75t_L g12606 ( 
.A(n_11460),
.Y(n_12606)
);

BUFx8_ASAP7_75t_L g12607 ( 
.A(n_11456),
.Y(n_12607)
);

AND2x2_ASAP7_75t_L g12608 ( 
.A(n_11985),
.B(n_10873),
.Y(n_12608)
);

AND2x4_ASAP7_75t_SL g12609 ( 
.A(n_11629),
.B(n_8052),
.Y(n_12609)
);

OR2x2_ASAP7_75t_L g12610 ( 
.A(n_11651),
.B(n_11353),
.Y(n_12610)
);

AND2x2_ASAP7_75t_L g12611 ( 
.A(n_12275),
.B(n_12288),
.Y(n_12611)
);

INVx1_ASAP7_75t_L g12612 ( 
.A(n_11685),
.Y(n_12612)
);

OR2x2_ASAP7_75t_L g12613 ( 
.A(n_11586),
.B(n_11354),
.Y(n_12613)
);

OR2x2_ASAP7_75t_L g12614 ( 
.A(n_11882),
.B(n_11364),
.Y(n_12614)
);

INVxp67_ASAP7_75t_SL g12615 ( 
.A(n_11790),
.Y(n_12615)
);

NAND2xp5_ASAP7_75t_L g12616 ( 
.A(n_11459),
.B(n_11366),
.Y(n_12616)
);

AND2x2_ASAP7_75t_L g12617 ( 
.A(n_12289),
.B(n_12172),
.Y(n_12617)
);

INVx3_ASAP7_75t_L g12618 ( 
.A(n_12127),
.Y(n_12618)
);

BUFx2_ASAP7_75t_L g12619 ( 
.A(n_11917),
.Y(n_12619)
);

NAND2xp5_ASAP7_75t_L g12620 ( 
.A(n_11489),
.B(n_11371),
.Y(n_12620)
);

AND2x2_ASAP7_75t_L g12621 ( 
.A(n_12172),
.B(n_10873),
.Y(n_12621)
);

INVx3_ASAP7_75t_L g12622 ( 
.A(n_12360),
.Y(n_12622)
);

INVx2_ASAP7_75t_L g12623 ( 
.A(n_12361),
.Y(n_12623)
);

INVx1_ASAP7_75t_L g12624 ( 
.A(n_11696),
.Y(n_12624)
);

HB1xp67_ASAP7_75t_L g12625 ( 
.A(n_12222),
.Y(n_12625)
);

INVx1_ASAP7_75t_L g12626 ( 
.A(n_11700),
.Y(n_12626)
);

AND2x2_ASAP7_75t_L g12627 ( 
.A(n_11678),
.B(n_11731),
.Y(n_12627)
);

INVx1_ASAP7_75t_L g12628 ( 
.A(n_11706),
.Y(n_12628)
);

INVxp67_ASAP7_75t_SL g12629 ( 
.A(n_11742),
.Y(n_12629)
);

AND2x2_ASAP7_75t_L g12630 ( 
.A(n_12112),
.B(n_10873),
.Y(n_12630)
);

INVx1_ASAP7_75t_L g12631 ( 
.A(n_11727),
.Y(n_12631)
);

INVx2_ASAP7_75t_L g12632 ( 
.A(n_12361),
.Y(n_12632)
);

INVx1_ASAP7_75t_L g12633 ( 
.A(n_11728),
.Y(n_12633)
);

OR2x2_ASAP7_75t_L g12634 ( 
.A(n_12223),
.B(n_11372),
.Y(n_12634)
);

AOI22xp33_ASAP7_75t_L g12635 ( 
.A1(n_11454),
.A2(n_10969),
.B1(n_10978),
.B2(n_10977),
.Y(n_12635)
);

AND2x2_ASAP7_75t_L g12636 ( 
.A(n_12112),
.B(n_10969),
.Y(n_12636)
);

HB1xp67_ASAP7_75t_L g12637 ( 
.A(n_12222),
.Y(n_12637)
);

INVx2_ASAP7_75t_L g12638 ( 
.A(n_11967),
.Y(n_12638)
);

INVx2_ASAP7_75t_L g12639 ( 
.A(n_11967),
.Y(n_12639)
);

BUFx2_ASAP7_75t_L g12640 ( 
.A(n_12203),
.Y(n_12640)
);

INVx2_ASAP7_75t_L g12641 ( 
.A(n_11967),
.Y(n_12641)
);

AND2x2_ASAP7_75t_L g12642 ( 
.A(n_12021),
.B(n_10969),
.Y(n_12642)
);

INVx1_ASAP7_75t_L g12643 ( 
.A(n_11758),
.Y(n_12643)
);

INVx2_ASAP7_75t_L g12644 ( 
.A(n_12402),
.Y(n_12644)
);

INVx1_ASAP7_75t_SL g12645 ( 
.A(n_11573),
.Y(n_12645)
);

NAND2xp5_ASAP7_75t_L g12646 ( 
.A(n_11462),
.B(n_11379),
.Y(n_12646)
);

OR2x2_ASAP7_75t_L g12647 ( 
.A(n_11816),
.B(n_11384),
.Y(n_12647)
);

INVx1_ASAP7_75t_L g12648 ( 
.A(n_11777),
.Y(n_12648)
);

INVx1_ASAP7_75t_L g12649 ( 
.A(n_11780),
.Y(n_12649)
);

BUFx2_ASAP7_75t_L g12650 ( 
.A(n_12202),
.Y(n_12650)
);

INVx1_ASAP7_75t_L g12651 ( 
.A(n_11800),
.Y(n_12651)
);

INVxp67_ASAP7_75t_L g12652 ( 
.A(n_12083),
.Y(n_12652)
);

AND2x2_ASAP7_75t_L g12653 ( 
.A(n_12027),
.B(n_10977),
.Y(n_12653)
);

BUFx3_ASAP7_75t_L g12654 ( 
.A(n_11460),
.Y(n_12654)
);

BUFx3_ASAP7_75t_L g12655 ( 
.A(n_11835),
.Y(n_12655)
);

AND2x2_ASAP7_75t_L g12656 ( 
.A(n_12154),
.B(n_10977),
.Y(n_12656)
);

AND2x2_ASAP7_75t_L g12657 ( 
.A(n_12154),
.B(n_10978),
.Y(n_12657)
);

INVx2_ASAP7_75t_L g12658 ( 
.A(n_12402),
.Y(n_12658)
);

NAND2xp5_ASAP7_75t_L g12659 ( 
.A(n_11660),
.B(n_11385),
.Y(n_12659)
);

AND2x2_ASAP7_75t_L g12660 ( 
.A(n_12292),
.B(n_10978),
.Y(n_12660)
);

INVx2_ASAP7_75t_L g12661 ( 
.A(n_11861),
.Y(n_12661)
);

INVx2_ASAP7_75t_L g12662 ( 
.A(n_11861),
.Y(n_12662)
);

HB1xp67_ASAP7_75t_L g12663 ( 
.A(n_12096),
.Y(n_12663)
);

INVx2_ASAP7_75t_L g12664 ( 
.A(n_11861),
.Y(n_12664)
);

INVx2_ASAP7_75t_L g12665 ( 
.A(n_11883),
.Y(n_12665)
);

INVx2_ASAP7_75t_L g12666 ( 
.A(n_11883),
.Y(n_12666)
);

INVx1_ASAP7_75t_L g12667 ( 
.A(n_11802),
.Y(n_12667)
);

BUFx3_ASAP7_75t_L g12668 ( 
.A(n_11890),
.Y(n_12668)
);

AND2x4_ASAP7_75t_L g12669 ( 
.A(n_11952),
.B(n_11955),
.Y(n_12669)
);

AND2x2_ASAP7_75t_L g12670 ( 
.A(n_11447),
.B(n_11068),
.Y(n_12670)
);

NAND2xp5_ASAP7_75t_L g12671 ( 
.A(n_11563),
.B(n_11386),
.Y(n_12671)
);

INVx1_ASAP7_75t_L g12672 ( 
.A(n_11809),
.Y(n_12672)
);

HB1xp67_ASAP7_75t_L g12673 ( 
.A(n_12179),
.Y(n_12673)
);

NAND2xp33_ASAP7_75t_R g12674 ( 
.A(n_11709),
.B(n_5175),
.Y(n_12674)
);

AND2x2_ASAP7_75t_L g12675 ( 
.A(n_11499),
.B(n_11068),
.Y(n_12675)
);

HB1xp67_ASAP7_75t_L g12676 ( 
.A(n_12308),
.Y(n_12676)
);

AND2x2_ASAP7_75t_L g12677 ( 
.A(n_11540),
.B(n_11068),
.Y(n_12677)
);

NAND2x1_ASAP7_75t_L g12678 ( 
.A(n_11865),
.B(n_11099),
.Y(n_12678)
);

INVx2_ASAP7_75t_L g12679 ( 
.A(n_11883),
.Y(n_12679)
);

AND2x2_ASAP7_75t_L g12680 ( 
.A(n_11549),
.B(n_11099),
.Y(n_12680)
);

INVx1_ASAP7_75t_L g12681 ( 
.A(n_11868),
.Y(n_12681)
);

INVx1_ASAP7_75t_L g12682 ( 
.A(n_11875),
.Y(n_12682)
);

INVx1_ASAP7_75t_L g12683 ( 
.A(n_11881),
.Y(n_12683)
);

INVx1_ASAP7_75t_L g12684 ( 
.A(n_11889),
.Y(n_12684)
);

AND2x2_ASAP7_75t_L g12685 ( 
.A(n_11597),
.B(n_11099),
.Y(n_12685)
);

INVx2_ASAP7_75t_L g12686 ( 
.A(n_12407),
.Y(n_12686)
);

NOR2xp33_ASAP7_75t_L g12687 ( 
.A(n_11732),
.B(n_6605),
.Y(n_12687)
);

AOI22xp33_ASAP7_75t_L g12688 ( 
.A1(n_11493),
.A2(n_11116),
.B1(n_11226),
.B2(n_11205),
.Y(n_12688)
);

INVx1_ASAP7_75t_L g12689 ( 
.A(n_11893),
.Y(n_12689)
);

INVx2_ASAP7_75t_L g12690 ( 
.A(n_12407),
.Y(n_12690)
);

INVx2_ASAP7_75t_L g12691 ( 
.A(n_12315),
.Y(n_12691)
);

NAND2xp5_ASAP7_75t_L g12692 ( 
.A(n_11500),
.B(n_11388),
.Y(n_12692)
);

INVx2_ASAP7_75t_L g12693 ( 
.A(n_11887),
.Y(n_12693)
);

AND2x2_ASAP7_75t_L g12694 ( 
.A(n_11612),
.B(n_11116),
.Y(n_12694)
);

AND2x2_ASAP7_75t_L g12695 ( 
.A(n_11622),
.B(n_11116),
.Y(n_12695)
);

INVx2_ASAP7_75t_L g12696 ( 
.A(n_11668),
.Y(n_12696)
);

INVxp67_ASAP7_75t_L g12697 ( 
.A(n_11901),
.Y(n_12697)
);

NAND2xp5_ASAP7_75t_L g12698 ( 
.A(n_11670),
.B(n_11609),
.Y(n_12698)
);

INVx2_ASAP7_75t_L g12699 ( 
.A(n_11668),
.Y(n_12699)
);

BUFx2_ASAP7_75t_L g12700 ( 
.A(n_12072),
.Y(n_12700)
);

AND2x2_ASAP7_75t_L g12701 ( 
.A(n_12122),
.B(n_11205),
.Y(n_12701)
);

INVx2_ASAP7_75t_L g12702 ( 
.A(n_11668),
.Y(n_12702)
);

INVx1_ASAP7_75t_L g12703 ( 
.A(n_11897),
.Y(n_12703)
);

INVx2_ASAP7_75t_L g12704 ( 
.A(n_11849),
.Y(n_12704)
);

AND2x2_ASAP7_75t_L g12705 ( 
.A(n_11553),
.B(n_11205),
.Y(n_12705)
);

INVx1_ASAP7_75t_L g12706 ( 
.A(n_11911),
.Y(n_12706)
);

NOR2x1_ASAP7_75t_L g12707 ( 
.A(n_11808),
.B(n_11226),
.Y(n_12707)
);

INVx2_ASAP7_75t_L g12708 ( 
.A(n_11849),
.Y(n_12708)
);

AND2x2_ASAP7_75t_L g12709 ( 
.A(n_11566),
.B(n_11226),
.Y(n_12709)
);

HB1xp67_ASAP7_75t_L g12710 ( 
.A(n_11973),
.Y(n_12710)
);

INVxp67_ASAP7_75t_SL g12711 ( 
.A(n_11568),
.Y(n_12711)
);

INVx1_ASAP7_75t_SL g12712 ( 
.A(n_12069),
.Y(n_12712)
);

AND2x4_ASAP7_75t_L g12713 ( 
.A(n_11952),
.B(n_11230),
.Y(n_12713)
);

AND2x2_ASAP7_75t_L g12714 ( 
.A(n_11570),
.B(n_11230),
.Y(n_12714)
);

INVx1_ASAP7_75t_L g12715 ( 
.A(n_11921),
.Y(n_12715)
);

INVx1_ASAP7_75t_L g12716 ( 
.A(n_11947),
.Y(n_12716)
);

INVx1_ASAP7_75t_L g12717 ( 
.A(n_11962),
.Y(n_12717)
);

HB1xp67_ASAP7_75t_L g12718 ( 
.A(n_11964),
.Y(n_12718)
);

INVxp67_ASAP7_75t_L g12719 ( 
.A(n_12236),
.Y(n_12719)
);

INVx2_ASAP7_75t_L g12720 ( 
.A(n_11849),
.Y(n_12720)
);

NAND2xp5_ASAP7_75t_L g12721 ( 
.A(n_11771),
.B(n_11389),
.Y(n_12721)
);

INVx5_ASAP7_75t_L g12722 ( 
.A(n_11629),
.Y(n_12722)
);

NAND2xp5_ASAP7_75t_L g12723 ( 
.A(n_11511),
.B(n_11390),
.Y(n_12723)
);

INVx2_ASAP7_75t_L g12724 ( 
.A(n_11850),
.Y(n_12724)
);

AND2x2_ASAP7_75t_L g12725 ( 
.A(n_11874),
.B(n_11230),
.Y(n_12725)
);

AOI22xp33_ASAP7_75t_L g12726 ( 
.A1(n_11481),
.A2(n_11290),
.B1(n_11331),
.B2(n_11293),
.Y(n_12726)
);

AND2x2_ASAP7_75t_L g12727 ( 
.A(n_11874),
.B(n_11290),
.Y(n_12727)
);

INVx2_ASAP7_75t_L g12728 ( 
.A(n_11850),
.Y(n_12728)
);

INVx1_ASAP7_75t_L g12729 ( 
.A(n_11963),
.Y(n_12729)
);

AND2x2_ASAP7_75t_L g12730 ( 
.A(n_11648),
.B(n_11290),
.Y(n_12730)
);

AND2x2_ASAP7_75t_L g12731 ( 
.A(n_11648),
.B(n_11293),
.Y(n_12731)
);

BUFx2_ASAP7_75t_L g12732 ( 
.A(n_12080),
.Y(n_12732)
);

AND2x2_ASAP7_75t_L g12733 ( 
.A(n_11955),
.B(n_12196),
.Y(n_12733)
);

NAND2xp5_ASAP7_75t_L g12734 ( 
.A(n_11442),
.B(n_11403),
.Y(n_12734)
);

AOI221xp5_ASAP7_75t_L g12735 ( 
.A1(n_11496),
.A2(n_11410),
.B1(n_11412),
.B2(n_11409),
.C(n_11404),
.Y(n_12735)
);

INVx2_ASAP7_75t_L g12736 ( 
.A(n_12327),
.Y(n_12736)
);

OAI22xp5_ASAP7_75t_L g12737 ( 
.A1(n_11490),
.A2(n_9310),
.B1(n_7798),
.B2(n_7811),
.Y(n_12737)
);

INVx2_ASAP7_75t_L g12738 ( 
.A(n_12327),
.Y(n_12738)
);

HB1xp67_ASAP7_75t_L g12739 ( 
.A(n_11948),
.Y(n_12739)
);

NAND2x1p5_ASAP7_75t_L g12740 ( 
.A(n_12095),
.B(n_11293),
.Y(n_12740)
);

INVxp67_ASAP7_75t_SL g12741 ( 
.A(n_11701),
.Y(n_12741)
);

AND2x2_ASAP7_75t_L g12742 ( 
.A(n_12196),
.B(n_11331),
.Y(n_12742)
);

INVx2_ASAP7_75t_L g12743 ( 
.A(n_12250),
.Y(n_12743)
);

NAND2xp5_ASAP7_75t_L g12744 ( 
.A(n_11607),
.B(n_11413),
.Y(n_12744)
);

INVx1_ASAP7_75t_L g12745 ( 
.A(n_11975),
.Y(n_12745)
);

AOI22xp33_ASAP7_75t_SL g12746 ( 
.A1(n_11453),
.A2(n_9310),
.B1(n_11336),
.B2(n_11331),
.Y(n_12746)
);

INVx2_ASAP7_75t_L g12747 ( 
.A(n_12250),
.Y(n_12747)
);

AND2x2_ASAP7_75t_L g12748 ( 
.A(n_11617),
.B(n_11336),
.Y(n_12748)
);

AND2x2_ASAP7_75t_L g12749 ( 
.A(n_12219),
.B(n_12225),
.Y(n_12749)
);

HB1xp67_ASAP7_75t_L g12750 ( 
.A(n_11987),
.Y(n_12750)
);

AND2x2_ASAP7_75t_L g12751 ( 
.A(n_11608),
.B(n_11336),
.Y(n_12751)
);

INVx2_ASAP7_75t_SL g12752 ( 
.A(n_11704),
.Y(n_12752)
);

INVx1_ASAP7_75t_L g12753 ( 
.A(n_11983),
.Y(n_12753)
);

INVx1_ASAP7_75t_L g12754 ( 
.A(n_12005),
.Y(n_12754)
);

INVx2_ASAP7_75t_L g12755 ( 
.A(n_11979),
.Y(n_12755)
);

BUFx3_ASAP7_75t_L g12756 ( 
.A(n_11965),
.Y(n_12756)
);

BUFx2_ASAP7_75t_L g12757 ( 
.A(n_12088),
.Y(n_12757)
);

INVx2_ASAP7_75t_L g12758 ( 
.A(n_11979),
.Y(n_12758)
);

INVx3_ASAP7_75t_L g12759 ( 
.A(n_12372),
.Y(n_12759)
);

INVx1_ASAP7_75t_L g12760 ( 
.A(n_12009),
.Y(n_12760)
);

HB1xp67_ASAP7_75t_L g12761 ( 
.A(n_11991),
.Y(n_12761)
);

AND2x2_ASAP7_75t_L g12762 ( 
.A(n_11608),
.B(n_11363),
.Y(n_12762)
);

INVx1_ASAP7_75t_L g12763 ( 
.A(n_12012),
.Y(n_12763)
);

INVxp67_ASAP7_75t_SL g12764 ( 
.A(n_11859),
.Y(n_12764)
);

BUFx3_ASAP7_75t_L g12765 ( 
.A(n_11801),
.Y(n_12765)
);

CKINVDCx14_ASAP7_75t_R g12766 ( 
.A(n_11828),
.Y(n_12766)
);

AND2x2_ASAP7_75t_L g12767 ( 
.A(n_11620),
.B(n_11363),
.Y(n_12767)
);

NAND2xp5_ASAP7_75t_L g12768 ( 
.A(n_11461),
.B(n_11417),
.Y(n_12768)
);

INVx1_ASAP7_75t_L g12769 ( 
.A(n_12036),
.Y(n_12769)
);

NAND2xp5_ASAP7_75t_L g12770 ( 
.A(n_11988),
.B(n_11418),
.Y(n_12770)
);

INVx1_ASAP7_75t_L g12771 ( 
.A(n_12040),
.Y(n_12771)
);

AND2x2_ASAP7_75t_L g12772 ( 
.A(n_11620),
.B(n_11363),
.Y(n_12772)
);

AND2x2_ASAP7_75t_L g12773 ( 
.A(n_11634),
.B(n_11378),
.Y(n_12773)
);

INVx1_ASAP7_75t_L g12774 ( 
.A(n_12043),
.Y(n_12774)
);

INVx2_ASAP7_75t_L g12775 ( 
.A(n_11808),
.Y(n_12775)
);

AND2x2_ASAP7_75t_L g12776 ( 
.A(n_11634),
.B(n_11378),
.Y(n_12776)
);

AND2x4_ASAP7_75t_L g12777 ( 
.A(n_11713),
.B(n_11378),
.Y(n_12777)
);

INVx2_ASAP7_75t_L g12778 ( 
.A(n_11832),
.Y(n_12778)
);

INVx3_ASAP7_75t_L g12779 ( 
.A(n_11832),
.Y(n_12779)
);

AND2x2_ASAP7_75t_L g12780 ( 
.A(n_11713),
.B(n_11430),
.Y(n_12780)
);

INVx1_ASAP7_75t_L g12781 ( 
.A(n_12049),
.Y(n_12781)
);

INVx1_ASAP7_75t_L g12782 ( 
.A(n_12052),
.Y(n_12782)
);

NAND2xp5_ASAP7_75t_L g12783 ( 
.A(n_11602),
.B(n_11436),
.Y(n_12783)
);

NAND2xp5_ASAP7_75t_L g12784 ( 
.A(n_11603),
.B(n_10567),
.Y(n_12784)
);

INVx1_ASAP7_75t_L g12785 ( 
.A(n_12056),
.Y(n_12785)
);

BUFx2_ASAP7_75t_L g12786 ( 
.A(n_11990),
.Y(n_12786)
);

HB1xp67_ASAP7_75t_L g12787 ( 
.A(n_11993),
.Y(n_12787)
);

INVx1_ASAP7_75t_L g12788 ( 
.A(n_12061),
.Y(n_12788)
);

INVx1_ASAP7_75t_L g12789 ( 
.A(n_12066),
.Y(n_12789)
);

AND2x2_ASAP7_75t_L g12790 ( 
.A(n_11785),
.B(n_7916),
.Y(n_12790)
);

BUFx6f_ASAP7_75t_L g12791 ( 
.A(n_11806),
.Y(n_12791)
);

AND2x2_ASAP7_75t_L g12792 ( 
.A(n_11785),
.B(n_7916),
.Y(n_12792)
);

HB1xp67_ASAP7_75t_L g12793 ( 
.A(n_11630),
.Y(n_12793)
);

INVx1_ASAP7_75t_L g12794 ( 
.A(n_12068),
.Y(n_12794)
);

AOI222xp33_ASAP7_75t_L g12795 ( 
.A1(n_11525),
.A2(n_9785),
.B1(n_9788),
.B2(n_9798),
.C1(n_9795),
.C2(n_9784),
.Y(n_12795)
);

INVx1_ASAP7_75t_L g12796 ( 
.A(n_12106),
.Y(n_12796)
);

INVx1_ASAP7_75t_L g12797 ( 
.A(n_12116),
.Y(n_12797)
);

HB1xp67_ASAP7_75t_L g12798 ( 
.A(n_12238),
.Y(n_12798)
);

NOR2x1_ASAP7_75t_SL g12799 ( 
.A(n_12031),
.B(n_6605),
.Y(n_12799)
);

INVx1_ASAP7_75t_L g12800 ( 
.A(n_12129),
.Y(n_12800)
);

INVx2_ASAP7_75t_L g12801 ( 
.A(n_11879),
.Y(n_12801)
);

INVx2_ASAP7_75t_L g12802 ( 
.A(n_11704),
.Y(n_12802)
);

NAND2xp5_ASAP7_75t_L g12803 ( 
.A(n_11494),
.B(n_10295),
.Y(n_12803)
);

AND2x4_ASAP7_75t_L g12804 ( 
.A(n_11812),
.B(n_7844),
.Y(n_12804)
);

AND2x2_ASAP7_75t_L g12805 ( 
.A(n_11812),
.B(n_7916),
.Y(n_12805)
);

AND2x2_ASAP7_75t_L g12806 ( 
.A(n_11825),
.B(n_7916),
.Y(n_12806)
);

BUFx3_ASAP7_75t_L g12807 ( 
.A(n_11945),
.Y(n_12807)
);

INVx2_ASAP7_75t_L g12808 ( 
.A(n_12398),
.Y(n_12808)
);

INVx1_ASAP7_75t_L g12809 ( 
.A(n_12134),
.Y(n_12809)
);

BUFx2_ASAP7_75t_L g12810 ( 
.A(n_11825),
.Y(n_12810)
);

INVx2_ASAP7_75t_L g12811 ( 
.A(n_12398),
.Y(n_12811)
);

INVx2_ASAP7_75t_L g12812 ( 
.A(n_12398),
.Y(n_12812)
);

INVx2_ASAP7_75t_L g12813 ( 
.A(n_12034),
.Y(n_12813)
);

NAND2xp5_ASAP7_75t_L g12814 ( 
.A(n_11624),
.B(n_10297),
.Y(n_12814)
);

INVx2_ASAP7_75t_L g12815 ( 
.A(n_12034),
.Y(n_12815)
);

BUFx3_ASAP7_75t_L g12816 ( 
.A(n_11610),
.Y(n_12816)
);

NAND2xp5_ASAP7_75t_L g12817 ( 
.A(n_11639),
.B(n_10301),
.Y(n_12817)
);

INVx1_ASAP7_75t_L g12818 ( 
.A(n_12139),
.Y(n_12818)
);

AND2x2_ASAP7_75t_L g12819 ( 
.A(n_12031),
.B(n_7939),
.Y(n_12819)
);

INVx1_ASAP7_75t_L g12820 ( 
.A(n_12143),
.Y(n_12820)
);

INVx2_ASAP7_75t_L g12821 ( 
.A(n_12045),
.Y(n_12821)
);

INVx2_ASAP7_75t_L g12822 ( 
.A(n_12045),
.Y(n_12822)
);

INVx1_ASAP7_75t_L g12823 ( 
.A(n_12144),
.Y(n_12823)
);

OR2x2_ASAP7_75t_L g12824 ( 
.A(n_12164),
.B(n_8512),
.Y(n_12824)
);

INVx2_ASAP7_75t_L g12825 ( 
.A(n_12071),
.Y(n_12825)
);

INVx1_ASAP7_75t_L g12826 ( 
.A(n_12145),
.Y(n_12826)
);

AND2x2_ASAP7_75t_L g12827 ( 
.A(n_12233),
.B(n_7939),
.Y(n_12827)
);

AND2x2_ASAP7_75t_L g12828 ( 
.A(n_11978),
.B(n_11524),
.Y(n_12828)
);

INVx1_ASAP7_75t_L g12829 ( 
.A(n_12161),
.Y(n_12829)
);

OR2x2_ASAP7_75t_L g12830 ( 
.A(n_12166),
.B(n_8512),
.Y(n_12830)
);

AND2x2_ASAP7_75t_L g12831 ( 
.A(n_11682),
.B(n_12047),
.Y(n_12831)
);

AND2x2_ASAP7_75t_L g12832 ( 
.A(n_11949),
.B(n_7939),
.Y(n_12832)
);

INVx2_ASAP7_75t_L g12833 ( 
.A(n_12071),
.Y(n_12833)
);

INVx1_ASAP7_75t_L g12834 ( 
.A(n_12180),
.Y(n_12834)
);

INVx4_ASAP7_75t_L g12835 ( 
.A(n_11674),
.Y(n_12835)
);

AND2x2_ASAP7_75t_L g12836 ( 
.A(n_11959),
.B(n_7944),
.Y(n_12836)
);

INVx2_ASAP7_75t_L g12837 ( 
.A(n_11950),
.Y(n_12837)
);

AO31x2_ASAP7_75t_L g12838 ( 
.A1(n_12076),
.A2(n_10312),
.A3(n_10313),
.B(n_10310),
.Y(n_12838)
);

OR2x2_ASAP7_75t_L g12839 ( 
.A(n_12168),
.B(n_8512),
.Y(n_12839)
);

INVx2_ASAP7_75t_L g12840 ( 
.A(n_11950),
.Y(n_12840)
);

OAI22xp5_ASAP7_75t_L g12841 ( 
.A1(n_11504),
.A2(n_7798),
.B1(n_7811),
.B2(n_7769),
.Y(n_12841)
);

INVx2_ASAP7_75t_L g12842 ( 
.A(n_11982),
.Y(n_12842)
);

AND2x2_ASAP7_75t_L g12843 ( 
.A(n_11674),
.B(n_7944),
.Y(n_12843)
);

AND2x2_ASAP7_75t_L g12844 ( 
.A(n_11694),
.B(n_7944),
.Y(n_12844)
);

INVx1_ASAP7_75t_L g12845 ( 
.A(n_12183),
.Y(n_12845)
);

AND2x2_ASAP7_75t_L g12846 ( 
.A(n_11694),
.B(n_7944),
.Y(n_12846)
);

INVx1_ASAP7_75t_SL g12847 ( 
.A(n_12406),
.Y(n_12847)
);

AND2x2_ASAP7_75t_L g12848 ( 
.A(n_12390),
.B(n_11671),
.Y(n_12848)
);

INVx2_ASAP7_75t_L g12849 ( 
.A(n_11982),
.Y(n_12849)
);

INVx2_ASAP7_75t_L g12850 ( 
.A(n_12404),
.Y(n_12850)
);

OR2x2_ASAP7_75t_L g12851 ( 
.A(n_12001),
.B(n_8512),
.Y(n_12851)
);

AND2x2_ASAP7_75t_L g12852 ( 
.A(n_11681),
.B(n_7958),
.Y(n_12852)
);

AND2x2_ASAP7_75t_L g12853 ( 
.A(n_12408),
.B(n_12410),
.Y(n_12853)
);

AND2x4_ASAP7_75t_L g12854 ( 
.A(n_11729),
.B(n_7844),
.Y(n_12854)
);

AND2x2_ASAP7_75t_L g12855 ( 
.A(n_11690),
.B(n_7958),
.Y(n_12855)
);

AND2x2_ASAP7_75t_L g12856 ( 
.A(n_11594),
.B(n_7958),
.Y(n_12856)
);

AND2x2_ASAP7_75t_L g12857 ( 
.A(n_11995),
.B(n_7958),
.Y(n_12857)
);

AND2x2_ASAP7_75t_L g12858 ( 
.A(n_12094),
.B(n_7958),
.Y(n_12858)
);

INVx1_ASAP7_75t_L g12859 ( 
.A(n_12188),
.Y(n_12859)
);

NAND2xp5_ASAP7_75t_L g12860 ( 
.A(n_11702),
.B(n_10314),
.Y(n_12860)
);

INVx1_ASAP7_75t_L g12861 ( 
.A(n_12192),
.Y(n_12861)
);

AND2x2_ASAP7_75t_L g12862 ( 
.A(n_12097),
.B(n_8115),
.Y(n_12862)
);

INVx1_ASAP7_75t_L g12863 ( 
.A(n_12205),
.Y(n_12863)
);

INVx2_ASAP7_75t_L g12864 ( 
.A(n_12404),
.Y(n_12864)
);

NAND2xp5_ASAP7_75t_L g12865 ( 
.A(n_11707),
.B(n_11721),
.Y(n_12865)
);

INVx2_ASAP7_75t_L g12866 ( 
.A(n_12358),
.Y(n_12866)
);

INVx2_ASAP7_75t_L g12867 ( 
.A(n_12401),
.Y(n_12867)
);

NAND2x1_ASAP7_75t_L g12868 ( 
.A(n_11824),
.B(n_8961),
.Y(n_12868)
);

AND2x4_ASAP7_75t_SL g12869 ( 
.A(n_11906),
.B(n_8052),
.Y(n_12869)
);

INVx3_ASAP7_75t_L g12870 ( 
.A(n_11908),
.Y(n_12870)
);

INVxp67_ASAP7_75t_L g12871 ( 
.A(n_11831),
.Y(n_12871)
);

INVx2_ASAP7_75t_L g12872 ( 
.A(n_12351),
.Y(n_12872)
);

OR2x2_ASAP7_75t_L g12873 ( 
.A(n_12091),
.B(n_8512),
.Y(n_12873)
);

AND2x2_ASAP7_75t_L g12874 ( 
.A(n_12100),
.B(n_8115),
.Y(n_12874)
);

AND2x2_ASAP7_75t_L g12875 ( 
.A(n_12111),
.B(n_8115),
.Y(n_12875)
);

INVxp67_ASAP7_75t_L g12876 ( 
.A(n_11650),
.Y(n_12876)
);

INVx1_ASAP7_75t_L g12877 ( 
.A(n_12207),
.Y(n_12877)
);

AND2x2_ASAP7_75t_L g12878 ( 
.A(n_12118),
.B(n_8115),
.Y(n_12878)
);

INVx2_ASAP7_75t_L g12879 ( 
.A(n_12373),
.Y(n_12879)
);

AND2x4_ASAP7_75t_L g12880 ( 
.A(n_11765),
.B(n_7908),
.Y(n_12880)
);

BUFx2_ASAP7_75t_L g12881 ( 
.A(n_12224),
.Y(n_12881)
);

INVx1_ASAP7_75t_L g12882 ( 
.A(n_12231),
.Y(n_12882)
);

AOI211xp5_ASAP7_75t_SL g12883 ( 
.A1(n_11565),
.A2(n_8997),
.B(n_9096),
.C(n_8974),
.Y(n_12883)
);

AND2x2_ASAP7_75t_L g12884 ( 
.A(n_11842),
.B(n_8115),
.Y(n_12884)
);

BUFx6f_ASAP7_75t_L g12885 ( 
.A(n_12038),
.Y(n_12885)
);

AOI22xp33_ASAP7_75t_SL g12886 ( 
.A1(n_11476),
.A2(n_7968),
.B1(n_7980),
.B2(n_7951),
.Y(n_12886)
);

BUFx3_ASAP7_75t_L g12887 ( 
.A(n_11725),
.Y(n_12887)
);

OR2x2_ASAP7_75t_L g12888 ( 
.A(n_12262),
.B(n_8512),
.Y(n_12888)
);

INVx1_ASAP7_75t_SL g12889 ( 
.A(n_12412),
.Y(n_12889)
);

BUFx2_ASAP7_75t_L g12890 ( 
.A(n_12325),
.Y(n_12890)
);

HB1xp67_ASAP7_75t_L g12891 ( 
.A(n_12329),
.Y(n_12891)
);

INVx1_ASAP7_75t_L g12892 ( 
.A(n_12237),
.Y(n_12892)
);

AOI22xp33_ASAP7_75t_L g12893 ( 
.A1(n_11477),
.A2(n_11793),
.B1(n_11527),
.B2(n_11530),
.Y(n_12893)
);

INVx1_ASAP7_75t_L g12894 ( 
.A(n_12242),
.Y(n_12894)
);

INVx2_ASAP7_75t_L g12895 ( 
.A(n_12105),
.Y(n_12895)
);

AND2x2_ASAP7_75t_L g12896 ( 
.A(n_11649),
.B(n_8160),
.Y(n_12896)
);

INVx2_ASAP7_75t_L g12897 ( 
.A(n_12133),
.Y(n_12897)
);

AND2x2_ASAP7_75t_L g12898 ( 
.A(n_12176),
.B(n_8160),
.Y(n_12898)
);

AND2x2_ASAP7_75t_L g12899 ( 
.A(n_11924),
.B(n_8160),
.Y(n_12899)
);

NAND2xp5_ASAP7_75t_L g12900 ( 
.A(n_11749),
.B(n_10316),
.Y(n_12900)
);

BUFx2_ASAP7_75t_L g12901 ( 
.A(n_12356),
.Y(n_12901)
);

INVx1_ASAP7_75t_L g12902 ( 
.A(n_12246),
.Y(n_12902)
);

AND2x2_ASAP7_75t_L g12903 ( 
.A(n_11933),
.B(n_11942),
.Y(n_12903)
);

NAND2x1p5_ASAP7_75t_L g12904 ( 
.A(n_11746),
.B(n_8351),
.Y(n_12904)
);

AND2x4_ASAP7_75t_L g12905 ( 
.A(n_11756),
.B(n_7908),
.Y(n_12905)
);

INVx1_ASAP7_75t_L g12906 ( 
.A(n_12251),
.Y(n_12906)
);

AND2x2_ASAP7_75t_L g12907 ( 
.A(n_11953),
.B(n_8160),
.Y(n_12907)
);

INVx1_ASAP7_75t_L g12908 ( 
.A(n_12271),
.Y(n_12908)
);

INVx3_ASAP7_75t_SL g12909 ( 
.A(n_11470),
.Y(n_12909)
);

AND2x2_ASAP7_75t_L g12910 ( 
.A(n_12103),
.B(n_8160),
.Y(n_12910)
);

AND2x2_ASAP7_75t_L g12911 ( 
.A(n_12107),
.B(n_8190),
.Y(n_12911)
);

NAND2xp5_ASAP7_75t_L g12912 ( 
.A(n_11768),
.B(n_10322),
.Y(n_12912)
);

INVx1_ASAP7_75t_L g12913 ( 
.A(n_12281),
.Y(n_12913)
);

AND2x2_ASAP7_75t_L g12914 ( 
.A(n_12108),
.B(n_8190),
.Y(n_12914)
);

INVx2_ASAP7_75t_L g12915 ( 
.A(n_12151),
.Y(n_12915)
);

INVx2_ASAP7_75t_L g12916 ( 
.A(n_12153),
.Y(n_12916)
);

INVx2_ASAP7_75t_L g12917 ( 
.A(n_12162),
.Y(n_12917)
);

AND2x2_ASAP7_75t_L g12918 ( 
.A(n_11692),
.B(n_8190),
.Y(n_12918)
);

AND2x2_ASAP7_75t_L g12919 ( 
.A(n_12313),
.B(n_8190),
.Y(n_12919)
);

AND2x4_ASAP7_75t_L g12920 ( 
.A(n_11787),
.B(n_8017),
.Y(n_12920)
);

AND2x2_ASAP7_75t_L g12921 ( 
.A(n_11564),
.B(n_8190),
.Y(n_12921)
);

INVx2_ASAP7_75t_L g12922 ( 
.A(n_12177),
.Y(n_12922)
);

BUFx2_ASAP7_75t_L g12923 ( 
.A(n_11840),
.Y(n_12923)
);

HB1xp67_ASAP7_75t_L g12924 ( 
.A(n_12248),
.Y(n_12924)
);

AND2x2_ASAP7_75t_L g12925 ( 
.A(n_11922),
.B(n_8215),
.Y(n_12925)
);

AND2x2_ASAP7_75t_L g12926 ( 
.A(n_12343),
.B(n_8215),
.Y(n_12926)
);

AND2x2_ASAP7_75t_L g12927 ( 
.A(n_12344),
.B(n_8215),
.Y(n_12927)
);

INVx1_ASAP7_75t_L g12928 ( 
.A(n_12293),
.Y(n_12928)
);

AND2x4_ASAP7_75t_L g12929 ( 
.A(n_11844),
.B(n_8017),
.Y(n_12929)
);

BUFx3_ASAP7_75t_L g12930 ( 
.A(n_11912),
.Y(n_12930)
);

BUFx2_ASAP7_75t_L g12931 ( 
.A(n_11846),
.Y(n_12931)
);

AND2x2_ASAP7_75t_L g12932 ( 
.A(n_11807),
.B(n_8215),
.Y(n_12932)
);

INVx2_ASAP7_75t_L g12933 ( 
.A(n_12267),
.Y(n_12933)
);

INVx1_ASAP7_75t_L g12934 ( 
.A(n_12302),
.Y(n_12934)
);

INVx2_ASAP7_75t_L g12935 ( 
.A(n_12269),
.Y(n_12935)
);

INVx2_ASAP7_75t_L g12936 ( 
.A(n_12279),
.Y(n_12936)
);

INVx1_ASAP7_75t_L g12937 ( 
.A(n_12312),
.Y(n_12937)
);

OR2x2_ASAP7_75t_L g12938 ( 
.A(n_12270),
.B(n_8512),
.Y(n_12938)
);

INVx1_ASAP7_75t_L g12939 ( 
.A(n_12317),
.Y(n_12939)
);

INVx2_ASAP7_75t_L g12940 ( 
.A(n_12334),
.Y(n_12940)
);

NAND2xp5_ASAP7_75t_L g12941 ( 
.A(n_11857),
.B(n_10329),
.Y(n_12941)
);

INVx1_ASAP7_75t_L g12942 ( 
.A(n_12328),
.Y(n_12942)
);

INVx1_ASAP7_75t_L g12943 ( 
.A(n_12330),
.Y(n_12943)
);

OR2x2_ASAP7_75t_L g12944 ( 
.A(n_12309),
.B(n_8512),
.Y(n_12944)
);

INVx4_ASAP7_75t_R g12945 ( 
.A(n_11584),
.Y(n_12945)
);

INVx2_ASAP7_75t_L g12946 ( 
.A(n_12387),
.Y(n_12946)
);

NAND2xp5_ASAP7_75t_L g12947 ( 
.A(n_11863),
.B(n_11864),
.Y(n_12947)
);

INVx1_ASAP7_75t_L g12948 ( 
.A(n_12331),
.Y(n_12948)
);

INVx1_ASAP7_75t_L g12949 ( 
.A(n_12363),
.Y(n_12949)
);

OR2x2_ASAP7_75t_L g12950 ( 
.A(n_11710),
.B(n_10331),
.Y(n_12950)
);

HB1xp67_ASAP7_75t_L g12951 ( 
.A(n_11871),
.Y(n_12951)
);

INVx1_ASAP7_75t_L g12952 ( 
.A(n_12369),
.Y(n_12952)
);

AND2x2_ASAP7_75t_L g12953 ( 
.A(n_12259),
.B(n_8215),
.Y(n_12953)
);

INVx1_ASAP7_75t_L g12954 ( 
.A(n_12374),
.Y(n_12954)
);

OR2x2_ASAP7_75t_L g12955 ( 
.A(n_12353),
.B(n_10332),
.Y(n_12955)
);

INVx1_ASAP7_75t_L g12956 ( 
.A(n_12380),
.Y(n_12956)
);

INVx1_ASAP7_75t_L g12957 ( 
.A(n_12397),
.Y(n_12957)
);

BUFx3_ASAP7_75t_L g12958 ( 
.A(n_11923),
.Y(n_12958)
);

OR2x2_ASAP7_75t_L g12959 ( 
.A(n_11537),
.B(n_10336),
.Y(n_12959)
);

NAND2xp5_ASAP7_75t_L g12960 ( 
.A(n_11880),
.B(n_11927),
.Y(n_12960)
);

OR2x2_ASAP7_75t_L g12961 ( 
.A(n_12388),
.B(n_10337),
.Y(n_12961)
);

INVx1_ASAP7_75t_L g12962 ( 
.A(n_12323),
.Y(n_12962)
);

INVx1_ASAP7_75t_L g12963 ( 
.A(n_12393),
.Y(n_12963)
);

INVx2_ASAP7_75t_L g12964 ( 
.A(n_11596),
.Y(n_12964)
);

NOR2x1_ASAP7_75t_SL g12965 ( 
.A(n_11501),
.B(n_6605),
.Y(n_12965)
);

BUFx3_ASAP7_75t_L g12966 ( 
.A(n_11986),
.Y(n_12966)
);

INVx2_ASAP7_75t_L g12967 ( 
.A(n_11596),
.Y(n_12967)
);

AND2x2_ASAP7_75t_L g12968 ( 
.A(n_12259),
.B(n_8235),
.Y(n_12968)
);

AND2x4_ASAP7_75t_L g12969 ( 
.A(n_11928),
.B(n_8185),
.Y(n_12969)
);

NAND2xp5_ASAP7_75t_L g12970 ( 
.A(n_11934),
.B(n_10339),
.Y(n_12970)
);

NAND2x1_ASAP7_75t_L g12971 ( 
.A(n_11824),
.B(n_11600),
.Y(n_12971)
);

INVx1_ASAP7_75t_L g12972 ( 
.A(n_11992),
.Y(n_12972)
);

INVx1_ASAP7_75t_L g12973 ( 
.A(n_11994),
.Y(n_12973)
);

INVx1_ASAP7_75t_L g12974 ( 
.A(n_12016),
.Y(n_12974)
);

INVx2_ASAP7_75t_L g12975 ( 
.A(n_11600),
.Y(n_12975)
);

AND2x2_ASAP7_75t_L g12976 ( 
.A(n_11532),
.B(n_8235),
.Y(n_12976)
);

INVx1_ASAP7_75t_L g12977 ( 
.A(n_12018),
.Y(n_12977)
);

INVx1_ASAP7_75t_L g12978 ( 
.A(n_12023),
.Y(n_12978)
);

BUFx3_ASAP7_75t_L g12979 ( 
.A(n_11803),
.Y(n_12979)
);

AND2x2_ASAP7_75t_L g12980 ( 
.A(n_11757),
.B(n_8235),
.Y(n_12980)
);

AND2x2_ASAP7_75t_L g12981 ( 
.A(n_11766),
.B(n_8235),
.Y(n_12981)
);

NAND2xp5_ASAP7_75t_L g12982 ( 
.A(n_12051),
.B(n_10341),
.Y(n_12982)
);

INVx1_ASAP7_75t_L g12983 ( 
.A(n_12053),
.Y(n_12983)
);

AND2x4_ASAP7_75t_L g12984 ( 
.A(n_12079),
.B(n_8185),
.Y(n_12984)
);

BUFx2_ASAP7_75t_L g12985 ( 
.A(n_11782),
.Y(n_12985)
);

INVx1_ASAP7_75t_L g12986 ( 
.A(n_12347),
.Y(n_12986)
);

AND2x2_ASAP7_75t_L g12987 ( 
.A(n_11773),
.B(n_8235),
.Y(n_12987)
);

AND2x2_ASAP7_75t_L g12988 ( 
.A(n_11774),
.B(n_8290),
.Y(n_12988)
);

NAND2xp5_ASAP7_75t_L g12989 ( 
.A(n_11518),
.B(n_10344),
.Y(n_12989)
);

HB1xp67_ASAP7_75t_L g12990 ( 
.A(n_12173),
.Y(n_12990)
);

INVx1_ASAP7_75t_L g12991 ( 
.A(n_12396),
.Y(n_12991)
);

BUFx6f_ASAP7_75t_L g12992 ( 
.A(n_11848),
.Y(n_12992)
);

INVxp67_ASAP7_75t_L g12993 ( 
.A(n_11920),
.Y(n_12993)
);

OR2x2_ASAP7_75t_L g12994 ( 
.A(n_11684),
.B(n_10345),
.Y(n_12994)
);

INVx1_ASAP7_75t_L g12995 ( 
.A(n_12039),
.Y(n_12995)
);

NOR2xp33_ASAP7_75t_L g12996 ( 
.A(n_12109),
.B(n_6605),
.Y(n_12996)
);

INVx2_ASAP7_75t_L g12997 ( 
.A(n_11611),
.Y(n_12997)
);

NOR2x1_ASAP7_75t_L g12998 ( 
.A(n_11937),
.B(n_8974),
.Y(n_12998)
);

BUFx6f_ASAP7_75t_L g12999 ( 
.A(n_11932),
.Y(n_12999)
);

INVx1_ASAP7_75t_L g13000 ( 
.A(n_12264),
.Y(n_13000)
);

INVx2_ASAP7_75t_L g13001 ( 
.A(n_11611),
.Y(n_13001)
);

BUFx4f_ASAP7_75t_SL g13002 ( 
.A(n_11656),
.Y(n_13002)
);

NAND2xp5_ASAP7_75t_L g13003 ( 
.A(n_11693),
.B(n_10347),
.Y(n_13003)
);

INVx1_ASAP7_75t_L g13004 ( 
.A(n_12266),
.Y(n_13004)
);

BUFx2_ASAP7_75t_L g13005 ( 
.A(n_11598),
.Y(n_13005)
);

AND2x2_ASAP7_75t_L g13006 ( 
.A(n_11775),
.B(n_8290),
.Y(n_13006)
);

NOR2x1_ASAP7_75t_L g13007 ( 
.A(n_11834),
.B(n_8974),
.Y(n_13007)
);

BUFx6f_ASAP7_75t_L g13008 ( 
.A(n_11656),
.Y(n_13008)
);

INVx3_ASAP7_75t_L g13009 ( 
.A(n_11661),
.Y(n_13009)
);

AND2x4_ASAP7_75t_L g13010 ( 
.A(n_11626),
.B(n_8356),
.Y(n_13010)
);

INVx1_ASAP7_75t_L g13011 ( 
.A(n_12089),
.Y(n_13011)
);

BUFx6f_ASAP7_75t_L g13012 ( 
.A(n_11661),
.Y(n_13012)
);

BUFx2_ASAP7_75t_L g13013 ( 
.A(n_11794),
.Y(n_13013)
);

INVx1_ASAP7_75t_L g13014 ( 
.A(n_12184),
.Y(n_13014)
);

HB1xp67_ASAP7_75t_L g13015 ( 
.A(n_12173),
.Y(n_13015)
);

INVx3_ASAP7_75t_L g13016 ( 
.A(n_11794),
.Y(n_13016)
);

OR2x2_ASAP7_75t_L g13017 ( 
.A(n_11745),
.B(n_10353),
.Y(n_13017)
);

INVx1_ASAP7_75t_L g13018 ( 
.A(n_12163),
.Y(n_13018)
);

HB1xp67_ASAP7_75t_L g13019 ( 
.A(n_11839),
.Y(n_13019)
);

AND2x2_ASAP7_75t_L g13020 ( 
.A(n_11783),
.B(n_8290),
.Y(n_13020)
);

INVx1_ASAP7_75t_L g13021 ( 
.A(n_12163),
.Y(n_13021)
);

INVx1_ASAP7_75t_L g13022 ( 
.A(n_12185),
.Y(n_13022)
);

INVx2_ASAP7_75t_L g13023 ( 
.A(n_11772),
.Y(n_13023)
);

AND2x4_ASAP7_75t_L g13024 ( 
.A(n_11733),
.B(n_8356),
.Y(n_13024)
);

INVxp67_ASAP7_75t_L g13025 ( 
.A(n_11632),
.Y(n_13025)
);

INVx2_ASAP7_75t_L g13026 ( 
.A(n_12255),
.Y(n_13026)
);

INVx2_ASAP7_75t_L g13027 ( 
.A(n_11545),
.Y(n_13027)
);

AND2x2_ASAP7_75t_L g13028 ( 
.A(n_11786),
.B(n_8290),
.Y(n_13028)
);

INVx2_ASAP7_75t_L g13029 ( 
.A(n_11613),
.Y(n_13029)
);

AND2x2_ASAP7_75t_L g13030 ( 
.A(n_11789),
.B(n_8290),
.Y(n_13030)
);

NAND2xp5_ASAP7_75t_L g13031 ( 
.A(n_11672),
.B(n_10354),
.Y(n_13031)
);

INVx1_ASAP7_75t_L g13032 ( 
.A(n_12185),
.Y(n_13032)
);

INVx2_ASAP7_75t_L g13033 ( 
.A(n_12249),
.Y(n_13033)
);

AND2x4_ASAP7_75t_L g13034 ( 
.A(n_12010),
.B(n_8451),
.Y(n_13034)
);

INVx1_ASAP7_75t_L g13035 ( 
.A(n_12297),
.Y(n_13035)
);

AND2x2_ASAP7_75t_L g13036 ( 
.A(n_11997),
.B(n_8340),
.Y(n_13036)
);

INVx1_ASAP7_75t_L g13037 ( 
.A(n_12249),
.Y(n_13037)
);

INVx3_ASAP7_75t_L g13038 ( 
.A(n_11913),
.Y(n_13038)
);

INVx2_ASAP7_75t_L g13039 ( 
.A(n_12307),
.Y(n_13039)
);

INVx2_ASAP7_75t_L g13040 ( 
.A(n_12307),
.Y(n_13040)
);

AND2x2_ASAP7_75t_L g13041 ( 
.A(n_11998),
.B(n_8340),
.Y(n_13041)
);

AND2x2_ASAP7_75t_L g13042 ( 
.A(n_12004),
.B(n_8340),
.Y(n_13042)
);

INVx2_ASAP7_75t_L g13043 ( 
.A(n_12339),
.Y(n_13043)
);

AND2x2_ASAP7_75t_L g13044 ( 
.A(n_12020),
.B(n_8340),
.Y(n_13044)
);

AND2x4_ASAP7_75t_L g13045 ( 
.A(n_11754),
.B(n_8451),
.Y(n_13045)
);

AND2x2_ASAP7_75t_L g13046 ( 
.A(n_12041),
.B(n_8340),
.Y(n_13046)
);

AND2x2_ASAP7_75t_L g13047 ( 
.A(n_12044),
.B(n_8443),
.Y(n_13047)
);

AND2x2_ASAP7_75t_L g13048 ( 
.A(n_12058),
.B(n_12333),
.Y(n_13048)
);

INVx2_ASAP7_75t_L g13049 ( 
.A(n_12339),
.Y(n_13049)
);

AND2x2_ASAP7_75t_L g13050 ( 
.A(n_11582),
.B(n_8443),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_12349),
.Y(n_13051)
);

INVx2_ASAP7_75t_L g13052 ( 
.A(n_12349),
.Y(n_13052)
);

INVx2_ASAP7_75t_L g13053 ( 
.A(n_12234),
.Y(n_13053)
);

INVx2_ASAP7_75t_L g13054 ( 
.A(n_12278),
.Y(n_13054)
);

INVx1_ASAP7_75t_L g13055 ( 
.A(n_12229),
.Y(n_13055)
);

AND2x2_ASAP7_75t_L g13056 ( 
.A(n_11989),
.B(n_8443),
.Y(n_13056)
);

NAND2xp5_ASAP7_75t_L g13057 ( 
.A(n_11507),
.B(n_10358),
.Y(n_13057)
);

AND2x2_ASAP7_75t_L g13058 ( 
.A(n_11588),
.B(n_11891),
.Y(n_13058)
);

BUFx6f_ASAP7_75t_L g13059 ( 
.A(n_11716),
.Y(n_13059)
);

INVx1_ASAP7_75t_L g13060 ( 
.A(n_12229),
.Y(n_13060)
);

NOR2x1_ASAP7_75t_L g13061 ( 
.A(n_11761),
.B(n_8997),
.Y(n_13061)
);

HB1xp67_ASAP7_75t_L g13062 ( 
.A(n_11905),
.Y(n_13062)
);

HB1xp67_ASAP7_75t_L g13063 ( 
.A(n_11516),
.Y(n_13063)
);

INVx2_ASAP7_75t_L g13064 ( 
.A(n_12278),
.Y(n_13064)
);

AND2x2_ASAP7_75t_L g13065 ( 
.A(n_11653),
.B(n_8443),
.Y(n_13065)
);

AND2x2_ASAP7_75t_L g13066 ( 
.A(n_11655),
.B(n_8443),
.Y(n_13066)
);

BUFx2_ASAP7_75t_L g13067 ( 
.A(n_11712),
.Y(n_13067)
);

AND2x2_ASAP7_75t_L g13068 ( 
.A(n_11738),
.B(n_8511),
.Y(n_13068)
);

NAND2xp5_ASAP7_75t_L g13069 ( 
.A(n_11579),
.B(n_10361),
.Y(n_13069)
);

NAND2xp5_ASAP7_75t_L g13070 ( 
.A(n_11554),
.B(n_10366),
.Y(n_13070)
);

AND2x2_ASAP7_75t_L g13071 ( 
.A(n_12227),
.B(n_8511),
.Y(n_13071)
);

BUFx3_ASAP7_75t_L g13072 ( 
.A(n_11956),
.Y(n_13072)
);

AND2x4_ASAP7_75t_L g13073 ( 
.A(n_11792),
.B(n_10372),
.Y(n_13073)
);

INVx3_ASAP7_75t_L g13074 ( 
.A(n_11913),
.Y(n_13074)
);

AND2x2_ASAP7_75t_L g13075 ( 
.A(n_12239),
.B(n_8511),
.Y(n_13075)
);

AND2x2_ASAP7_75t_L g13076 ( 
.A(n_12243),
.B(n_8511),
.Y(n_13076)
);

BUFx2_ASAP7_75t_L g13077 ( 
.A(n_11941),
.Y(n_13077)
);

INVx1_ASAP7_75t_L g13078 ( 
.A(n_12278),
.Y(n_13078)
);

INVx2_ASAP7_75t_L g13079 ( 
.A(n_11976),
.Y(n_13079)
);

INVxp67_ASAP7_75t_SL g13080 ( 
.A(n_11614),
.Y(n_13080)
);

INVxp67_ASAP7_75t_L g13081 ( 
.A(n_11506),
.Y(n_13081)
);

NAND2xp5_ASAP7_75t_L g13082 ( 
.A(n_11559),
.B(n_10373),
.Y(n_13082)
);

OR2x2_ASAP7_75t_L g13083 ( 
.A(n_11778),
.B(n_10379),
.Y(n_13083)
);

INVx2_ASAP7_75t_L g13084 ( 
.A(n_11516),
.Y(n_13084)
);

INVx2_ASAP7_75t_L g13085 ( 
.A(n_12138),
.Y(n_13085)
);

AND2x2_ASAP7_75t_L g13086 ( 
.A(n_12252),
.B(n_8511),
.Y(n_13086)
);

INVx2_ASAP7_75t_L g13087 ( 
.A(n_11841),
.Y(n_13087)
);

AND2x2_ASAP7_75t_L g13088 ( 
.A(n_12256),
.B(n_8625),
.Y(n_13088)
);

OR2x2_ASAP7_75t_L g13089 ( 
.A(n_11555),
.B(n_10383),
.Y(n_13089)
);

AND2x2_ASAP7_75t_L g13090 ( 
.A(n_12277),
.B(n_8625),
.Y(n_13090)
);

AND2x4_ASAP7_75t_L g13091 ( 
.A(n_11877),
.B(n_10384),
.Y(n_13091)
);

AND2x2_ASAP7_75t_L g13092 ( 
.A(n_12287),
.B(n_8625),
.Y(n_13092)
);

AND2x2_ASAP7_75t_L g13093 ( 
.A(n_12291),
.B(n_8625),
.Y(n_13093)
);

AND2x2_ASAP7_75t_L g13094 ( 
.A(n_11830),
.B(n_8625),
.Y(n_13094)
);

BUFx2_ASAP7_75t_L g13095 ( 
.A(n_11957),
.Y(n_13095)
);

BUFx3_ASAP7_75t_L g13096 ( 
.A(n_11667),
.Y(n_13096)
);

AND2x2_ASAP7_75t_L g13097 ( 
.A(n_11838),
.B(n_11853),
.Y(n_13097)
);

INVx2_ASAP7_75t_L g13098 ( 
.A(n_11748),
.Y(n_13098)
);

HB1xp67_ASAP7_75t_L g13099 ( 
.A(n_11958),
.Y(n_13099)
);

AND2x2_ASAP7_75t_L g13100 ( 
.A(n_11855),
.B(n_11899),
.Y(n_13100)
);

NAND2xp5_ASAP7_75t_L g13101 ( 
.A(n_11539),
.B(n_10387),
.Y(n_13101)
);

AND2x2_ASAP7_75t_L g13102 ( 
.A(n_11750),
.B(n_8677),
.Y(n_13102)
);

AND2x4_ASAP7_75t_L g13103 ( 
.A(n_12007),
.B(n_10389),
.Y(n_13103)
);

INVx1_ASAP7_75t_L g13104 ( 
.A(n_12218),
.Y(n_13104)
);

INVx2_ASAP7_75t_L g13105 ( 
.A(n_11748),
.Y(n_13105)
);

INVx2_ASAP7_75t_L g13106 ( 
.A(n_11981),
.Y(n_13106)
);

NAND2xp5_ASAP7_75t_L g13107 ( 
.A(n_11467),
.B(n_10390),
.Y(n_13107)
);

BUFx2_ASAP7_75t_L g13108 ( 
.A(n_11961),
.Y(n_13108)
);

INVx1_ASAP7_75t_L g13109 ( 
.A(n_12218),
.Y(n_13109)
);

AND2x2_ASAP7_75t_L g13110 ( 
.A(n_12019),
.B(n_8677),
.Y(n_13110)
);

INVx1_ASAP7_75t_L g13111 ( 
.A(n_12272),
.Y(n_13111)
);

INVx1_ASAP7_75t_L g13112 ( 
.A(n_11938),
.Y(n_13112)
);

AND2x4_ASAP7_75t_L g13113 ( 
.A(n_12060),
.B(n_10408),
.Y(n_13113)
);

INVx2_ASAP7_75t_L g13114 ( 
.A(n_12160),
.Y(n_13114)
);

AND2x2_ASAP7_75t_L g13115 ( 
.A(n_12067),
.B(n_12226),
.Y(n_13115)
);

HB1xp67_ASAP7_75t_L g13116 ( 
.A(n_11996),
.Y(n_13116)
);

AND2x2_ASAP7_75t_L g13117 ( 
.A(n_12204),
.B(n_8677),
.Y(n_13117)
);

INVx4_ASAP7_75t_L g13118 ( 
.A(n_11815),
.Y(n_13118)
);

AND2x2_ASAP7_75t_L g13119 ( 
.A(n_12211),
.B(n_8677),
.Y(n_13119)
);

INVx1_ASAP7_75t_L g13120 ( 
.A(n_11938),
.Y(n_13120)
);

INVx1_ASAP7_75t_L g13121 ( 
.A(n_12367),
.Y(n_13121)
);

AND2x2_ASAP7_75t_L g13122 ( 
.A(n_12221),
.B(n_8677),
.Y(n_13122)
);

INVx2_ASAP7_75t_L g13123 ( 
.A(n_12141),
.Y(n_13123)
);

AND2x2_ASAP7_75t_L g13124 ( 
.A(n_12300),
.B(n_8689),
.Y(n_13124)
);

BUFx2_ASAP7_75t_L g13125 ( 
.A(n_11730),
.Y(n_13125)
);

INVx2_ASAP7_75t_L g13126 ( 
.A(n_11631),
.Y(n_13126)
);

INVx1_ASAP7_75t_L g13127 ( 
.A(n_12326),
.Y(n_13127)
);

AND2x4_ASAP7_75t_L g13128 ( 
.A(n_11675),
.B(n_10409),
.Y(n_13128)
);

NOR3xp33_ASAP7_75t_L g13129 ( 
.A(n_11854),
.B(n_9096),
.C(n_8997),
.Y(n_13129)
);

NAND2xp5_ASAP7_75t_L g13130 ( 
.A(n_11464),
.B(n_11531),
.Y(n_13130)
);

INVx2_ASAP7_75t_L g13131 ( 
.A(n_12159),
.Y(n_13131)
);

INVx1_ASAP7_75t_L g13132 ( 
.A(n_12311),
.Y(n_13132)
);

INVx2_ASAP7_75t_L g13133 ( 
.A(n_12159),
.Y(n_13133)
);

INVx1_ASAP7_75t_L g13134 ( 
.A(n_12320),
.Y(n_13134)
);

NAND2xp5_ASAP7_75t_L g13135 ( 
.A(n_11581),
.B(n_10413),
.Y(n_13135)
);

BUFx2_ASAP7_75t_L g13136 ( 
.A(n_11473),
.Y(n_13136)
);

INVx1_ASAP7_75t_L g13137 ( 
.A(n_12316),
.Y(n_13137)
);

BUFx2_ASAP7_75t_L g13138 ( 
.A(n_11551),
.Y(n_13138)
);

INVx2_ASAP7_75t_SL g13139 ( 
.A(n_12055),
.Y(n_13139)
);

HB1xp67_ASAP7_75t_L g13140 ( 
.A(n_11900),
.Y(n_13140)
);

INVx1_ASAP7_75t_L g13141 ( 
.A(n_11954),
.Y(n_13141)
);

HB1xp67_ASAP7_75t_L g13142 ( 
.A(n_11898),
.Y(n_13142)
);

BUFx2_ASAP7_75t_L g13143 ( 
.A(n_11760),
.Y(n_13143)
);

BUFx3_ASAP7_75t_L g13144 ( 
.A(n_11763),
.Y(n_13144)
);

INVx3_ASAP7_75t_L g13145 ( 
.A(n_11813),
.Y(n_13145)
);

INVx3_ASAP7_75t_L g13146 ( 
.A(n_11488),
.Y(n_13146)
);

INVx2_ASAP7_75t_L g13147 ( 
.A(n_12379),
.Y(n_13147)
);

AO31x2_ASAP7_75t_L g13148 ( 
.A1(n_11907),
.A2(n_10418),
.A3(n_10424),
.B(n_10416),
.Y(n_13148)
);

AND2x4_ASAP7_75t_L g13149 ( 
.A(n_11677),
.B(n_11686),
.Y(n_13149)
);

AND2x2_ASAP7_75t_L g13150 ( 
.A(n_11711),
.B(n_8689),
.Y(n_13150)
);

INVx1_ASAP7_75t_L g13151 ( 
.A(n_11896),
.Y(n_13151)
);

AND2x2_ASAP7_75t_L g13152 ( 
.A(n_12314),
.B(n_8689),
.Y(n_13152)
);

INVx1_ASAP7_75t_L g13153 ( 
.A(n_11915),
.Y(n_13153)
);

INVx1_ASAP7_75t_L g13154 ( 
.A(n_11925),
.Y(n_13154)
);

AND2x2_ASAP7_75t_L g13155 ( 
.A(n_11485),
.B(n_8689),
.Y(n_13155)
);

INVx1_ASAP7_75t_L g13156 ( 
.A(n_11966),
.Y(n_13156)
);

AND2x2_ASAP7_75t_L g13157 ( 
.A(n_11776),
.B(n_8689),
.Y(n_13157)
);

INVx1_ASAP7_75t_L g13158 ( 
.A(n_11676),
.Y(n_13158)
);

NOR2xp33_ASAP7_75t_L g13159 ( 
.A(n_11483),
.B(n_6259),
.Y(n_13159)
);

AND2x4_ASAP7_75t_L g13160 ( 
.A(n_12155),
.B(n_10438),
.Y(n_13160)
);

INVx1_ASAP7_75t_L g13161 ( 
.A(n_11699),
.Y(n_13161)
);

NAND2xp5_ASAP7_75t_L g13162 ( 
.A(n_11449),
.B(n_10439),
.Y(n_13162)
);

INVx2_ASAP7_75t_L g13163 ( 
.A(n_12301),
.Y(n_13163)
);

INVx1_ASAP7_75t_L g13164 ( 
.A(n_11781),
.Y(n_13164)
);

INVx2_ASAP7_75t_L g13165 ( 
.A(n_12132),
.Y(n_13165)
);

INVx1_ASAP7_75t_L g13166 ( 
.A(n_11856),
.Y(n_13166)
);

BUFx6f_ASAP7_75t_L g13167 ( 
.A(n_11815),
.Y(n_13167)
);

INVxp67_ASAP7_75t_L g13168 ( 
.A(n_11627),
.Y(n_13168)
);

INVx1_ASAP7_75t_L g13169 ( 
.A(n_11909),
.Y(n_13169)
);

OR2x2_ASAP7_75t_L g13170 ( 
.A(n_11495),
.B(n_10442),
.Y(n_13170)
);

HB1xp67_ASAP7_75t_L g13171 ( 
.A(n_11903),
.Y(n_13171)
);

HB1xp67_ASAP7_75t_L g13172 ( 
.A(n_12104),
.Y(n_13172)
);

INVx2_ASAP7_75t_L g13173 ( 
.A(n_12132),
.Y(n_13173)
);

AND2x2_ASAP7_75t_L g13174 ( 
.A(n_11486),
.B(n_8702),
.Y(n_13174)
);

CKINVDCx8_ASAP7_75t_R g13175 ( 
.A(n_12336),
.Y(n_13175)
);

INVx3_ASAP7_75t_L g13176 ( 
.A(n_11885),
.Y(n_13176)
);

NAND2xp5_ASAP7_75t_L g13177 ( 
.A(n_11822),
.B(n_11526),
.Y(n_13177)
);

INVx2_ASAP7_75t_L g13178 ( 
.A(n_11885),
.Y(n_13178)
);

INVx2_ASAP7_75t_SL g13179 ( 
.A(n_12057),
.Y(n_13179)
);

INVx2_ASAP7_75t_L g13180 ( 
.A(n_11811),
.Y(n_13180)
);

OR2x2_ASAP7_75t_L g13181 ( 
.A(n_11571),
.B(n_10445),
.Y(n_13181)
);

INVx1_ASAP7_75t_L g13182 ( 
.A(n_11862),
.Y(n_13182)
);

INVx2_ASAP7_75t_L g13183 ( 
.A(n_11870),
.Y(n_13183)
);

BUFx6f_ASAP7_75t_L g13184 ( 
.A(n_12059),
.Y(n_13184)
);

AND2x2_ASAP7_75t_L g13185 ( 
.A(n_12324),
.B(n_8702),
.Y(n_13185)
);

AND2x2_ASAP7_75t_L g13186 ( 
.A(n_12194),
.B(n_8702),
.Y(n_13186)
);

BUFx2_ASAP7_75t_L g13187 ( 
.A(n_11575),
.Y(n_13187)
);

AND2x2_ASAP7_75t_L g13188 ( 
.A(n_11589),
.B(n_8702),
.Y(n_13188)
);

AND2x2_ASAP7_75t_L g13189 ( 
.A(n_11604),
.B(n_8702),
.Y(n_13189)
);

AND2x2_ASAP7_75t_L g13190 ( 
.A(n_11606),
.B(n_8703),
.Y(n_13190)
);

INVx2_ASAP7_75t_L g13191 ( 
.A(n_12286),
.Y(n_13191)
);

INVx1_ASAP7_75t_L g13192 ( 
.A(n_11940),
.Y(n_13192)
);

INVx1_ASAP7_75t_L g13193 ( 
.A(n_11791),
.Y(n_13193)
);

INVx1_ASAP7_75t_L g13194 ( 
.A(n_11804),
.Y(n_13194)
);

NAND2xp5_ASAP7_75t_L g13195 ( 
.A(n_11444),
.B(n_10450),
.Y(n_13195)
);

AND2x2_ASAP7_75t_L g13196 ( 
.A(n_12282),
.B(n_8703),
.Y(n_13196)
);

AND2x2_ASAP7_75t_L g13197 ( 
.A(n_12191),
.B(n_8703),
.Y(n_13197)
);

AND2x2_ASAP7_75t_L g13198 ( 
.A(n_12193),
.B(n_8703),
.Y(n_13198)
);

AND2x2_ASAP7_75t_L g13199 ( 
.A(n_12209),
.B(n_8703),
.Y(n_13199)
);

BUFx6f_ASAP7_75t_L g13200 ( 
.A(n_12077),
.Y(n_13200)
);

AND2x2_ASAP7_75t_L g13201 ( 
.A(n_11740),
.B(n_8831),
.Y(n_13201)
);

INVx1_ASAP7_75t_L g13202 ( 
.A(n_11843),
.Y(n_13202)
);

AND2x2_ASAP7_75t_L g13203 ( 
.A(n_11592),
.B(n_8831),
.Y(n_13203)
);

BUFx2_ASAP7_75t_L g13204 ( 
.A(n_11818),
.Y(n_13204)
);

INVxp67_ASAP7_75t_SL g13205 ( 
.A(n_12013),
.Y(n_13205)
);

AND2x2_ASAP7_75t_L g13206 ( 
.A(n_12149),
.B(n_8831),
.Y(n_13206)
);

INVx1_ASAP7_75t_L g13207 ( 
.A(n_11919),
.Y(n_13207)
);

NAND2xp5_ASAP7_75t_L g13208 ( 
.A(n_11910),
.B(n_10454),
.Y(n_13208)
);

INVx1_ASAP7_75t_L g13209 ( 
.A(n_12355),
.Y(n_13209)
);

BUFx3_ASAP7_75t_L g13210 ( 
.A(n_12063),
.Y(n_13210)
);

BUFx2_ASAP7_75t_L g13211 ( 
.A(n_11751),
.Y(n_13211)
);

HB1xp67_ASAP7_75t_L g13212 ( 
.A(n_12006),
.Y(n_13212)
);

INVx1_ASAP7_75t_L g13213 ( 
.A(n_12285),
.Y(n_13213)
);

INVx2_ASAP7_75t_SL g13214 ( 
.A(n_12017),
.Y(n_13214)
);

NAND2xp5_ASAP7_75t_L g13215 ( 
.A(n_12113),
.B(n_10455),
.Y(n_13215)
);

BUFx6f_ASAP7_75t_L g13216 ( 
.A(n_12142),
.Y(n_13216)
);

OR2x2_ASAP7_75t_L g13217 ( 
.A(n_11587),
.B(n_10456),
.Y(n_13217)
);

AND2x2_ASAP7_75t_SL g13218 ( 
.A(n_11508),
.B(n_8291),
.Y(n_13218)
);

AND2x2_ASAP7_75t_L g13219 ( 
.A(n_11590),
.B(n_11829),
.Y(n_13219)
);

AND2x2_ASAP7_75t_L g13220 ( 
.A(n_12025),
.B(n_8831),
.Y(n_13220)
);

NOR2xp33_ASAP7_75t_L g13221 ( 
.A(n_11708),
.B(n_6368),
.Y(n_13221)
);

INVx1_ASAP7_75t_L g13222 ( 
.A(n_12081),
.Y(n_13222)
);

AND2x2_ASAP7_75t_L g13223 ( 
.A(n_12029),
.B(n_12054),
.Y(n_13223)
);

AND2x2_ASAP7_75t_L g13224 ( 
.A(n_11715),
.B(n_8831),
.Y(n_13224)
);

OR2x2_ASAP7_75t_L g13225 ( 
.A(n_11502),
.B(n_10457),
.Y(n_13225)
);

INVx1_ASAP7_75t_L g13226 ( 
.A(n_12241),
.Y(n_13226)
);

AND2x2_ASAP7_75t_L g13227 ( 
.A(n_11482),
.B(n_8910),
.Y(n_13227)
);

INVx2_ASAP7_75t_SL g13228 ( 
.A(n_12206),
.Y(n_13228)
);

INVx1_ASAP7_75t_L g13229 ( 
.A(n_12136),
.Y(n_13229)
);

HB1xp67_ASAP7_75t_L g13230 ( 
.A(n_12073),
.Y(n_13230)
);

HB1xp67_ASAP7_75t_L g13231 ( 
.A(n_11762),
.Y(n_13231)
);

INVx4_ASAP7_75t_R g13232 ( 
.A(n_12400),
.Y(n_13232)
);

NOR2xp33_ASAP7_75t_L g13233 ( 
.A(n_11472),
.B(n_6368),
.Y(n_13233)
);

AND2x2_ASAP7_75t_L g13234 ( 
.A(n_12150),
.B(n_8910),
.Y(n_13234)
);

INVx2_ASAP7_75t_L g13235 ( 
.A(n_12286),
.Y(n_13235)
);

INVx1_ASAP7_75t_L g13236 ( 
.A(n_12208),
.Y(n_13236)
);

NAND2x1p5_ASAP7_75t_L g13237 ( 
.A(n_12098),
.B(n_8417),
.Y(n_13237)
);

OR2x2_ASAP7_75t_L g13238 ( 
.A(n_11683),
.B(n_10459),
.Y(n_13238)
);

NAND2xp5_ASAP7_75t_L g13239 ( 
.A(n_11515),
.B(n_10465),
.Y(n_13239)
);

INVx1_ASAP7_75t_L g13240 ( 
.A(n_12210),
.Y(n_13240)
);

BUFx3_ASAP7_75t_L g13241 ( 
.A(n_12304),
.Y(n_13241)
);

INVx1_ASAP7_75t_L g13242 ( 
.A(n_11719),
.Y(n_13242)
);

AND2x2_ASAP7_75t_L g13243 ( 
.A(n_12310),
.B(n_12322),
.Y(n_13243)
);

AND2x4_ASAP7_75t_L g13244 ( 
.A(n_12378),
.B(n_12384),
.Y(n_13244)
);

INVx1_ASAP7_75t_L g13245 ( 
.A(n_11796),
.Y(n_13245)
);

INVx2_ASAP7_75t_L g13246 ( 
.A(n_12148),
.Y(n_13246)
);

AND2x4_ASAP7_75t_L g13247 ( 
.A(n_12385),
.B(n_10466),
.Y(n_13247)
);

AOI22xp33_ASAP7_75t_SL g13248 ( 
.A1(n_11647),
.A2(n_7968),
.B1(n_7980),
.B2(n_7951),
.Y(n_13248)
);

BUFx6f_ASAP7_75t_L g13249 ( 
.A(n_12085),
.Y(n_13249)
);

AND2x2_ASAP7_75t_L g13250 ( 
.A(n_12140),
.B(n_8910),
.Y(n_13250)
);

AND2x4_ASAP7_75t_L g13251 ( 
.A(n_12399),
.B(n_10467),
.Y(n_13251)
);

OR2x2_ASAP7_75t_L g13252 ( 
.A(n_11658),
.B(n_10470),
.Y(n_13252)
);

OR2x2_ASAP7_75t_L g13253 ( 
.A(n_11574),
.B(n_11591),
.Y(n_13253)
);

AND2x4_ASAP7_75t_L g13254 ( 
.A(n_11930),
.B(n_10471),
.Y(n_13254)
);

INVx1_ASAP7_75t_L g13255 ( 
.A(n_11736),
.Y(n_13255)
);

OR2x2_ASAP7_75t_L g13256 ( 
.A(n_12190),
.B(n_10472),
.Y(n_13256)
);

NAND2xp5_ASAP7_75t_L g13257 ( 
.A(n_11561),
.B(n_10473),
.Y(n_13257)
);

AND2x2_ASAP7_75t_L g13258 ( 
.A(n_12170),
.B(n_8910),
.Y(n_13258)
);

BUFx2_ASAP7_75t_L g13259 ( 
.A(n_11743),
.Y(n_13259)
);

INVx1_ASAP7_75t_L g13260 ( 
.A(n_11739),
.Y(n_13260)
);

INVx2_ASAP7_75t_L g13261 ( 
.A(n_11814),
.Y(n_13261)
);

INVx3_ASAP7_75t_L g13262 ( 
.A(n_12319),
.Y(n_13262)
);

AND2x2_ASAP7_75t_L g13263 ( 
.A(n_12175),
.B(n_8910),
.Y(n_13263)
);

BUFx3_ASAP7_75t_L g13264 ( 
.A(n_12247),
.Y(n_13264)
);

INVx2_ASAP7_75t_L g13265 ( 
.A(n_11819),
.Y(n_13265)
);

OR2x2_ASAP7_75t_L g13266 ( 
.A(n_11469),
.B(n_10476),
.Y(n_13266)
);

BUFx3_ASAP7_75t_L g13267 ( 
.A(n_12280),
.Y(n_13267)
);

OR2x2_ASAP7_75t_L g13268 ( 
.A(n_11635),
.B(n_10480),
.Y(n_13268)
);

INVx2_ASAP7_75t_L g13269 ( 
.A(n_12137),
.Y(n_13269)
);

INVx2_ASAP7_75t_L g13270 ( 
.A(n_12146),
.Y(n_13270)
);

OR2x6_ASAP7_75t_SL g13271 ( 
.A(n_11717),
.B(n_5222),
.Y(n_13271)
);

AND2x4_ASAP7_75t_L g13272 ( 
.A(n_12178),
.B(n_10482),
.Y(n_13272)
);

AND2x2_ASAP7_75t_L g13273 ( 
.A(n_12186),
.B(n_10484),
.Y(n_13273)
);

AND2x2_ASAP7_75t_L g13274 ( 
.A(n_11652),
.B(n_10486),
.Y(n_13274)
);

AND2x2_ASAP7_75t_L g13275 ( 
.A(n_12156),
.B(n_10489),
.Y(n_13275)
);

INVxp67_ASAP7_75t_L g13276 ( 
.A(n_11972),
.Y(n_13276)
);

INVx1_ASAP7_75t_L g13277 ( 
.A(n_11817),
.Y(n_13277)
);

INVx2_ASAP7_75t_L g13278 ( 
.A(n_12189),
.Y(n_13278)
);

NOR2xp33_ASAP7_75t_L g13279 ( 
.A(n_12400),
.B(n_6368),
.Y(n_13279)
);

OAI22xp5_ASAP7_75t_L g13280 ( 
.A1(n_11542),
.A2(n_7798),
.B1(n_7811),
.B2(n_7769),
.Y(n_13280)
);

INVx1_ASAP7_75t_L g13281 ( 
.A(n_11827),
.Y(n_13281)
);

AND2x2_ASAP7_75t_L g13282 ( 
.A(n_11852),
.B(n_10494),
.Y(n_13282)
);

INVx1_ASAP7_75t_L g13283 ( 
.A(n_11645),
.Y(n_13283)
);

INVxp67_ASAP7_75t_SL g13284 ( 
.A(n_11595),
.Y(n_13284)
);

OR2x2_ASAP7_75t_L g13285 ( 
.A(n_11644),
.B(n_10495),
.Y(n_13285)
);

AND2x4_ASAP7_75t_L g13286 ( 
.A(n_12411),
.B(n_10496),
.Y(n_13286)
);

INVx2_ASAP7_75t_R g13287 ( 
.A(n_11914),
.Y(n_13287)
);

HB1xp67_ASAP7_75t_L g13288 ( 
.A(n_11665),
.Y(n_13288)
);

NOR2x1_ASAP7_75t_L g13289 ( 
.A(n_11946),
.B(n_9096),
.Y(n_13289)
);

OR2x2_ASAP7_75t_L g13290 ( 
.A(n_11747),
.B(n_10497),
.Y(n_13290)
);

INVx1_ASAP7_75t_L g13291 ( 
.A(n_12403),
.Y(n_13291)
);

NAND2xp5_ASAP7_75t_L g13292 ( 
.A(n_11536),
.B(n_11866),
.Y(n_13292)
);

INVx1_ASAP7_75t_L g13293 ( 
.A(n_12375),
.Y(n_13293)
);

NAND2x1p5_ASAP7_75t_SL g13294 ( 
.A(n_11560),
.B(n_7720),
.Y(n_13294)
);

NAND2xp5_ASAP7_75t_L g13295 ( 
.A(n_11552),
.B(n_10498),
.Y(n_13295)
);

NAND2xp5_ASAP7_75t_L g13296 ( 
.A(n_11847),
.B(n_10502),
.Y(n_13296)
);

INVx3_ASAP7_75t_L g13297 ( 
.A(n_12261),
.Y(n_13297)
);

INVx1_ASAP7_75t_L g13298 ( 
.A(n_12165),
.Y(n_13298)
);

BUFx3_ASAP7_75t_L g13299 ( 
.A(n_12086),
.Y(n_13299)
);

INVx1_ASAP7_75t_L g13300 ( 
.A(n_12389),
.Y(n_13300)
);

INVx2_ASAP7_75t_L g13301 ( 
.A(n_12394),
.Y(n_13301)
);

INVx1_ASAP7_75t_L g13302 ( 
.A(n_11679),
.Y(n_13302)
);

OR2x2_ASAP7_75t_L g13303 ( 
.A(n_11769),
.B(n_11583),
.Y(n_13303)
);

BUFx2_ASAP7_75t_L g13304 ( 
.A(n_11578),
.Y(n_13304)
);

INVxp67_ASAP7_75t_L g13305 ( 
.A(n_12048),
.Y(n_13305)
);

BUFx3_ASAP7_75t_L g13306 ( 
.A(n_12011),
.Y(n_13306)
);

NAND2xp5_ASAP7_75t_L g13307 ( 
.A(n_12099),
.B(n_10509),
.Y(n_13307)
);

OR2x2_ASAP7_75t_L g13308 ( 
.A(n_11884),
.B(n_10510),
.Y(n_13308)
);

BUFx3_ASAP7_75t_L g13309 ( 
.A(n_11562),
.Y(n_13309)
);

INVx1_ASAP7_75t_SL g13310 ( 
.A(n_11487),
.Y(n_13310)
);

BUFx2_ASAP7_75t_L g13311 ( 
.A(n_12078),
.Y(n_13311)
);

AND2x2_ASAP7_75t_L g13312 ( 
.A(n_12131),
.B(n_10512),
.Y(n_13312)
);

OR2x2_ASAP7_75t_L g13313 ( 
.A(n_11688),
.B(n_10513),
.Y(n_13313)
);

AND2x2_ASAP7_75t_L g13314 ( 
.A(n_11576),
.B(n_10517),
.Y(n_13314)
);

BUFx3_ASAP7_75t_L g13315 ( 
.A(n_12382),
.Y(n_13315)
);

AND2x2_ASAP7_75t_L g13316 ( 
.A(n_11577),
.B(n_10518),
.Y(n_13316)
);

INVx2_ASAP7_75t_L g13317 ( 
.A(n_11833),
.Y(n_13317)
);

HB1xp67_ASAP7_75t_L g13318 ( 
.A(n_11969),
.Y(n_13318)
);

HB1xp67_ASAP7_75t_L g13319 ( 
.A(n_11886),
.Y(n_13319)
);

NAND2xp5_ASAP7_75t_L g13320 ( 
.A(n_11892),
.B(n_10521),
.Y(n_13320)
);

NAND2xp5_ASAP7_75t_L g13321 ( 
.A(n_11753),
.B(n_10527),
.Y(n_13321)
);

NAND2xp5_ASAP7_75t_L g13322 ( 
.A(n_12090),
.B(n_11916),
.Y(n_13322)
);

INVx1_ASAP7_75t_L g13323 ( 
.A(n_12434),
.Y(n_13323)
);

AND2x2_ASAP7_75t_L g13324 ( 
.A(n_12457),
.B(n_11623),
.Y(n_13324)
);

AND2x2_ASAP7_75t_L g13325 ( 
.A(n_12693),
.B(n_12187),
.Y(n_13325)
);

AND2x2_ASAP7_75t_L g13326 ( 
.A(n_12786),
.B(n_12124),
.Y(n_13326)
);

NAND2xp5_ASAP7_75t_L g13327 ( 
.A(n_12645),
.B(n_11572),
.Y(n_13327)
);

OR2x2_ASAP7_75t_L g13328 ( 
.A(n_12467),
.B(n_12093),
.Y(n_13328)
);

INVx3_ASAP7_75t_L g13329 ( 
.A(n_12527),
.Y(n_13329)
);

NAND2xp5_ASAP7_75t_L g13330 ( 
.A(n_13262),
.B(n_11723),
.Y(n_13330)
);

INVx2_ASAP7_75t_L g13331 ( 
.A(n_12584),
.Y(n_13331)
);

AND2x2_ASAP7_75t_L g13332 ( 
.A(n_12700),
.B(n_12348),
.Y(n_13332)
);

AND2x2_ASAP7_75t_L g13333 ( 
.A(n_12640),
.B(n_11943),
.Y(n_13333)
);

INVx1_ASAP7_75t_L g13334 ( 
.A(n_12439),
.Y(n_13334)
);

OR2x2_ASAP7_75t_L g13335 ( 
.A(n_12482),
.B(n_11558),
.Y(n_13335)
);

NAND2xp5_ASAP7_75t_L g13336 ( 
.A(n_13262),
.B(n_12065),
.Y(n_13336)
);

BUFx3_ASAP7_75t_L g13337 ( 
.A(n_12607),
.Y(n_13337)
);

AND2x2_ASAP7_75t_L g13338 ( 
.A(n_12558),
.B(n_12130),
.Y(n_13338)
);

AND2x2_ASAP7_75t_L g13339 ( 
.A(n_12483),
.B(n_11858),
.Y(n_13339)
);

AND2x2_ASAP7_75t_L g13340 ( 
.A(n_12615),
.B(n_12392),
.Y(n_13340)
);

AND2x2_ASAP7_75t_L g13341 ( 
.A(n_12487),
.B(n_11823),
.Y(n_13341)
);

AND2x2_ASAP7_75t_L g13342 ( 
.A(n_12516),
.B(n_12084),
.Y(n_13342)
);

INVx1_ASAP7_75t_SL g13343 ( 
.A(n_12599),
.Y(n_13343)
);

AND2x4_ASAP7_75t_L g13344 ( 
.A(n_12491),
.B(n_10622),
.Y(n_13344)
);

AND2x2_ASAP7_75t_L g13345 ( 
.A(n_12546),
.B(n_12128),
.Y(n_13345)
);

INVx2_ASAP7_75t_L g13346 ( 
.A(n_12550),
.Y(n_13346)
);

INVx2_ASAP7_75t_L g13347 ( 
.A(n_12607),
.Y(n_13347)
);

NOR2xp67_ASAP7_75t_L g13348 ( 
.A(n_12722),
.B(n_12022),
.Y(n_13348)
);

OAI22xp5_ASAP7_75t_L g13349 ( 
.A1(n_12893),
.A2(n_12213),
.B1(n_12216),
.B2(n_12214),
.Y(n_13349)
);

NAND2xp5_ASAP7_75t_L g13350 ( 
.A(n_13136),
.B(n_12087),
.Y(n_13350)
);

NOR2xp33_ASAP7_75t_SL g13351 ( 
.A(n_12565),
.B(n_11935),
.Y(n_13351)
);

BUFx8_ASAP7_75t_SL g13352 ( 
.A(n_12606),
.Y(n_13352)
);

INVx2_ASAP7_75t_L g13353 ( 
.A(n_12501),
.Y(n_13353)
);

AND2x2_ASAP7_75t_L g13354 ( 
.A(n_12650),
.B(n_11836),
.Y(n_13354)
);

HB1xp67_ASAP7_75t_L g13355 ( 
.A(n_12421),
.Y(n_13355)
);

INVx2_ASAP7_75t_L g13356 ( 
.A(n_12501),
.Y(n_13356)
);

INVxp67_ASAP7_75t_L g13357 ( 
.A(n_12440),
.Y(n_13357)
);

INVx2_ASAP7_75t_L g13358 ( 
.A(n_12622),
.Y(n_13358)
);

INVxp67_ASAP7_75t_L g13359 ( 
.A(n_12810),
.Y(n_13359)
);

INVx1_ASAP7_75t_L g13360 ( 
.A(n_12449),
.Y(n_13360)
);

INVx4_ASAP7_75t_L g13361 ( 
.A(n_12606),
.Y(n_13361)
);

INVx1_ASAP7_75t_L g13362 ( 
.A(n_12476),
.Y(n_13362)
);

OR2x2_ASAP7_75t_L g13363 ( 
.A(n_12479),
.B(n_11735),
.Y(n_13363)
);

AND2x2_ASAP7_75t_L g13364 ( 
.A(n_12462),
.B(n_12464),
.Y(n_13364)
);

AND2x2_ASAP7_75t_L g13365 ( 
.A(n_12801),
.B(n_11873),
.Y(n_13365)
);

OAI22xp5_ASAP7_75t_L g13366 ( 
.A1(n_13038),
.A2(n_12258),
.B1(n_12296),
.B2(n_11918),
.Y(n_13366)
);

NAND2x1_ASAP7_75t_L g13367 ( 
.A(n_12945),
.B(n_12240),
.Y(n_13367)
);

AOI22xp33_ASAP7_75t_SL g13368 ( 
.A1(n_13138),
.A2(n_11888),
.B1(n_12014),
.B2(n_11845),
.Y(n_13368)
);

INVx3_ASAP7_75t_L g13369 ( 
.A(n_12491),
.Y(n_13369)
);

AOI22xp33_ASAP7_75t_SL g13370 ( 
.A1(n_13187),
.A2(n_11664),
.B1(n_11902),
.B2(n_12119),
.Y(n_13370)
);

INVx1_ASAP7_75t_L g13371 ( 
.A(n_12891),
.Y(n_13371)
);

INVx2_ASAP7_75t_SL g13372 ( 
.A(n_12722),
.Y(n_13372)
);

INVx2_ASAP7_75t_L g13373 ( 
.A(n_12622),
.Y(n_13373)
);

INVx1_ASAP7_75t_L g13374 ( 
.A(n_12416),
.Y(n_13374)
);

INVx1_ASAP7_75t_L g13375 ( 
.A(n_12416),
.Y(n_13375)
);

INVx1_ASAP7_75t_L g13376 ( 
.A(n_12420),
.Y(n_13376)
);

AND2x2_ASAP7_75t_L g13377 ( 
.A(n_12506),
.B(n_12028),
.Y(n_13377)
);

INVx2_ASAP7_75t_L g13378 ( 
.A(n_12759),
.Y(n_13378)
);

INVx2_ASAP7_75t_L g13379 ( 
.A(n_12759),
.Y(n_13379)
);

INVx2_ASAP7_75t_L g13380 ( 
.A(n_12722),
.Y(n_13380)
);

NAND2xp5_ASAP7_75t_L g13381 ( 
.A(n_12507),
.B(n_11867),
.Y(n_13381)
);

OR2x2_ASAP7_75t_L g13382 ( 
.A(n_12430),
.B(n_12415),
.Y(n_13382)
);

AOI21xp33_ASAP7_75t_L g13383 ( 
.A1(n_12784),
.A2(n_11669),
.B(n_11795),
.Y(n_13383)
);

INVx2_ASAP7_75t_L g13384 ( 
.A(n_12791),
.Y(n_13384)
);

NOR2xp33_ASAP7_75t_L g13385 ( 
.A(n_12519),
.B(n_5019),
.Y(n_13385)
);

BUFx3_ASAP7_75t_L g13386 ( 
.A(n_12494),
.Y(n_13386)
);

NAND2xp5_ASAP7_75t_L g13387 ( 
.A(n_12718),
.B(n_11718),
.Y(n_13387)
);

INVx1_ASAP7_75t_L g13388 ( 
.A(n_12420),
.Y(n_13388)
);

AND2x2_ASAP7_75t_L g13389 ( 
.A(n_12419),
.B(n_12050),
.Y(n_13389)
);

INVx1_ASAP7_75t_L g13390 ( 
.A(n_12425),
.Y(n_13390)
);

AND2x2_ASAP7_75t_L g13391 ( 
.A(n_12428),
.B(n_12376),
.Y(n_13391)
);

NAND2xp5_ASAP7_75t_L g13392 ( 
.A(n_12521),
.B(n_11936),
.Y(n_13392)
);

HB1xp67_ASAP7_75t_L g13393 ( 
.A(n_12663),
.Y(n_13393)
);

AND2x2_ASAP7_75t_L g13394 ( 
.A(n_12732),
.B(n_12391),
.Y(n_13394)
);

AND2x2_ASAP7_75t_L g13395 ( 
.A(n_12757),
.B(n_12125),
.Y(n_13395)
);

AND2x2_ASAP7_75t_L g13396 ( 
.A(n_12563),
.B(n_10534),
.Y(n_13396)
);

INVx1_ASAP7_75t_L g13397 ( 
.A(n_12425),
.Y(n_13397)
);

INVx3_ASAP7_75t_L g13398 ( 
.A(n_12791),
.Y(n_13398)
);

INVxp67_ASAP7_75t_L g13399 ( 
.A(n_12543),
.Y(n_13399)
);

AOI22xp33_ASAP7_75t_SL g13400 ( 
.A1(n_13038),
.A2(n_12230),
.B1(n_12120),
.B2(n_12215),
.Y(n_13400)
);

AOI22xp33_ASAP7_75t_L g13401 ( 
.A1(n_13287),
.A2(n_12000),
.B1(n_12220),
.B2(n_12200),
.Y(n_13401)
);

INVx1_ASAP7_75t_L g13402 ( 
.A(n_12436),
.Y(n_13402)
);

AND2x4_ASAP7_75t_L g13403 ( 
.A(n_12484),
.B(n_12438),
.Y(n_13403)
);

HB1xp67_ASAP7_75t_L g13404 ( 
.A(n_12990),
.Y(n_13404)
);

INVx1_ASAP7_75t_L g13405 ( 
.A(n_12436),
.Y(n_13405)
);

NAND2xp5_ASAP7_75t_L g13406 ( 
.A(n_12876),
.B(n_12345),
.Y(n_13406)
);

AND2x2_ASAP7_75t_L g13407 ( 
.A(n_12564),
.B(n_10542),
.Y(n_13407)
);

OR2x2_ASAP7_75t_L g13408 ( 
.A(n_12535),
.B(n_12492),
.Y(n_13408)
);

INVx1_ASAP7_75t_L g13409 ( 
.A(n_12437),
.Y(n_13409)
);

BUFx2_ASAP7_75t_L g13410 ( 
.A(n_13015),
.Y(n_13410)
);

INVx1_ASAP7_75t_L g13411 ( 
.A(n_12437),
.Y(n_13411)
);

OAI211xp5_ASAP7_75t_SL g13412 ( 
.A1(n_13177),
.A2(n_13130),
.B(n_13025),
.C(n_13081),
.Y(n_13412)
);

BUFx3_ASAP7_75t_L g13413 ( 
.A(n_12495),
.Y(n_13413)
);

AND2x2_ASAP7_75t_L g13414 ( 
.A(n_12567),
.B(n_10546),
.Y(n_13414)
);

INVx1_ASAP7_75t_SL g13415 ( 
.A(n_12596),
.Y(n_13415)
);

AND2x2_ASAP7_75t_L g13416 ( 
.A(n_12733),
.B(n_10553),
.Y(n_13416)
);

AND2x2_ASAP7_75t_L g13417 ( 
.A(n_12435),
.B(n_10559),
.Y(n_13417)
);

INVx2_ASAP7_75t_L g13418 ( 
.A(n_12791),
.Y(n_13418)
);

INVx1_ASAP7_75t_L g13419 ( 
.A(n_12441),
.Y(n_13419)
);

INVx2_ASAP7_75t_L g13420 ( 
.A(n_12442),
.Y(n_13420)
);

AND2x4_ASAP7_75t_L g13421 ( 
.A(n_12578),
.B(n_10622),
.Y(n_13421)
);

AND2x2_ASAP7_75t_L g13422 ( 
.A(n_12443),
.B(n_10562),
.Y(n_13422)
);

AND2x2_ASAP7_75t_L g13423 ( 
.A(n_12485),
.B(n_10569),
.Y(n_13423)
);

INVx2_ASAP7_75t_L g13424 ( 
.A(n_12442),
.Y(n_13424)
);

AND2x2_ASAP7_75t_L g13425 ( 
.A(n_12445),
.B(n_10574),
.Y(n_13425)
);

INVx1_ASAP7_75t_L g13426 ( 
.A(n_12441),
.Y(n_13426)
);

AND2x2_ASAP7_75t_L g13427 ( 
.A(n_12448),
.B(n_10582),
.Y(n_13427)
);

AOI22xp33_ASAP7_75t_L g13428 ( 
.A1(n_13204),
.A2(n_12024),
.B1(n_12199),
.B2(n_12157),
.Y(n_13428)
);

OR2x2_ASAP7_75t_L g13429 ( 
.A(n_13107),
.B(n_10622),
.Y(n_13429)
);

AND2x2_ASAP7_75t_L g13430 ( 
.A(n_12452),
.B(n_10584),
.Y(n_13430)
);

AND2x2_ASAP7_75t_L g13431 ( 
.A(n_12454),
.B(n_10586),
.Y(n_13431)
);

AND2x2_ASAP7_75t_L g13432 ( 
.A(n_12414),
.B(n_10590),
.Y(n_13432)
);

NOR2xp33_ASAP7_75t_L g13433 ( 
.A(n_12606),
.B(n_12424),
.Y(n_13433)
);

INVx1_ASAP7_75t_L g13434 ( 
.A(n_12446),
.Y(n_13434)
);

CKINVDCx20_ASAP7_75t_R g13435 ( 
.A(n_12766),
.Y(n_13435)
);

AND2x2_ASAP7_75t_L g13436 ( 
.A(n_12423),
.B(n_10592),
.Y(n_13436)
);

AND2x2_ASAP7_75t_L g13437 ( 
.A(n_12542),
.B(n_10594),
.Y(n_13437)
);

AND2x2_ASAP7_75t_L g13438 ( 
.A(n_12542),
.B(n_10597),
.Y(n_13438)
);

INVxp67_ASAP7_75t_L g13439 ( 
.A(n_12560),
.Y(n_13439)
);

INVx2_ASAP7_75t_L g13440 ( 
.A(n_12765),
.Y(n_13440)
);

NAND2xp5_ASAP7_75t_L g13441 ( 
.A(n_13074),
.B(n_12350),
.Y(n_13441)
);

INVx1_ASAP7_75t_L g13442 ( 
.A(n_12446),
.Y(n_13442)
);

HB1xp67_ASAP7_75t_L g13443 ( 
.A(n_13063),
.Y(n_13443)
);

AND2x2_ASAP7_75t_L g13444 ( 
.A(n_12512),
.B(n_10598),
.Y(n_13444)
);

INVx1_ASAP7_75t_L g13445 ( 
.A(n_12451),
.Y(n_13445)
);

NAND2xp5_ASAP7_75t_L g13446 ( 
.A(n_13074),
.B(n_11643),
.Y(n_13446)
);

INVx1_ASAP7_75t_L g13447 ( 
.A(n_12451),
.Y(n_13447)
);

HB1xp67_ASAP7_75t_L g13448 ( 
.A(n_12697),
.Y(n_13448)
);

NAND2xp5_ASAP7_75t_L g13449 ( 
.A(n_13231),
.B(n_12352),
.Y(n_13449)
);

OAI22xp5_ASAP7_75t_L g13450 ( 
.A1(n_13304),
.A2(n_12158),
.B1(n_12362),
.B2(n_12354),
.Y(n_13450)
);

NAND2xp5_ASAP7_75t_L g13451 ( 
.A(n_13019),
.B(n_12115),
.Y(n_13451)
);

OR2x2_ASAP7_75t_L g13452 ( 
.A(n_13225),
.B(n_10622),
.Y(n_13452)
);

INVxp33_ASAP7_75t_L g13453 ( 
.A(n_12687),
.Y(n_13453)
);

INVxp67_ASAP7_75t_SL g13454 ( 
.A(n_12461),
.Y(n_13454)
);

INVx1_ASAP7_75t_L g13455 ( 
.A(n_12456),
.Y(n_13455)
);

INVx1_ASAP7_75t_L g13456 ( 
.A(n_12456),
.Y(n_13456)
);

INVx2_ASAP7_75t_L g13457 ( 
.A(n_12756),
.Y(n_13457)
);

AND2x4_ASAP7_75t_L g13458 ( 
.A(n_12588),
.B(n_11066),
.Y(n_13458)
);

HB1xp67_ASAP7_75t_L g13459 ( 
.A(n_12798),
.Y(n_13459)
);

INVx1_ASAP7_75t_L g13460 ( 
.A(n_12458),
.Y(n_13460)
);

AND2x2_ASAP7_75t_L g13461 ( 
.A(n_12523),
.B(n_10604),
.Y(n_13461)
);

INVx2_ASAP7_75t_L g13462 ( 
.A(n_12618),
.Y(n_13462)
);

INVx1_ASAP7_75t_L g13463 ( 
.A(n_12458),
.Y(n_13463)
);

AND2x4_ASAP7_75t_L g13464 ( 
.A(n_12669),
.B(n_11066),
.Y(n_13464)
);

HB1xp67_ASAP7_75t_L g13465 ( 
.A(n_12710),
.Y(n_13465)
);

AND2x2_ASAP7_75t_L g13466 ( 
.A(n_12529),
.B(n_10606),
.Y(n_13466)
);

AND2x2_ASAP7_75t_L g13467 ( 
.A(n_12712),
.B(n_10607),
.Y(n_13467)
);

INVx1_ASAP7_75t_L g13468 ( 
.A(n_12468),
.Y(n_13468)
);

NAND2xp5_ASAP7_75t_L g13469 ( 
.A(n_12525),
.B(n_12147),
.Y(n_13469)
);

INVx3_ASAP7_75t_L g13470 ( 
.A(n_12777),
.Y(n_13470)
);

INVx2_ASAP7_75t_L g13471 ( 
.A(n_12618),
.Y(n_13471)
);

INVx1_ASAP7_75t_L g13472 ( 
.A(n_12468),
.Y(n_13472)
);

AOI22xp33_ASAP7_75t_L g13473 ( 
.A1(n_13143),
.A2(n_11636),
.B1(n_11695),
.B2(n_11697),
.Y(n_13473)
);

NAND2xp5_ASAP7_75t_L g13474 ( 
.A(n_12652),
.B(n_12386),
.Y(n_13474)
);

BUFx2_ASAP7_75t_L g13475 ( 
.A(n_12576),
.Y(n_13475)
);

INVx1_ASAP7_75t_L g13476 ( 
.A(n_12469),
.Y(n_13476)
);

AND2x4_ASAP7_75t_L g13477 ( 
.A(n_12669),
.B(n_11066),
.Y(n_13477)
);

INVx1_ASAP7_75t_L g13478 ( 
.A(n_12469),
.Y(n_13478)
);

INVx1_ASAP7_75t_L g13479 ( 
.A(n_12472),
.Y(n_13479)
);

INVx4_ASAP7_75t_L g13480 ( 
.A(n_12496),
.Y(n_13480)
);

INVx1_ASAP7_75t_SL g13481 ( 
.A(n_12496),
.Y(n_13481)
);

AND2x2_ASAP7_75t_L g13482 ( 
.A(n_12466),
.B(n_10612),
.Y(n_13482)
);

OR2x2_ASAP7_75t_L g13483 ( 
.A(n_12602),
.B(n_10614),
.Y(n_13483)
);

INVx2_ASAP7_75t_L g13484 ( 
.A(n_12779),
.Y(n_13484)
);

INVx1_ASAP7_75t_L g13485 ( 
.A(n_12472),
.Y(n_13485)
);

NAND2xp5_ASAP7_75t_L g13486 ( 
.A(n_12627),
.B(n_12764),
.Y(n_13486)
);

INVx1_ASAP7_75t_L g13487 ( 
.A(n_12473),
.Y(n_13487)
);

INVx2_ASAP7_75t_L g13488 ( 
.A(n_12779),
.Y(n_13488)
);

OR2x2_ASAP7_75t_L g13489 ( 
.A(n_13170),
.B(n_10618),
.Y(n_13489)
);

HB1xp67_ASAP7_75t_L g13490 ( 
.A(n_12625),
.Y(n_13490)
);

AND2x2_ASAP7_75t_L g13491 ( 
.A(n_12466),
.B(n_10621),
.Y(n_13491)
);

INVx3_ASAP7_75t_L g13492 ( 
.A(n_12777),
.Y(n_13492)
);

INVx1_ASAP7_75t_L g13493 ( 
.A(n_12473),
.Y(n_13493)
);

INVx1_ASAP7_75t_L g13494 ( 
.A(n_12474),
.Y(n_13494)
);

NAND2xp5_ASAP7_75t_L g13495 ( 
.A(n_13116),
.B(n_10624),
.Y(n_13495)
);

AND2x4_ASAP7_75t_SL g13496 ( 
.A(n_12471),
.B(n_8052),
.Y(n_13496)
);

AND2x2_ASAP7_75t_L g13497 ( 
.A(n_12429),
.B(n_10629),
.Y(n_13497)
);

OR2x2_ASAP7_75t_L g13498 ( 
.A(n_13268),
.B(n_10641),
.Y(n_13498)
);

NOR2x1_ASAP7_75t_L g13499 ( 
.A(n_13121),
.B(n_12126),
.Y(n_13499)
);

OR2x2_ASAP7_75t_L g13500 ( 
.A(n_13285),
.B(n_10652),
.Y(n_13500)
);

INVx1_ASAP7_75t_L g13501 ( 
.A(n_12474),
.Y(n_13501)
);

AND2x4_ASAP7_75t_L g13502 ( 
.A(n_12522),
.B(n_11066),
.Y(n_13502)
);

INVx2_ASAP7_75t_L g13503 ( 
.A(n_12816),
.Y(n_13503)
);

AND2x2_ASAP7_75t_L g13504 ( 
.A(n_12431),
.B(n_10655),
.Y(n_13504)
);

AND2x2_ASAP7_75t_L g13505 ( 
.A(n_12617),
.B(n_10656),
.Y(n_13505)
);

AOI22xp33_ASAP7_75t_L g13506 ( 
.A1(n_13297),
.A2(n_12092),
.B1(n_12181),
.B2(n_11659),
.Y(n_13506)
);

INVx1_ASAP7_75t_L g13507 ( 
.A(n_12480),
.Y(n_13507)
);

INVx1_ASAP7_75t_L g13508 ( 
.A(n_12480),
.Y(n_13508)
);

OR2x2_ASAP7_75t_L g13509 ( 
.A(n_13238),
.B(n_10657),
.Y(n_13509)
);

BUFx3_ASAP7_75t_L g13510 ( 
.A(n_12557),
.Y(n_13510)
);

INVx2_ASAP7_75t_L g13511 ( 
.A(n_12655),
.Y(n_13511)
);

HB1xp67_ASAP7_75t_L g13512 ( 
.A(n_12637),
.Y(n_13512)
);

INVx1_ASAP7_75t_L g13513 ( 
.A(n_12432),
.Y(n_13513)
);

OR2x2_ASAP7_75t_L g13514 ( 
.A(n_13132),
.B(n_10661),
.Y(n_13514)
);

AND2x2_ASAP7_75t_L g13515 ( 
.A(n_12561),
.B(n_10665),
.Y(n_13515)
);

AND2x2_ASAP7_75t_L g13516 ( 
.A(n_12566),
.B(n_10666),
.Y(n_13516)
);

INVx1_ASAP7_75t_L g13517 ( 
.A(n_12450),
.Y(n_13517)
);

INVx2_ASAP7_75t_L g13518 ( 
.A(n_12668),
.Y(n_13518)
);

OR2x2_ASAP7_75t_L g13519 ( 
.A(n_13132),
.B(n_10669),
.Y(n_13519)
);

INVx1_ASAP7_75t_SL g13520 ( 
.A(n_12909),
.Y(n_13520)
);

AND2x2_ASAP7_75t_L g13521 ( 
.A(n_12568),
.B(n_10671),
.Y(n_13521)
);

INVx1_ASAP7_75t_L g13522 ( 
.A(n_12453),
.Y(n_13522)
);

INVx1_ASAP7_75t_L g13523 ( 
.A(n_12497),
.Y(n_13523)
);

INVx3_ASAP7_75t_L g13524 ( 
.A(n_12654),
.Y(n_13524)
);

OR2x2_ASAP7_75t_L g13525 ( 
.A(n_13134),
.B(n_10673),
.Y(n_13525)
);

NAND2xp5_ASAP7_75t_L g13526 ( 
.A(n_13062),
.B(n_10679),
.Y(n_13526)
);

INVx2_ASAP7_75t_L g13527 ( 
.A(n_12505),
.Y(n_13527)
);

INVx1_ASAP7_75t_L g13528 ( 
.A(n_12497),
.Y(n_13528)
);

AND2x2_ASAP7_75t_L g13529 ( 
.A(n_12847),
.B(n_10687),
.Y(n_13529)
);

INVx1_ASAP7_75t_L g13530 ( 
.A(n_12498),
.Y(n_13530)
);

AND2x2_ASAP7_75t_L g13531 ( 
.A(n_12889),
.B(n_10689),
.Y(n_13531)
);

OR2x2_ASAP7_75t_L g13532 ( 
.A(n_13134),
.B(n_12413),
.Y(n_13532)
);

AND2x2_ASAP7_75t_L g13533 ( 
.A(n_12488),
.B(n_10690),
.Y(n_13533)
);

INVx2_ASAP7_75t_L g13534 ( 
.A(n_12505),
.Y(n_13534)
);

OR2x2_ASAP7_75t_L g13535 ( 
.A(n_13181),
.B(n_10691),
.Y(n_13535)
);

AND2x2_ASAP7_75t_L g13536 ( 
.A(n_12490),
.B(n_10700),
.Y(n_13536)
);

AND2x2_ASAP7_75t_L g13537 ( 
.A(n_12594),
.B(n_12619),
.Y(n_13537)
);

OR2x2_ASAP7_75t_L g13538 ( 
.A(n_13217),
.B(n_10702),
.Y(n_13538)
);

AND2x2_ASAP7_75t_L g13539 ( 
.A(n_12537),
.B(n_10703),
.Y(n_13539)
);

AND2x4_ASAP7_75t_L g13540 ( 
.A(n_12534),
.B(n_10705),
.Y(n_13540)
);

OR2x2_ASAP7_75t_L g13541 ( 
.A(n_13083),
.B(n_10710),
.Y(n_13541)
);

NAND2x1p5_ASAP7_75t_L g13542 ( 
.A(n_12835),
.B(n_6628),
.Y(n_13542)
);

BUFx3_ASAP7_75t_L g13543 ( 
.A(n_12557),
.Y(n_13543)
);

INVx1_ASAP7_75t_L g13544 ( 
.A(n_12498),
.Y(n_13544)
);

INVx1_ASAP7_75t_L g13545 ( 
.A(n_12499),
.Y(n_13545)
);

INVx1_ASAP7_75t_L g13546 ( 
.A(n_12499),
.Y(n_13546)
);

OR2x2_ASAP7_75t_L g13547 ( 
.A(n_12601),
.B(n_10711),
.Y(n_13547)
);

INVx1_ASAP7_75t_L g13548 ( 
.A(n_12500),
.Y(n_13548)
);

INVx1_ASAP7_75t_L g13549 ( 
.A(n_12500),
.Y(n_13549)
);

INVx1_ASAP7_75t_L g13550 ( 
.A(n_12502),
.Y(n_13550)
);

INVx2_ASAP7_75t_L g13551 ( 
.A(n_12537),
.Y(n_13551)
);

INVx1_ASAP7_75t_L g13552 ( 
.A(n_12502),
.Y(n_13552)
);

INVx1_ASAP7_75t_L g13553 ( 
.A(n_12612),
.Y(n_13553)
);

INVx2_ASAP7_75t_L g13554 ( 
.A(n_12433),
.Y(n_13554)
);

AOI22xp33_ASAP7_75t_SL g13555 ( 
.A1(n_13297),
.A2(n_11984),
.B1(n_12110),
.B2(n_12121),
.Y(n_13555)
);

INVx1_ASAP7_75t_L g13556 ( 
.A(n_12612),
.Y(n_13556)
);

INVx3_ASAP7_75t_R g13557 ( 
.A(n_12985),
.Y(n_13557)
);

OR2x2_ASAP7_75t_L g13558 ( 
.A(n_13193),
.B(n_13194),
.Y(n_13558)
);

OR2x2_ASAP7_75t_L g13559 ( 
.A(n_13193),
.B(n_10717),
.Y(n_13559)
);

NOR2xp33_ASAP7_75t_L g13560 ( 
.A(n_12489),
.B(n_5037),
.Y(n_13560)
);

NAND2xp5_ASAP7_75t_L g13561 ( 
.A(n_12426),
.B(n_12427),
.Y(n_13561)
);

INVx1_ASAP7_75t_L g13562 ( 
.A(n_12624),
.Y(n_13562)
);

INVx1_ASAP7_75t_L g13563 ( 
.A(n_12624),
.Y(n_13563)
);

AOI21x1_ASAP7_75t_L g13564 ( 
.A1(n_13084),
.A2(n_12338),
.B(n_12276),
.Y(n_13564)
);

NAND2xp5_ASAP7_75t_L g13565 ( 
.A(n_12444),
.B(n_10720),
.Y(n_13565)
);

AND2x4_ASAP7_75t_L g13566 ( 
.A(n_12736),
.B(n_12738),
.Y(n_13566)
);

HB1xp67_ASAP7_75t_L g13567 ( 
.A(n_12838),
.Y(n_13567)
);

INVx1_ASAP7_75t_L g13568 ( 
.A(n_12626),
.Y(n_13568)
);

INVx2_ASAP7_75t_L g13569 ( 
.A(n_12433),
.Y(n_13569)
);

OR2x2_ASAP7_75t_L g13570 ( 
.A(n_13194),
.B(n_10722),
.Y(n_13570)
);

AND2x2_ASAP7_75t_L g13571 ( 
.A(n_12611),
.B(n_10733),
.Y(n_13571)
);

INVx1_ASAP7_75t_L g13572 ( 
.A(n_12626),
.Y(n_13572)
);

INVx2_ASAP7_75t_L g13573 ( 
.A(n_12885),
.Y(n_13573)
);

OR2x2_ASAP7_75t_L g13574 ( 
.A(n_13252),
.B(n_10734),
.Y(n_13574)
);

INVx2_ASAP7_75t_L g13575 ( 
.A(n_12885),
.Y(n_13575)
);

INVx1_ASAP7_75t_L g13576 ( 
.A(n_12667),
.Y(n_13576)
);

INVx1_ASAP7_75t_L g13577 ( 
.A(n_12667),
.Y(n_13577)
);

INVx1_ASAP7_75t_L g13578 ( 
.A(n_12672),
.Y(n_13578)
);

INVx2_ASAP7_75t_L g13579 ( 
.A(n_12885),
.Y(n_13579)
);

NAND2xp5_ASAP7_75t_L g13580 ( 
.A(n_12447),
.B(n_10735),
.Y(n_13580)
);

INVx1_ASAP7_75t_L g13581 ( 
.A(n_12672),
.Y(n_13581)
);

HB1xp67_ASAP7_75t_L g13582 ( 
.A(n_12838),
.Y(n_13582)
);

INVx1_ASAP7_75t_L g13583 ( 
.A(n_12681),
.Y(n_13583)
);

INVx1_ASAP7_75t_L g13584 ( 
.A(n_12681),
.Y(n_13584)
);

NAND2xp5_ASAP7_75t_L g13585 ( 
.A(n_12459),
.B(n_10738),
.Y(n_13585)
);

OR2x2_ASAP7_75t_L g13586 ( 
.A(n_13209),
.B(n_10748),
.Y(n_13586)
);

INVx3_ASAP7_75t_L g13587 ( 
.A(n_12605),
.Y(n_13587)
);

NAND2xp5_ASAP7_75t_L g13588 ( 
.A(n_12465),
.B(n_10751),
.Y(n_13588)
);

INVx1_ASAP7_75t_L g13589 ( 
.A(n_12682),
.Y(n_13589)
);

AND2x2_ASAP7_75t_L g13590 ( 
.A(n_12630),
.B(n_10756),
.Y(n_13590)
);

OR2x6_ASAP7_75t_L g13591 ( 
.A(n_12807),
.B(n_5222),
.Y(n_13591)
);

NOR2x1_ASAP7_75t_L g13592 ( 
.A(n_13121),
.B(n_12174),
.Y(n_13592)
);

BUFx3_ASAP7_75t_L g13593 ( 
.A(n_12881),
.Y(n_13593)
);

INVxp67_ASAP7_75t_L g13594 ( 
.A(n_12629),
.Y(n_13594)
);

INVx2_ASAP7_75t_L g13595 ( 
.A(n_12477),
.Y(n_13595)
);

INVx1_ASAP7_75t_L g13596 ( 
.A(n_12682),
.Y(n_13596)
);

NAND2xp5_ASAP7_75t_L g13597 ( 
.A(n_12638),
.B(n_10758),
.Y(n_13597)
);

AND2x2_ASAP7_75t_L g13598 ( 
.A(n_12636),
.B(n_10759),
.Y(n_13598)
);

OR2x2_ASAP7_75t_L g13599 ( 
.A(n_13209),
.B(n_12768),
.Y(n_13599)
);

AND2x2_ASAP7_75t_L g13600 ( 
.A(n_12670),
.B(n_10761),
.Y(n_13600)
);

NOR2xp33_ASAP7_75t_L g13601 ( 
.A(n_12475),
.B(n_5037),
.Y(n_13601)
);

INVx2_ASAP7_75t_L g13602 ( 
.A(n_12481),
.Y(n_13602)
);

HB1xp67_ASAP7_75t_L g13603 ( 
.A(n_12838),
.Y(n_13603)
);

AND2x4_ASAP7_75t_L g13604 ( 
.A(n_12743),
.B(n_12747),
.Y(n_13604)
);

INVxp67_ASAP7_75t_SL g13605 ( 
.A(n_12676),
.Y(n_13605)
);

NAND2xp5_ASAP7_75t_L g13606 ( 
.A(n_12639),
.B(n_10770),
.Y(n_13606)
);

NAND2x1_ASAP7_75t_L g13607 ( 
.A(n_13232),
.B(n_10771),
.Y(n_13607)
);

AOI22xp33_ASAP7_75t_L g13608 ( 
.A1(n_13309),
.A2(n_11860),
.B1(n_11939),
.B2(n_11931),
.Y(n_13608)
);

AND2x2_ASAP7_75t_L g13609 ( 
.A(n_12478),
.B(n_10774),
.Y(n_13609)
);

INVx1_ASAP7_75t_L g13610 ( 
.A(n_12683),
.Y(n_13610)
);

INVx1_ASAP7_75t_L g13611 ( 
.A(n_12683),
.Y(n_13611)
);

NAND2xp5_ASAP7_75t_SL g13612 ( 
.A(n_12503),
.B(n_12381),
.Y(n_13612)
);

INVx1_ASAP7_75t_L g13613 ( 
.A(n_12684),
.Y(n_13613)
);

INVx1_ASAP7_75t_L g13614 ( 
.A(n_12684),
.Y(n_13614)
);

INVx1_ASAP7_75t_L g13615 ( 
.A(n_12689),
.Y(n_13615)
);

INVx1_ASAP7_75t_L g13616 ( 
.A(n_12689),
.Y(n_13616)
);

NOR2xp33_ASAP7_75t_L g13617 ( 
.A(n_12890),
.B(n_5071),
.Y(n_13617)
);

AND2x2_ASAP7_75t_L g13618 ( 
.A(n_12621),
.B(n_10779),
.Y(n_13618)
);

AND2x2_ASAP7_75t_L g13619 ( 
.A(n_12901),
.B(n_10783),
.Y(n_13619)
);

AND2x4_ASAP7_75t_L g13620 ( 
.A(n_12510),
.B(n_10786),
.Y(n_13620)
);

INVx2_ASAP7_75t_L g13621 ( 
.A(n_12418),
.Y(n_13621)
);

CKINVDCx14_ASAP7_75t_R g13622 ( 
.A(n_12828),
.Y(n_13622)
);

INVx1_ASAP7_75t_L g13623 ( 
.A(n_12703),
.Y(n_13623)
);

NOR2xp33_ASAP7_75t_R g13624 ( 
.A(n_12674),
.B(n_5257),
.Y(n_13624)
);

INVx2_ASAP7_75t_L g13625 ( 
.A(n_12740),
.Y(n_13625)
);

NAND2xp5_ASAP7_75t_L g13626 ( 
.A(n_12641),
.B(n_10791),
.Y(n_13626)
);

OAI22xp5_ASAP7_75t_L g13627 ( 
.A1(n_13292),
.A2(n_12182),
.B1(n_12364),
.B2(n_12365),
.Y(n_13627)
);

INVxp67_ASAP7_75t_SL g13628 ( 
.A(n_13061),
.Y(n_13628)
);

INVx2_ASAP7_75t_L g13629 ( 
.A(n_12530),
.Y(n_13629)
);

INVx2_ASAP7_75t_L g13630 ( 
.A(n_12531),
.Y(n_13630)
);

AOI22xp33_ASAP7_75t_L g13631 ( 
.A1(n_12979),
.A2(n_12332),
.B1(n_12198),
.B2(n_12201),
.Y(n_13631)
);

AND2x2_ASAP7_75t_L g13632 ( 
.A(n_12540),
.B(n_10792),
.Y(n_13632)
);

INVx1_ASAP7_75t_L g13633 ( 
.A(n_12703),
.Y(n_13633)
);

INVx2_ASAP7_75t_L g13634 ( 
.A(n_12544),
.Y(n_13634)
);

HB1xp67_ASAP7_75t_L g13635 ( 
.A(n_12673),
.Y(n_13635)
);

NOR2x1_ASAP7_75t_SL g13636 ( 
.A(n_13059),
.B(n_12359),
.Y(n_13636)
);

NOR2xp67_ASAP7_75t_L g13637 ( 
.A(n_13009),
.B(n_12395),
.Y(n_13637)
);

AND2x4_ASAP7_75t_L g13638 ( 
.A(n_12696),
.B(n_10797),
.Y(n_13638)
);

INVx2_ASAP7_75t_L g13639 ( 
.A(n_12545),
.Y(n_13639)
);

OR2x2_ASAP7_75t_L g13640 ( 
.A(n_13308),
.B(n_10798),
.Y(n_13640)
);

BUFx3_ASAP7_75t_L g13641 ( 
.A(n_12755),
.Y(n_13641)
);

AND2x4_ASAP7_75t_L g13642 ( 
.A(n_12699),
.B(n_10799),
.Y(n_13642)
);

INVx2_ASAP7_75t_L g13643 ( 
.A(n_12555),
.Y(n_13643)
);

INVx2_ASAP7_75t_L g13644 ( 
.A(n_13008),
.Y(n_13644)
);

AND2x2_ASAP7_75t_L g13645 ( 
.A(n_12742),
.B(n_12591),
.Y(n_13645)
);

OR2x2_ASAP7_75t_L g13646 ( 
.A(n_13281),
.B(n_10800),
.Y(n_13646)
);

BUFx2_ASAP7_75t_L g13647 ( 
.A(n_13111),
.Y(n_13647)
);

INVx1_ASAP7_75t_L g13648 ( 
.A(n_12706),
.Y(n_13648)
);

INVx2_ASAP7_75t_L g13649 ( 
.A(n_13008),
.Y(n_13649)
);

NOR2xp67_ASAP7_75t_L g13650 ( 
.A(n_13009),
.B(n_12346),
.Y(n_13650)
);

AOI22xp33_ASAP7_75t_SL g13651 ( 
.A1(n_13259),
.A2(n_12357),
.B1(n_12377),
.B2(n_12370),
.Y(n_13651)
);

AND2x2_ASAP7_75t_L g13652 ( 
.A(n_12592),
.B(n_12598),
.Y(n_13652)
);

OR2x2_ASAP7_75t_L g13653 ( 
.A(n_12646),
.B(n_10809),
.Y(n_13653)
);

NOR2xp33_ASAP7_75t_L g13654 ( 
.A(n_12719),
.B(n_5071),
.Y(n_13654)
);

AND2x2_ASAP7_75t_L g13655 ( 
.A(n_12603),
.B(n_10815),
.Y(n_13655)
);

INVx1_ASAP7_75t_L g13656 ( 
.A(n_12706),
.Y(n_13656)
);

INVx1_ASAP7_75t_L g13657 ( 
.A(n_12716),
.Y(n_13657)
);

AND2x2_ASAP7_75t_L g13658 ( 
.A(n_12749),
.B(n_10817),
.Y(n_13658)
);

AND2x2_ASAP7_75t_L g13659 ( 
.A(n_12751),
.B(n_10818),
.Y(n_13659)
);

HB1xp67_ASAP7_75t_L g13660 ( 
.A(n_12924),
.Y(n_13660)
);

BUFx2_ASAP7_75t_L g13661 ( 
.A(n_13111),
.Y(n_13661)
);

INVx1_ASAP7_75t_L g13662 ( 
.A(n_12716),
.Y(n_13662)
);

AND2x2_ASAP7_75t_L g13663 ( 
.A(n_12762),
.B(n_10819),
.Y(n_13663)
);

HB1xp67_ASAP7_75t_L g13664 ( 
.A(n_12923),
.Y(n_13664)
);

OR2x2_ASAP7_75t_L g13665 ( 
.A(n_13313),
.B(n_10820),
.Y(n_13665)
);

AND2x4_ASAP7_75t_L g13666 ( 
.A(n_12702),
.B(n_12704),
.Y(n_13666)
);

INVx1_ASAP7_75t_L g13667 ( 
.A(n_12717),
.Y(n_13667)
);

INVx2_ASAP7_75t_L g13668 ( 
.A(n_13008),
.Y(n_13668)
);

INVx5_ASAP7_75t_L g13669 ( 
.A(n_12708),
.Y(n_13669)
);

INVx1_ASAP7_75t_L g13670 ( 
.A(n_12717),
.Y(n_13670)
);

AOI22xp33_ASAP7_75t_L g13671 ( 
.A1(n_13299),
.A2(n_12245),
.B1(n_12306),
.B2(n_12295),
.Y(n_13671)
);

INVx1_ASAP7_75t_L g13672 ( 
.A(n_12729),
.Y(n_13672)
);

INVx1_ASAP7_75t_L g13673 ( 
.A(n_12729),
.Y(n_13673)
);

INVx1_ASAP7_75t_L g13674 ( 
.A(n_12745),
.Y(n_13674)
);

HB1xp67_ASAP7_75t_L g13675 ( 
.A(n_12931),
.Y(n_13675)
);

AND2x2_ASAP7_75t_L g13676 ( 
.A(n_12767),
.B(n_10826),
.Y(n_13676)
);

AND2x2_ASAP7_75t_L g13677 ( 
.A(n_12772),
.B(n_10827),
.Y(n_13677)
);

NAND2xp5_ASAP7_75t_L g13678 ( 
.A(n_13230),
.B(n_13099),
.Y(n_13678)
);

INVx1_ASAP7_75t_L g13679 ( 
.A(n_12745),
.Y(n_13679)
);

INVx2_ASAP7_75t_L g13680 ( 
.A(n_13012),
.Y(n_13680)
);

INVx1_ASAP7_75t_L g13681 ( 
.A(n_12753),
.Y(n_13681)
);

INVx2_ASAP7_75t_L g13682 ( 
.A(n_13012),
.Y(n_13682)
);

INVx1_ASAP7_75t_L g13683 ( 
.A(n_12753),
.Y(n_13683)
);

INVx2_ASAP7_75t_L g13684 ( 
.A(n_13012),
.Y(n_13684)
);

HB1xp67_ASAP7_75t_L g13685 ( 
.A(n_12951),
.Y(n_13685)
);

INVx1_ASAP7_75t_L g13686 ( 
.A(n_12754),
.Y(n_13686)
);

INVx2_ASAP7_75t_L g13687 ( 
.A(n_12720),
.Y(n_13687)
);

AND2x2_ASAP7_75t_L g13688 ( 
.A(n_12773),
.B(n_10830),
.Y(n_13688)
);

NAND2xp5_ASAP7_75t_L g13689 ( 
.A(n_12661),
.B(n_10832),
.Y(n_13689)
);

INVx2_ASAP7_75t_L g13690 ( 
.A(n_12644),
.Y(n_13690)
);

AND2x2_ASAP7_75t_L g13691 ( 
.A(n_12776),
.B(n_10845),
.Y(n_13691)
);

INVx1_ASAP7_75t_L g13692 ( 
.A(n_12754),
.Y(n_13692)
);

INVx1_ASAP7_75t_L g13693 ( 
.A(n_12760),
.Y(n_13693)
);

INVx1_ASAP7_75t_L g13694 ( 
.A(n_12760),
.Y(n_13694)
);

INVxp67_ASAP7_75t_SL g13695 ( 
.A(n_13237),
.Y(n_13695)
);

INVx1_ASAP7_75t_L g13696 ( 
.A(n_12763),
.Y(n_13696)
);

AND2x2_ASAP7_75t_L g13697 ( 
.A(n_12658),
.B(n_10849),
.Y(n_13697)
);

AND2x4_ASAP7_75t_L g13698 ( 
.A(n_12539),
.B(n_10851),
.Y(n_13698)
);

INVx2_ASAP7_75t_L g13699 ( 
.A(n_12686),
.Y(n_13699)
);

AND2x2_ASAP7_75t_L g13700 ( 
.A(n_12690),
.B(n_12709),
.Y(n_13700)
);

AOI22xp33_ASAP7_75t_L g13701 ( 
.A1(n_13300),
.A2(n_12257),
.B1(n_12273),
.B2(n_12260),
.Y(n_13701)
);

OR2x2_ASAP7_75t_L g13702 ( 
.A(n_12770),
.B(n_10854),
.Y(n_13702)
);

INVx4_ASAP7_75t_L g13703 ( 
.A(n_12724),
.Y(n_13703)
);

AND2x2_ASAP7_75t_L g13704 ( 
.A(n_12714),
.B(n_10856),
.Y(n_13704)
);

INVx1_ASAP7_75t_SL g13705 ( 
.A(n_13002),
.Y(n_13705)
);

HB1xp67_ASAP7_75t_L g13706 ( 
.A(n_13023),
.Y(n_13706)
);

AOI22xp33_ASAP7_75t_L g13707 ( 
.A1(n_13226),
.A2(n_12117),
.B1(n_12042),
.B2(n_12046),
.Y(n_13707)
);

NAND2x1p5_ASAP7_75t_SL g13708 ( 
.A(n_13214),
.B(n_7720),
.Y(n_13708)
);

INVx2_ASAP7_75t_L g13709 ( 
.A(n_12713),
.Y(n_13709)
);

AND2x2_ASAP7_75t_L g13710 ( 
.A(n_12705),
.B(n_10869),
.Y(n_13710)
);

NOR2xp33_ASAP7_75t_L g13711 ( 
.A(n_13175),
.B(n_5257),
.Y(n_13711)
);

INVx2_ASAP7_75t_L g13712 ( 
.A(n_12713),
.Y(n_13712)
);

INVx1_ASAP7_75t_L g13713 ( 
.A(n_12763),
.Y(n_13713)
);

AND2x2_ASAP7_75t_L g13714 ( 
.A(n_12832),
.B(n_10877),
.Y(n_13714)
);

NAND2xp5_ASAP7_75t_L g13715 ( 
.A(n_12662),
.B(n_10879),
.Y(n_13715)
);

OR2x2_ASAP7_75t_L g13716 ( 
.A(n_12593),
.B(n_10883),
.Y(n_13716)
);

AOI22xp33_ASAP7_75t_SL g13717 ( 
.A1(n_13322),
.A2(n_12340),
.B1(n_7730),
.B2(n_7968),
.Y(n_13717)
);

NAND2xp5_ASAP7_75t_L g13718 ( 
.A(n_12664),
.B(n_10886),
.Y(n_13718)
);

OR2x2_ASAP7_75t_L g13719 ( 
.A(n_12803),
.B(n_10887),
.Y(n_13719)
);

NAND2xp5_ASAP7_75t_L g13720 ( 
.A(n_12665),
.B(n_12666),
.Y(n_13720)
);

AND2x2_ASAP7_75t_L g13721 ( 
.A(n_13157),
.B(n_7610),
.Y(n_13721)
);

OR2x2_ASAP7_75t_L g13722 ( 
.A(n_13212),
.B(n_8470),
.Y(n_13722)
);

AND2x2_ASAP7_75t_L g13723 ( 
.A(n_12848),
.B(n_7610),
.Y(n_13723)
);

INVx2_ASAP7_75t_L g13724 ( 
.A(n_13016),
.Y(n_13724)
);

INVx2_ASAP7_75t_L g13725 ( 
.A(n_13016),
.Y(n_13725)
);

AND2x2_ASAP7_75t_L g13726 ( 
.A(n_13210),
.B(n_7610),
.Y(n_13726)
);

AND2x2_ASAP7_75t_L g13727 ( 
.A(n_12748),
.B(n_7610),
.Y(n_13727)
);

INVx1_ASAP7_75t_L g13728 ( 
.A(n_12769),
.Y(n_13728)
);

INVx2_ASAP7_75t_L g13729 ( 
.A(n_12678),
.Y(n_13729)
);

HB1xp67_ASAP7_75t_L g13730 ( 
.A(n_12679),
.Y(n_13730)
);

INVx2_ASAP7_75t_L g13731 ( 
.A(n_12605),
.Y(n_13731)
);

INVx2_ASAP7_75t_L g13732 ( 
.A(n_12790),
.Y(n_13732)
);

INVx2_ASAP7_75t_L g13733 ( 
.A(n_12792),
.Y(n_13733)
);

INVx1_ASAP7_75t_L g13734 ( 
.A(n_12769),
.Y(n_13734)
);

NAND2xp5_ASAP7_75t_L g13735 ( 
.A(n_13311),
.B(n_11951),
.Y(n_13735)
);

INVx1_ASAP7_75t_L g13736 ( 
.A(n_12771),
.Y(n_13736)
);

INVx1_ASAP7_75t_SL g13737 ( 
.A(n_13077),
.Y(n_13737)
);

INVx2_ASAP7_75t_L g13738 ( 
.A(n_12805),
.Y(n_13738)
);

NAND2xp5_ASAP7_75t_L g13739 ( 
.A(n_13288),
.B(n_11968),
.Y(n_13739)
);

OR2x2_ASAP7_75t_L g13740 ( 
.A(n_13266),
.B(n_8483),
.Y(n_13740)
);

INVx3_ASAP7_75t_L g13741 ( 
.A(n_12804),
.Y(n_13741)
);

INVx1_ASAP7_75t_L g13742 ( 
.A(n_12771),
.Y(n_13742)
);

AND2x2_ASAP7_75t_L g13743 ( 
.A(n_12701),
.B(n_7610),
.Y(n_13743)
);

INVx1_ASAP7_75t_L g13744 ( 
.A(n_12774),
.Y(n_13744)
);

AND2x2_ASAP7_75t_L g13745 ( 
.A(n_12691),
.B(n_7622),
.Y(n_13745)
);

AND2x2_ASAP7_75t_L g13746 ( 
.A(n_13223),
.B(n_7622),
.Y(n_13746)
);

AND2x2_ASAP7_75t_L g13747 ( 
.A(n_12806),
.B(n_7622),
.Y(n_13747)
);

AND2x2_ASAP7_75t_L g13748 ( 
.A(n_12741),
.B(n_13095),
.Y(n_13748)
);

AND2x4_ASAP7_75t_L g13749 ( 
.A(n_12549),
.B(n_12551),
.Y(n_13749)
);

INVx2_ASAP7_75t_L g13750 ( 
.A(n_12758),
.Y(n_13750)
);

INVx4_ASAP7_75t_L g13751 ( 
.A(n_12728),
.Y(n_13751)
);

AND2x2_ASAP7_75t_L g13752 ( 
.A(n_13108),
.B(n_7622),
.Y(n_13752)
);

OR2x2_ASAP7_75t_L g13753 ( 
.A(n_13003),
.B(n_8483),
.Y(n_13753)
);

HB1xp67_ASAP7_75t_L g13754 ( 
.A(n_13013),
.Y(n_13754)
);

AND2x2_ASAP7_75t_L g13755 ( 
.A(n_12730),
.B(n_7622),
.Y(n_13755)
);

NAND2xp5_ASAP7_75t_L g13756 ( 
.A(n_13168),
.B(n_11971),
.Y(n_13756)
);

INVx1_ASAP7_75t_L g13757 ( 
.A(n_12774),
.Y(n_13757)
);

INVx1_ASAP7_75t_L g13758 ( 
.A(n_12781),
.Y(n_13758)
);

INVx2_ASAP7_75t_L g13759 ( 
.A(n_12574),
.Y(n_13759)
);

BUFx2_ASAP7_75t_L g13760 ( 
.A(n_12517),
.Y(n_13760)
);

INVx1_ASAP7_75t_L g13761 ( 
.A(n_12781),
.Y(n_13761)
);

OR2x2_ASAP7_75t_L g13762 ( 
.A(n_12455),
.B(n_8491),
.Y(n_13762)
);

NAND2xp5_ASAP7_75t_L g13763 ( 
.A(n_13080),
.B(n_12003),
.Y(n_13763)
);

INVx2_ASAP7_75t_SL g13764 ( 
.A(n_12971),
.Y(n_13764)
);

INVx1_ASAP7_75t_L g13765 ( 
.A(n_12782),
.Y(n_13765)
);

NAND2x1p5_ASAP7_75t_L g13766 ( 
.A(n_12835),
.B(n_12707),
.Y(n_13766)
);

OR2x2_ASAP7_75t_L g13767 ( 
.A(n_13239),
.B(n_8491),
.Y(n_13767)
);

AND2x2_ASAP7_75t_SL g13768 ( 
.A(n_13233),
.B(n_8291),
.Y(n_13768)
);

AND2x2_ASAP7_75t_L g13769 ( 
.A(n_12731),
.B(n_7632),
.Y(n_13769)
);

AND2x2_ASAP7_75t_L g13770 ( 
.A(n_12604),
.B(n_12608),
.Y(n_13770)
);

AND2x2_ASAP7_75t_L g13771 ( 
.A(n_12656),
.B(n_7632),
.Y(n_13771)
);

NOR2xp67_ASAP7_75t_L g13772 ( 
.A(n_13139),
.B(n_9096),
.Y(n_13772)
);

NOR2xp67_ASAP7_75t_L g13773 ( 
.A(n_13179),
.B(n_9100),
.Y(n_13773)
);

NAND2xp5_ASAP7_75t_L g13774 ( 
.A(n_13318),
.B(n_12026),
.Y(n_13774)
);

NAND2xp5_ASAP7_75t_L g13775 ( 
.A(n_13156),
.B(n_12033),
.Y(n_13775)
);

INVx2_ASAP7_75t_L g13776 ( 
.A(n_12575),
.Y(n_13776)
);

INVx1_ASAP7_75t_L g13777 ( 
.A(n_12782),
.Y(n_13777)
);

NAND2xp5_ASAP7_75t_L g13778 ( 
.A(n_13156),
.B(n_13305),
.Y(n_13778)
);

HB1xp67_ASAP7_75t_L g13779 ( 
.A(n_12463),
.Y(n_13779)
);

INVx1_ASAP7_75t_L g13780 ( 
.A(n_12785),
.Y(n_13780)
);

NOR2x1_ASAP7_75t_L g13781 ( 
.A(n_13146),
.B(n_12335),
.Y(n_13781)
);

NAND4xp25_ASAP7_75t_L g13782 ( 
.A(n_12688),
.B(n_11999),
.C(n_12366),
.D(n_12409),
.Y(n_13782)
);

INVx2_ASAP7_75t_L g13783 ( 
.A(n_12585),
.Y(n_13783)
);

HB1xp67_ASAP7_75t_L g13784 ( 
.A(n_12470),
.Y(n_13784)
);

INVx1_ASAP7_75t_L g13785 ( 
.A(n_12785),
.Y(n_13785)
);

INVx1_ASAP7_75t_L g13786 ( 
.A(n_12859),
.Y(n_13786)
);

AND2x2_ASAP7_75t_L g13787 ( 
.A(n_12657),
.B(n_12836),
.Y(n_13787)
);

HB1xp67_ASAP7_75t_L g13788 ( 
.A(n_12595),
.Y(n_13788)
);

INVx1_ASAP7_75t_L g13789 ( 
.A(n_12859),
.Y(n_13789)
);

INVx4_ASAP7_75t_L g13790 ( 
.A(n_12775),
.Y(n_13790)
);

AND2x2_ASAP7_75t_L g13791 ( 
.A(n_12831),
.B(n_7632),
.Y(n_13791)
);

INVx1_ASAP7_75t_L g13792 ( 
.A(n_12861),
.Y(n_13792)
);

HB1xp67_ASAP7_75t_L g13793 ( 
.A(n_12597),
.Y(n_13793)
);

NOR2xp33_ASAP7_75t_L g13794 ( 
.A(n_12887),
.B(n_5285),
.Y(n_13794)
);

NAND2xp5_ASAP7_75t_L g13795 ( 
.A(n_13192),
.B(n_12037),
.Y(n_13795)
);

AOI22xp33_ASAP7_75t_L g13796 ( 
.A1(n_13140),
.A2(n_12265),
.B1(n_12290),
.B2(n_12284),
.Y(n_13796)
);

INVx3_ASAP7_75t_L g13797 ( 
.A(n_12804),
.Y(n_13797)
);

INVx2_ASAP7_75t_L g13798 ( 
.A(n_12600),
.Y(n_13798)
);

INVx1_ASAP7_75t_L g13799 ( 
.A(n_12861),
.Y(n_13799)
);

AOI22xp5_ASAP7_75t_L g13800 ( 
.A1(n_13283),
.A2(n_12299),
.B1(n_12368),
.B2(n_12318),
.Y(n_13800)
);

INVx2_ASAP7_75t_L g13801 ( 
.A(n_12623),
.Y(n_13801)
);

INVx1_ASAP7_75t_L g13802 ( 
.A(n_12948),
.Y(n_13802)
);

AND2x2_ASAP7_75t_L g13803 ( 
.A(n_12417),
.B(n_7632),
.Y(n_13803)
);

NAND2xp5_ASAP7_75t_L g13804 ( 
.A(n_13192),
.B(n_10259),
.Y(n_13804)
);

OR2x2_ASAP7_75t_L g13805 ( 
.A(n_12739),
.B(n_8499),
.Y(n_13805)
);

INVx1_ASAP7_75t_L g13806 ( 
.A(n_12948),
.Y(n_13806)
);

AND2x2_ASAP7_75t_L g13807 ( 
.A(n_12675),
.B(n_7632),
.Y(n_13807)
);

INVx2_ASAP7_75t_L g13808 ( 
.A(n_12632),
.Y(n_13808)
);

INVx1_ASAP7_75t_L g13809 ( 
.A(n_12614),
.Y(n_13809)
);

NAND2xp5_ASAP7_75t_L g13810 ( 
.A(n_12422),
.B(n_10260),
.Y(n_13810)
);

INVxp67_ASAP7_75t_SL g13811 ( 
.A(n_12904),
.Y(n_13811)
);

INVx1_ASAP7_75t_L g13812 ( 
.A(n_12659),
.Y(n_13812)
);

BUFx5_ASAP7_75t_L g13813 ( 
.A(n_13018),
.Y(n_13813)
);

INVx2_ASAP7_75t_L g13814 ( 
.A(n_12868),
.Y(n_13814)
);

INVx1_ASAP7_75t_L g13815 ( 
.A(n_12508),
.Y(n_13815)
);

INVx1_ASAP7_75t_L g13816 ( 
.A(n_12513),
.Y(n_13816)
);

OR2x2_ASAP7_75t_L g13817 ( 
.A(n_12750),
.B(n_8499),
.Y(n_13817)
);

AND2x2_ASAP7_75t_L g13818 ( 
.A(n_12677),
.B(n_7674),
.Y(n_13818)
);

OR2x2_ASAP7_75t_L g13819 ( 
.A(n_12761),
.B(n_8125),
.Y(n_13819)
);

AND2x2_ASAP7_75t_L g13820 ( 
.A(n_12680),
.B(n_7674),
.Y(n_13820)
);

AND2x2_ASAP7_75t_L g13821 ( 
.A(n_12685),
.B(n_12694),
.Y(n_13821)
);

OR2x2_ASAP7_75t_L g13822 ( 
.A(n_12787),
.B(n_8125),
.Y(n_13822)
);

AND2x2_ASAP7_75t_L g13823 ( 
.A(n_12695),
.B(n_7674),
.Y(n_13823)
);

AND2x2_ASAP7_75t_L g13824 ( 
.A(n_12966),
.B(n_7674),
.Y(n_13824)
);

BUFx2_ASAP7_75t_L g13825 ( 
.A(n_12514),
.Y(n_13825)
);

INVx2_ASAP7_75t_L g13826 ( 
.A(n_12752),
.Y(n_13826)
);

INVxp67_ASAP7_75t_SL g13827 ( 
.A(n_12556),
.Y(n_13827)
);

INVx3_ASAP7_75t_L g13828 ( 
.A(n_12609),
.Y(n_13828)
);

INVx2_ASAP7_75t_L g13829 ( 
.A(n_12552),
.Y(n_13829)
);

INVxp67_ASAP7_75t_SL g13830 ( 
.A(n_12998),
.Y(n_13830)
);

AND2x2_ASAP7_75t_L g13831 ( 
.A(n_13097),
.B(n_7674),
.Y(n_13831)
);

BUFx2_ASAP7_75t_L g13832 ( 
.A(n_13059),
.Y(n_13832)
);

INVx2_ASAP7_75t_L g13833 ( 
.A(n_12559),
.Y(n_13833)
);

AND2x4_ASAP7_75t_L g13834 ( 
.A(n_12562),
.B(n_9100),
.Y(n_13834)
);

INVx1_ASAP7_75t_L g13835 ( 
.A(n_12515),
.Y(n_13835)
);

AND2x2_ASAP7_75t_L g13836 ( 
.A(n_12725),
.B(n_7708),
.Y(n_13836)
);

INVx3_ASAP7_75t_L g13837 ( 
.A(n_13010),
.Y(n_13837)
);

AND2x2_ASAP7_75t_L g13838 ( 
.A(n_12727),
.B(n_7708),
.Y(n_13838)
);

INVx1_ASAP7_75t_L g13839 ( 
.A(n_12518),
.Y(n_13839)
);

AND2x2_ASAP7_75t_L g13840 ( 
.A(n_12884),
.B(n_7708),
.Y(n_13840)
);

INVx2_ASAP7_75t_L g13841 ( 
.A(n_12778),
.Y(n_13841)
);

AND2x2_ASAP7_75t_L g13842 ( 
.A(n_13243),
.B(n_7708),
.Y(n_13842)
);

INVx3_ASAP7_75t_L g13843 ( 
.A(n_13010),
.Y(n_13843)
);

AND2x2_ASAP7_75t_L g13844 ( 
.A(n_12867),
.B(n_7708),
.Y(n_13844)
);

AND2x2_ASAP7_75t_L g13845 ( 
.A(n_12872),
.B(n_7784),
.Y(n_13845)
);

INVx1_ASAP7_75t_L g13846 ( 
.A(n_12520),
.Y(n_13846)
);

AND2x2_ASAP7_75t_L g13847 ( 
.A(n_12879),
.B(n_7784),
.Y(n_13847)
);

INVx1_ASAP7_75t_L g13848 ( 
.A(n_12524),
.Y(n_13848)
);

NAND2xp5_ASAP7_75t_L g13849 ( 
.A(n_13211),
.B(n_10262),
.Y(n_13849)
);

OR2x2_ASAP7_75t_SL g13850 ( 
.A(n_13172),
.B(n_10277),
.Y(n_13850)
);

AND2x2_ASAP7_75t_L g13851 ( 
.A(n_13067),
.B(n_7784),
.Y(n_13851)
);

NAND2xp5_ASAP7_75t_L g13852 ( 
.A(n_13142),
.B(n_10262),
.Y(n_13852)
);

HB1xp67_ASAP7_75t_L g13853 ( 
.A(n_12992),
.Y(n_13853)
);

BUFx2_ASAP7_75t_L g13854 ( 
.A(n_13059),
.Y(n_13854)
);

INVx2_ASAP7_75t_L g13855 ( 
.A(n_12569),
.Y(n_13855)
);

AND2x2_ASAP7_75t_L g13856 ( 
.A(n_13125),
.B(n_13100),
.Y(n_13856)
);

AND2x4_ASAP7_75t_L g13857 ( 
.A(n_12486),
.B(n_9100),
.Y(n_13857)
);

NAND2xp5_ASAP7_75t_L g13858 ( 
.A(n_13171),
.B(n_10263),
.Y(n_13858)
);

AND2x2_ASAP7_75t_L g13859 ( 
.A(n_13115),
.B(n_12930),
.Y(n_13859)
);

INVx1_ASAP7_75t_L g13860 ( 
.A(n_12532),
.Y(n_13860)
);

OR2x2_ASAP7_75t_L g13861 ( 
.A(n_13302),
.B(n_8135),
.Y(n_13861)
);

INVx2_ASAP7_75t_L g13862 ( 
.A(n_12570),
.Y(n_13862)
);

INVx1_ASAP7_75t_L g13863 ( 
.A(n_12533),
.Y(n_13863)
);

OR2x2_ASAP7_75t_L g13864 ( 
.A(n_12734),
.B(n_8135),
.Y(n_13864)
);

AND2x4_ASAP7_75t_SL g13865 ( 
.A(n_12992),
.B(n_8547),
.Y(n_13865)
);

NOR2x1_ASAP7_75t_L g13866 ( 
.A(n_13146),
.B(n_9100),
.Y(n_13866)
);

AND2x2_ASAP7_75t_L g13867 ( 
.A(n_12958),
.B(n_7784),
.Y(n_13867)
);

INVx1_ASAP7_75t_L g13868 ( 
.A(n_12536),
.Y(n_13868)
);

AND2x4_ASAP7_75t_L g13869 ( 
.A(n_12493),
.B(n_9124),
.Y(n_13869)
);

INVx2_ASAP7_75t_L g13870 ( 
.A(n_12571),
.Y(n_13870)
);

INVx1_ASAP7_75t_L g13871 ( 
.A(n_12538),
.Y(n_13871)
);

OR2x2_ASAP7_75t_L g13872 ( 
.A(n_13307),
.B(n_8146),
.Y(n_13872)
);

AND2x2_ASAP7_75t_L g13873 ( 
.A(n_12996),
.B(n_7784),
.Y(n_13873)
);

AND2x4_ASAP7_75t_L g13874 ( 
.A(n_12504),
.B(n_9124),
.Y(n_13874)
);

NAND2xp5_ASAP7_75t_L g13875 ( 
.A(n_13276),
.B(n_10263),
.Y(n_13875)
);

AND2x2_ASAP7_75t_L g13876 ( 
.A(n_13048),
.B(n_8729),
.Y(n_13876)
);

NAND2xp5_ASAP7_75t_L g13877 ( 
.A(n_13284),
.B(n_10265),
.Y(n_13877)
);

AND2x2_ASAP7_75t_L g13878 ( 
.A(n_13241),
.B(n_10265),
.Y(n_13878)
);

AND2x2_ASAP7_75t_L g13879 ( 
.A(n_13163),
.B(n_13141),
.Y(n_13879)
);

INVx1_ASAP7_75t_L g13880 ( 
.A(n_12541),
.Y(n_13880)
);

INVx2_ASAP7_75t_L g13881 ( 
.A(n_12572),
.Y(n_13881)
);

OR2x2_ASAP7_75t_L g13882 ( 
.A(n_13215),
.B(n_8146),
.Y(n_13882)
);

NOR2x1_ASAP7_75t_L g13883 ( 
.A(n_13145),
.B(n_9124),
.Y(n_13883)
);

INVx1_ASAP7_75t_L g13884 ( 
.A(n_12548),
.Y(n_13884)
);

INVx2_ASAP7_75t_L g13885 ( 
.A(n_12581),
.Y(n_13885)
);

HB1xp67_ASAP7_75t_L g13886 ( 
.A(n_12992),
.Y(n_13886)
);

AND2x2_ASAP7_75t_L g13887 ( 
.A(n_13141),
.B(n_10269),
.Y(n_13887)
);

AND2x2_ASAP7_75t_L g13888 ( 
.A(n_12711),
.B(n_12660),
.Y(n_13888)
);

AND2x2_ASAP7_75t_L g13889 ( 
.A(n_13114),
.B(n_10269),
.Y(n_13889)
);

NAND2xp5_ASAP7_75t_L g13890 ( 
.A(n_12972),
.B(n_10270),
.Y(n_13890)
);

INVx1_ASAP7_75t_L g13891 ( 
.A(n_12554),
.Y(n_13891)
);

INVx1_ASAP7_75t_SL g13892 ( 
.A(n_12780),
.Y(n_13892)
);

INVx1_ASAP7_75t_L g13893 ( 
.A(n_12573),
.Y(n_13893)
);

OR2x2_ASAP7_75t_L g13894 ( 
.A(n_12783),
.B(n_8336),
.Y(n_13894)
);

NAND2xp5_ASAP7_75t_L g13895 ( 
.A(n_12973),
.B(n_10270),
.Y(n_13895)
);

INVx1_ASAP7_75t_L g13896 ( 
.A(n_12577),
.Y(n_13896)
);

NOR2xp33_ASAP7_75t_L g13897 ( 
.A(n_13159),
.B(n_5285),
.Y(n_13897)
);

OR2x2_ASAP7_75t_L g13898 ( 
.A(n_13057),
.B(n_8336),
.Y(n_13898)
);

AND2x2_ASAP7_75t_L g13899 ( 
.A(n_13207),
.B(n_12586),
.Y(n_13899)
);

HB1xp67_ASAP7_75t_L g13900 ( 
.A(n_12999),
.Y(n_13900)
);

INVx1_ASAP7_75t_L g13901 ( 
.A(n_12579),
.Y(n_13901)
);

INVx1_ASAP7_75t_L g13902 ( 
.A(n_12582),
.Y(n_13902)
);

HB1xp67_ASAP7_75t_L g13903 ( 
.A(n_12999),
.Y(n_13903)
);

INVxp67_ASAP7_75t_SL g13904 ( 
.A(n_12965),
.Y(n_13904)
);

AOI22xp33_ASAP7_75t_L g13905 ( 
.A1(n_13213),
.A2(n_8225),
.B1(n_8386),
.B2(n_7800),
.Y(n_13905)
);

AND2x2_ASAP7_75t_L g13906 ( 
.A(n_13207),
.B(n_10274),
.Y(n_13906)
);

OAI222xp33_ASAP7_75t_L g13907 ( 
.A1(n_13289),
.A2(n_12074),
.B1(n_11820),
.B2(n_9153),
.C1(n_9128),
.C2(n_9154),
.Y(n_13907)
);

NAND2xp5_ASAP7_75t_L g13908 ( 
.A(n_12974),
.B(n_10274),
.Y(n_13908)
);

OR2x2_ASAP7_75t_L g13909 ( 
.A(n_13035),
.B(n_8375),
.Y(n_13909)
);

AND2x2_ASAP7_75t_L g13910 ( 
.A(n_12589),
.B(n_10287),
.Y(n_13910)
);

AND2x2_ASAP7_75t_L g13911 ( 
.A(n_13158),
.B(n_10287),
.Y(n_13911)
);

INVx1_ASAP7_75t_L g13912 ( 
.A(n_12587),
.Y(n_13912)
);

HB1xp67_ASAP7_75t_L g13913 ( 
.A(n_12999),
.Y(n_13913)
);

INVx1_ASAP7_75t_L g13914 ( 
.A(n_12590),
.Y(n_13914)
);

AND2x2_ASAP7_75t_L g13915 ( 
.A(n_13158),
.B(n_13161),
.Y(n_13915)
);

INVx1_ASAP7_75t_L g13916 ( 
.A(n_12628),
.Y(n_13916)
);

INVx1_ASAP7_75t_L g13917 ( 
.A(n_12631),
.Y(n_13917)
);

NAND2xp5_ASAP7_75t_L g13918 ( 
.A(n_12977),
.B(n_9822),
.Y(n_13918)
);

AND2x2_ASAP7_75t_L g13919 ( 
.A(n_13161),
.B(n_9124),
.Y(n_13919)
);

INVx1_ASAP7_75t_L g13920 ( 
.A(n_12633),
.Y(n_13920)
);

INVx1_ASAP7_75t_L g13921 ( 
.A(n_12643),
.Y(n_13921)
);

INVx2_ASAP7_75t_L g13922 ( 
.A(n_12642),
.Y(n_13922)
);

INVx1_ASAP7_75t_L g13923 ( 
.A(n_12648),
.Y(n_13923)
);

BUFx3_ASAP7_75t_L g13924 ( 
.A(n_12802),
.Y(n_13924)
);

AND2x4_ASAP7_75t_L g13925 ( 
.A(n_12837),
.B(n_9128),
.Y(n_13925)
);

INVx1_ASAP7_75t_L g13926 ( 
.A(n_12649),
.Y(n_13926)
);

INVx5_ASAP7_75t_L g13927 ( 
.A(n_13167),
.Y(n_13927)
);

INVx3_ASAP7_75t_L g13928 ( 
.A(n_13024),
.Y(n_13928)
);

AND2x4_ASAP7_75t_L g13929 ( 
.A(n_12840),
.B(n_9128),
.Y(n_13929)
);

BUFx6f_ASAP7_75t_L g13930 ( 
.A(n_12813),
.Y(n_13930)
);

OAI22xp5_ASAP7_75t_L g13931 ( 
.A1(n_12726),
.A2(n_12371),
.B1(n_7798),
.B2(n_7811),
.Y(n_13931)
);

INVx1_ASAP7_75t_L g13932 ( 
.A(n_12651),
.Y(n_13932)
);

AOI22xp33_ASAP7_75t_L g13933 ( 
.A1(n_13213),
.A2(n_8225),
.B1(n_8386),
.B2(n_7800),
.Y(n_13933)
);

NAND2xp5_ASAP7_75t_L g13934 ( 
.A(n_12978),
.B(n_9822),
.Y(n_13934)
);

INVx1_ASAP7_75t_L g13935 ( 
.A(n_12715),
.Y(n_13935)
);

INVx2_ASAP7_75t_L g13936 ( 
.A(n_12653),
.Y(n_13936)
);

INVx1_ASAP7_75t_L g13937 ( 
.A(n_12788),
.Y(n_13937)
);

AND2x2_ASAP7_75t_L g13938 ( 
.A(n_12856),
.B(n_9128),
.Y(n_13938)
);

INVx1_ASAP7_75t_L g13939 ( 
.A(n_12789),
.Y(n_13939)
);

HB1xp67_ASAP7_75t_L g13940 ( 
.A(n_12793),
.Y(n_13940)
);

INVx1_ASAP7_75t_L g13941 ( 
.A(n_12794),
.Y(n_13941)
);

OR2x2_ASAP7_75t_L g13942 ( 
.A(n_13035),
.B(n_8375),
.Y(n_13942)
);

INVx2_ASAP7_75t_L g13943 ( 
.A(n_12850),
.Y(n_13943)
);

NAND2xp5_ASAP7_75t_L g13944 ( 
.A(n_12983),
.B(n_9825),
.Y(n_13944)
);

BUFx2_ASAP7_75t_L g13945 ( 
.A(n_13148),
.Y(n_13945)
);

AND2x2_ASAP7_75t_L g13946 ( 
.A(n_12898),
.B(n_9139),
.Y(n_13946)
);

BUFx3_ASAP7_75t_L g13947 ( 
.A(n_12815),
.Y(n_13947)
);

BUFx3_ASAP7_75t_L g13948 ( 
.A(n_12821),
.Y(n_13948)
);

INVx1_ASAP7_75t_L g13949 ( 
.A(n_12796),
.Y(n_13949)
);

NAND2xp5_ASAP7_75t_L g13950 ( 
.A(n_12822),
.B(n_9825),
.Y(n_13950)
);

OR2x2_ASAP7_75t_L g13951 ( 
.A(n_12721),
.B(n_8377),
.Y(n_13951)
);

AND2x2_ASAP7_75t_L g13952 ( 
.A(n_13279),
.B(n_9139),
.Y(n_13952)
);

NAND2xp5_ASAP7_75t_L g13953 ( 
.A(n_12825),
.B(n_9833),
.Y(n_13953)
);

INVx1_ASAP7_75t_L g13954 ( 
.A(n_12797),
.Y(n_13954)
);

INVx2_ASAP7_75t_L g13955 ( 
.A(n_12864),
.Y(n_13955)
);

INVx1_ASAP7_75t_L g13956 ( 
.A(n_12800),
.Y(n_13956)
);

INVx1_ASAP7_75t_L g13957 ( 
.A(n_12809),
.Y(n_13957)
);

NAND2xp5_ASAP7_75t_L g13958 ( 
.A(n_12833),
.B(n_9833),
.Y(n_13958)
);

AND2x2_ASAP7_75t_L g13959 ( 
.A(n_13164),
.B(n_13166),
.Y(n_13959)
);

INVx1_ASAP7_75t_L g13960 ( 
.A(n_12818),
.Y(n_13960)
);

NAND2xp5_ASAP7_75t_L g13961 ( 
.A(n_13283),
.B(n_9842),
.Y(n_13961)
);

OR2x2_ASAP7_75t_L g13962 ( 
.A(n_13089),
.B(n_8377),
.Y(n_13962)
);

INVx1_ASAP7_75t_L g13963 ( 
.A(n_12820),
.Y(n_13963)
);

INVx1_ASAP7_75t_L g13964 ( 
.A(n_12823),
.Y(n_13964)
);

OR2x2_ASAP7_75t_L g13965 ( 
.A(n_13011),
.B(n_8380),
.Y(n_13965)
);

AND2x4_ASAP7_75t_L g13966 ( 
.A(n_12842),
.B(n_9139),
.Y(n_13966)
);

AND2x2_ASAP7_75t_L g13967 ( 
.A(n_13164),
.B(n_9139),
.Y(n_13967)
);

INVx2_ASAP7_75t_L g13968 ( 
.A(n_12854),
.Y(n_13968)
);

INVx2_ASAP7_75t_L g13969 ( 
.A(n_12854),
.Y(n_13969)
);

INVx2_ASAP7_75t_L g13970 ( 
.A(n_12870),
.Y(n_13970)
);

INVx2_ASAP7_75t_L g13971 ( 
.A(n_12870),
.Y(n_13971)
);

NAND2xp5_ASAP7_75t_L g13972 ( 
.A(n_13222),
.B(n_9842),
.Y(n_13972)
);

INVx2_ASAP7_75t_L g13973 ( 
.A(n_12849),
.Y(n_13973)
);

AND2x4_ASAP7_75t_L g13974 ( 
.A(n_12808),
.B(n_9153),
.Y(n_13974)
);

HB1xp67_ASAP7_75t_L g13975 ( 
.A(n_13148),
.Y(n_13975)
);

AND2x2_ASAP7_75t_L g13976 ( 
.A(n_13166),
.B(n_9153),
.Y(n_13976)
);

BUFx2_ASAP7_75t_L g13977 ( 
.A(n_13148),
.Y(n_13977)
);

AND2x4_ASAP7_75t_L g13978 ( 
.A(n_12811),
.B(n_9153),
.Y(n_13978)
);

INVx1_ASAP7_75t_L g13979 ( 
.A(n_12826),
.Y(n_13979)
);

NOR2xp33_ASAP7_75t_L g13980 ( 
.A(n_12871),
.B(n_5301),
.Y(n_13980)
);

AND2x4_ASAP7_75t_L g13981 ( 
.A(n_12812),
.B(n_9154),
.Y(n_13981)
);

OAI22xp5_ASAP7_75t_L g13982 ( 
.A1(n_13253),
.A2(n_7798),
.B1(n_7811),
.B2(n_7769),
.Y(n_13982)
);

INVx1_ASAP7_75t_L g13983 ( 
.A(n_12829),
.Y(n_13983)
);

INVx2_ASAP7_75t_SL g13984 ( 
.A(n_12869),
.Y(n_13984)
);

AND2x4_ASAP7_75t_L g13985 ( 
.A(n_12866),
.B(n_9154),
.Y(n_13985)
);

OR2x2_ASAP7_75t_L g13986 ( 
.A(n_13011),
.B(n_8380),
.Y(n_13986)
);

AND2x2_ASAP7_75t_L g13987 ( 
.A(n_13182),
.B(n_9154),
.Y(n_13987)
);

AND2x2_ASAP7_75t_L g13988 ( 
.A(n_13182),
.B(n_9155),
.Y(n_13988)
);

AND2x2_ASAP7_75t_L g13989 ( 
.A(n_13169),
.B(n_12853),
.Y(n_13989)
);

AND2x4_ASAP7_75t_L g13990 ( 
.A(n_12799),
.B(n_9155),
.Y(n_13990)
);

INVx1_ASAP7_75t_L g13991 ( 
.A(n_12834),
.Y(n_13991)
);

NAND2xp5_ASAP7_75t_L g13992 ( 
.A(n_13137),
.B(n_9849),
.Y(n_13992)
);

NAND2xp33_ASAP7_75t_SL g13993 ( 
.A(n_13216),
.B(n_5301),
.Y(n_13993)
);

INVx2_ASAP7_75t_L g13994 ( 
.A(n_13026),
.Y(n_13994)
);

HB1xp67_ASAP7_75t_L g13995 ( 
.A(n_13014),
.Y(n_13995)
);

OR2x6_ASAP7_75t_SL g13996 ( 
.A(n_12698),
.B(n_5128),
.Y(n_13996)
);

INVx3_ASAP7_75t_L g13997 ( 
.A(n_13024),
.Y(n_13997)
);

HB1xp67_ASAP7_75t_L g13998 ( 
.A(n_13014),
.Y(n_13998)
);

AND2x2_ASAP7_75t_L g13999 ( 
.A(n_13149),
.B(n_9155),
.Y(n_13999)
);

NOR2x1_ASAP7_75t_SL g14000 ( 
.A(n_13216),
.B(n_8168),
.Y(n_14000)
);

AND2x4_ASAP7_75t_L g14001 ( 
.A(n_12799),
.B(n_9155),
.Y(n_14001)
);

AND2x2_ASAP7_75t_L g14002 ( 
.A(n_13149),
.B(n_9183),
.Y(n_14002)
);

NAND2xp5_ASAP7_75t_L g14003 ( 
.A(n_13137),
.B(n_9849),
.Y(n_14003)
);

OAI221xp5_ASAP7_75t_L g14004 ( 
.A1(n_12746),
.A2(n_12254),
.B1(n_7767),
.B2(n_7845),
.C(n_7755),
.Y(n_14004)
);

INVx1_ASAP7_75t_L g14005 ( 
.A(n_12845),
.Y(n_14005)
);

INVx3_ASAP7_75t_L g14006 ( 
.A(n_13045),
.Y(n_14006)
);

INVx2_ASAP7_75t_L g14007 ( 
.A(n_12953),
.Y(n_14007)
);

INVx1_ASAP7_75t_L g14008 ( 
.A(n_12863),
.Y(n_14008)
);

NAND2xp5_ASAP7_75t_L g14009 ( 
.A(n_13205),
.B(n_13202),
.Y(n_14009)
);

INVx1_ASAP7_75t_L g14010 ( 
.A(n_12877),
.Y(n_14010)
);

INVx2_ASAP7_75t_R g14011 ( 
.A(n_13037),
.Y(n_14011)
);

INVx1_ASAP7_75t_L g14012 ( 
.A(n_12882),
.Y(n_14012)
);

INVx3_ASAP7_75t_L g14013 ( 
.A(n_13045),
.Y(n_14013)
);

AND2x4_ASAP7_75t_L g14014 ( 
.A(n_13073),
.B(n_9183),
.Y(n_14014)
);

AND2x2_ASAP7_75t_L g14015 ( 
.A(n_13264),
.B(n_9183),
.Y(n_14015)
);

AND2x2_ASAP7_75t_L g14016 ( 
.A(n_13267),
.B(n_9183),
.Y(n_14016)
);

INVx2_ASAP7_75t_L g14017 ( 
.A(n_12968),
.Y(n_14017)
);

INVx1_ASAP7_75t_L g14018 ( 
.A(n_12892),
.Y(n_14018)
);

AND2x2_ASAP7_75t_L g14019 ( 
.A(n_12903),
.B(n_9194),
.Y(n_14019)
);

INVx1_ASAP7_75t_L g14020 ( 
.A(n_12894),
.Y(n_14020)
);

AND2x2_ASAP7_75t_L g14021 ( 
.A(n_13242),
.B(n_9194),
.Y(n_14021)
);

AND2x2_ASAP7_75t_L g14022 ( 
.A(n_13255),
.B(n_9194),
.Y(n_14022)
);

INVx1_ASAP7_75t_L g14023 ( 
.A(n_12902),
.Y(n_14023)
);

NAND2xp5_ASAP7_75t_L g14024 ( 
.A(n_13202),
.B(n_9861),
.Y(n_14024)
);

BUFx6f_ASAP7_75t_L g14025 ( 
.A(n_12865),
.Y(n_14025)
);

OR2x2_ASAP7_75t_L g14026 ( 
.A(n_13290),
.B(n_8189),
.Y(n_14026)
);

AND2x2_ASAP7_75t_L g14027 ( 
.A(n_13260),
.B(n_9194),
.Y(n_14027)
);

BUFx2_ASAP7_75t_L g14028 ( 
.A(n_13118),
.Y(n_14028)
);

INVx1_ASAP7_75t_L g14029 ( 
.A(n_12906),
.Y(n_14029)
);

NAND2xp5_ASAP7_75t_L g14030 ( 
.A(n_12989),
.B(n_9861),
.Y(n_14030)
);

AND2x4_ASAP7_75t_L g14031 ( 
.A(n_13073),
.B(n_9229),
.Y(n_14031)
);

AND2x2_ASAP7_75t_L g14032 ( 
.A(n_13269),
.B(n_9229),
.Y(n_14032)
);

OAI22xp5_ASAP7_75t_L g14033 ( 
.A1(n_12744),
.A2(n_7798),
.B1(n_7769),
.B2(n_8247),
.Y(n_14033)
);

OR2x2_ASAP7_75t_L g14034 ( 
.A(n_13162),
.B(n_8200),
.Y(n_14034)
);

INVx1_ASAP7_75t_L g14035 ( 
.A(n_12908),
.Y(n_14035)
);

OR2x2_ASAP7_75t_L g14036 ( 
.A(n_13195),
.B(n_8200),
.Y(n_14036)
);

HB1xp67_ASAP7_75t_L g14037 ( 
.A(n_13113),
.Y(n_14037)
);

NAND2xp5_ASAP7_75t_L g14038 ( 
.A(n_13245),
.B(n_13277),
.Y(n_14038)
);

OAI21xp5_ASAP7_75t_SL g14039 ( 
.A1(n_12883),
.A2(n_8236),
.B(n_8057),
.Y(n_14039)
);

AND2x4_ASAP7_75t_L g14040 ( 
.A(n_13103),
.B(n_9229),
.Y(n_14040)
);

INVx1_ASAP7_75t_L g14041 ( 
.A(n_12913),
.Y(n_14041)
);

OR2x2_ASAP7_75t_L g14042 ( 
.A(n_13256),
.B(n_8536),
.Y(n_14042)
);

INVx2_ASAP7_75t_L g14043 ( 
.A(n_12964),
.Y(n_14043)
);

NOR2xp67_ASAP7_75t_L g14044 ( 
.A(n_12553),
.B(n_9229),
.Y(n_14044)
);

INVx1_ASAP7_75t_L g14045 ( 
.A(n_12928),
.Y(n_14045)
);

AND2x2_ASAP7_75t_L g14046 ( 
.A(n_13270),
.B(n_9245),
.Y(n_14046)
);

INVx1_ASAP7_75t_L g14047 ( 
.A(n_12934),
.Y(n_14047)
);

OAI22xp5_ASAP7_75t_L g14048 ( 
.A1(n_13221),
.A2(n_7769),
.B1(n_8247),
.B2(n_8416),
.Y(n_14048)
);

INVx1_ASAP7_75t_L g14049 ( 
.A(n_12937),
.Y(n_14049)
);

OAI22xp5_ASAP7_75t_SL g14050 ( 
.A1(n_13245),
.A2(n_6894),
.B1(n_6922),
.B2(n_6772),
.Y(n_14050)
);

NOR2xp33_ASAP7_75t_L g14051 ( 
.A(n_13096),
.B(n_9864),
.Y(n_14051)
);

AND2x2_ASAP7_75t_L g14052 ( 
.A(n_13228),
.B(n_9245),
.Y(n_14052)
);

AND2x2_ASAP7_75t_L g14053 ( 
.A(n_13315),
.B(n_13190),
.Y(n_14053)
);

AND2x2_ASAP7_75t_L g14054 ( 
.A(n_12976),
.B(n_9245),
.Y(n_14054)
);

NOR2x1_ASAP7_75t_SL g14055 ( 
.A(n_13216),
.B(n_8168),
.Y(n_14055)
);

INVx2_ASAP7_75t_L g14056 ( 
.A(n_12967),
.Y(n_14056)
);

INVx1_ASAP7_75t_L g14057 ( 
.A(n_12939),
.Y(n_14057)
);

AND2x2_ASAP7_75t_L g14058 ( 
.A(n_13301),
.B(n_9245),
.Y(n_14058)
);

NAND2xp5_ASAP7_75t_L g14059 ( 
.A(n_13277),
.B(n_9864),
.Y(n_14059)
);

NOR2x1p5_ASAP7_75t_L g14060 ( 
.A(n_13144),
.B(n_13072),
.Y(n_14060)
);

AND2x2_ASAP7_75t_L g14061 ( 
.A(n_12855),
.B(n_9262),
.Y(n_14061)
);

INVx2_ASAP7_75t_L g14062 ( 
.A(n_12975),
.Y(n_14062)
);

INVx4_ASAP7_75t_L g14063 ( 
.A(n_12962),
.Y(n_14063)
);

AND2x2_ASAP7_75t_L g14064 ( 
.A(n_12896),
.B(n_9262),
.Y(n_14064)
);

INVx2_ASAP7_75t_L g14065 ( 
.A(n_12997),
.Y(n_14065)
);

AND2x4_ASAP7_75t_L g14066 ( 
.A(n_13103),
.B(n_9262),
.Y(n_14066)
);

AND2x2_ASAP7_75t_L g14067 ( 
.A(n_13218),
.B(n_9262),
.Y(n_14067)
);

NOR2x1_ASAP7_75t_L g14068 ( 
.A(n_13145),
.B(n_13104),
.Y(n_14068)
);

NAND2xp5_ASAP7_75t_L g14069 ( 
.A(n_12993),
.B(n_9874),
.Y(n_14069)
);

INVx2_ASAP7_75t_L g14070 ( 
.A(n_13001),
.Y(n_14070)
);

INVx1_ASAP7_75t_L g14071 ( 
.A(n_12942),
.Y(n_14071)
);

AND2x4_ASAP7_75t_L g14072 ( 
.A(n_12895),
.B(n_9299),
.Y(n_14072)
);

AND2x2_ASAP7_75t_L g14073 ( 
.A(n_12965),
.B(n_9299),
.Y(n_14073)
);

INVx2_ASAP7_75t_L g14074 ( 
.A(n_13196),
.Y(n_14074)
);

HB1xp67_ASAP7_75t_L g14075 ( 
.A(n_13113),
.Y(n_14075)
);

OR2x2_ASAP7_75t_L g14076 ( 
.A(n_12616),
.B(n_8536),
.Y(n_14076)
);

INVx1_ASAP7_75t_L g14077 ( 
.A(n_12943),
.Y(n_14077)
);

AOI22xp33_ASAP7_75t_L g14078 ( 
.A1(n_13082),
.A2(n_8225),
.B1(n_8386),
.B2(n_7800),
.Y(n_14078)
);

INVx2_ASAP7_75t_L g14079 ( 
.A(n_12899),
.Y(n_14079)
);

AND2x2_ASAP7_75t_L g14080 ( 
.A(n_13189),
.B(n_9299),
.Y(n_14080)
);

INVx2_ASAP7_75t_L g14081 ( 
.A(n_13036),
.Y(n_14081)
);

INVx2_ASAP7_75t_L g14082 ( 
.A(n_13041),
.Y(n_14082)
);

INVx2_ASAP7_75t_L g14083 ( 
.A(n_13042),
.Y(n_14083)
);

NAND2xp5_ASAP7_75t_L g14084 ( 
.A(n_13058),
.B(n_9874),
.Y(n_14084)
);

INVx2_ASAP7_75t_L g14085 ( 
.A(n_13044),
.Y(n_14085)
);

INVx1_ASAP7_75t_L g14086 ( 
.A(n_12949),
.Y(n_14086)
);

BUFx2_ASAP7_75t_L g14087 ( 
.A(n_13118),
.Y(n_14087)
);

AND2x2_ASAP7_75t_L g14088 ( 
.A(n_13278),
.B(n_9299),
.Y(n_14088)
);

AND2x2_ASAP7_75t_L g14089 ( 
.A(n_13091),
.B(n_13065),
.Y(n_14089)
);

INVx1_ASAP7_75t_L g14090 ( 
.A(n_12952),
.Y(n_14090)
);

AND2x2_ASAP7_75t_L g14091 ( 
.A(n_13091),
.B(n_9300),
.Y(n_14091)
);

AND2x4_ASAP7_75t_L g14092 ( 
.A(n_12897),
.B(n_9300),
.Y(n_14092)
);

NOR2xp33_ASAP7_75t_L g14093 ( 
.A(n_12963),
.B(n_9875),
.Y(n_14093)
);

INVx3_ASAP7_75t_L g14094 ( 
.A(n_13034),
.Y(n_14094)
);

AND2x2_ASAP7_75t_L g14095 ( 
.A(n_13066),
.B(n_9300),
.Y(n_14095)
);

AOI22xp33_ASAP7_75t_L g14096 ( 
.A1(n_13336),
.A2(n_13306),
.B1(n_13219),
.B2(n_13291),
.Y(n_14096)
);

INVx1_ASAP7_75t_L g14097 ( 
.A(n_13355),
.Y(n_14097)
);

OR2x2_ASAP7_75t_L g14098 ( 
.A(n_13554),
.B(n_12620),
.Y(n_14098)
);

NAND3xp33_ASAP7_75t_L g14099 ( 
.A(n_13401),
.B(n_12735),
.C(n_13319),
.Y(n_14099)
);

NAND2xp5_ASAP7_75t_L g14100 ( 
.A(n_13454),
.B(n_13106),
.Y(n_14100)
);

AND2x4_ASAP7_75t_L g14101 ( 
.A(n_13337),
.B(n_12947),
.Y(n_14101)
);

INVx4_ASAP7_75t_L g14102 ( 
.A(n_13480),
.Y(n_14102)
);

INVx2_ASAP7_75t_SL g14103 ( 
.A(n_13669),
.Y(n_14103)
);

INVx1_ASAP7_75t_L g14104 ( 
.A(n_13465),
.Y(n_14104)
);

INVx2_ASAP7_75t_L g14105 ( 
.A(n_13927),
.Y(n_14105)
);

AND2x2_ASAP7_75t_L g14106 ( 
.A(n_13537),
.B(n_13298),
.Y(n_14106)
);

INVx1_ASAP7_75t_SL g14107 ( 
.A(n_13352),
.Y(n_14107)
);

OR2x2_ASAP7_75t_L g14108 ( 
.A(n_13569),
.B(n_13000),
.Y(n_14108)
);

NAND2xp5_ASAP7_75t_SL g14109 ( 
.A(n_13368),
.B(n_13254),
.Y(n_14109)
);

INVx2_ASAP7_75t_L g14110 ( 
.A(n_13927),
.Y(n_14110)
);

INVx2_ASAP7_75t_L g14111 ( 
.A(n_13927),
.Y(n_14111)
);

AOI22xp33_ASAP7_75t_L g14112 ( 
.A1(n_13330),
.A2(n_13229),
.B1(n_13254),
.B2(n_12723),
.Y(n_14112)
);

AND2x2_ASAP7_75t_L g14113 ( 
.A(n_13347),
.B(n_13236),
.Y(n_14113)
);

INVx2_ASAP7_75t_L g14114 ( 
.A(n_13386),
.Y(n_14114)
);

OR2x2_ASAP7_75t_L g14115 ( 
.A(n_13737),
.B(n_13004),
.Y(n_14115)
);

OR2x2_ASAP7_75t_L g14116 ( 
.A(n_14037),
.B(n_13031),
.Y(n_14116)
);

INVx1_ASAP7_75t_L g14117 ( 
.A(n_13393),
.Y(n_14117)
);

BUFx3_ASAP7_75t_L g14118 ( 
.A(n_13413),
.Y(n_14118)
);

INVx1_ASAP7_75t_L g14119 ( 
.A(n_13685),
.Y(n_14119)
);

INVx1_ASAP7_75t_L g14120 ( 
.A(n_13660),
.Y(n_14120)
);

AND2x2_ASAP7_75t_L g14121 ( 
.A(n_13415),
.B(n_13240),
.Y(n_14121)
);

AND2x2_ASAP7_75t_L g14122 ( 
.A(n_13888),
.B(n_13180),
.Y(n_14122)
);

AND2x4_ASAP7_75t_L g14123 ( 
.A(n_13481),
.B(n_12960),
.Y(n_14123)
);

AND2x2_ASAP7_75t_L g14124 ( 
.A(n_13343),
.B(n_13183),
.Y(n_14124)
);

NAND2xp5_ASAP7_75t_L g14125 ( 
.A(n_13856),
.B(n_13127),
.Y(n_14125)
);

INVx1_ASAP7_75t_L g14126 ( 
.A(n_14028),
.Y(n_14126)
);

INVx1_ASAP7_75t_L g14127 ( 
.A(n_14028),
.Y(n_14127)
);

INVx5_ASAP7_75t_L g14128 ( 
.A(n_13361),
.Y(n_14128)
);

INVx2_ASAP7_75t_L g14129 ( 
.A(n_13369),
.Y(n_14129)
);

CKINVDCx5p33_ASAP7_75t_R g14130 ( 
.A(n_13624),
.Y(n_14130)
);

BUFx6f_ASAP7_75t_L g14131 ( 
.A(n_13510),
.Y(n_14131)
);

INVx1_ASAP7_75t_L g14132 ( 
.A(n_14087),
.Y(n_14132)
);

AND2x2_ASAP7_75t_L g14133 ( 
.A(n_13705),
.B(n_13261),
.Y(n_14133)
);

INVx5_ASAP7_75t_L g14134 ( 
.A(n_13372),
.Y(n_14134)
);

AND2x2_ASAP7_75t_L g14135 ( 
.A(n_13329),
.B(n_13265),
.Y(n_14135)
);

INVx2_ASAP7_75t_L g14136 ( 
.A(n_13587),
.Y(n_14136)
);

BUFx2_ASAP7_75t_L g14137 ( 
.A(n_13475),
.Y(n_14137)
);

NAND2xp5_ASAP7_75t_L g14138 ( 
.A(n_13748),
.B(n_13127),
.Y(n_14138)
);

AND2x2_ASAP7_75t_L g14139 ( 
.A(n_13520),
.B(n_12986),
.Y(n_14139)
);

HB1xp67_ASAP7_75t_L g14140 ( 
.A(n_13475),
.Y(n_14140)
);

INVx1_ASAP7_75t_L g14141 ( 
.A(n_14087),
.Y(n_14141)
);

AND2x2_ASAP7_75t_L g14142 ( 
.A(n_13652),
.B(n_12991),
.Y(n_14142)
);

INVx2_ASAP7_75t_L g14143 ( 
.A(n_13766),
.Y(n_14143)
);

INVx2_ASAP7_75t_L g14144 ( 
.A(n_13470),
.Y(n_14144)
);

NAND2xp5_ASAP7_75t_L g14145 ( 
.A(n_13827),
.B(n_12692),
.Y(n_14145)
);

AND2x4_ASAP7_75t_L g14146 ( 
.A(n_13543),
.B(n_12995),
.Y(n_14146)
);

INVx1_ASAP7_75t_L g14147 ( 
.A(n_13995),
.Y(n_14147)
);

AND2x2_ASAP7_75t_L g14148 ( 
.A(n_13395),
.B(n_13312),
.Y(n_14148)
);

INVx1_ASAP7_75t_L g14149 ( 
.A(n_13998),
.Y(n_14149)
);

INVx2_ASAP7_75t_L g14150 ( 
.A(n_13492),
.Y(n_14150)
);

INVx4_ASAP7_75t_L g14151 ( 
.A(n_13398),
.Y(n_14151)
);

OR2x2_ASAP7_75t_L g14152 ( 
.A(n_14075),
.B(n_12583),
.Y(n_14152)
);

NAND2xp5_ASAP7_75t_L g14153 ( 
.A(n_13754),
.B(n_13310),
.Y(n_14153)
);

INVx1_ASAP7_75t_L g14154 ( 
.A(n_13664),
.Y(n_14154)
);

BUFx2_ASAP7_75t_L g14155 ( 
.A(n_13945),
.Y(n_14155)
);

INVx1_ASAP7_75t_L g14156 ( 
.A(n_13675),
.Y(n_14156)
);

INVx2_ASAP7_75t_SL g14157 ( 
.A(n_13669),
.Y(n_14157)
);

AND2x2_ASAP7_75t_L g14158 ( 
.A(n_13770),
.B(n_13246),
.Y(n_14158)
);

OAI22xp5_ASAP7_75t_L g14159 ( 
.A1(n_13428),
.A2(n_13101),
.B1(n_13303),
.B2(n_13208),
.Y(n_14159)
);

AND2x2_ASAP7_75t_L g14160 ( 
.A(n_13364),
.B(n_13005),
.Y(n_14160)
);

INVx2_ASAP7_75t_L g14161 ( 
.A(n_13764),
.Y(n_14161)
);

NAND2xp5_ASAP7_75t_L g14162 ( 
.A(n_13825),
.B(n_13666),
.Y(n_14162)
);

BUFx2_ASAP7_75t_L g14163 ( 
.A(n_13591),
.Y(n_14163)
);

AND2x2_ASAP7_75t_L g14164 ( 
.A(n_13645),
.B(n_13275),
.Y(n_14164)
);

OR2x2_ASAP7_75t_L g14165 ( 
.A(n_13357),
.B(n_13070),
.Y(n_14165)
);

AND2x4_ASAP7_75t_L g14166 ( 
.A(n_13593),
.B(n_13128),
.Y(n_14166)
);

INVxp67_ASAP7_75t_L g14167 ( 
.A(n_13832),
.Y(n_14167)
);

AND2x4_ASAP7_75t_L g14168 ( 
.A(n_13331),
.B(n_13128),
.Y(n_14168)
);

AOI22xp33_ASAP7_75t_L g14169 ( 
.A1(n_13412),
.A2(n_13244),
.B1(n_13295),
.B2(n_13200),
.Y(n_14169)
);

AND2x2_ASAP7_75t_L g14170 ( 
.A(n_13524),
.B(n_13273),
.Y(n_14170)
);

INVx1_ASAP7_75t_SL g14171 ( 
.A(n_13825),
.Y(n_14171)
);

BUFx2_ASAP7_75t_L g14172 ( 
.A(n_13591),
.Y(n_14172)
);

AO21x2_ASAP7_75t_L g14173 ( 
.A1(n_13567),
.A2(n_13021),
.B(n_13018),
.Y(n_14173)
);

AND2x2_ASAP7_75t_L g14174 ( 
.A(n_13899),
.B(n_13314),
.Y(n_14174)
);

AND2x2_ASAP7_75t_L g14175 ( 
.A(n_13384),
.B(n_13316),
.Y(n_14175)
);

INVx2_ASAP7_75t_L g14176 ( 
.A(n_13760),
.Y(n_14176)
);

NAND2xp5_ASAP7_75t_L g14177 ( 
.A(n_13666),
.B(n_13069),
.Y(n_14177)
);

INVx2_ASAP7_75t_L g14178 ( 
.A(n_13760),
.Y(n_14178)
);

AOI22xp33_ASAP7_75t_L g14179 ( 
.A1(n_13350),
.A2(n_13244),
.B1(n_13200),
.B2(n_13184),
.Y(n_14179)
);

AND2x2_ASAP7_75t_L g14180 ( 
.A(n_13418),
.B(n_12857),
.Y(n_14180)
);

HB1xp67_ASAP7_75t_L g14181 ( 
.A(n_13832),
.Y(n_14181)
);

AND2x2_ASAP7_75t_L g14182 ( 
.A(n_13440),
.B(n_12858),
.Y(n_14182)
);

AND2x2_ASAP7_75t_L g14183 ( 
.A(n_13700),
.B(n_12862),
.Y(n_14183)
);

OR2x2_ASAP7_75t_L g14184 ( 
.A(n_13532),
.B(n_12955),
.Y(n_14184)
);

HB1xp67_ASAP7_75t_L g14185 ( 
.A(n_13854),
.Y(n_14185)
);

INVx1_ASAP7_75t_L g14186 ( 
.A(n_13448),
.Y(n_14186)
);

INVx1_ASAP7_75t_L g14187 ( 
.A(n_13459),
.Y(n_14187)
);

INVx2_ASAP7_75t_L g14188 ( 
.A(n_13420),
.Y(n_14188)
);

INVx4_ASAP7_75t_L g14189 ( 
.A(n_13669),
.Y(n_14189)
);

INVx2_ASAP7_75t_L g14190 ( 
.A(n_13424),
.Y(n_14190)
);

AND2x2_ASAP7_75t_L g14191 ( 
.A(n_13821),
.B(n_12874),
.Y(n_14191)
);

INVxp67_ASAP7_75t_SL g14192 ( 
.A(n_13607),
.Y(n_14192)
);

AND2x2_ASAP7_75t_L g14193 ( 
.A(n_13324),
.B(n_12635),
.Y(n_14193)
);

AND2x2_ASAP7_75t_L g14194 ( 
.A(n_13503),
.B(n_13068),
.Y(n_14194)
);

AND2x2_ASAP7_75t_L g14195 ( 
.A(n_13527),
.B(n_12875),
.Y(n_14195)
);

INVx1_ASAP7_75t_SL g14196 ( 
.A(n_13854),
.Y(n_14196)
);

NAND2xp5_ASAP7_75t_L g14197 ( 
.A(n_13647),
.B(n_13135),
.Y(n_14197)
);

INVx1_ASAP7_75t_L g14198 ( 
.A(n_13779),
.Y(n_14198)
);

INVx2_ASAP7_75t_L g14199 ( 
.A(n_13731),
.Y(n_14199)
);

AND2x2_ASAP7_75t_L g14200 ( 
.A(n_13534),
.B(n_13551),
.Y(n_14200)
);

INVx1_ASAP7_75t_SL g14201 ( 
.A(n_13647),
.Y(n_14201)
);

AND2x4_ASAP7_75t_L g14202 ( 
.A(n_13403),
.B(n_12580),
.Y(n_14202)
);

INVx3_ASAP7_75t_L g14203 ( 
.A(n_13703),
.Y(n_14203)
);

INVx2_ASAP7_75t_L g14204 ( 
.A(n_13924),
.Y(n_14204)
);

INVx2_ASAP7_75t_L g14205 ( 
.A(n_13729),
.Y(n_14205)
);

BUFx3_ASAP7_75t_L g14206 ( 
.A(n_13403),
.Y(n_14206)
);

AND2x2_ASAP7_75t_L g14207 ( 
.A(n_13354),
.B(n_12878),
.Y(n_14207)
);

AND2x2_ASAP7_75t_L g14208 ( 
.A(n_14089),
.B(n_13174),
.Y(n_14208)
);

OR2x6_ASAP7_75t_L g14209 ( 
.A(n_13399),
.B(n_13104),
.Y(n_14209)
);

INVx2_ASAP7_75t_L g14210 ( 
.A(n_13947),
.Y(n_14210)
);

INVx1_ASAP7_75t_L g14211 ( 
.A(n_13784),
.Y(n_14211)
);

INVx2_ASAP7_75t_L g14212 ( 
.A(n_13948),
.Y(n_14212)
);

INVx1_ASAP7_75t_L g14213 ( 
.A(n_13490),
.Y(n_14213)
);

INVx1_ASAP7_75t_L g14214 ( 
.A(n_13512),
.Y(n_14214)
);

INVx2_ASAP7_75t_L g14215 ( 
.A(n_13930),
.Y(n_14215)
);

INVx2_ASAP7_75t_SL g14216 ( 
.A(n_13853),
.Y(n_14216)
);

INVx1_ASAP7_75t_L g14217 ( 
.A(n_13945),
.Y(n_14217)
);

OR2x6_ASAP7_75t_L g14218 ( 
.A(n_13439),
.B(n_13109),
.Y(n_14218)
);

NOR2xp33_ASAP7_75t_SL g14219 ( 
.A(n_13794),
.B(n_13617),
.Y(n_14219)
);

AND2x2_ASAP7_75t_L g14220 ( 
.A(n_13346),
.B(n_12910),
.Y(n_14220)
);

OR2x2_ASAP7_75t_SL g14221 ( 
.A(n_13408),
.B(n_13184),
.Y(n_14221)
);

NAND2xp5_ASAP7_75t_SL g14222 ( 
.A(n_13370),
.B(n_13184),
.Y(n_14222)
);

INVx4_ASAP7_75t_L g14223 ( 
.A(n_13930),
.Y(n_14223)
);

INVx2_ASAP7_75t_L g14224 ( 
.A(n_13641),
.Y(n_14224)
);

INVx1_ASAP7_75t_L g14225 ( 
.A(n_13977),
.Y(n_14225)
);

AND2x6_ASAP7_75t_L g14226 ( 
.A(n_13380),
.B(n_13109),
.Y(n_14226)
);

BUFx3_ASAP7_75t_L g14227 ( 
.A(n_13749),
.Y(n_14227)
);

AND2x4_ASAP7_75t_SL g14228 ( 
.A(n_14063),
.B(n_12843),
.Y(n_14228)
);

AND2x4_ASAP7_75t_SL g14229 ( 
.A(n_13828),
.B(n_12844),
.Y(n_14229)
);

OR2x2_ASAP7_75t_L g14230 ( 
.A(n_13382),
.B(n_12634),
.Y(n_14230)
);

INVxp67_ASAP7_75t_SL g14231 ( 
.A(n_13772),
.Y(n_14231)
);

AO21x2_ASAP7_75t_L g14232 ( 
.A1(n_13582),
.A2(n_13022),
.B(n_13021),
.Y(n_14232)
);

AND2x2_ASAP7_75t_L g14233 ( 
.A(n_13811),
.B(n_12911),
.Y(n_14233)
);

INVx1_ASAP7_75t_L g14234 ( 
.A(n_13977),
.Y(n_14234)
);

AOI22xp33_ASAP7_75t_L g14235 ( 
.A1(n_13622),
.A2(n_13200),
.B1(n_13249),
.B2(n_12886),
.Y(n_14235)
);

OR2x6_ASAP7_75t_L g14236 ( 
.A(n_13457),
.B(n_13160),
.Y(n_14236)
);

AO21x2_ASAP7_75t_L g14237 ( 
.A1(n_13603),
.A2(n_13032),
.B(n_13022),
.Y(n_14237)
);

NOR2x1_ASAP7_75t_SL g14238 ( 
.A(n_13573),
.B(n_13249),
.Y(n_14238)
);

INVx1_ASAP7_75t_L g14239 ( 
.A(n_13940),
.Y(n_14239)
);

AND2x4_ASAP7_75t_L g14240 ( 
.A(n_13566),
.B(n_12915),
.Y(n_14240)
);

HB1xp67_ASAP7_75t_L g14241 ( 
.A(n_13661),
.Y(n_14241)
);

OAI33xp33_ASAP7_75t_L g14242 ( 
.A1(n_13446),
.A2(n_13296),
.A3(n_13320),
.B1(n_13321),
.B2(n_13257),
.B3(n_12956),
.Y(n_14242)
);

AND2x2_ASAP7_75t_L g14243 ( 
.A(n_13787),
.B(n_14053),
.Y(n_14243)
);

INVx2_ASAP7_75t_L g14244 ( 
.A(n_13358),
.Y(n_14244)
);

AND2x2_ASAP7_75t_L g14245 ( 
.A(n_13989),
.B(n_12914),
.Y(n_14245)
);

INVx1_ASAP7_75t_L g14246 ( 
.A(n_13813),
.Y(n_14246)
);

INVx2_ASAP7_75t_L g14247 ( 
.A(n_13373),
.Y(n_14247)
);

AND2x2_ASAP7_75t_L g14248 ( 
.A(n_13394),
.B(n_12907),
.Y(n_14248)
);

OR2x2_ASAP7_75t_L g14249 ( 
.A(n_13362),
.B(n_13363),
.Y(n_14249)
);

INVx2_ASAP7_75t_L g14250 ( 
.A(n_13378),
.Y(n_14250)
);

INVx1_ASAP7_75t_L g14251 ( 
.A(n_13813),
.Y(n_14251)
);

INVx2_ASAP7_75t_L g14252 ( 
.A(n_13379),
.Y(n_14252)
);

OR2x2_ASAP7_75t_L g14253 ( 
.A(n_13678),
.B(n_12526),
.Y(n_14253)
);

AND2x4_ASAP7_75t_L g14254 ( 
.A(n_13566),
.B(n_12916),
.Y(n_14254)
);

AOI22xp33_ASAP7_75t_L g14255 ( 
.A1(n_13349),
.A2(n_13249),
.B1(n_13224),
.B2(n_12460),
.Y(n_14255)
);

HB1xp67_ASAP7_75t_L g14256 ( 
.A(n_13661),
.Y(n_14256)
);

NAND2x1_ASAP7_75t_L g14257 ( 
.A(n_13344),
.B(n_13007),
.Y(n_14257)
);

AND2x2_ASAP7_75t_L g14258 ( 
.A(n_13826),
.B(n_12921),
.Y(n_14258)
);

AND2x2_ASAP7_75t_L g14259 ( 
.A(n_13709),
.B(n_12846),
.Y(n_14259)
);

BUFx3_ASAP7_75t_L g14260 ( 
.A(n_13749),
.Y(n_14260)
);

NOR2x1_ASAP7_75t_L g14261 ( 
.A(n_13435),
.B(n_13032),
.Y(n_14261)
);

AND2x2_ASAP7_75t_L g14262 ( 
.A(n_13712),
.B(n_13433),
.Y(n_14262)
);

AND2x2_ASAP7_75t_L g14263 ( 
.A(n_13325),
.B(n_13317),
.Y(n_14263)
);

INVx2_ASAP7_75t_L g14264 ( 
.A(n_13866),
.Y(n_14264)
);

INVx2_ASAP7_75t_L g14265 ( 
.A(n_13883),
.Y(n_14265)
);

AND2x2_ASAP7_75t_L g14266 ( 
.A(n_13575),
.B(n_13155),
.Y(n_14266)
);

INVx2_ASAP7_75t_L g14267 ( 
.A(n_13579),
.Y(n_14267)
);

OAI22xp33_ASAP7_75t_L g14268 ( 
.A1(n_13351),
.A2(n_13271),
.B1(n_13293),
.B2(n_13280),
.Y(n_14268)
);

INVx1_ASAP7_75t_L g14269 ( 
.A(n_13813),
.Y(n_14269)
);

INVx2_ASAP7_75t_L g14270 ( 
.A(n_14000),
.Y(n_14270)
);

BUFx2_ASAP7_75t_L g14271 ( 
.A(n_13830),
.Y(n_14271)
);

AND2x2_ASAP7_75t_L g14272 ( 
.A(n_13342),
.B(n_13339),
.Y(n_14272)
);

NOR3xp33_ASAP7_75t_L g14273 ( 
.A(n_13486),
.B(n_13126),
.C(n_13274),
.Y(n_14273)
);

HB1xp67_ASAP7_75t_L g14274 ( 
.A(n_13886),
.Y(n_14274)
);

BUFx2_ASAP7_75t_L g14275 ( 
.A(n_13410),
.Y(n_14275)
);

NAND2xp5_ASAP7_75t_SL g14276 ( 
.A(n_13348),
.B(n_13160),
.Y(n_14276)
);

INVx1_ASAP7_75t_L g14277 ( 
.A(n_13813),
.Y(n_14277)
);

AND2x4_ASAP7_75t_L g14278 ( 
.A(n_13604),
.B(n_12917),
.Y(n_14278)
);

AND2x2_ASAP7_75t_L g14279 ( 
.A(n_13332),
.B(n_12925),
.Y(n_14279)
);

INVx1_ASAP7_75t_L g14280 ( 
.A(n_13410),
.Y(n_14280)
);

INVx2_ASAP7_75t_L g14281 ( 
.A(n_14055),
.Y(n_14281)
);

AND2x2_ASAP7_75t_L g14282 ( 
.A(n_13340),
.B(n_13695),
.Y(n_14282)
);

OR2x2_ASAP7_75t_L g14283 ( 
.A(n_13359),
.B(n_12613),
.Y(n_14283)
);

AND2x2_ASAP7_75t_L g14284 ( 
.A(n_13892),
.B(n_13046),
.Y(n_14284)
);

NAND2xp5_ASAP7_75t_L g14285 ( 
.A(n_13594),
.B(n_12922),
.Y(n_14285)
);

INVx1_ASAP7_75t_L g14286 ( 
.A(n_13975),
.Y(n_14286)
);

NAND2xp5_ASAP7_75t_L g14287 ( 
.A(n_13404),
.B(n_12933),
.Y(n_14287)
);

AOI22xp33_ASAP7_75t_SL g14288 ( 
.A1(n_13366),
.A2(n_12841),
.B1(n_12737),
.B2(n_13282),
.Y(n_14288)
);

INVx1_ASAP7_75t_L g14289 ( 
.A(n_13371),
.Y(n_14289)
);

INVx2_ASAP7_75t_SL g14290 ( 
.A(n_13900),
.Y(n_14290)
);

INVx3_ASAP7_75t_L g14291 ( 
.A(n_13751),
.Y(n_14291)
);

INVx2_ASAP7_75t_L g14292 ( 
.A(n_13353),
.Y(n_14292)
);

AND2x2_ASAP7_75t_L g14293 ( 
.A(n_13922),
.B(n_13936),
.Y(n_14293)
);

NAND2xp5_ASAP7_75t_L g14294 ( 
.A(n_13706),
.B(n_12935),
.Y(n_14294)
);

INVx1_ASAP7_75t_L g14295 ( 
.A(n_13443),
.Y(n_14295)
);

INVx1_ASAP7_75t_L g14296 ( 
.A(n_13323),
.Y(n_14296)
);

AND2x2_ASAP7_75t_L g14297 ( 
.A(n_13604),
.B(n_13047),
.Y(n_14297)
);

AOI211xp5_ASAP7_75t_L g14298 ( 
.A1(n_13383),
.A2(n_13129),
.B(n_13105),
.C(n_13098),
.Y(n_14298)
);

AND2x2_ASAP7_75t_L g14299 ( 
.A(n_13365),
.B(n_13150),
.Y(n_14299)
);

BUFx3_ASAP7_75t_L g14300 ( 
.A(n_13542),
.Y(n_14300)
);

INVx5_ASAP7_75t_SL g14301 ( 
.A(n_14025),
.Y(n_14301)
);

CKINVDCx20_ASAP7_75t_R g14302 ( 
.A(n_13993),
.Y(n_14302)
);

NOR2xp67_ASAP7_75t_L g14303 ( 
.A(n_13903),
.B(n_12959),
.Y(n_14303)
);

INVx2_ASAP7_75t_L g14304 ( 
.A(n_13356),
.Y(n_14304)
);

OR2x2_ASAP7_75t_L g14305 ( 
.A(n_13558),
.B(n_12647),
.Y(n_14305)
);

AND2x4_ASAP7_75t_L g14306 ( 
.A(n_13511),
.B(n_12936),
.Y(n_14306)
);

OR2x6_ASAP7_75t_SL g14307 ( 
.A(n_13599),
.B(n_12940),
.Y(n_14307)
);

HB1xp67_ASAP7_75t_L g14308 ( 
.A(n_13913),
.Y(n_14308)
);

INVx2_ASAP7_75t_L g14309 ( 
.A(n_13724),
.Y(n_14309)
);

INVx2_ASAP7_75t_L g14310 ( 
.A(n_13725),
.Y(n_14310)
);

AND2x2_ASAP7_75t_L g14311 ( 
.A(n_13595),
.B(n_12819),
.Y(n_14311)
);

AND2x2_ASAP7_75t_L g14312 ( 
.A(n_13333),
.B(n_12919),
.Y(n_14312)
);

AND2x4_ASAP7_75t_L g14313 ( 
.A(n_13518),
.B(n_12946),
.Y(n_14313)
);

OR2x2_ASAP7_75t_SL g14314 ( 
.A(n_13635),
.B(n_12954),
.Y(n_14314)
);

INVx1_ASAP7_75t_L g14315 ( 
.A(n_13334),
.Y(n_14315)
);

AND2x2_ASAP7_75t_SL g14316 ( 
.A(n_13859),
.B(n_12671),
.Y(n_14316)
);

INVx3_ASAP7_75t_L g14317 ( 
.A(n_13790),
.Y(n_14317)
);

AOI22xp33_ASAP7_75t_L g14318 ( 
.A1(n_13592),
.A2(n_13203),
.B1(n_13248),
.B2(n_13188),
.Y(n_14318)
);

OR2x2_ASAP7_75t_L g14319 ( 
.A(n_13722),
.B(n_12950),
.Y(n_14319)
);

HB1xp67_ASAP7_75t_L g14320 ( 
.A(n_13773),
.Y(n_14320)
);

BUFx2_ASAP7_75t_L g14321 ( 
.A(n_13628),
.Y(n_14321)
);

OR2x2_ASAP7_75t_L g14322 ( 
.A(n_13778),
.B(n_12509),
.Y(n_14322)
);

OR2x2_ASAP7_75t_L g14323 ( 
.A(n_13360),
.B(n_12511),
.Y(n_14323)
);

HB1xp67_ASAP7_75t_L g14324 ( 
.A(n_14068),
.Y(n_14324)
);

AND2x2_ASAP7_75t_L g14325 ( 
.A(n_13915),
.B(n_13050),
.Y(n_14325)
);

INVx1_ASAP7_75t_L g14326 ( 
.A(n_13374),
.Y(n_14326)
);

NAND2xp5_ASAP7_75t_L g14327 ( 
.A(n_13730),
.B(n_12957),
.Y(n_14327)
);

OR2x2_ASAP7_75t_L g14328 ( 
.A(n_14026),
.B(n_12528),
.Y(n_14328)
);

INVx3_ASAP7_75t_L g14329 ( 
.A(n_14040),
.Y(n_14329)
);

AND2x4_ASAP7_75t_L g14330 ( 
.A(n_13462),
.B(n_13110),
.Y(n_14330)
);

AND2x2_ASAP7_75t_L g14331 ( 
.A(n_13959),
.B(n_13629),
.Y(n_14331)
);

AND2x2_ASAP7_75t_L g14332 ( 
.A(n_13630),
.B(n_13102),
.Y(n_14332)
);

INVx1_ASAP7_75t_L g14333 ( 
.A(n_13375),
.Y(n_14333)
);

OR2x2_ASAP7_75t_L g14334 ( 
.A(n_13687),
.B(n_12961),
.Y(n_14334)
);

INVx1_ASAP7_75t_L g14335 ( 
.A(n_13376),
.Y(n_14335)
);

BUFx2_ASAP7_75t_L g14336 ( 
.A(n_13904),
.Y(n_14336)
);

INVx1_ASAP7_75t_L g14337 ( 
.A(n_13388),
.Y(n_14337)
);

INVx2_ASAP7_75t_SL g14338 ( 
.A(n_13865),
.Y(n_14338)
);

INVx2_ASAP7_75t_L g14339 ( 
.A(n_13741),
.Y(n_14339)
);

OR2x2_ASAP7_75t_L g14340 ( 
.A(n_13690),
.B(n_12547),
.Y(n_14340)
);

INVx1_ASAP7_75t_SL g14341 ( 
.A(n_13999),
.Y(n_14341)
);

INVx1_ASAP7_75t_L g14342 ( 
.A(n_13390),
.Y(n_14342)
);

INVx4_ASAP7_75t_L g14343 ( 
.A(n_13471),
.Y(n_14343)
);

INVx2_ASAP7_75t_L g14344 ( 
.A(n_13797),
.Y(n_14344)
);

BUFx2_ASAP7_75t_L g14345 ( 
.A(n_13708),
.Y(n_14345)
);

HB1xp67_ASAP7_75t_L g14346 ( 
.A(n_13788),
.Y(n_14346)
);

INVx2_ASAP7_75t_L g14347 ( 
.A(n_13814),
.Y(n_14347)
);

INVx2_ASAP7_75t_L g14348 ( 
.A(n_14040),
.Y(n_14348)
);

AND2x2_ASAP7_75t_L g14349 ( 
.A(n_13634),
.B(n_12980),
.Y(n_14349)
);

AND2x2_ASAP7_75t_L g14350 ( 
.A(n_13639),
.B(n_12981),
.Y(n_14350)
);

INVx2_ASAP7_75t_L g14351 ( 
.A(n_14066),
.Y(n_14351)
);

BUFx2_ASAP7_75t_L g14352 ( 
.A(n_13793),
.Y(n_14352)
);

INVx2_ASAP7_75t_SL g14353 ( 
.A(n_14014),
.Y(n_14353)
);

INVx4_ASAP7_75t_L g14354 ( 
.A(n_13484),
.Y(n_14354)
);

AND2x2_ASAP7_75t_L g14355 ( 
.A(n_13643),
.B(n_12987),
.Y(n_14355)
);

BUFx2_ASAP7_75t_L g14356 ( 
.A(n_13644),
.Y(n_14356)
);

BUFx6f_ASAP7_75t_L g14357 ( 
.A(n_13649),
.Y(n_14357)
);

INVx2_ASAP7_75t_L g14358 ( 
.A(n_14066),
.Y(n_14358)
);

INVx1_ASAP7_75t_L g14359 ( 
.A(n_13397),
.Y(n_14359)
);

AND2x2_ASAP7_75t_L g14360 ( 
.A(n_13602),
.B(n_12988),
.Y(n_14360)
);

AND2x2_ASAP7_75t_L g14361 ( 
.A(n_13621),
.B(n_13326),
.Y(n_14361)
);

INVx2_ASAP7_75t_L g14362 ( 
.A(n_13837),
.Y(n_14362)
);

INVxp67_ASAP7_75t_SL g14363 ( 
.A(n_13636),
.Y(n_14363)
);

NOR2xp33_ASAP7_75t_L g14364 ( 
.A(n_13453),
.B(n_12610),
.Y(n_14364)
);

HB1xp67_ASAP7_75t_L g14365 ( 
.A(n_13557),
.Y(n_14365)
);

INVx3_ASAP7_75t_L g14366 ( 
.A(n_14014),
.Y(n_14366)
);

AND2x2_ASAP7_75t_L g14367 ( 
.A(n_13338),
.B(n_13768),
.Y(n_14367)
);

AND2x2_ASAP7_75t_L g14368 ( 
.A(n_13711),
.B(n_13006),
.Y(n_14368)
);

HB1xp67_ASAP7_75t_L g14369 ( 
.A(n_13668),
.Y(n_14369)
);

INVx1_ASAP7_75t_L g14370 ( 
.A(n_13402),
.Y(n_14370)
);

OR2x6_ASAP7_75t_L g14371 ( 
.A(n_14060),
.B(n_12814),
.Y(n_14371)
);

HB1xp67_ASAP7_75t_L g14372 ( 
.A(n_13680),
.Y(n_14372)
);

INVx1_ASAP7_75t_L g14373 ( 
.A(n_13405),
.Y(n_14373)
);

BUFx2_ASAP7_75t_L g14374 ( 
.A(n_13682),
.Y(n_14374)
);

OR2x2_ASAP7_75t_L g14375 ( 
.A(n_13699),
.B(n_12994),
.Y(n_14375)
);

BUFx2_ASAP7_75t_L g14376 ( 
.A(n_13684),
.Y(n_14376)
);

OR2x6_ASAP7_75t_L g14377 ( 
.A(n_14025),
.B(n_12817),
.Y(n_14377)
);

AOI22xp33_ASAP7_75t_L g14378 ( 
.A1(n_13555),
.A2(n_13028),
.B1(n_13030),
.B2(n_13020),
.Y(n_14378)
);

INVxp67_ASAP7_75t_SL g14379 ( 
.A(n_13367),
.Y(n_14379)
);

INVx1_ASAP7_75t_L g14380 ( 
.A(n_13409),
.Y(n_14380)
);

INVx1_ASAP7_75t_L g14381 ( 
.A(n_13411),
.Y(n_14381)
);

INVx1_ASAP7_75t_L g14382 ( 
.A(n_13419),
.Y(n_14382)
);

INVx1_ASAP7_75t_L g14383 ( 
.A(n_13426),
.Y(n_14383)
);

NAND2xp5_ASAP7_75t_L g14384 ( 
.A(n_13879),
.B(n_13272),
.Y(n_14384)
);

INVx2_ASAP7_75t_SL g14385 ( 
.A(n_14031),
.Y(n_14385)
);

AO21x2_ASAP7_75t_L g14386 ( 
.A1(n_13605),
.A2(n_13120),
.B(n_13112),
.Y(n_14386)
);

AND2x4_ASAP7_75t_L g14387 ( 
.A(n_13750),
.B(n_13094),
.Y(n_14387)
);

AND2x2_ASAP7_75t_L g14388 ( 
.A(n_13855),
.B(n_12926),
.Y(n_14388)
);

INVx1_ASAP7_75t_L g14389 ( 
.A(n_13434),
.Y(n_14389)
);

NAND2xp5_ASAP7_75t_L g14390 ( 
.A(n_13488),
.B(n_13272),
.Y(n_14390)
);

INVx2_ASAP7_75t_L g14391 ( 
.A(n_13843),
.Y(n_14391)
);

AND2x2_ASAP7_75t_L g14392 ( 
.A(n_13862),
.B(n_12927),
.Y(n_14392)
);

BUFx2_ASAP7_75t_L g14393 ( 
.A(n_13499),
.Y(n_14393)
);

INVx1_ASAP7_75t_L g14394 ( 
.A(n_13442),
.Y(n_14394)
);

INVx1_ASAP7_75t_L g14395 ( 
.A(n_13445),
.Y(n_14395)
);

AND2x2_ASAP7_75t_L g14396 ( 
.A(n_13870),
.B(n_12932),
.Y(n_14396)
);

INVx1_ASAP7_75t_L g14397 ( 
.A(n_13447),
.Y(n_14397)
);

BUFx2_ASAP7_75t_SL g14398 ( 
.A(n_13973),
.Y(n_14398)
);

NOR2xp33_ASAP7_75t_L g14399 ( 
.A(n_13385),
.B(n_13017),
.Y(n_14399)
);

INVx2_ASAP7_75t_L g14400 ( 
.A(n_13928),
.Y(n_14400)
);

INVx1_ASAP7_75t_L g14401 ( 
.A(n_13455),
.Y(n_14401)
);

INVx1_ASAP7_75t_L g14402 ( 
.A(n_13456),
.Y(n_14402)
);

INVx1_ASAP7_75t_L g14403 ( 
.A(n_13460),
.Y(n_14403)
);

INVx3_ASAP7_75t_L g14404 ( 
.A(n_14031),
.Y(n_14404)
);

INVx1_ASAP7_75t_L g14405 ( 
.A(n_13463),
.Y(n_14405)
);

INVx1_ASAP7_75t_L g14406 ( 
.A(n_13468),
.Y(n_14406)
);

INVx2_ASAP7_75t_L g14407 ( 
.A(n_13997),
.Y(n_14407)
);

INVx2_ASAP7_75t_L g14408 ( 
.A(n_14094),
.Y(n_14408)
);

OR2x2_ASAP7_75t_L g14409 ( 
.A(n_13740),
.B(n_12860),
.Y(n_14409)
);

HB1xp67_ASAP7_75t_L g14410 ( 
.A(n_13344),
.Y(n_14410)
);

INVx1_ASAP7_75t_L g14411 ( 
.A(n_13472),
.Y(n_14411)
);

AND2x2_ASAP7_75t_L g14412 ( 
.A(n_13881),
.B(n_13885),
.Y(n_14412)
);

INVx2_ASAP7_75t_SL g14413 ( 
.A(n_13990),
.Y(n_14413)
);

INVx2_ASAP7_75t_L g14414 ( 
.A(n_14006),
.Y(n_14414)
);

NAND2xp5_ASAP7_75t_L g14415 ( 
.A(n_13529),
.B(n_12900),
.Y(n_14415)
);

INVx1_ASAP7_75t_L g14416 ( 
.A(n_13476),
.Y(n_14416)
);

INVx2_ASAP7_75t_L g14417 ( 
.A(n_14013),
.Y(n_14417)
);

INVx3_ASAP7_75t_L g14418 ( 
.A(n_13990),
.Y(n_14418)
);

AND2x2_ASAP7_75t_L g14419 ( 
.A(n_13531),
.B(n_13071),
.Y(n_14419)
);

INVx1_ASAP7_75t_L g14420 ( 
.A(n_13478),
.Y(n_14420)
);

AOI22xp5_ASAP7_75t_L g14421 ( 
.A1(n_13450),
.A2(n_13735),
.B1(n_13774),
.B2(n_13763),
.Y(n_14421)
);

INVx1_ASAP7_75t_L g14422 ( 
.A(n_13479),
.Y(n_14422)
);

INVx1_ASAP7_75t_L g14423 ( 
.A(n_13485),
.Y(n_14423)
);

INVx1_ASAP7_75t_L g14424 ( 
.A(n_13487),
.Y(n_14424)
);

HB1xp67_ASAP7_75t_L g14425 ( 
.A(n_13970),
.Y(n_14425)
);

INVx1_ASAP7_75t_L g14426 ( 
.A(n_13493),
.Y(n_14426)
);

INVx1_ASAP7_75t_L g14427 ( 
.A(n_13494),
.Y(n_14427)
);

INVx1_ASAP7_75t_L g14428 ( 
.A(n_13501),
.Y(n_14428)
);

AND2x2_ASAP7_75t_L g14429 ( 
.A(n_14002),
.B(n_13075),
.Y(n_14429)
);

INVx2_ASAP7_75t_L g14430 ( 
.A(n_13464),
.Y(n_14430)
);

BUFx3_ASAP7_75t_L g14431 ( 
.A(n_13560),
.Y(n_14431)
);

HB1xp67_ASAP7_75t_L g14432 ( 
.A(n_13971),
.Y(n_14432)
);

AND2x2_ASAP7_75t_L g14433 ( 
.A(n_13876),
.B(n_13076),
.Y(n_14433)
);

OR2x2_ASAP7_75t_L g14434 ( 
.A(n_13561),
.B(n_12912),
.Y(n_14434)
);

INVx1_ASAP7_75t_L g14435 ( 
.A(n_13507),
.Y(n_14435)
);

BUFx3_ASAP7_75t_L g14436 ( 
.A(n_13620),
.Y(n_14436)
);

INVx2_ASAP7_75t_L g14437 ( 
.A(n_13464),
.Y(n_14437)
);

INVx1_ASAP7_75t_L g14438 ( 
.A(n_13508),
.Y(n_14438)
);

OR2x2_ASAP7_75t_L g14439 ( 
.A(n_14009),
.B(n_12941),
.Y(n_14439)
);

BUFx2_ASAP7_75t_L g14440 ( 
.A(n_13638),
.Y(n_14440)
);

HB1xp67_ASAP7_75t_L g14441 ( 
.A(n_13638),
.Y(n_14441)
);

NAND4xp25_ASAP7_75t_L g14442 ( 
.A(n_13335),
.B(n_13201),
.C(n_13087),
.D(n_12982),
.Y(n_14442)
);

AND2x2_ASAP7_75t_L g14443 ( 
.A(n_14079),
.B(n_13086),
.Y(n_14443)
);

BUFx3_ASAP7_75t_L g14444 ( 
.A(n_13620),
.Y(n_14444)
);

HB1xp67_ASAP7_75t_L g14445 ( 
.A(n_13642),
.Y(n_14445)
);

OR2x2_ASAP7_75t_L g14446 ( 
.A(n_13720),
.B(n_12970),
.Y(n_14446)
);

BUFx2_ASAP7_75t_L g14447 ( 
.A(n_13642),
.Y(n_14447)
);

INVx1_ASAP7_75t_L g14448 ( 
.A(n_13513),
.Y(n_14448)
);

INVx2_ASAP7_75t_L g14449 ( 
.A(n_13477),
.Y(n_14449)
);

AND2x2_ASAP7_75t_L g14450 ( 
.A(n_14081),
.B(n_13088),
.Y(n_14450)
);

INVx1_ASAP7_75t_L g14451 ( 
.A(n_13517),
.Y(n_14451)
);

INVx1_ASAP7_75t_SL g14452 ( 
.A(n_14073),
.Y(n_14452)
);

OR2x2_ASAP7_75t_L g14453 ( 
.A(n_13849),
.B(n_12851),
.Y(n_14453)
);

INVx1_ASAP7_75t_L g14454 ( 
.A(n_13522),
.Y(n_14454)
);

INVxp67_ASAP7_75t_SL g14455 ( 
.A(n_13781),
.Y(n_14455)
);

AND2x2_ASAP7_75t_L g14456 ( 
.A(n_14082),
.B(n_13090),
.Y(n_14456)
);

AND2x2_ASAP7_75t_L g14457 ( 
.A(n_14083),
.B(n_13092),
.Y(n_14457)
);

INVx1_ASAP7_75t_L g14458 ( 
.A(n_13523),
.Y(n_14458)
);

BUFx6f_ASAP7_75t_L g14459 ( 
.A(n_13841),
.Y(n_14459)
);

INVx1_ASAP7_75t_L g14460 ( 
.A(n_13528),
.Y(n_14460)
);

AND2x2_ASAP7_75t_L g14461 ( 
.A(n_14085),
.B(n_13093),
.Y(n_14461)
);

INVx1_ASAP7_75t_L g14462 ( 
.A(n_13530),
.Y(n_14462)
);

AO21x2_ASAP7_75t_L g14463 ( 
.A1(n_14038),
.A2(n_13120),
.B(n_13112),
.Y(n_14463)
);

AND2x2_ASAP7_75t_L g14464 ( 
.A(n_14019),
.B(n_13247),
.Y(n_14464)
);

AND2x4_ASAP7_75t_L g14465 ( 
.A(n_13829),
.B(n_12852),
.Y(n_14465)
);

AND2x4_ASAP7_75t_L g14466 ( 
.A(n_13833),
.B(n_13034),
.Y(n_14466)
);

INVx2_ASAP7_75t_L g14467 ( 
.A(n_13477),
.Y(n_14467)
);

BUFx6f_ASAP7_75t_L g14468 ( 
.A(n_13943),
.Y(n_14468)
);

OR2x2_ASAP7_75t_L g14469 ( 
.A(n_13955),
.B(n_12873),
.Y(n_14469)
);

AOI22xp33_ASAP7_75t_L g14470 ( 
.A1(n_13473),
.A2(n_13227),
.B1(n_13220),
.B2(n_12918),
.Y(n_14470)
);

INVx2_ASAP7_75t_L g14471 ( 
.A(n_13752),
.Y(n_14471)
);

INVx2_ASAP7_75t_L g14472 ( 
.A(n_13625),
.Y(n_14472)
);

INVx4_ASAP7_75t_L g14473 ( 
.A(n_13467),
.Y(n_14473)
);

AND2x2_ASAP7_75t_L g14474 ( 
.A(n_14074),
.B(n_13247),
.Y(n_14474)
);

INVx2_ASAP7_75t_L g14475 ( 
.A(n_13968),
.Y(n_14475)
);

AND2x2_ASAP7_75t_L g14476 ( 
.A(n_14021),
.B(n_13251),
.Y(n_14476)
);

BUFx3_ASAP7_75t_L g14477 ( 
.A(n_13619),
.Y(n_14477)
);

INVx2_ASAP7_75t_SL g14478 ( 
.A(n_14001),
.Y(n_14478)
);

INVx1_ASAP7_75t_SL g14479 ( 
.A(n_14015),
.Y(n_14479)
);

AND2x2_ASAP7_75t_L g14480 ( 
.A(n_14022),
.B(n_14027),
.Y(n_14480)
);

AND2x2_ASAP7_75t_L g14481 ( 
.A(n_14016),
.B(n_13251),
.Y(n_14481)
);

INVx1_ASAP7_75t_L g14482 ( 
.A(n_13544),
.Y(n_14482)
);

AO21x2_ASAP7_75t_L g14483 ( 
.A1(n_13650),
.A2(n_13060),
.B(n_13055),
.Y(n_14483)
);

OAI21xp5_ASAP7_75t_L g14484 ( 
.A1(n_13701),
.A2(n_13053),
.B(n_12880),
.Y(n_14484)
);

AND2x2_ASAP7_75t_L g14485 ( 
.A(n_14007),
.B(n_13056),
.Y(n_14485)
);

INVx2_ASAP7_75t_L g14486 ( 
.A(n_13969),
.Y(n_14486)
);

INVx2_ASAP7_75t_L g14487 ( 
.A(n_13746),
.Y(n_14487)
);

AND2x2_ASAP7_75t_L g14488 ( 
.A(n_14017),
.B(n_13423),
.Y(n_14488)
);

INVx2_ASAP7_75t_L g14489 ( 
.A(n_13925),
.Y(n_14489)
);

INVx1_ASAP7_75t_L g14490 ( 
.A(n_13545),
.Y(n_14490)
);

BUFx3_ASAP7_75t_L g14491 ( 
.A(n_13601),
.Y(n_14491)
);

INVx2_ASAP7_75t_L g14492 ( 
.A(n_13925),
.Y(n_14492)
);

INVx2_ASAP7_75t_L g14493 ( 
.A(n_13929),
.Y(n_14493)
);

BUFx2_ASAP7_75t_L g14494 ( 
.A(n_14001),
.Y(n_14494)
);

AND2x2_ASAP7_75t_L g14495 ( 
.A(n_13732),
.B(n_13152),
.Y(n_14495)
);

HB1xp67_ASAP7_75t_L g14496 ( 
.A(n_13539),
.Y(n_14496)
);

INVx5_ASAP7_75t_L g14497 ( 
.A(n_13437),
.Y(n_14497)
);

INVx1_ASAP7_75t_L g14498 ( 
.A(n_13546),
.Y(n_14498)
);

INVx1_ASAP7_75t_L g14499 ( 
.A(n_13548),
.Y(n_14499)
);

AND2x4_ASAP7_75t_L g14500 ( 
.A(n_13984),
.B(n_13117),
.Y(n_14500)
);

OR2x2_ASAP7_75t_L g14501 ( 
.A(n_13392),
.B(n_12888),
.Y(n_14501)
);

INVx2_ASAP7_75t_L g14502 ( 
.A(n_13929),
.Y(n_14502)
);

OR2x2_ASAP7_75t_SL g14503 ( 
.A(n_13328),
.B(n_13167),
.Y(n_14503)
);

INVx1_ASAP7_75t_L g14504 ( 
.A(n_13549),
.Y(n_14504)
);

BUFx2_ASAP7_75t_L g14505 ( 
.A(n_14052),
.Y(n_14505)
);

BUFx3_ASAP7_75t_L g14506 ( 
.A(n_13482),
.Y(n_14506)
);

AND2x2_ASAP7_75t_L g14507 ( 
.A(n_13733),
.B(n_13119),
.Y(n_14507)
);

INVx1_ASAP7_75t_L g14508 ( 
.A(n_13550),
.Y(n_14508)
);

INVxp67_ASAP7_75t_SL g14509 ( 
.A(n_13637),
.Y(n_14509)
);

AND2x2_ASAP7_75t_L g14510 ( 
.A(n_13738),
.B(n_13122),
.Y(n_14510)
);

HB1xp67_ASAP7_75t_L g14511 ( 
.A(n_13421),
.Y(n_14511)
);

INVx1_ASAP7_75t_L g14512 ( 
.A(n_13552),
.Y(n_14512)
);

AND2x2_ASAP7_75t_L g14513 ( 
.A(n_14032),
.B(n_13124),
.Y(n_14513)
);

AND2x4_ASAP7_75t_L g14514 ( 
.A(n_13491),
.B(n_13286),
.Y(n_14514)
);

INVx1_ASAP7_75t_L g14515 ( 
.A(n_13553),
.Y(n_14515)
);

AND2x2_ASAP7_75t_L g14516 ( 
.A(n_14046),
.B(n_13185),
.Y(n_14516)
);

INVx1_ASAP7_75t_L g14517 ( 
.A(n_13556),
.Y(n_14517)
);

NAND2xp5_ASAP7_75t_SL g14518 ( 
.A(n_14044),
.B(n_12880),
.Y(n_14518)
);

NOR2xp33_ASAP7_75t_L g14519 ( 
.A(n_13996),
.B(n_13286),
.Y(n_14519)
);

NAND2xp5_ASAP7_75t_L g14520 ( 
.A(n_13438),
.B(n_13294),
.Y(n_14520)
);

INVx1_ASAP7_75t_L g14521 ( 
.A(n_13562),
.Y(n_14521)
);

INVx3_ASAP7_75t_L g14522 ( 
.A(n_13985),
.Y(n_14522)
);

INVx2_ASAP7_75t_L g14523 ( 
.A(n_13966),
.Y(n_14523)
);

NAND2xp5_ASAP7_75t_L g14524 ( 
.A(n_13994),
.B(n_12938),
.Y(n_14524)
);

OR2x2_ASAP7_75t_L g14525 ( 
.A(n_13767),
.B(n_12824),
.Y(n_14525)
);

NOR2xp33_ASAP7_75t_SL g14526 ( 
.A(n_13654),
.B(n_13079),
.Y(n_14526)
);

AND2x2_ASAP7_75t_L g14527 ( 
.A(n_13345),
.B(n_13197),
.Y(n_14527)
);

AND2x2_ASAP7_75t_L g14528 ( 
.A(n_13919),
.B(n_13198),
.Y(n_14528)
);

AND2x2_ASAP7_75t_L g14529 ( 
.A(n_13967),
.B(n_13199),
.Y(n_14529)
);

HB1xp67_ASAP7_75t_L g14530 ( 
.A(n_13421),
.Y(n_14530)
);

INVx1_ASAP7_75t_L g14531 ( 
.A(n_13563),
.Y(n_14531)
);

AND2x2_ASAP7_75t_L g14532 ( 
.A(n_13976),
.B(n_13206),
.Y(n_14532)
);

AND2x4_ASAP7_75t_L g14533 ( 
.A(n_13571),
.B(n_13186),
.Y(n_14533)
);

OR2x6_ASAP7_75t_L g14534 ( 
.A(n_13980),
.B(n_13055),
.Y(n_14534)
);

AND2x4_ASAP7_75t_L g14535 ( 
.A(n_14043),
.B(n_13250),
.Y(n_14535)
);

NAND2x1p5_ASAP7_75t_L g14536 ( 
.A(n_14056),
.B(n_12905),
.Y(n_14536)
);

AND2x4_ASAP7_75t_L g14537 ( 
.A(n_14062),
.B(n_12827),
.Y(n_14537)
);

INVx1_ASAP7_75t_L g14538 ( 
.A(n_13568),
.Y(n_14538)
);

NAND2xp5_ASAP7_75t_L g14539 ( 
.A(n_14065),
.B(n_12830),
.Y(n_14539)
);

INVx3_ASAP7_75t_L g14540 ( 
.A(n_13985),
.Y(n_14540)
);

NOR2xp33_ASAP7_75t_L g14541 ( 
.A(n_13897),
.B(n_13327),
.Y(n_14541)
);

OR2x2_ASAP7_75t_L g14542 ( 
.A(n_13805),
.B(n_13817),
.Y(n_14542)
);

OR2x2_ASAP7_75t_L g14543 ( 
.A(n_13753),
.B(n_12839),
.Y(n_14543)
);

HB1xp67_ASAP7_75t_L g14544 ( 
.A(n_13878),
.Y(n_14544)
);

AOI22xp33_ASAP7_75t_L g14545 ( 
.A1(n_13756),
.A2(n_13234),
.B1(n_13263),
.B2(n_13258),
.Y(n_14545)
);

INVx3_ASAP7_75t_L g14546 ( 
.A(n_13966),
.Y(n_14546)
);

OR2x2_ASAP7_75t_L g14547 ( 
.A(n_14084),
.B(n_12944),
.Y(n_14547)
);

HB1xp67_ASAP7_75t_L g14548 ( 
.A(n_13489),
.Y(n_14548)
);

AND2x4_ASAP7_75t_L g14549 ( 
.A(n_14070),
.B(n_12905),
.Y(n_14549)
);

OR2x2_ASAP7_75t_L g14550 ( 
.A(n_13762),
.B(n_13151),
.Y(n_14550)
);

INVx1_ASAP7_75t_L g14551 ( 
.A(n_13572),
.Y(n_14551)
);

INVx3_ASAP7_75t_L g14552 ( 
.A(n_13834),
.Y(n_14552)
);

INVx1_ASAP7_75t_L g14553 ( 
.A(n_13576),
.Y(n_14553)
);

INVx2_ASAP7_75t_L g14554 ( 
.A(n_13726),
.Y(n_14554)
);

INVx2_ASAP7_75t_L g14555 ( 
.A(n_13851),
.Y(n_14555)
);

INVx1_ASAP7_75t_L g14556 ( 
.A(n_13577),
.Y(n_14556)
);

NAND2xp5_ASAP7_75t_L g14557 ( 
.A(n_13416),
.B(n_13151),
.Y(n_14557)
);

HB1xp67_ASAP7_75t_L g14558 ( 
.A(n_13640),
.Y(n_14558)
);

INVx2_ASAP7_75t_L g14559 ( 
.A(n_13987),
.Y(n_14559)
);

HB1xp67_ASAP7_75t_L g14560 ( 
.A(n_14011),
.Y(n_14560)
);

INVx1_ASAP7_75t_L g14561 ( 
.A(n_13578),
.Y(n_14561)
);

HB1xp67_ASAP7_75t_L g14562 ( 
.A(n_13509),
.Y(n_14562)
);

AND2x4_ASAP7_75t_L g14563 ( 
.A(n_13432),
.B(n_12920),
.Y(n_14563)
);

BUFx3_ASAP7_75t_L g14564 ( 
.A(n_13809),
.Y(n_14564)
);

NAND2x1_ASAP7_75t_L g14565 ( 
.A(n_13458),
.B(n_13176),
.Y(n_14565)
);

AOI22xp33_ASAP7_75t_L g14566 ( 
.A1(n_13377),
.A2(n_13029),
.B1(n_13027),
.B2(n_13167),
.Y(n_14566)
);

NAND2xp5_ASAP7_75t_L g14567 ( 
.A(n_13759),
.B(n_13153),
.Y(n_14567)
);

AND2x2_ASAP7_75t_L g14568 ( 
.A(n_13988),
.B(n_13341),
.Y(n_14568)
);

AND2x4_ASAP7_75t_L g14569 ( 
.A(n_13436),
.B(n_12920),
.Y(n_14569)
);

BUFx3_ASAP7_75t_L g14570 ( 
.A(n_13776),
.Y(n_14570)
);

INVx2_ASAP7_75t_L g14571 ( 
.A(n_14091),
.Y(n_14571)
);

INVx2_ASAP7_75t_L g14572 ( 
.A(n_13723),
.Y(n_14572)
);

HB1xp67_ASAP7_75t_L g14573 ( 
.A(n_13498),
.Y(n_14573)
);

AO21x2_ASAP7_75t_L g14574 ( 
.A1(n_13441),
.A2(n_13060),
.B(n_13051),
.Y(n_14574)
);

INVx5_ASAP7_75t_L g14575 ( 
.A(n_13698),
.Y(n_14575)
);

AND2x4_ASAP7_75t_L g14576 ( 
.A(n_13783),
.B(n_12929),
.Y(n_14576)
);

BUFx2_ASAP7_75t_L g14577 ( 
.A(n_13540),
.Y(n_14577)
);

OR2x2_ASAP7_75t_L g14578 ( 
.A(n_13547),
.B(n_13153),
.Y(n_14578)
);

HB1xp67_ASAP7_75t_L g14579 ( 
.A(n_13500),
.Y(n_14579)
);

NOR2xp33_ASAP7_75t_L g14580 ( 
.A(n_13812),
.B(n_13085),
.Y(n_14580)
);

INVx2_ASAP7_75t_L g14581 ( 
.A(n_13857),
.Y(n_14581)
);

AND2x4_ASAP7_75t_L g14582 ( 
.A(n_13798),
.B(n_13801),
.Y(n_14582)
);

AND2x2_ASAP7_75t_L g14583 ( 
.A(n_13600),
.B(n_12929),
.Y(n_14583)
);

NAND2xp5_ASAP7_75t_L g14584 ( 
.A(n_13808),
.B(n_13154),
.Y(n_14584)
);

INVx2_ASAP7_75t_L g14585 ( 
.A(n_13857),
.Y(n_14585)
);

INVx1_ASAP7_75t_L g14586 ( 
.A(n_13581),
.Y(n_14586)
);

AND2x2_ASAP7_75t_L g14587 ( 
.A(n_14088),
.B(n_12969),
.Y(n_14587)
);

AND2x2_ASAP7_75t_L g14588 ( 
.A(n_13658),
.B(n_12969),
.Y(n_14588)
);

INVx1_ASAP7_75t_L g14589 ( 
.A(n_13583),
.Y(n_14589)
);

OR2x2_ASAP7_75t_L g14590 ( 
.A(n_13898),
.B(n_13154),
.Y(n_14590)
);

NOR2x1_ASAP7_75t_SL g14591 ( 
.A(n_13612),
.B(n_13131),
.Y(n_14591)
);

INVx3_ASAP7_75t_L g14592 ( 
.A(n_13834),
.Y(n_14592)
);

OAI221xp5_ASAP7_75t_L g14593 ( 
.A1(n_13400),
.A2(n_12795),
.B1(n_13123),
.B2(n_13147),
.C(n_13037),
.Y(n_14593)
);

AOI22xp33_ASAP7_75t_L g14594 ( 
.A1(n_13739),
.A2(n_12984),
.B1(n_13235),
.B2(n_13191),
.Y(n_14594)
);

AND2x2_ASAP7_75t_SL g14595 ( 
.A(n_13381),
.B(n_12984),
.Y(n_14595)
);

INVx1_ASAP7_75t_L g14596 ( 
.A(n_13584),
.Y(n_14596)
);

INVx1_ASAP7_75t_L g14597 ( 
.A(n_13589),
.Y(n_14597)
);

AND2x2_ASAP7_75t_L g14598 ( 
.A(n_13704),
.B(n_13133),
.Y(n_14598)
);

AND2x2_ASAP7_75t_L g14599 ( 
.A(n_13497),
.B(n_13178),
.Y(n_14599)
);

AND2x2_ASAP7_75t_L g14600 ( 
.A(n_13504),
.B(n_13033),
.Y(n_14600)
);

INVx2_ASAP7_75t_L g14601 ( 
.A(n_13869),
.Y(n_14601)
);

AOI221xp5_ASAP7_75t_L g14602 ( 
.A1(n_13506),
.A2(n_13387),
.B1(n_13474),
.B2(n_13406),
.C(n_13795),
.Y(n_14602)
);

INVx1_ASAP7_75t_L g14603 ( 
.A(n_13596),
.Y(n_14603)
);

AND2x2_ASAP7_75t_L g14604 ( 
.A(n_13710),
.B(n_13039),
.Y(n_14604)
);

AND2x2_ASAP7_75t_L g14605 ( 
.A(n_13444),
.B(n_13040),
.Y(n_14605)
);

INVx1_ASAP7_75t_L g14606 ( 
.A(n_13610),
.Y(n_14606)
);

AND2x2_ASAP7_75t_L g14607 ( 
.A(n_13461),
.B(n_13043),
.Y(n_14607)
);

OR2x6_ASAP7_75t_L g14608 ( 
.A(n_14050),
.B(n_13049),
.Y(n_14608)
);

INVx1_ASAP7_75t_L g14609 ( 
.A(n_13611),
.Y(n_14609)
);

INVx2_ASAP7_75t_L g14610 ( 
.A(n_13869),
.Y(n_14610)
);

BUFx6f_ASAP7_75t_L g14611 ( 
.A(n_13698),
.Y(n_14611)
);

BUFx3_ASAP7_75t_L g14612 ( 
.A(n_13609),
.Y(n_14612)
);

INVx1_ASAP7_75t_L g14613 ( 
.A(n_13613),
.Y(n_14613)
);

INVx1_ASAP7_75t_L g14614 ( 
.A(n_13614),
.Y(n_14614)
);

INVx2_ASAP7_75t_L g14615 ( 
.A(n_13874),
.Y(n_14615)
);

AND2x2_ASAP7_75t_L g14616 ( 
.A(n_13466),
.B(n_13515),
.Y(n_14616)
);

AND2x2_ASAP7_75t_L g14617 ( 
.A(n_13516),
.B(n_13052),
.Y(n_14617)
);

INVx1_ASAP7_75t_L g14618 ( 
.A(n_13615),
.Y(n_14618)
);

NAND2xp5_ASAP7_75t_L g14619 ( 
.A(n_13505),
.B(n_13165),
.Y(n_14619)
);

INVx1_ASAP7_75t_L g14620 ( 
.A(n_13616),
.Y(n_14620)
);

BUFx2_ASAP7_75t_L g14621 ( 
.A(n_13540),
.Y(n_14621)
);

AND2x2_ASAP7_75t_L g14622 ( 
.A(n_13521),
.B(n_13173),
.Y(n_14622)
);

AND2x2_ASAP7_75t_L g14623 ( 
.A(n_13417),
.B(n_13176),
.Y(n_14623)
);

INVx1_ASAP7_75t_L g14624 ( 
.A(n_13623),
.Y(n_14624)
);

INVx2_ASAP7_75t_L g14625 ( 
.A(n_13874),
.Y(n_14625)
);

NOR2xp33_ASAP7_75t_L g14626 ( 
.A(n_13882),
.B(n_9875),
.Y(n_14626)
);

INVx2_ASAP7_75t_L g14627 ( 
.A(n_13974),
.Y(n_14627)
);

INVx1_ASAP7_75t_L g14628 ( 
.A(n_13633),
.Y(n_14628)
);

NAND2xp5_ASAP7_75t_L g14629 ( 
.A(n_14051),
.B(n_9879),
.Y(n_14629)
);

OR2x2_ASAP7_75t_L g14630 ( 
.A(n_13894),
.B(n_13051),
.Y(n_14630)
);

BUFx3_ASAP7_75t_L g14631 ( 
.A(n_13396),
.Y(n_14631)
);

NOR2x1_ASAP7_75t_L g14632 ( 
.A(n_13429),
.B(n_13078),
.Y(n_14632)
);

INVx1_ASAP7_75t_L g14633 ( 
.A(n_13648),
.Y(n_14633)
);

INVx1_ASAP7_75t_L g14634 ( 
.A(n_13656),
.Y(n_14634)
);

INVx1_ASAP7_75t_L g14635 ( 
.A(n_13657),
.Y(n_14635)
);

NOR2xp67_ASAP7_75t_L g14636 ( 
.A(n_13574),
.B(n_13078),
.Y(n_14636)
);

OR2x2_ASAP7_75t_L g14637 ( 
.A(n_14034),
.B(n_13054),
.Y(n_14637)
);

HB1xp67_ASAP7_75t_L g14638 ( 
.A(n_13665),
.Y(n_14638)
);

INVx1_ASAP7_75t_L g14639 ( 
.A(n_13662),
.Y(n_14639)
);

INVx1_ASAP7_75t_L g14640 ( 
.A(n_13667),
.Y(n_14640)
);

INVx4_ASAP7_75t_L g14641 ( 
.A(n_13407),
.Y(n_14641)
);

INVx2_ASAP7_75t_L g14642 ( 
.A(n_13974),
.Y(n_14642)
);

INVx2_ASAP7_75t_L g14643 ( 
.A(n_13978),
.Y(n_14643)
);

HB1xp67_ASAP7_75t_L g14644 ( 
.A(n_13535),
.Y(n_14644)
);

INVx1_ASAP7_75t_L g14645 ( 
.A(n_13670),
.Y(n_14645)
);

INVx1_ASAP7_75t_L g14646 ( 
.A(n_13672),
.Y(n_14646)
);

OAI33xp33_ASAP7_75t_L g14647 ( 
.A1(n_13775),
.A2(n_13064),
.A3(n_9795),
.B1(n_9785),
.B2(n_9798),
.B3(n_9788),
.Y(n_14647)
);

AND2x4_ASAP7_75t_L g14648 ( 
.A(n_13414),
.B(n_7663),
.Y(n_14648)
);

INVx1_ASAP7_75t_L g14649 ( 
.A(n_13673),
.Y(n_14649)
);

AND2x2_ASAP7_75t_L g14650 ( 
.A(n_13422),
.B(n_9300),
.Y(n_14650)
);

INVx1_ASAP7_75t_L g14651 ( 
.A(n_13674),
.Y(n_14651)
);

INVx1_ASAP7_75t_L g14652 ( 
.A(n_13679),
.Y(n_14652)
);

INVx1_ASAP7_75t_L g14653 ( 
.A(n_13681),
.Y(n_14653)
);

AND2x4_ASAP7_75t_L g14654 ( 
.A(n_13590),
.B(n_7663),
.Y(n_14654)
);

AND2x2_ASAP7_75t_L g14655 ( 
.A(n_13425),
.B(n_9309),
.Y(n_14655)
);

INVx5_ASAP7_75t_SL g14656 ( 
.A(n_13978),
.Y(n_14656)
);

INVx2_ASAP7_75t_SL g14657 ( 
.A(n_13496),
.Y(n_14657)
);

AND2x2_ASAP7_75t_L g14658 ( 
.A(n_13427),
.B(n_9309),
.Y(n_14658)
);

NAND2xp5_ASAP7_75t_L g14659 ( 
.A(n_13906),
.B(n_13887),
.Y(n_14659)
);

HB1xp67_ASAP7_75t_L g14660 ( 
.A(n_13538),
.Y(n_14660)
);

INVxp67_ASAP7_75t_L g14661 ( 
.A(n_13469),
.Y(n_14661)
);

OAI21xp5_ASAP7_75t_L g14662 ( 
.A1(n_13707),
.A2(n_9218),
.B(n_10178),
.Y(n_14662)
);

OR2x2_ASAP7_75t_L g14663 ( 
.A(n_14036),
.B(n_8411),
.Y(n_14663)
);

BUFx2_ASAP7_75t_L g14664 ( 
.A(n_13850),
.Y(n_14664)
);

AOI22xp5_ASAP7_75t_L g14665 ( 
.A1(n_13627),
.A2(n_8175),
.B1(n_8207),
.B2(n_8168),
.Y(n_14665)
);

INVxp67_ASAP7_75t_SL g14666 ( 
.A(n_13877),
.Y(n_14666)
);

NAND2xp5_ASAP7_75t_L g14667 ( 
.A(n_13911),
.B(n_9879),
.Y(n_14667)
);

INVx2_ASAP7_75t_L g14668 ( 
.A(n_13981),
.Y(n_14668)
);

AND2x2_ASAP7_75t_L g14669 ( 
.A(n_13430),
.B(n_13431),
.Y(n_14669)
);

NOR2x1_ASAP7_75t_SL g14670 ( 
.A(n_13514),
.B(n_8175),
.Y(n_14670)
);

INVx4_ASAP7_75t_L g14671 ( 
.A(n_13981),
.Y(n_14671)
);

NOR2xp33_ASAP7_75t_R g14672 ( 
.A(n_13495),
.B(n_5075),
.Y(n_14672)
);

AND2x2_ASAP7_75t_L g14673 ( 
.A(n_13533),
.B(n_9309),
.Y(n_14673)
);

AND2x2_ASAP7_75t_L g14674 ( 
.A(n_13536),
.B(n_9309),
.Y(n_14674)
);

INVx1_ASAP7_75t_L g14675 ( 
.A(n_13683),
.Y(n_14675)
);

INVx1_ASAP7_75t_L g14676 ( 
.A(n_13686),
.Y(n_14676)
);

NAND2xp5_ASAP7_75t_L g14677 ( 
.A(n_13598),
.B(n_9885),
.Y(n_14677)
);

INVx1_ASAP7_75t_L g14678 ( 
.A(n_13692),
.Y(n_14678)
);

BUFx2_ASAP7_75t_L g14679 ( 
.A(n_13693),
.Y(n_14679)
);

INVx1_ASAP7_75t_L g14680 ( 
.A(n_13694),
.Y(n_14680)
);

INVx1_ASAP7_75t_L g14681 ( 
.A(n_13696),
.Y(n_14681)
);

OR2x6_ASAP7_75t_L g14682 ( 
.A(n_13526),
.B(n_6628),
.Y(n_14682)
);

OA21x2_ASAP7_75t_L g14683 ( 
.A1(n_13907),
.A2(n_10296),
.B(n_10292),
.Y(n_14683)
);

INVx1_ASAP7_75t_L g14684 ( 
.A(n_13713),
.Y(n_14684)
);

AND2x2_ASAP7_75t_L g14685 ( 
.A(n_13632),
.B(n_9318),
.Y(n_14685)
);

OAI21xp5_ASAP7_75t_L g14686 ( 
.A1(n_13631),
.A2(n_9040),
.B(n_9019),
.Y(n_14686)
);

INVx3_ASAP7_75t_L g14687 ( 
.A(n_14072),
.Y(n_14687)
);

INVx2_ASAP7_75t_L g14688 ( 
.A(n_14067),
.Y(n_14688)
);

AND2x2_ASAP7_75t_L g14689 ( 
.A(n_14058),
.B(n_13618),
.Y(n_14689)
);

AND2x2_ASAP7_75t_L g14690 ( 
.A(n_13389),
.B(n_9318),
.Y(n_14690)
);

INVx1_ASAP7_75t_L g14691 ( 
.A(n_13728),
.Y(n_14691)
);

INVx1_ASAP7_75t_L g14692 ( 
.A(n_13734),
.Y(n_14692)
);

INVx1_ASAP7_75t_L g14693 ( 
.A(n_13736),
.Y(n_14693)
);

INVx2_ASAP7_75t_L g14694 ( 
.A(n_13842),
.Y(n_14694)
);

AND2x2_ASAP7_75t_L g14695 ( 
.A(n_13659),
.B(n_9318),
.Y(n_14695)
);

INVx1_ASAP7_75t_L g14696 ( 
.A(n_13742),
.Y(n_14696)
);

INVx1_ASAP7_75t_L g14697 ( 
.A(n_13744),
.Y(n_14697)
);

INVx3_ASAP7_75t_L g14698 ( 
.A(n_14072),
.Y(n_14698)
);

INVx2_ASAP7_75t_L g14699 ( 
.A(n_14092),
.Y(n_14699)
);

AOI222xp33_ASAP7_75t_L g14700 ( 
.A1(n_13449),
.A2(n_9795),
.B1(n_9785),
.B2(n_9798),
.C1(n_9788),
.C2(n_9784),
.Y(n_14700)
);

AND2x2_ASAP7_75t_L g14701 ( 
.A(n_13663),
.B(n_9318),
.Y(n_14701)
);

OR2x2_ASAP7_75t_L g14702 ( 
.A(n_14030),
.B(n_8411),
.Y(n_14702)
);

AOI22xp33_ASAP7_75t_L g14703 ( 
.A1(n_13451),
.A2(n_9930),
.B1(n_9941),
.B2(n_8225),
.Y(n_14703)
);

INVx2_ASAP7_75t_L g14704 ( 
.A(n_14092),
.Y(n_14704)
);

AND2x2_ASAP7_75t_L g14705 ( 
.A(n_13676),
.B(n_9352),
.Y(n_14705)
);

HB1xp67_ASAP7_75t_L g14706 ( 
.A(n_13819),
.Y(n_14706)
);

AO21x2_ASAP7_75t_L g14707 ( 
.A1(n_13452),
.A2(n_10296),
.B(n_10292),
.Y(n_14707)
);

INVx2_ASAP7_75t_L g14708 ( 
.A(n_13727),
.Y(n_14708)
);

INVx1_ASAP7_75t_L g14709 ( 
.A(n_13757),
.Y(n_14709)
);

INVx3_ASAP7_75t_L g14710 ( 
.A(n_13867),
.Y(n_14710)
);

AND2x6_ASAP7_75t_L g14711 ( 
.A(n_13758),
.B(n_8175),
.Y(n_14711)
);

AND2x4_ASAP7_75t_L g14712 ( 
.A(n_13677),
.B(n_7663),
.Y(n_14712)
);

BUFx2_ASAP7_75t_L g14713 ( 
.A(n_13761),
.Y(n_14713)
);

INVx2_ASAP7_75t_L g14714 ( 
.A(n_13824),
.Y(n_14714)
);

INVx2_ASAP7_75t_L g14715 ( 
.A(n_14064),
.Y(n_14715)
);

NAND2xp5_ASAP7_75t_L g14716 ( 
.A(n_13697),
.B(n_9885),
.Y(n_14716)
);

AOI22xp5_ASAP7_75t_L g14717 ( 
.A1(n_13796),
.A2(n_8207),
.B1(n_8618),
.B2(n_8175),
.Y(n_14717)
);

INVx2_ASAP7_75t_L g14718 ( 
.A(n_13938),
.Y(n_14718)
);

INVx2_ASAP7_75t_L g14719 ( 
.A(n_14095),
.Y(n_14719)
);

AND2x2_ASAP7_75t_L g14720 ( 
.A(n_13688),
.B(n_9352),
.Y(n_14720)
);

BUFx2_ASAP7_75t_L g14721 ( 
.A(n_13765),
.Y(n_14721)
);

OR2x2_ASAP7_75t_L g14722 ( 
.A(n_13864),
.B(n_13483),
.Y(n_14722)
);

HB1xp67_ASAP7_75t_L g14723 ( 
.A(n_13822),
.Y(n_14723)
);

OR2x2_ASAP7_75t_L g14724 ( 
.A(n_13719),
.B(n_13861),
.Y(n_14724)
);

INVx2_ASAP7_75t_L g14725 ( 
.A(n_13831),
.Y(n_14725)
);

AND2x2_ASAP7_75t_L g14726 ( 
.A(n_13691),
.B(n_9352),
.Y(n_14726)
);

INVx4_ASAP7_75t_L g14727 ( 
.A(n_13815),
.Y(n_14727)
);

INVx2_ASAP7_75t_L g14728 ( 
.A(n_13791),
.Y(n_14728)
);

INVx1_ASAP7_75t_L g14729 ( 
.A(n_13777),
.Y(n_14729)
);

BUFx3_ASAP7_75t_L g14730 ( 
.A(n_13565),
.Y(n_14730)
);

INVx1_ASAP7_75t_L g14731 ( 
.A(n_13780),
.Y(n_14731)
);

BUFx3_ASAP7_75t_L g14732 ( 
.A(n_13580),
.Y(n_14732)
);

INVx1_ASAP7_75t_L g14733 ( 
.A(n_13785),
.Y(n_14733)
);

BUFx3_ASAP7_75t_L g14734 ( 
.A(n_13585),
.Y(n_14734)
);

INVx1_ASAP7_75t_L g14735 ( 
.A(n_13786),
.Y(n_14735)
);

INVx4_ASAP7_75t_L g14736 ( 
.A(n_13816),
.Y(n_14736)
);

INVx1_ASAP7_75t_L g14737 ( 
.A(n_13789),
.Y(n_14737)
);

INVx1_ASAP7_75t_SL g14738 ( 
.A(n_13586),
.Y(n_14738)
);

INVx1_ASAP7_75t_L g14739 ( 
.A(n_13792),
.Y(n_14739)
);

AND2x2_ASAP7_75t_L g14740 ( 
.A(n_13714),
.B(n_9352),
.Y(n_14740)
);

NOR2xp33_ASAP7_75t_L g14741 ( 
.A(n_13951),
.B(n_9892),
.Y(n_14741)
);

NAND2xp5_ASAP7_75t_L g14742 ( 
.A(n_13889),
.B(n_14093),
.Y(n_14742)
);

INVx2_ASAP7_75t_L g14743 ( 
.A(n_14080),
.Y(n_14743)
);

AND2x2_ASAP7_75t_L g14744 ( 
.A(n_13655),
.B(n_9438),
.Y(n_14744)
);

NAND2xp5_ASAP7_75t_L g14745 ( 
.A(n_13810),
.B(n_9892),
.Y(n_14745)
);

AND2x2_ASAP7_75t_L g14746 ( 
.A(n_13952),
.B(n_9438),
.Y(n_14746)
);

INVx1_ASAP7_75t_L g14747 ( 
.A(n_13799),
.Y(n_14747)
);

INVx2_ASAP7_75t_L g14748 ( 
.A(n_13743),
.Y(n_14748)
);

INVx2_ASAP7_75t_L g14749 ( 
.A(n_13502),
.Y(n_14749)
);

AND2x2_ASAP7_75t_L g14750 ( 
.A(n_13391),
.B(n_9438),
.Y(n_14750)
);

INVx2_ASAP7_75t_L g14751 ( 
.A(n_13502),
.Y(n_14751)
);

INVx1_ASAP7_75t_L g14752 ( 
.A(n_13802),
.Y(n_14752)
);

INVx1_ASAP7_75t_L g14753 ( 
.A(n_13806),
.Y(n_14753)
);

INVxp67_ASAP7_75t_SL g14754 ( 
.A(n_13852),
.Y(n_14754)
);

INVx2_ASAP7_75t_L g14755 ( 
.A(n_14054),
.Y(n_14755)
);

INVx2_ASAP7_75t_L g14756 ( 
.A(n_13458),
.Y(n_14756)
);

INVx2_ASAP7_75t_L g14757 ( 
.A(n_13721),
.Y(n_14757)
);

AND2x4_ASAP7_75t_L g14758 ( 
.A(n_13646),
.B(n_7663),
.Y(n_14758)
);

INVx1_ASAP7_75t_L g14759 ( 
.A(n_13519),
.Y(n_14759)
);

OR2x2_ASAP7_75t_L g14760 ( 
.A(n_14042),
.B(n_8412),
.Y(n_14760)
);

BUFx3_ASAP7_75t_L g14761 ( 
.A(n_13588),
.Y(n_14761)
);

INVx2_ASAP7_75t_L g14762 ( 
.A(n_13946),
.Y(n_14762)
);

INVx1_ASAP7_75t_L g14763 ( 
.A(n_13525),
.Y(n_14763)
);

AND2x2_ASAP7_75t_L g14764 ( 
.A(n_13873),
.B(n_9438),
.Y(n_14764)
);

AND2x2_ASAP7_75t_L g14765 ( 
.A(n_13745),
.B(n_9449),
.Y(n_14765)
);

AND2x4_ASAP7_75t_L g14766 ( 
.A(n_13597),
.B(n_7663),
.Y(n_14766)
);

AND2x2_ASAP7_75t_L g14767 ( 
.A(n_13836),
.B(n_9449),
.Y(n_14767)
);

INVx1_ASAP7_75t_L g14768 ( 
.A(n_13890),
.Y(n_14768)
);

AND2x2_ASAP7_75t_L g14769 ( 
.A(n_13838),
.B(n_9449),
.Y(n_14769)
);

BUFx3_ASAP7_75t_L g14770 ( 
.A(n_13606),
.Y(n_14770)
);

OR2x2_ASAP7_75t_L g14771 ( 
.A(n_13541),
.B(n_8412),
.Y(n_14771)
);

AOI221xp5_ASAP7_75t_L g14772 ( 
.A1(n_13782),
.A2(n_9814),
.B1(n_9816),
.B2(n_9811),
.C(n_9807),
.Y(n_14772)
);

HB1xp67_ASAP7_75t_L g14773 ( 
.A(n_13858),
.Y(n_14773)
);

INVx1_ASAP7_75t_L g14774 ( 
.A(n_13895),
.Y(n_14774)
);

AND2x2_ASAP7_75t_SL g14775 ( 
.A(n_14393),
.B(n_13653),
.Y(n_14775)
);

AND2x4_ASAP7_75t_L g14776 ( 
.A(n_14575),
.B(n_13835),
.Y(n_14776)
);

NAND2xp5_ASAP7_75t_L g14777 ( 
.A(n_14201),
.B(n_13626),
.Y(n_14777)
);

INVx2_ASAP7_75t_L g14778 ( 
.A(n_14575),
.Y(n_14778)
);

OAI22xp5_ASAP7_75t_L g14779 ( 
.A1(n_14455),
.A2(n_14393),
.B1(n_14099),
.B2(n_14421),
.Y(n_14779)
);

AND2x2_ASAP7_75t_L g14780 ( 
.A(n_14107),
.B(n_13875),
.Y(n_14780)
);

NAND2xp5_ASAP7_75t_L g14781 ( 
.A(n_14171),
.B(n_13992),
.Y(n_14781)
);

HB1xp67_ASAP7_75t_L g14782 ( 
.A(n_14560),
.Y(n_14782)
);

AND2x2_ASAP7_75t_L g14783 ( 
.A(n_14243),
.B(n_13771),
.Y(n_14783)
);

INVxp67_ASAP7_75t_SL g14784 ( 
.A(n_14241),
.Y(n_14784)
);

INVx1_ASAP7_75t_L g14785 ( 
.A(n_14275),
.Y(n_14785)
);

INVx2_ASAP7_75t_L g14786 ( 
.A(n_14575),
.Y(n_14786)
);

AND2x4_ASAP7_75t_L g14787 ( 
.A(n_14440),
.B(n_13839),
.Y(n_14787)
);

INVx1_ASAP7_75t_L g14788 ( 
.A(n_14275),
.Y(n_14788)
);

OR2x2_ASAP7_75t_L g14789 ( 
.A(n_14196),
.B(n_13804),
.Y(n_14789)
);

INVx1_ASAP7_75t_L g14790 ( 
.A(n_14140),
.Y(n_14790)
);

INVx2_ASAP7_75t_L g14791 ( 
.A(n_14440),
.Y(n_14791)
);

AND2x4_ASAP7_75t_L g14792 ( 
.A(n_14227),
.B(n_13846),
.Y(n_14792)
);

INVx2_ASAP7_75t_L g14793 ( 
.A(n_14447),
.Y(n_14793)
);

INVx1_ASAP7_75t_L g14794 ( 
.A(n_14137),
.Y(n_14794)
);

NAND2xp5_ASAP7_75t_L g14795 ( 
.A(n_14106),
.B(n_14003),
.Y(n_14795)
);

NOR2xp67_ASAP7_75t_L g14796 ( 
.A(n_14256),
.B(n_13716),
.Y(n_14796)
);

BUFx2_ASAP7_75t_L g14797 ( 
.A(n_14324),
.Y(n_14797)
);

OR2x2_ASAP7_75t_L g14798 ( 
.A(n_14108),
.B(n_13972),
.Y(n_14798)
);

INVx2_ASAP7_75t_L g14799 ( 
.A(n_14447),
.Y(n_14799)
);

AND2x2_ASAP7_75t_L g14800 ( 
.A(n_14282),
.B(n_13755),
.Y(n_14800)
);

NAND2xp5_ASAP7_75t_L g14801 ( 
.A(n_14148),
.B(n_13689),
.Y(n_14801)
);

INVx2_ASAP7_75t_L g14802 ( 
.A(n_14189),
.Y(n_14802)
);

NOR2xp67_ASAP7_75t_L g14803 ( 
.A(n_14497),
.B(n_13559),
.Y(n_14803)
);

INVx2_ASAP7_75t_L g14804 ( 
.A(n_14577),
.Y(n_14804)
);

AND2x2_ASAP7_75t_L g14805 ( 
.A(n_14568),
.B(n_13769),
.Y(n_14805)
);

INVx1_ASAP7_75t_L g14806 ( 
.A(n_14155),
.Y(n_14806)
);

OAI221xp5_ASAP7_75t_SL g14807 ( 
.A1(n_14318),
.A2(n_13608),
.B1(n_13800),
.B2(n_14004),
.C(n_14078),
.Y(n_14807)
);

INVx2_ASAP7_75t_L g14808 ( 
.A(n_14577),
.Y(n_14808)
);

AND2x2_ASAP7_75t_L g14809 ( 
.A(n_14160),
.B(n_13910),
.Y(n_14809)
);

INVxp67_ASAP7_75t_L g14810 ( 
.A(n_14192),
.Y(n_14810)
);

OR2x2_ASAP7_75t_L g14811 ( 
.A(n_14116),
.B(n_13570),
.Y(n_14811)
);

NOR3x1_ASAP7_75t_L g14812 ( 
.A(n_14222),
.B(n_13718),
.C(n_13715),
.Y(n_14812)
);

AND2x2_ASAP7_75t_L g14813 ( 
.A(n_14206),
.B(n_14061),
.Y(n_14813)
);

HB1xp67_ASAP7_75t_L g14814 ( 
.A(n_14621),
.Y(n_14814)
);

NAND2xp5_ASAP7_75t_L g14815 ( 
.A(n_14336),
.B(n_13848),
.Y(n_14815)
);

INVx1_ASAP7_75t_L g14816 ( 
.A(n_14155),
.Y(n_14816)
);

AND2x2_ASAP7_75t_L g14817 ( 
.A(n_14118),
.B(n_13651),
.Y(n_14817)
);

OR2x2_ASAP7_75t_L g14818 ( 
.A(n_14162),
.B(n_13702),
.Y(n_14818)
);

INVx1_ASAP7_75t_L g14819 ( 
.A(n_14621),
.Y(n_14819)
);

NAND2x1_ASAP7_75t_L g14820 ( 
.A(n_14226),
.B(n_13860),
.Y(n_14820)
);

INVx1_ASAP7_75t_L g14821 ( 
.A(n_14181),
.Y(n_14821)
);

NAND2xp5_ASAP7_75t_L g14822 ( 
.A(n_14260),
.B(n_13863),
.Y(n_14822)
);

AND2x2_ASAP7_75t_L g14823 ( 
.A(n_14207),
.B(n_13807),
.Y(n_14823)
);

AND2x2_ASAP7_75t_L g14824 ( 
.A(n_14297),
.B(n_13818),
.Y(n_14824)
);

INVx1_ASAP7_75t_L g14825 ( 
.A(n_14185),
.Y(n_14825)
);

INVx2_ASAP7_75t_L g14826 ( 
.A(n_14565),
.Y(n_14826)
);

NAND2x1p5_ASAP7_75t_L g14827 ( 
.A(n_14128),
.B(n_13868),
.Y(n_14827)
);

INVx1_ASAP7_75t_L g14828 ( 
.A(n_14511),
.Y(n_14828)
);

INVx1_ASAP7_75t_L g14829 ( 
.A(n_14530),
.Y(n_14829)
);

INVx1_ASAP7_75t_L g14830 ( 
.A(n_14441),
.Y(n_14830)
);

NAND2xp5_ASAP7_75t_L g14831 ( 
.A(n_14365),
.B(n_13871),
.Y(n_14831)
);

INVx3_ASAP7_75t_L g14832 ( 
.A(n_14102),
.Y(n_14832)
);

AND2x2_ASAP7_75t_L g14833 ( 
.A(n_14124),
.B(n_13820),
.Y(n_14833)
);

AND2x2_ASAP7_75t_L g14834 ( 
.A(n_14170),
.B(n_13823),
.Y(n_14834)
);

INVx1_ASAP7_75t_L g14835 ( 
.A(n_14445),
.Y(n_14835)
);

NAND2xp5_ASAP7_75t_L g14836 ( 
.A(n_14174),
.B(n_13880),
.Y(n_14836)
);

OR2x2_ASAP7_75t_L g14837 ( 
.A(n_14152),
.B(n_13962),
.Y(n_14837)
);

INVx1_ASAP7_75t_L g14838 ( 
.A(n_14346),
.Y(n_14838)
);

INVx1_ASAP7_75t_L g14839 ( 
.A(n_14679),
.Y(n_14839)
);

INVx1_ASAP7_75t_L g14840 ( 
.A(n_14679),
.Y(n_14840)
);

AND2x2_ASAP7_75t_L g14841 ( 
.A(n_14464),
.B(n_13840),
.Y(n_14841)
);

INVx2_ASAP7_75t_L g14842 ( 
.A(n_14103),
.Y(n_14842)
);

NAND2xp5_ASAP7_75t_L g14843 ( 
.A(n_14303),
.B(n_13884),
.Y(n_14843)
);

AND2x2_ASAP7_75t_L g14844 ( 
.A(n_14248),
.B(n_13891),
.Y(n_14844)
);

INVx1_ASAP7_75t_L g14845 ( 
.A(n_14713),
.Y(n_14845)
);

AOI211xp5_ASAP7_75t_L g14846 ( 
.A1(n_14109),
.A2(n_13931),
.B(n_13961),
.C(n_14059),
.Y(n_14846)
);

OR2x2_ASAP7_75t_L g14847 ( 
.A(n_14098),
.B(n_13872),
.Y(n_14847)
);

AND2x2_ASAP7_75t_L g14848 ( 
.A(n_14299),
.B(n_13893),
.Y(n_14848)
);

AND2x2_ASAP7_75t_L g14849 ( 
.A(n_14164),
.B(n_13896),
.Y(n_14849)
);

OR2x2_ASAP7_75t_L g14850 ( 
.A(n_14197),
.B(n_13909),
.Y(n_14850)
);

INVx1_ASAP7_75t_L g14851 ( 
.A(n_14713),
.Y(n_14851)
);

AND2x2_ASAP7_75t_L g14852 ( 
.A(n_14114),
.B(n_13901),
.Y(n_14852)
);

BUFx3_ASAP7_75t_L g14853 ( 
.A(n_14203),
.Y(n_14853)
);

AND2x2_ASAP7_75t_L g14854 ( 
.A(n_14121),
.B(n_13902),
.Y(n_14854)
);

OR2x2_ASAP7_75t_L g14855 ( 
.A(n_14221),
.B(n_13942),
.Y(n_14855)
);

AND2x2_ASAP7_75t_L g14856 ( 
.A(n_14476),
.B(n_13912),
.Y(n_14856)
);

HB1xp67_ASAP7_75t_L g14857 ( 
.A(n_14134),
.Y(n_14857)
);

AND2x2_ASAP7_75t_L g14858 ( 
.A(n_14262),
.B(n_14233),
.Y(n_14858)
);

AND2x2_ASAP7_75t_L g14859 ( 
.A(n_14183),
.B(n_13914),
.Y(n_14859)
);

INVx4_ASAP7_75t_L g14860 ( 
.A(n_14128),
.Y(n_14860)
);

NAND2xp5_ASAP7_75t_L g14861 ( 
.A(n_14509),
.B(n_13916),
.Y(n_14861)
);

AND2x4_ASAP7_75t_L g14862 ( 
.A(n_14166),
.B(n_13917),
.Y(n_14862)
);

HB1xp67_ASAP7_75t_L g14863 ( 
.A(n_14134),
.Y(n_14863)
);

INVx1_ASAP7_75t_L g14864 ( 
.A(n_14721),
.Y(n_14864)
);

AND2x2_ASAP7_75t_L g14865 ( 
.A(n_14325),
.B(n_13920),
.Y(n_14865)
);

NAND2xp5_ASAP7_75t_L g14866 ( 
.A(n_14123),
.B(n_13921),
.Y(n_14866)
);

AND2x2_ASAP7_75t_L g14867 ( 
.A(n_14229),
.B(n_13923),
.Y(n_14867)
);

INVxp67_ASAP7_75t_SL g14868 ( 
.A(n_14379),
.Y(n_14868)
);

AND2x2_ASAP7_75t_L g14869 ( 
.A(n_14208),
.B(n_13926),
.Y(n_14869)
);

INVx1_ASAP7_75t_L g14870 ( 
.A(n_14721),
.Y(n_14870)
);

INVx2_ASAP7_75t_L g14871 ( 
.A(n_14157),
.Y(n_14871)
);

AND2x2_ASAP7_75t_L g14872 ( 
.A(n_14301),
.B(n_13932),
.Y(n_14872)
);

AND2x2_ASAP7_75t_L g14873 ( 
.A(n_14301),
.B(n_13935),
.Y(n_14873)
);

AND2x2_ASAP7_75t_L g14874 ( 
.A(n_14291),
.B(n_14317),
.Y(n_14874)
);

AND2x2_ASAP7_75t_L g14875 ( 
.A(n_14481),
.B(n_13937),
.Y(n_14875)
);

INVx2_ASAP7_75t_L g14876 ( 
.A(n_14128),
.Y(n_14876)
);

AND2x2_ASAP7_75t_L g14877 ( 
.A(n_14331),
.B(n_13939),
.Y(n_14877)
);

HB1xp67_ASAP7_75t_L g14878 ( 
.A(n_14134),
.Y(n_14878)
);

INVx1_ASAP7_75t_L g14879 ( 
.A(n_14352),
.Y(n_14879)
);

OR2x2_ASAP7_75t_L g14880 ( 
.A(n_14221),
.B(n_14503),
.Y(n_14880)
);

AND2x2_ASAP7_75t_L g14881 ( 
.A(n_14168),
.B(n_13941),
.Y(n_14881)
);

INVx2_ASAP7_75t_L g14882 ( 
.A(n_14497),
.Y(n_14882)
);

AND2x2_ASAP7_75t_L g14883 ( 
.A(n_14101),
.B(n_13949),
.Y(n_14883)
);

INVx1_ASAP7_75t_L g14884 ( 
.A(n_14410),
.Y(n_14884)
);

AND2x2_ASAP7_75t_L g14885 ( 
.A(n_14175),
.B(n_13954),
.Y(n_14885)
);

INVx2_ASAP7_75t_L g14886 ( 
.A(n_14497),
.Y(n_14886)
);

INVx2_ASAP7_75t_L g14887 ( 
.A(n_14611),
.Y(n_14887)
);

AND2x2_ASAP7_75t_L g14888 ( 
.A(n_14419),
.B(n_13956),
.Y(n_14888)
);

INVx1_ASAP7_75t_SL g14889 ( 
.A(n_14271),
.Y(n_14889)
);

NAND2xp5_ASAP7_75t_L g14890 ( 
.A(n_14122),
.B(n_13957),
.Y(n_14890)
);

INVx2_ASAP7_75t_L g14891 ( 
.A(n_14611),
.Y(n_14891)
);

OR2x2_ASAP7_75t_L g14892 ( 
.A(n_14503),
.B(n_13965),
.Y(n_14892)
);

AND2x2_ASAP7_75t_L g14893 ( 
.A(n_14113),
.B(n_13960),
.Y(n_14893)
);

INVx1_ASAP7_75t_L g14894 ( 
.A(n_14274),
.Y(n_14894)
);

AND2x4_ASAP7_75t_L g14895 ( 
.A(n_14477),
.B(n_13963),
.Y(n_14895)
);

AND2x4_ASAP7_75t_L g14896 ( 
.A(n_14431),
.B(n_13964),
.Y(n_14896)
);

INVx1_ASAP7_75t_L g14897 ( 
.A(n_14308),
.Y(n_14897)
);

INVx1_ASAP7_75t_L g14898 ( 
.A(n_14280),
.Y(n_14898)
);

AND2x2_ASAP7_75t_L g14899 ( 
.A(n_14158),
.B(n_13979),
.Y(n_14899)
);

OR2x2_ASAP7_75t_L g14900 ( 
.A(n_14249),
.B(n_13986),
.Y(n_14900)
);

INVx1_ASAP7_75t_L g14901 ( 
.A(n_14126),
.Y(n_14901)
);

NOR2xp33_ASAP7_75t_L g14902 ( 
.A(n_14151),
.B(n_13983),
.Y(n_14902)
);

AND2x2_ASAP7_75t_SL g14903 ( 
.A(n_14316),
.B(n_13991),
.Y(n_14903)
);

NAND2xp33_ASAP7_75t_R g14904 ( 
.A(n_14130),
.B(n_14005),
.Y(n_14904)
);

NOR3xp33_ASAP7_75t_L g14905 ( 
.A(n_14602),
.B(n_14159),
.C(n_14242),
.Y(n_14905)
);

NAND2xp5_ASAP7_75t_L g14906 ( 
.A(n_14167),
.B(n_14008),
.Y(n_14906)
);

HB1xp67_ASAP7_75t_L g14907 ( 
.A(n_14636),
.Y(n_14907)
);

INVx2_ASAP7_75t_SL g14908 ( 
.A(n_14494),
.Y(n_14908)
);

INVx1_ASAP7_75t_L g14909 ( 
.A(n_14127),
.Y(n_14909)
);

INVx2_ASAP7_75t_L g14910 ( 
.A(n_14236),
.Y(n_14910)
);

AND2x2_ASAP7_75t_L g14911 ( 
.A(n_14133),
.B(n_14010),
.Y(n_14911)
);

INVx1_ASAP7_75t_L g14912 ( 
.A(n_14132),
.Y(n_14912)
);

INVx1_ASAP7_75t_L g14913 ( 
.A(n_14141),
.Y(n_14913)
);

AND2x2_ASAP7_75t_L g14914 ( 
.A(n_14367),
.B(n_14012),
.Y(n_14914)
);

HB1xp67_ASAP7_75t_L g14915 ( 
.A(n_14236),
.Y(n_14915)
);

NAND3xp33_ASAP7_75t_L g14916 ( 
.A(n_14261),
.B(n_14024),
.C(n_14020),
.Y(n_14916)
);

INVx1_ASAP7_75t_L g14917 ( 
.A(n_14548),
.Y(n_14917)
);

INVx2_ASAP7_75t_L g14918 ( 
.A(n_14131),
.Y(n_14918)
);

INVx1_ASAP7_75t_L g14919 ( 
.A(n_14558),
.Y(n_14919)
);

INVx1_ASAP7_75t_L g14920 ( 
.A(n_14562),
.Y(n_14920)
);

AND2x2_ASAP7_75t_L g14921 ( 
.A(n_14129),
.B(n_14163),
.Y(n_14921)
);

NAND2xp5_ASAP7_75t_SL g14922 ( 
.A(n_14473),
.B(n_13564),
.Y(n_14922)
);

AND2x2_ASAP7_75t_L g14923 ( 
.A(n_14172),
.B(n_14204),
.Y(n_14923)
);

INVx2_ASAP7_75t_L g14924 ( 
.A(n_14131),
.Y(n_14924)
);

INVx1_ASAP7_75t_L g14925 ( 
.A(n_14573),
.Y(n_14925)
);

AND2x2_ASAP7_75t_L g14926 ( 
.A(n_14245),
.B(n_14018),
.Y(n_14926)
);

AND2x2_ASAP7_75t_L g14927 ( 
.A(n_14139),
.B(n_14023),
.Y(n_14927)
);

AND2x2_ASAP7_75t_L g14928 ( 
.A(n_14200),
.B(n_14474),
.Y(n_14928)
);

INVx1_ASAP7_75t_L g14929 ( 
.A(n_14579),
.Y(n_14929)
);

NOR2xp33_ASAP7_75t_L g14930 ( 
.A(n_14219),
.B(n_14029),
.Y(n_14930)
);

NAND2xp5_ASAP7_75t_L g14931 ( 
.A(n_14240),
.B(n_14035),
.Y(n_14931)
);

AND2x4_ASAP7_75t_SL g14932 ( 
.A(n_14223),
.B(n_14041),
.Y(n_14932)
);

NAND2xp5_ASAP7_75t_L g14933 ( 
.A(n_14254),
.B(n_14045),
.Y(n_14933)
);

NAND2xp5_ASAP7_75t_L g14934 ( 
.A(n_14278),
.B(n_14047),
.Y(n_14934)
);

NAND2xp5_ASAP7_75t_L g14935 ( 
.A(n_14321),
.B(n_14049),
.Y(n_14935)
);

INVx2_ASAP7_75t_L g14936 ( 
.A(n_14656),
.Y(n_14936)
);

NAND2xp5_ASAP7_75t_L g14937 ( 
.A(n_14210),
.B(n_14057),
.Y(n_14937)
);

NAND2x1_ASAP7_75t_L g14938 ( 
.A(n_14226),
.B(n_14071),
.Y(n_14938)
);

NAND2x1p5_ASAP7_75t_L g14939 ( 
.A(n_14491),
.B(n_14077),
.Y(n_14939)
);

AND2x2_ASAP7_75t_L g14940 ( 
.A(n_14362),
.B(n_14086),
.Y(n_14940)
);

INVx1_ASAP7_75t_L g14941 ( 
.A(n_14638),
.Y(n_14941)
);

OR2x2_ASAP7_75t_L g14942 ( 
.A(n_14216),
.B(n_14076),
.Y(n_14942)
);

INVxp67_ASAP7_75t_SL g14943 ( 
.A(n_14238),
.Y(n_14943)
);

NAND2xp5_ASAP7_75t_L g14944 ( 
.A(n_14212),
.B(n_14090),
.Y(n_14944)
);

NAND2xp5_ASAP7_75t_L g14945 ( 
.A(n_14224),
.B(n_13950),
.Y(n_14945)
);

INVx1_ASAP7_75t_L g14946 ( 
.A(n_14644),
.Y(n_14946)
);

OAI21xp5_ASAP7_75t_SL g14947 ( 
.A1(n_14288),
.A2(n_14112),
.B(n_14169),
.Y(n_14947)
);

OR2x2_ASAP7_75t_L g14948 ( 
.A(n_14290),
.B(n_13953),
.Y(n_14948)
);

INVx1_ASAP7_75t_L g14949 ( 
.A(n_14660),
.Y(n_14949)
);

AND2x2_ASAP7_75t_L g14950 ( 
.A(n_14391),
.B(n_13803),
.Y(n_14950)
);

OR2x2_ASAP7_75t_L g14951 ( 
.A(n_14153),
.B(n_13958),
.Y(n_14951)
);

INVx1_ASAP7_75t_L g14952 ( 
.A(n_14213),
.Y(n_14952)
);

CKINVDCx5p33_ASAP7_75t_R g14953 ( 
.A(n_14302),
.Y(n_14953)
);

AND2x2_ASAP7_75t_L g14954 ( 
.A(n_14400),
.B(n_13747),
.Y(n_14954)
);

OR2x2_ASAP7_75t_L g14955 ( 
.A(n_14138),
.B(n_14069),
.Y(n_14955)
);

NAND2xp5_ASAP7_75t_L g14956 ( 
.A(n_14407),
.B(n_13908),
.Y(n_14956)
);

NOR2xp33_ASAP7_75t_R g14957 ( 
.A(n_14198),
.B(n_13918),
.Y(n_14957)
);

INVx1_ASAP7_75t_L g14958 ( 
.A(n_14214),
.Y(n_14958)
);

AND2x2_ASAP7_75t_L g14959 ( 
.A(n_14408),
.B(n_13844),
.Y(n_14959)
);

AND2x2_ASAP7_75t_L g14960 ( 
.A(n_14414),
.B(n_13845),
.Y(n_14960)
);

AND2x4_ASAP7_75t_SL g14961 ( 
.A(n_14146),
.B(n_13847),
.Y(n_14961)
);

AND2x2_ASAP7_75t_L g14962 ( 
.A(n_14417),
.B(n_13982),
.Y(n_14962)
);

NAND2x1p5_ASAP7_75t_L g14963 ( 
.A(n_14436),
.B(n_13934),
.Y(n_14963)
);

INVx1_ASAP7_75t_L g14964 ( 
.A(n_14217),
.Y(n_14964)
);

AND2x2_ASAP7_75t_L g14965 ( 
.A(n_14284),
.B(n_13944),
.Y(n_14965)
);

INVx1_ASAP7_75t_L g14966 ( 
.A(n_14225),
.Y(n_14966)
);

AND2x2_ASAP7_75t_L g14967 ( 
.A(n_14191),
.B(n_14144),
.Y(n_14967)
);

INVx1_ASAP7_75t_L g14968 ( 
.A(n_14234),
.Y(n_14968)
);

AND2x2_ASAP7_75t_SL g14969 ( 
.A(n_14273),
.B(n_14272),
.Y(n_14969)
);

AND2x2_ASAP7_75t_L g14970 ( 
.A(n_14150),
.B(n_14033),
.Y(n_14970)
);

INVx1_ASAP7_75t_L g14971 ( 
.A(n_14544),
.Y(n_14971)
);

INVx2_ASAP7_75t_L g14972 ( 
.A(n_14656),
.Y(n_14972)
);

INVx1_ASAP7_75t_L g14973 ( 
.A(n_14271),
.Y(n_14973)
);

OR2x2_ASAP7_75t_L g14974 ( 
.A(n_14184),
.B(n_13905),
.Y(n_14974)
);

AND2x2_ASAP7_75t_L g14975 ( 
.A(n_14136),
.B(n_14339),
.Y(n_14975)
);

INVx1_ASAP7_75t_L g14976 ( 
.A(n_14115),
.Y(n_14976)
);

AND2x2_ASAP7_75t_L g14977 ( 
.A(n_14344),
.B(n_14039),
.Y(n_14977)
);

INVx2_ASAP7_75t_L g14978 ( 
.A(n_14418),
.Y(n_14978)
);

AND2x2_ASAP7_75t_L g14979 ( 
.A(n_14142),
.B(n_13717),
.Y(n_14979)
);

INVx3_ASAP7_75t_L g14980 ( 
.A(n_14671),
.Y(n_14980)
);

HB1xp67_ASAP7_75t_L g14981 ( 
.A(n_14320),
.Y(n_14981)
);

INVx1_ASAP7_75t_L g14982 ( 
.A(n_14154),
.Y(n_14982)
);

AND2x4_ASAP7_75t_SL g14983 ( 
.A(n_14209),
.B(n_8547),
.Y(n_14983)
);

BUFx2_ASAP7_75t_L g14984 ( 
.A(n_14314),
.Y(n_14984)
);

INVxp33_ASAP7_75t_L g14985 ( 
.A(n_14591),
.Y(n_14985)
);

BUFx3_ASAP7_75t_L g14986 ( 
.A(n_14444),
.Y(n_14986)
);

INVx1_ASAP7_75t_L g14987 ( 
.A(n_14156),
.Y(n_14987)
);

INVx1_ASAP7_75t_L g14988 ( 
.A(n_14187),
.Y(n_14988)
);

AND2x2_ASAP7_75t_L g14989 ( 
.A(n_14480),
.B(n_14048),
.Y(n_14989)
);

HB1xp67_ASAP7_75t_L g14990 ( 
.A(n_14209),
.Y(n_14990)
);

OR2x2_ASAP7_75t_L g14991 ( 
.A(n_14314),
.B(n_13933),
.Y(n_14991)
);

INVx1_ASAP7_75t_L g14992 ( 
.A(n_14496),
.Y(n_14992)
);

NAND2xp5_ASAP7_75t_L g14993 ( 
.A(n_14343),
.B(n_13671),
.Y(n_14993)
);

INVx1_ASAP7_75t_L g14994 ( 
.A(n_14369),
.Y(n_14994)
);

AND2x2_ASAP7_75t_L g14995 ( 
.A(n_14135),
.B(n_9449),
.Y(n_14995)
);

AND2x2_ASAP7_75t_L g14996 ( 
.A(n_14279),
.B(n_9472),
.Y(n_14996)
);

NAND2xp5_ASAP7_75t_L g14997 ( 
.A(n_14354),
.B(n_9894),
.Y(n_14997)
);

OR2x2_ASAP7_75t_L g14998 ( 
.A(n_14177),
.B(n_10304),
.Y(n_14998)
);

AND2x2_ASAP7_75t_L g14999 ( 
.A(n_14514),
.B(n_9472),
.Y(n_14999)
);

INVx1_ASAP7_75t_L g15000 ( 
.A(n_14372),
.Y(n_15000)
);

INVx1_ASAP7_75t_L g15001 ( 
.A(n_14097),
.Y(n_15001)
);

INVx2_ASAP7_75t_L g15002 ( 
.A(n_14218),
.Y(n_15002)
);

INVxp67_ASAP7_75t_SL g15003 ( 
.A(n_14363),
.Y(n_15003)
);

OR2x2_ASAP7_75t_L g15004 ( 
.A(n_14125),
.B(n_14100),
.Y(n_15004)
);

NAND2xp5_ASAP7_75t_L g15005 ( 
.A(n_14263),
.B(n_9894),
.Y(n_15005)
);

NAND2xp5_ASAP7_75t_L g15006 ( 
.A(n_14356),
.B(n_9899),
.Y(n_15006)
);

OR2x2_ASAP7_75t_L g15007 ( 
.A(n_14230),
.B(n_10304),
.Y(n_15007)
);

OAI22xp33_ASAP7_75t_L g15008 ( 
.A1(n_14717),
.A2(n_8207),
.B1(n_8618),
.B2(n_8175),
.Y(n_15008)
);

INVx1_ASAP7_75t_L g15009 ( 
.A(n_14117),
.Y(n_15009)
);

NOR2x1_ASAP7_75t_L g15010 ( 
.A(n_14483),
.B(n_9472),
.Y(n_15010)
);

INVx1_ASAP7_75t_L g15011 ( 
.A(n_14104),
.Y(n_15011)
);

BUFx2_ASAP7_75t_L g15012 ( 
.A(n_14307),
.Y(n_15012)
);

OR2x2_ASAP7_75t_L g15013 ( 
.A(n_14305),
.B(n_10306),
.Y(n_15013)
);

AND2x2_ASAP7_75t_L g15014 ( 
.A(n_14228),
.B(n_9472),
.Y(n_15014)
);

INVx1_ASAP7_75t_L g15015 ( 
.A(n_14211),
.Y(n_15015)
);

AND2x2_ASAP7_75t_L g15016 ( 
.A(n_14361),
.B(n_9665),
.Y(n_15016)
);

HB1xp67_ASAP7_75t_L g15017 ( 
.A(n_14218),
.Y(n_15017)
);

AND2x2_ASAP7_75t_L g15018 ( 
.A(n_14266),
.B(n_9665),
.Y(n_15018)
);

HB1xp67_ASAP7_75t_L g15019 ( 
.A(n_14377),
.Y(n_15019)
);

AND2x4_ASAP7_75t_L g15020 ( 
.A(n_14506),
.B(n_9665),
.Y(n_15020)
);

NAND2xp5_ASAP7_75t_L g15021 ( 
.A(n_14374),
.B(n_9899),
.Y(n_15021)
);

INVx2_ASAP7_75t_L g15022 ( 
.A(n_14329),
.Y(n_15022)
);

INVx1_ASAP7_75t_SL g15023 ( 
.A(n_14542),
.Y(n_15023)
);

INVx2_ASAP7_75t_L g15024 ( 
.A(n_14552),
.Y(n_15024)
);

OR2x2_ASAP7_75t_L g15025 ( 
.A(n_14328),
.B(n_10306),
.Y(n_15025)
);

AND2x2_ASAP7_75t_L g15026 ( 
.A(n_14616),
.B(n_9665),
.Y(n_15026)
);

INVx1_ASAP7_75t_L g15027 ( 
.A(n_14756),
.Y(n_15027)
);

AND2x4_ASAP7_75t_L g15028 ( 
.A(n_14631),
.B(n_9674),
.Y(n_15028)
);

HB1xp67_ASAP7_75t_L g15029 ( 
.A(n_14377),
.Y(n_15029)
);

HB1xp67_ASAP7_75t_L g15030 ( 
.A(n_14706),
.Y(n_15030)
);

INVx2_ASAP7_75t_L g15031 ( 
.A(n_14592),
.Y(n_15031)
);

OR2x2_ASAP7_75t_L g15032 ( 
.A(n_14186),
.B(n_10318),
.Y(n_15032)
);

NAND2xp5_ASAP7_75t_L g15033 ( 
.A(n_14376),
.B(n_9902),
.Y(n_15033)
);

INVx2_ASAP7_75t_L g15034 ( 
.A(n_14522),
.Y(n_15034)
);

INVx1_ASAP7_75t_L g15035 ( 
.A(n_14147),
.Y(n_15035)
);

INVx1_ASAP7_75t_L g15036 ( 
.A(n_14149),
.Y(n_15036)
);

HB1xp67_ASAP7_75t_L g15037 ( 
.A(n_14723),
.Y(n_15037)
);

INVxp67_ASAP7_75t_SL g15038 ( 
.A(n_14276),
.Y(n_15038)
);

AND2x2_ASAP7_75t_L g15039 ( 
.A(n_14669),
.B(n_9674),
.Y(n_15039)
);

NAND2xp5_ASAP7_75t_SL g15040 ( 
.A(n_14202),
.B(n_14268),
.Y(n_15040)
);

AND2x2_ASAP7_75t_L g15041 ( 
.A(n_14312),
.B(n_9674),
.Y(n_15041)
);

NAND2xp5_ASAP7_75t_L g15042 ( 
.A(n_14505),
.B(n_14341),
.Y(n_15042)
);

AND2x2_ASAP7_75t_L g15043 ( 
.A(n_14182),
.B(n_9674),
.Y(n_15043)
);

INVx2_ASAP7_75t_L g15044 ( 
.A(n_14540),
.Y(n_15044)
);

INVx1_ASAP7_75t_L g15045 ( 
.A(n_14287),
.Y(n_15045)
);

AND2x2_ASAP7_75t_L g15046 ( 
.A(n_14195),
.B(n_9685),
.Y(n_15046)
);

INVx1_ASAP7_75t_L g15047 ( 
.A(n_14119),
.Y(n_15047)
);

INVxp67_ASAP7_75t_L g15048 ( 
.A(n_14526),
.Y(n_15048)
);

INVx1_ASAP7_75t_L g15049 ( 
.A(n_14120),
.Y(n_15049)
);

OR2x2_ASAP7_75t_L g15050 ( 
.A(n_14145),
.B(n_10318),
.Y(n_15050)
);

INVx1_ASAP7_75t_L g15051 ( 
.A(n_14239),
.Y(n_15051)
);

INVx1_ASAP7_75t_L g15052 ( 
.A(n_14323),
.Y(n_15052)
);

INVx1_ASAP7_75t_L g15053 ( 
.A(n_14749),
.Y(n_15053)
);

NAND2xp5_ASAP7_75t_L g15054 ( 
.A(n_14413),
.B(n_9902),
.Y(n_15054)
);

AND2x2_ASAP7_75t_L g15055 ( 
.A(n_14258),
.B(n_9685),
.Y(n_15055)
);

AND2x2_ASAP7_75t_L g15056 ( 
.A(n_14220),
.B(n_9685),
.Y(n_15056)
);

AND2x4_ASAP7_75t_L g15057 ( 
.A(n_14612),
.B(n_9685),
.Y(n_15057)
);

INVx1_ASAP7_75t_L g15058 ( 
.A(n_14751),
.Y(n_15058)
);

AND2x2_ASAP7_75t_L g15059 ( 
.A(n_14194),
.B(n_9734),
.Y(n_15059)
);

NAND2xp5_ASAP7_75t_L g15060 ( 
.A(n_14478),
.B(n_9903),
.Y(n_15060)
);

OR2x2_ASAP7_75t_L g15061 ( 
.A(n_14475),
.B(n_10326),
.Y(n_15061)
);

NAND2xp5_ASAP7_75t_L g15062 ( 
.A(n_14179),
.B(n_9903),
.Y(n_15062)
);

INVx1_ASAP7_75t_L g15063 ( 
.A(n_14286),
.Y(n_15063)
);

AND2x2_ASAP7_75t_L g15064 ( 
.A(n_14259),
.B(n_9734),
.Y(n_15064)
);

AND2x4_ASAP7_75t_L g15065 ( 
.A(n_14231),
.B(n_9734),
.Y(n_15065)
);

NAND2xp5_ASAP7_75t_L g15066 ( 
.A(n_14226),
.B(n_9904),
.Y(n_15066)
);

NAND2xp5_ASAP7_75t_L g15067 ( 
.A(n_14357),
.B(n_9904),
.Y(n_15067)
);

NAND2x1_ASAP7_75t_L g15068 ( 
.A(n_14641),
.B(n_9734),
.Y(n_15068)
);

OR2x2_ASAP7_75t_L g15069 ( 
.A(n_14486),
.B(n_10326),
.Y(n_15069)
);

AND2x2_ASAP7_75t_L g15070 ( 
.A(n_14500),
.B(n_9755),
.Y(n_15070)
);

AND2x2_ASAP7_75t_L g15071 ( 
.A(n_14583),
.B(n_14368),
.Y(n_15071)
);

NAND2xp5_ASAP7_75t_L g15072 ( 
.A(n_14357),
.B(n_9911),
.Y(n_15072)
);

NAND2xp5_ASAP7_75t_L g15073 ( 
.A(n_14161),
.B(n_9911),
.Y(n_15073)
);

INVx1_ASAP7_75t_L g15074 ( 
.A(n_14283),
.Y(n_15074)
);

INVx1_ASAP7_75t_L g15075 ( 
.A(n_14425),
.Y(n_15075)
);

AND2x4_ASAP7_75t_L g15076 ( 
.A(n_14105),
.B(n_9755),
.Y(n_15076)
);

INVx2_ASAP7_75t_L g15077 ( 
.A(n_14670),
.Y(n_15077)
);

NAND2x1_ASAP7_75t_SL g15078 ( 
.A(n_14546),
.B(n_9755),
.Y(n_15078)
);

NAND2xp5_ASAP7_75t_L g15079 ( 
.A(n_14479),
.B(n_9917),
.Y(n_15079)
);

INVx2_ASAP7_75t_L g15080 ( 
.A(n_14536),
.Y(n_15080)
);

INVx1_ASAP7_75t_L g15081 ( 
.A(n_14432),
.Y(n_15081)
);

NAND2xp33_ASAP7_75t_SL g15082 ( 
.A(n_14257),
.B(n_6772),
.Y(n_15082)
);

INVx2_ASAP7_75t_L g15083 ( 
.A(n_14366),
.Y(n_15083)
);

INVx2_ASAP7_75t_SL g15084 ( 
.A(n_14687),
.Y(n_15084)
);

NAND2xp5_ASAP7_75t_L g15085 ( 
.A(n_14452),
.B(n_9917),
.Y(n_15085)
);

INVx1_ASAP7_75t_L g15086 ( 
.A(n_14564),
.Y(n_15086)
);

AND2x4_ASAP7_75t_SL g15087 ( 
.A(n_14306),
.B(n_8547),
.Y(n_15087)
);

INVx1_ASAP7_75t_L g15088 ( 
.A(n_14340),
.Y(n_15088)
);

NAND2x1_ASAP7_75t_L g15089 ( 
.A(n_14698),
.B(n_9755),
.Y(n_15089)
);

OAI21xp33_ASAP7_75t_L g15090 ( 
.A1(n_14255),
.A2(n_9019),
.B(n_8962),
.Y(n_15090)
);

OR2x2_ASAP7_75t_L g15091 ( 
.A(n_14659),
.B(n_10330),
.Y(n_15091)
);

AND2x2_ASAP7_75t_L g15092 ( 
.A(n_14689),
.B(n_9761),
.Y(n_15092)
);

AND2x2_ASAP7_75t_L g15093 ( 
.A(n_14349),
.B(n_9761),
.Y(n_15093)
);

NAND2xp5_ASAP7_75t_L g15094 ( 
.A(n_14598),
.B(n_9924),
.Y(n_15094)
);

AND2x4_ASAP7_75t_L g15095 ( 
.A(n_14143),
.B(n_14215),
.Y(n_15095)
);

AND2x2_ASAP7_75t_L g15096 ( 
.A(n_14350),
.B(n_9761),
.Y(n_15096)
);

NAND2xp5_ASAP7_75t_SL g15097 ( 
.A(n_14459),
.B(n_8175),
.Y(n_15097)
);

AND2x4_ASAP7_75t_L g15098 ( 
.A(n_14199),
.B(n_9761),
.Y(n_15098)
);

AND2x2_ASAP7_75t_L g15099 ( 
.A(n_14355),
.B(n_14360),
.Y(n_15099)
);

AND2x2_ASAP7_75t_L g15100 ( 
.A(n_14332),
.B(n_9767),
.Y(n_15100)
);

BUFx2_ASAP7_75t_L g15101 ( 
.A(n_14664),
.Y(n_15101)
);

AND2x4_ASAP7_75t_L g15102 ( 
.A(n_14188),
.B(n_9767),
.Y(n_15102)
);

AND2x4_ASAP7_75t_SL g15103 ( 
.A(n_14313),
.B(n_8547),
.Y(n_15103)
);

INVx2_ASAP7_75t_L g15104 ( 
.A(n_14404),
.Y(n_15104)
);

INVx1_ASAP7_75t_L g15105 ( 
.A(n_14375),
.Y(n_15105)
);

INVx3_ASAP7_75t_L g15106 ( 
.A(n_14300),
.Y(n_15106)
);

AND2x2_ASAP7_75t_L g15107 ( 
.A(n_14396),
.B(n_9767),
.Y(n_15107)
);

INVx1_ASAP7_75t_L g15108 ( 
.A(n_14173),
.Y(n_15108)
);

INVx1_ASAP7_75t_L g15109 ( 
.A(n_14232),
.Y(n_15109)
);

AND2x2_ASAP7_75t_L g15110 ( 
.A(n_14330),
.B(n_14527),
.Y(n_15110)
);

AND2x2_ASAP7_75t_L g15111 ( 
.A(n_14180),
.B(n_9767),
.Y(n_15111)
);

NOR3xp33_ASAP7_75t_L g15112 ( 
.A(n_14541),
.B(n_14442),
.C(n_14661),
.Y(n_15112)
);

INVx3_ASAP7_75t_R g15113 ( 
.A(n_14176),
.Y(n_15113)
);

AND2x2_ASAP7_75t_L g15114 ( 
.A(n_14488),
.B(n_9782),
.Y(n_15114)
);

INVx2_ASAP7_75t_L g15115 ( 
.A(n_14707),
.Y(n_15115)
);

INVx2_ASAP7_75t_L g15116 ( 
.A(n_14430),
.Y(n_15116)
);

AND2x4_ASAP7_75t_SL g15117 ( 
.A(n_14459),
.B(n_8547),
.Y(n_15117)
);

INVx1_ASAP7_75t_L g15118 ( 
.A(n_14237),
.Y(n_15118)
);

NOR2xp67_ASAP7_75t_L g15119 ( 
.A(n_14178),
.B(n_9782),
.Y(n_15119)
);

NOR2xp67_ASAP7_75t_L g15120 ( 
.A(n_14264),
.B(n_9782),
.Y(n_15120)
);

INVx1_ASAP7_75t_L g15121 ( 
.A(n_14386),
.Y(n_15121)
);

INVx2_ASAP7_75t_L g15122 ( 
.A(n_14437),
.Y(n_15122)
);

AND2x2_ASAP7_75t_L g15123 ( 
.A(n_14443),
.B(n_9782),
.Y(n_15123)
);

INVx2_ASAP7_75t_L g15124 ( 
.A(n_14449),
.Y(n_15124)
);

AND2x2_ASAP7_75t_L g15125 ( 
.A(n_14450),
.B(n_9909),
.Y(n_15125)
);

AND2x2_ASAP7_75t_L g15126 ( 
.A(n_14456),
.B(n_9909),
.Y(n_15126)
);

NOR2xp67_ASAP7_75t_L g15127 ( 
.A(n_14265),
.B(n_9909),
.Y(n_15127)
);

INVx1_ASAP7_75t_L g15128 ( 
.A(n_14295),
.Y(n_15128)
);

OR2x2_ASAP7_75t_L g15129 ( 
.A(n_14253),
.B(n_10330),
.Y(n_15129)
);

INVx1_ASAP7_75t_L g15130 ( 
.A(n_14557),
.Y(n_15130)
);

OR2x2_ASAP7_75t_L g15131 ( 
.A(n_14294),
.B(n_10342),
.Y(n_15131)
);

OR2x2_ASAP7_75t_L g15132 ( 
.A(n_14165),
.B(n_14319),
.Y(n_15132)
);

AOI211xp5_ASAP7_75t_L g15133 ( 
.A1(n_14593),
.A2(n_6894),
.B(n_6922),
.C(n_6772),
.Y(n_15133)
);

INVx1_ASAP7_75t_L g15134 ( 
.A(n_14327),
.Y(n_15134)
);

INVx1_ASAP7_75t_L g15135 ( 
.A(n_14632),
.Y(n_15135)
);

AND2x2_ASAP7_75t_L g15136 ( 
.A(n_14457),
.B(n_9909),
.Y(n_15136)
);

AND2x4_ASAP7_75t_L g15137 ( 
.A(n_14110),
.B(n_9918),
.Y(n_15137)
);

HB1xp67_ASAP7_75t_L g15138 ( 
.A(n_14664),
.Y(n_15138)
);

INVx2_ASAP7_75t_L g15139 ( 
.A(n_14467),
.Y(n_15139)
);

AND2x2_ASAP7_75t_L g15140 ( 
.A(n_14461),
.B(n_9918),
.Y(n_15140)
);

NAND2x1_ASAP7_75t_SL g15141 ( 
.A(n_14270),
.B(n_9918),
.Y(n_15141)
);

AND2x2_ASAP7_75t_L g15142 ( 
.A(n_14588),
.B(n_9918),
.Y(n_15142)
);

AND2x2_ASAP7_75t_L g15143 ( 
.A(n_14495),
.B(n_9997),
.Y(n_15143)
);

INVx2_ASAP7_75t_L g15144 ( 
.A(n_14111),
.Y(n_15144)
);

NAND2xp5_ASAP7_75t_L g15145 ( 
.A(n_14205),
.B(n_9924),
.Y(n_15145)
);

INVx1_ASAP7_75t_L g15146 ( 
.A(n_14334),
.Y(n_15146)
);

INVx1_ASAP7_75t_L g15147 ( 
.A(n_14285),
.Y(n_15147)
);

AND2x4_ASAP7_75t_L g15148 ( 
.A(n_14353),
.B(n_14385),
.Y(n_15148)
);

NAND2xp5_ASAP7_75t_L g15149 ( 
.A(n_14096),
.B(n_9997),
.Y(n_15149)
);

NAND2xp5_ASAP7_75t_SL g15150 ( 
.A(n_14468),
.B(n_8175),
.Y(n_15150)
);

AND2x2_ASAP7_75t_L g15151 ( 
.A(n_14532),
.B(n_9997),
.Y(n_15151)
);

AND2x2_ASAP7_75t_L g15152 ( 
.A(n_14528),
.B(n_9997),
.Y(n_15152)
);

INVx1_ASAP7_75t_L g15153 ( 
.A(n_14759),
.Y(n_15153)
);

AND2x4_ASAP7_75t_L g15154 ( 
.A(n_14190),
.B(n_10005),
.Y(n_15154)
);

INVx1_ASAP7_75t_SL g15155 ( 
.A(n_14345),
.Y(n_15155)
);

AND2x2_ASAP7_75t_L g15156 ( 
.A(n_14529),
.B(n_10005),
.Y(n_15156)
);

INVx1_ASAP7_75t_SL g15157 ( 
.A(n_14398),
.Y(n_15157)
);

INVxp67_ASAP7_75t_SL g15158 ( 
.A(n_14519),
.Y(n_15158)
);

AND2x2_ASAP7_75t_L g15159 ( 
.A(n_14429),
.B(n_14485),
.Y(n_15159)
);

INVx1_ASAP7_75t_L g15160 ( 
.A(n_14763),
.Y(n_15160)
);

INVx2_ASAP7_75t_L g15161 ( 
.A(n_14623),
.Y(n_15161)
);

INVx3_ASAP7_75t_L g15162 ( 
.A(n_14468),
.Y(n_15162)
);

NAND2xp5_ASAP7_75t_L g15163 ( 
.A(n_14738),
.B(n_10005),
.Y(n_15163)
);

INVx1_ASAP7_75t_L g15164 ( 
.A(n_14412),
.Y(n_15164)
);

HB1xp67_ASAP7_75t_L g15165 ( 
.A(n_14682),
.Y(n_15165)
);

NOR2x1p5_ASAP7_75t_L g15166 ( 
.A(n_14384),
.B(n_5370),
.Y(n_15166)
);

AND2x2_ASAP7_75t_L g15167 ( 
.A(n_14388),
.B(n_10005),
.Y(n_15167)
);

OR2x2_ASAP7_75t_L g15168 ( 
.A(n_14439),
.B(n_10342),
.Y(n_15168)
);

AND2x4_ASAP7_75t_L g15169 ( 
.A(n_14570),
.B(n_10084),
.Y(n_15169)
);

INVx2_ASAP7_75t_SL g15170 ( 
.A(n_14581),
.Y(n_15170)
);

AND2x2_ASAP7_75t_L g15171 ( 
.A(n_14392),
.B(n_10084),
.Y(n_15171)
);

INVx1_ASAP7_75t_L g15172 ( 
.A(n_14293),
.Y(n_15172)
);

NAND2xp5_ASAP7_75t_L g15173 ( 
.A(n_14347),
.B(n_10084),
.Y(n_15173)
);

NAND2xp5_ASAP7_75t_L g15174 ( 
.A(n_14594),
.B(n_10084),
.Y(n_15174)
);

AND2x2_ASAP7_75t_L g15175 ( 
.A(n_14311),
.B(n_10089),
.Y(n_15175)
);

AND2x2_ASAP7_75t_L g15176 ( 
.A(n_14587),
.B(n_10089),
.Y(n_15176)
);

OR2x2_ASAP7_75t_L g15177 ( 
.A(n_14292),
.B(n_10369),
.Y(n_15177)
);

AND2x6_ASAP7_75t_SL g15178 ( 
.A(n_14534),
.B(n_7769),
.Y(n_15178)
);

AND2x2_ASAP7_75t_L g15179 ( 
.A(n_14387),
.B(n_10089),
.Y(n_15179)
);

INVx2_ASAP7_75t_L g15180 ( 
.A(n_14348),
.Y(n_15180)
);

OR2x2_ASAP7_75t_L g15181 ( 
.A(n_14304),
.B(n_10369),
.Y(n_15181)
);

AND2x2_ASAP7_75t_L g15182 ( 
.A(n_14533),
.B(n_10089),
.Y(n_15182)
);

INVx2_ASAP7_75t_SL g15183 ( 
.A(n_14585),
.Y(n_15183)
);

AND2x4_ASAP7_75t_L g15184 ( 
.A(n_14559),
.B(n_10138),
.Y(n_15184)
);

BUFx3_ASAP7_75t_L g15185 ( 
.A(n_14466),
.Y(n_15185)
);

AND2x2_ASAP7_75t_L g15186 ( 
.A(n_14193),
.B(n_10138),
.Y(n_15186)
);

INVxp33_ASAP7_75t_SL g15187 ( 
.A(n_14364),
.Y(n_15187)
);

AND2x2_ASAP7_75t_L g15188 ( 
.A(n_14507),
.B(n_10138),
.Y(n_15188)
);

OR2x2_ASAP7_75t_L g15189 ( 
.A(n_14724),
.B(n_14322),
.Y(n_15189)
);

INVxp67_ASAP7_75t_L g15190 ( 
.A(n_14390),
.Y(n_15190)
);

AOI22xp33_ASAP7_75t_L g15191 ( 
.A1(n_14235),
.A2(n_9941),
.B1(n_9930),
.B2(n_7823),
.Y(n_15191)
);

AND2x2_ASAP7_75t_L g15192 ( 
.A(n_14510),
.B(n_10138),
.Y(n_15192)
);

INVx1_ASAP7_75t_L g15193 ( 
.A(n_14578),
.Y(n_15193)
);

INVx1_ASAP7_75t_L g15194 ( 
.A(n_14599),
.Y(n_15194)
);

AND2x4_ASAP7_75t_L g15195 ( 
.A(n_14267),
.B(n_10151),
.Y(n_15195)
);

OR2x2_ASAP7_75t_L g15196 ( 
.A(n_14309),
.B(n_10374),
.Y(n_15196)
);

INVx1_ASAP7_75t_L g15197 ( 
.A(n_14622),
.Y(n_15197)
);

INVx1_ASAP7_75t_L g15198 ( 
.A(n_14600),
.Y(n_15198)
);

INVx1_ASAP7_75t_L g15199 ( 
.A(n_14605),
.Y(n_15199)
);

NAND2xp5_ASAP7_75t_L g15200 ( 
.A(n_14351),
.B(n_14358),
.Y(n_15200)
);

AND2x2_ASAP7_75t_L g15201 ( 
.A(n_14371),
.B(n_10151),
.Y(n_15201)
);

NAND2xp5_ASAP7_75t_L g15202 ( 
.A(n_14601),
.B(n_10151),
.Y(n_15202)
);

NAND2xp5_ASAP7_75t_L g15203 ( 
.A(n_14610),
.B(n_10151),
.Y(n_15203)
);

NAND2xp5_ASAP7_75t_L g15204 ( 
.A(n_14615),
.B(n_10205),
.Y(n_15204)
);

INVx2_ASAP7_75t_L g15205 ( 
.A(n_14625),
.Y(n_15205)
);

AND2x2_ASAP7_75t_SL g15206 ( 
.A(n_14595),
.B(n_8291),
.Y(n_15206)
);

INVx2_ASAP7_75t_L g15207 ( 
.A(n_14627),
.Y(n_15207)
);

AND2x2_ASAP7_75t_L g15208 ( 
.A(n_14371),
.B(n_10205),
.Y(n_15208)
);

INVx1_ASAP7_75t_L g15209 ( 
.A(n_14607),
.Y(n_15209)
);

AND2x2_ASAP7_75t_L g15210 ( 
.A(n_14465),
.B(n_10205),
.Y(n_15210)
);

INVx2_ASAP7_75t_L g15211 ( 
.A(n_14642),
.Y(n_15211)
);

NAND2xp5_ASAP7_75t_L g15212 ( 
.A(n_14643),
.B(n_10205),
.Y(n_15212)
);

INVx1_ASAP7_75t_L g15213 ( 
.A(n_14617),
.Y(n_15213)
);

INVx1_ASAP7_75t_L g15214 ( 
.A(n_14567),
.Y(n_15214)
);

NAND2xp5_ASAP7_75t_L g15215 ( 
.A(n_14668),
.B(n_10217),
.Y(n_15215)
);

AND2x2_ASAP7_75t_L g15216 ( 
.A(n_14516),
.B(n_10217),
.Y(n_15216)
);

INVx1_ASAP7_75t_L g15217 ( 
.A(n_14584),
.Y(n_15217)
);

NAND2xp5_ASAP7_75t_L g15218 ( 
.A(n_14566),
.B(n_10217),
.Y(n_15218)
);

OR2x6_ASAP7_75t_L g15219 ( 
.A(n_14534),
.B(n_6628),
.Y(n_15219)
);

INVx2_ASAP7_75t_L g15220 ( 
.A(n_14489),
.Y(n_15220)
);

NAND2xp5_ASAP7_75t_L g15221 ( 
.A(n_14244),
.B(n_10217),
.Y(n_15221)
);

INVx1_ASAP7_75t_L g15222 ( 
.A(n_14289),
.Y(n_15222)
);

OR2x2_ASAP7_75t_L g15223 ( 
.A(n_14310),
.B(n_10374),
.Y(n_15223)
);

NAND2x1p5_ASAP7_75t_L g15224 ( 
.A(n_14338),
.B(n_14727),
.Y(n_15224)
);

HB1xp67_ASAP7_75t_L g15225 ( 
.A(n_14682),
.Y(n_15225)
);

NAND2xp5_ASAP7_75t_L g15226 ( 
.A(n_14247),
.B(n_10288),
.Y(n_15226)
);

INVxp67_ASAP7_75t_SL g15227 ( 
.A(n_14520),
.Y(n_15227)
);

INVx1_ASAP7_75t_L g15228 ( 
.A(n_14296),
.Y(n_15228)
);

INVx1_ASAP7_75t_L g15229 ( 
.A(n_14315),
.Y(n_15229)
);

INVx1_ASAP7_75t_L g15230 ( 
.A(n_14448),
.Y(n_15230)
);

INVx1_ASAP7_75t_SL g15231 ( 
.A(n_14722),
.Y(n_15231)
);

NAND2xp5_ASAP7_75t_L g15232 ( 
.A(n_14250),
.B(n_10288),
.Y(n_15232)
);

INVx1_ASAP7_75t_L g15233 ( 
.A(n_14451),
.Y(n_15233)
);

INVxp67_ASAP7_75t_L g15234 ( 
.A(n_14399),
.Y(n_15234)
);

HB1xp67_ASAP7_75t_L g15235 ( 
.A(n_14608),
.Y(n_15235)
);

NAND2xp5_ASAP7_75t_L g15236 ( 
.A(n_14252),
.B(n_10288),
.Y(n_15236)
);

AND2x2_ASAP7_75t_L g15237 ( 
.A(n_14688),
.B(n_10288),
.Y(n_15237)
);

AND2x4_ASAP7_75t_L g15238 ( 
.A(n_14472),
.B(n_14657),
.Y(n_15238)
);

AND2x2_ASAP7_75t_L g15239 ( 
.A(n_14433),
.B(n_8783),
.Y(n_15239)
);

AND2x2_ASAP7_75t_L g15240 ( 
.A(n_14535),
.B(n_8783),
.Y(n_15240)
);

INVx3_ASAP7_75t_L g15241 ( 
.A(n_14563),
.Y(n_15241)
);

INVx2_ASAP7_75t_L g15242 ( 
.A(n_14492),
.Y(n_15242)
);

INVx1_ASAP7_75t_L g15243 ( 
.A(n_14454),
.Y(n_15243)
);

INVx1_ASAP7_75t_SL g15244 ( 
.A(n_14409),
.Y(n_15244)
);

NAND2xp5_ASAP7_75t_L g15245 ( 
.A(n_14493),
.B(n_9252),
.Y(n_15245)
);

INVx2_ASAP7_75t_L g15246 ( 
.A(n_14502),
.Y(n_15246)
);

OR2x2_ASAP7_75t_L g15247 ( 
.A(n_14619),
.B(n_10377),
.Y(n_15247)
);

INVx1_ASAP7_75t_L g15248 ( 
.A(n_14590),
.Y(n_15248)
);

AND2x2_ASAP7_75t_L g15249 ( 
.A(n_14725),
.B(n_8783),
.Y(n_15249)
);

AND2x4_ASAP7_75t_SL g15250 ( 
.A(n_14569),
.B(n_8861),
.Y(n_15250)
);

AND2x2_ASAP7_75t_L g15251 ( 
.A(n_14513),
.B(n_14471),
.Y(n_15251)
);

NAND2xp5_ASAP7_75t_L g15252 ( 
.A(n_14523),
.B(n_9252),
.Y(n_15252)
);

INVx2_ASAP7_75t_L g15253 ( 
.A(n_14281),
.Y(n_15253)
);

AND2x2_ASAP7_75t_L g15254 ( 
.A(n_14555),
.B(n_8921),
.Y(n_15254)
);

OR2x2_ASAP7_75t_L g15255 ( 
.A(n_14742),
.B(n_10377),
.Y(n_15255)
);

NOR2xp67_ASAP7_75t_L g15256 ( 
.A(n_14736),
.B(n_10385),
.Y(n_15256)
);

AND2x4_ASAP7_75t_L g15257 ( 
.A(n_14571),
.B(n_7720),
.Y(n_15257)
);

HB1xp67_ASAP7_75t_L g15258 ( 
.A(n_14608),
.Y(n_15258)
);

OR2x2_ASAP7_75t_L g15259 ( 
.A(n_14415),
.B(n_10385),
.Y(n_15259)
);

OR2x2_ASAP7_75t_L g15260 ( 
.A(n_14434),
.B(n_10391),
.Y(n_15260)
);

NAND2xp5_ASAP7_75t_L g15261 ( 
.A(n_14582),
.B(n_9263),
.Y(n_15261)
);

AND2x2_ASAP7_75t_L g15262 ( 
.A(n_14537),
.B(n_8921),
.Y(n_15262)
);

INVx1_ASAP7_75t_L g15263 ( 
.A(n_14550),
.Y(n_15263)
);

AND2x2_ASAP7_75t_L g15264 ( 
.A(n_14715),
.B(n_8921),
.Y(n_15264)
);

AND2x4_ASAP7_75t_L g15265 ( 
.A(n_14554),
.B(n_14714),
.Y(n_15265)
);

AND2x2_ASAP7_75t_L g15266 ( 
.A(n_14718),
.B(n_8777),
.Y(n_15266)
);

AND2x2_ASAP7_75t_L g15267 ( 
.A(n_14719),
.B(n_8777),
.Y(n_15267)
);

AND2x2_ASAP7_75t_L g15268 ( 
.A(n_14487),
.B(n_8777),
.Y(n_15268)
);

AND2x2_ASAP7_75t_L g15269 ( 
.A(n_14694),
.B(n_8793),
.Y(n_15269)
);

INVx1_ASAP7_75t_L g15270 ( 
.A(n_14604),
.Y(n_15270)
);

AND2x2_ASAP7_75t_L g15271 ( 
.A(n_14743),
.B(n_8793),
.Y(n_15271)
);

INVx1_ASAP7_75t_L g15272 ( 
.A(n_14326),
.Y(n_15272)
);

BUFx2_ASAP7_75t_L g15273 ( 
.A(n_14463),
.Y(n_15273)
);

NAND2xp5_ASAP7_75t_L g15274 ( 
.A(n_14666),
.B(n_9263),
.Y(n_15274)
);

AND2x2_ASAP7_75t_L g15275 ( 
.A(n_14755),
.B(n_8793),
.Y(n_15275)
);

OR2x2_ASAP7_75t_L g15276 ( 
.A(n_14446),
.B(n_10391),
.Y(n_15276)
);

AND2x2_ASAP7_75t_L g15277 ( 
.A(n_14762),
.B(n_8794),
.Y(n_15277)
);

INVx2_ASAP7_75t_L g15278 ( 
.A(n_14699),
.Y(n_15278)
);

NAND2xp5_ASAP7_75t_L g15279 ( 
.A(n_14704),
.B(n_9265),
.Y(n_15279)
);

AND2x4_ASAP7_75t_L g15280 ( 
.A(n_14730),
.B(n_7755),
.Y(n_15280)
);

INVx2_ASAP7_75t_L g15281 ( 
.A(n_14690),
.Y(n_15281)
);

INVx1_ASAP7_75t_L g15282 ( 
.A(n_14333),
.Y(n_15282)
);

OAI221xp5_ASAP7_75t_SL g15283 ( 
.A1(n_14378),
.A2(n_9814),
.B1(n_9816),
.B2(n_9811),
.C(n_9807),
.Y(n_15283)
);

AND2x2_ASAP7_75t_L g15284 ( 
.A(n_14572),
.B(n_8794),
.Y(n_15284)
);

NAND2xp5_ASAP7_75t_L g15285 ( 
.A(n_14549),
.B(n_9265),
.Y(n_15285)
);

OR2x2_ASAP7_75t_L g15286 ( 
.A(n_14469),
.B(n_10393),
.Y(n_15286)
);

INVx1_ASAP7_75t_L g15287 ( 
.A(n_14335),
.Y(n_15287)
);

OR2x2_ASAP7_75t_L g15288 ( 
.A(n_14543),
.B(n_10393),
.Y(n_15288)
);

INVxp67_ASAP7_75t_L g15289 ( 
.A(n_14518),
.Y(n_15289)
);

NAND2xp5_ASAP7_75t_L g15290 ( 
.A(n_14576),
.B(n_9270),
.Y(n_15290)
);

AND2x2_ASAP7_75t_L g15291 ( 
.A(n_14728),
.B(n_8794),
.Y(n_15291)
);

AND2x2_ASAP7_75t_L g15292 ( 
.A(n_14708),
.B(n_14710),
.Y(n_15292)
);

OR2x2_ASAP7_75t_L g15293 ( 
.A(n_14525),
.B(n_10400),
.Y(n_15293)
);

OR2x2_ASAP7_75t_L g15294 ( 
.A(n_14453),
.B(n_14524),
.Y(n_15294)
);

NOR2xp33_ASAP7_75t_L g15295 ( 
.A(n_14732),
.B(n_8450),
.Y(n_15295)
);

NAND2xp5_ASAP7_75t_L g15296 ( 
.A(n_14754),
.B(n_9270),
.Y(n_15296)
);

OR2x2_ASAP7_75t_L g15297 ( 
.A(n_14547),
.B(n_14501),
.Y(n_15297)
);

OR2x2_ASAP7_75t_L g15298 ( 
.A(n_14771),
.B(n_10400),
.Y(n_15298)
);

INVx2_ASAP7_75t_L g15299 ( 
.A(n_14750),
.Y(n_15299)
);

INVx1_ASAP7_75t_L g15300 ( 
.A(n_14337),
.Y(n_15300)
);

INVx1_ASAP7_75t_SL g15301 ( 
.A(n_14672),
.Y(n_15301)
);

INVx1_ASAP7_75t_L g15302 ( 
.A(n_14342),
.Y(n_15302)
);

AND2x2_ASAP7_75t_L g15303 ( 
.A(n_14748),
.B(n_14757),
.Y(n_15303)
);

NAND2xp5_ASAP7_75t_L g15304 ( 
.A(n_14298),
.B(n_9280),
.Y(n_15304)
);

AND2x2_ASAP7_75t_L g15305 ( 
.A(n_14734),
.B(n_8802),
.Y(n_15305)
);

AND2x2_ASAP7_75t_L g15306 ( 
.A(n_14761),
.B(n_8802),
.Y(n_15306)
);

AND2x2_ASAP7_75t_L g15307 ( 
.A(n_14770),
.B(n_8802),
.Y(n_15307)
);

AND2x2_ASAP7_75t_L g15308 ( 
.A(n_14484),
.B(n_14545),
.Y(n_15308)
);

AND2x2_ASAP7_75t_L g15309 ( 
.A(n_14773),
.B(n_8873),
.Y(n_15309)
);

INVxp67_ASAP7_75t_SL g15310 ( 
.A(n_14630),
.Y(n_15310)
);

AND2x2_ASAP7_75t_L g15311 ( 
.A(n_14470),
.B(n_8873),
.Y(n_15311)
);

AND2x2_ASAP7_75t_L g15312 ( 
.A(n_14648),
.B(n_8873),
.Y(n_15312)
);

AND2x2_ASAP7_75t_L g15313 ( 
.A(n_14654),
.B(n_8874),
.Y(n_15313)
);

AND2x4_ASAP7_75t_L g15314 ( 
.A(n_14359),
.B(n_7755),
.Y(n_15314)
);

OR2x2_ASAP7_75t_L g15315 ( 
.A(n_14539),
.B(n_14702),
.Y(n_15315)
);

INVx2_ASAP7_75t_L g15316 ( 
.A(n_14712),
.Y(n_15316)
);

NAND2xp5_ASAP7_75t_L g15317 ( 
.A(n_14580),
.B(n_9280),
.Y(n_15317)
);

INVx1_ASAP7_75t_L g15318 ( 
.A(n_14370),
.Y(n_15318)
);

AND2x2_ASAP7_75t_L g15319 ( 
.A(n_14758),
.B(n_8874),
.Y(n_15319)
);

NAND2xp5_ASAP7_75t_L g15320 ( 
.A(n_14768),
.B(n_9296),
.Y(n_15320)
);

INVx1_ASAP7_75t_L g15321 ( 
.A(n_14373),
.Y(n_15321)
);

NAND2xp5_ASAP7_75t_L g15322 ( 
.A(n_14774),
.B(n_9296),
.Y(n_15322)
);

INVx2_ASAP7_75t_L g15323 ( 
.A(n_14740),
.Y(n_15323)
);

OR2x2_ASAP7_75t_L g15324 ( 
.A(n_14663),
.B(n_10405),
.Y(n_15324)
);

INVx1_ASAP7_75t_L g15325 ( 
.A(n_14380),
.Y(n_15325)
);

NAND2xp5_ASAP7_75t_L g15326 ( 
.A(n_14741),
.B(n_9297),
.Y(n_15326)
);

AND2x4_ASAP7_75t_L g15327 ( 
.A(n_14381),
.B(n_10570),
.Y(n_15327)
);

AOI22xp33_ASAP7_75t_L g15328 ( 
.A1(n_14686),
.A2(n_9941),
.B1(n_9930),
.B2(n_7823),
.Y(n_15328)
);

INVx2_ASAP7_75t_L g15329 ( 
.A(n_14695),
.Y(n_15329)
);

INVx1_ASAP7_75t_L g15330 ( 
.A(n_14382),
.Y(n_15330)
);

NAND2xp5_ASAP7_75t_L g15331 ( 
.A(n_14626),
.B(n_9297),
.Y(n_15331)
);

AND2x2_ASAP7_75t_L g15332 ( 
.A(n_14766),
.B(n_8874),
.Y(n_15332)
);

INVx4_ASAP7_75t_L g15333 ( 
.A(n_14246),
.Y(n_15333)
);

INVx2_ASAP7_75t_L g15334 ( 
.A(n_14701),
.Y(n_15334)
);

INVx1_ASAP7_75t_SL g15335 ( 
.A(n_14637),
.Y(n_15335)
);

INVx2_ASAP7_75t_L g15336 ( 
.A(n_14705),
.Y(n_15336)
);

HB1xp67_ASAP7_75t_L g15337 ( 
.A(n_14251),
.Y(n_15337)
);

INVx1_ASAP7_75t_L g15338 ( 
.A(n_14383),
.Y(n_15338)
);

AND2x4_ASAP7_75t_L g15339 ( 
.A(n_14389),
.B(n_11118),
.Y(n_15339)
);

OR2x2_ASAP7_75t_L g15340 ( 
.A(n_14760),
.B(n_14677),
.Y(n_15340)
);

AND2x2_ASAP7_75t_L g15341 ( 
.A(n_14746),
.B(n_8879),
.Y(n_15341)
);

INVx2_ASAP7_75t_SL g15342 ( 
.A(n_14720),
.Y(n_15342)
);

INVx1_ASAP7_75t_L g15343 ( 
.A(n_14394),
.Y(n_15343)
);

OR2x2_ASAP7_75t_L g15344 ( 
.A(n_14629),
.B(n_10405),
.Y(n_15344)
);

AND2x2_ASAP7_75t_L g15345 ( 
.A(n_14726),
.B(n_8879),
.Y(n_15345)
);

OR2x2_ASAP7_75t_L g15346 ( 
.A(n_14716),
.B(n_14395),
.Y(n_15346)
);

NAND2x1p5_ASAP7_75t_L g15347 ( 
.A(n_14397),
.B(n_8057),
.Y(n_15347)
);

INVx1_ASAP7_75t_L g15348 ( 
.A(n_14401),
.Y(n_15348)
);

AND2x2_ASAP7_75t_L g15349 ( 
.A(n_14744),
.B(n_8879),
.Y(n_15349)
);

INVx1_ASAP7_75t_L g15350 ( 
.A(n_14402),
.Y(n_15350)
);

INVx1_ASAP7_75t_L g15351 ( 
.A(n_14403),
.Y(n_15351)
);

AND2x4_ASAP7_75t_SL g15352 ( 
.A(n_14405),
.B(n_8861),
.Y(n_15352)
);

INVx2_ASAP7_75t_L g15353 ( 
.A(n_14650),
.Y(n_15353)
);

NAND2xp5_ASAP7_75t_L g15354 ( 
.A(n_14406),
.B(n_9311),
.Y(n_15354)
);

BUFx2_ASAP7_75t_L g15355 ( 
.A(n_14574),
.Y(n_15355)
);

AND2x2_ASAP7_75t_L g15356 ( 
.A(n_14655),
.B(n_8952),
.Y(n_15356)
);

INVx1_ASAP7_75t_L g15357 ( 
.A(n_14411),
.Y(n_15357)
);

INVx1_ASAP7_75t_L g15358 ( 
.A(n_14416),
.Y(n_15358)
);

INVx1_ASAP7_75t_L g15359 ( 
.A(n_14420),
.Y(n_15359)
);

INVx1_ASAP7_75t_L g15360 ( 
.A(n_14422),
.Y(n_15360)
);

INVx1_ASAP7_75t_L g15361 ( 
.A(n_14423),
.Y(n_15361)
);

INVx1_ASAP7_75t_L g15362 ( 
.A(n_14424),
.Y(n_15362)
);

NAND3xp33_ASAP7_75t_L g15363 ( 
.A(n_14683),
.B(n_9941),
.C(n_9930),
.Y(n_15363)
);

AND2x2_ASAP7_75t_L g15364 ( 
.A(n_14658),
.B(n_8952),
.Y(n_15364)
);

INVx2_ASAP7_75t_SL g15365 ( 
.A(n_14673),
.Y(n_15365)
);

INVx2_ASAP7_75t_L g15366 ( 
.A(n_14674),
.Y(n_15366)
);

HB1xp67_ASAP7_75t_L g15367 ( 
.A(n_14269),
.Y(n_15367)
);

INVx2_ASAP7_75t_L g15368 ( 
.A(n_14685),
.Y(n_15368)
);

INVx2_ASAP7_75t_L g15369 ( 
.A(n_14767),
.Y(n_15369)
);

AND2x4_ASAP7_75t_L g15370 ( 
.A(n_14426),
.B(n_7767),
.Y(n_15370)
);

INVx2_ASAP7_75t_L g15371 ( 
.A(n_14769),
.Y(n_15371)
);

INVx2_ASAP7_75t_L g15372 ( 
.A(n_14711),
.Y(n_15372)
);

INVx1_ASAP7_75t_L g15373 ( 
.A(n_14427),
.Y(n_15373)
);

NAND2xp5_ASAP7_75t_L g15374 ( 
.A(n_14428),
.B(n_9311),
.Y(n_15374)
);

INVx2_ASAP7_75t_L g15375 ( 
.A(n_14711),
.Y(n_15375)
);

NAND2xp5_ASAP7_75t_L g15376 ( 
.A(n_14435),
.B(n_9312),
.Y(n_15376)
);

NOR2x1_ASAP7_75t_R g15377 ( 
.A(n_14438),
.B(n_6628),
.Y(n_15377)
);

AND2x2_ASAP7_75t_L g15378 ( 
.A(n_14764),
.B(n_14765),
.Y(n_15378)
);

AND2x4_ASAP7_75t_L g15379 ( 
.A(n_14277),
.B(n_11118),
.Y(n_15379)
);

AND2x4_ASAP7_75t_L g15380 ( 
.A(n_14458),
.B(n_11134),
.Y(n_15380)
);

NAND2xp5_ASAP7_75t_L g15381 ( 
.A(n_14460),
.B(n_9312),
.Y(n_15381)
);

AOI221xp5_ASAP7_75t_L g15382 ( 
.A1(n_14662),
.A2(n_9814),
.B1(n_9816),
.B2(n_9811),
.C(n_9807),
.Y(n_15382)
);

INVx2_ASAP7_75t_L g15383 ( 
.A(n_14711),
.Y(n_15383)
);

OR2x2_ASAP7_75t_L g15384 ( 
.A(n_14667),
.B(n_10411),
.Y(n_15384)
);

INVx1_ASAP7_75t_L g15385 ( 
.A(n_14462),
.Y(n_15385)
);

INVx1_ASAP7_75t_SL g15386 ( 
.A(n_14880),
.Y(n_15386)
);

NOR2xp67_ASAP7_75t_L g15387 ( 
.A(n_14857),
.B(n_14482),
.Y(n_15387)
);

AND2x2_ASAP7_75t_L g15388 ( 
.A(n_14858),
.B(n_14490),
.Y(n_15388)
);

AND2x2_ASAP7_75t_L g15389 ( 
.A(n_14928),
.B(n_14498),
.Y(n_15389)
);

INVx1_ASAP7_75t_L g15390 ( 
.A(n_15355),
.Y(n_15390)
);

INVx2_ASAP7_75t_L g15391 ( 
.A(n_14820),
.Y(n_15391)
);

NOR3xp33_ASAP7_75t_SL g15392 ( 
.A(n_14953),
.B(n_14504),
.C(n_14499),
.Y(n_15392)
);

INVx1_ASAP7_75t_L g15393 ( 
.A(n_15355),
.Y(n_15393)
);

INVx1_ASAP7_75t_L g15394 ( 
.A(n_15273),
.Y(n_15394)
);

INVx2_ASAP7_75t_L g15395 ( 
.A(n_14938),
.Y(n_15395)
);

INVx3_ASAP7_75t_L g15396 ( 
.A(n_15148),
.Y(n_15396)
);

AND2x2_ASAP7_75t_L g15397 ( 
.A(n_15110),
.B(n_14508),
.Y(n_15397)
);

INVx2_ASAP7_75t_L g15398 ( 
.A(n_14860),
.Y(n_15398)
);

NAND2xp5_ASAP7_75t_L g15399 ( 
.A(n_14868),
.B(n_14512),
.Y(n_15399)
);

BUFx3_ASAP7_75t_L g15400 ( 
.A(n_15148),
.Y(n_15400)
);

AND2x2_ASAP7_75t_L g15401 ( 
.A(n_14809),
.B(n_14515),
.Y(n_15401)
);

AND2x4_ASAP7_75t_L g15402 ( 
.A(n_14943),
.B(n_14517),
.Y(n_15402)
);

AND2x2_ASAP7_75t_L g15403 ( 
.A(n_15071),
.B(n_14521),
.Y(n_15403)
);

AND2x2_ASAP7_75t_L g15404 ( 
.A(n_14874),
.B(n_14531),
.Y(n_15404)
);

INVx2_ASAP7_75t_L g15405 ( 
.A(n_15078),
.Y(n_15405)
);

INVx1_ASAP7_75t_L g15406 ( 
.A(n_15273),
.Y(n_15406)
);

OR2x2_ASAP7_75t_L g15407 ( 
.A(n_15012),
.B(n_14745),
.Y(n_15407)
);

AND2x2_ASAP7_75t_L g15408 ( 
.A(n_15159),
.B(n_14538),
.Y(n_15408)
);

NAND2xp5_ASAP7_75t_L g15409 ( 
.A(n_15003),
.B(n_14551),
.Y(n_15409)
);

AND2x2_ASAP7_75t_L g15410 ( 
.A(n_14800),
.B(n_14553),
.Y(n_15410)
);

INVx2_ASAP7_75t_L g15411 ( 
.A(n_14863),
.Y(n_15411)
);

INVx1_ASAP7_75t_SL g15412 ( 
.A(n_14903),
.Y(n_15412)
);

AND2x2_ASAP7_75t_L g15413 ( 
.A(n_15038),
.B(n_14556),
.Y(n_15413)
);

AND2x2_ASAP7_75t_L g15414 ( 
.A(n_15157),
.B(n_14561),
.Y(n_15414)
);

NAND2xp5_ASAP7_75t_L g15415 ( 
.A(n_14810),
.B(n_14586),
.Y(n_15415)
);

INVx1_ASAP7_75t_L g15416 ( 
.A(n_14814),
.Y(n_15416)
);

NAND2xp5_ASAP7_75t_L g15417 ( 
.A(n_14908),
.B(n_14589),
.Y(n_15417)
);

INVxp67_ASAP7_75t_L g15418 ( 
.A(n_14878),
.Y(n_15418)
);

OR2x2_ASAP7_75t_L g15419 ( 
.A(n_15012),
.B(n_14596),
.Y(n_15419)
);

INVx1_ASAP7_75t_L g15420 ( 
.A(n_14782),
.Y(n_15420)
);

INVx1_ASAP7_75t_L g15421 ( 
.A(n_15121),
.Y(n_15421)
);

NAND2xp5_ASAP7_75t_L g15422 ( 
.A(n_14990),
.B(n_14597),
.Y(n_15422)
);

INVx1_ASAP7_75t_L g15423 ( 
.A(n_15108),
.Y(n_15423)
);

INVx1_ASAP7_75t_L g15424 ( 
.A(n_15109),
.Y(n_15424)
);

AND2x2_ASAP7_75t_L g15425 ( 
.A(n_14813),
.B(n_14603),
.Y(n_15425)
);

NOR4xp25_ASAP7_75t_SL g15426 ( 
.A(n_14984),
.B(n_14609),
.C(n_14613),
.D(n_14606),
.Y(n_15426)
);

NAND2xp5_ASAP7_75t_L g15427 ( 
.A(n_15017),
.B(n_14614),
.Y(n_15427)
);

AND2x2_ASAP7_75t_L g15428 ( 
.A(n_14967),
.B(n_14618),
.Y(n_15428)
);

INVx2_ASAP7_75t_L g15429 ( 
.A(n_14827),
.Y(n_15429)
);

INVx1_ASAP7_75t_L g15430 ( 
.A(n_15118),
.Y(n_15430)
);

AND2x2_ASAP7_75t_L g15431 ( 
.A(n_15099),
.B(n_14620),
.Y(n_15431)
);

AND2x4_ASAP7_75t_L g15432 ( 
.A(n_15185),
.B(n_14624),
.Y(n_15432)
);

AND2x2_ASAP7_75t_L g15433 ( 
.A(n_15002),
.B(n_14628),
.Y(n_15433)
);

BUFx3_ASAP7_75t_L g15434 ( 
.A(n_15224),
.Y(n_15434)
);

AND2x2_ASAP7_75t_L g15435 ( 
.A(n_14921),
.B(n_14633),
.Y(n_15435)
);

NAND3xp33_ASAP7_75t_SL g15436 ( 
.A(n_14985),
.B(n_14665),
.C(n_14635),
.Y(n_15436)
);

AND2x2_ASAP7_75t_L g15437 ( 
.A(n_15155),
.B(n_14634),
.Y(n_15437)
);

INVxp67_ASAP7_75t_L g15438 ( 
.A(n_15030),
.Y(n_15438)
);

NAND2xp5_ASAP7_75t_L g15439 ( 
.A(n_14889),
.B(n_14639),
.Y(n_15439)
);

OAI33xp33_ASAP7_75t_L g15440 ( 
.A1(n_14779),
.A2(n_14649),
.A3(n_14645),
.B1(n_14651),
.B2(n_14646),
.B3(n_14640),
.Y(n_15440)
);

INVx3_ASAP7_75t_L g15441 ( 
.A(n_14986),
.Y(n_15441)
);

HB1xp67_ASAP7_75t_L g15442 ( 
.A(n_14803),
.Y(n_15442)
);

INVx1_ASAP7_75t_L g15443 ( 
.A(n_15037),
.Y(n_15443)
);

NAND2xp5_ASAP7_75t_L g15444 ( 
.A(n_14915),
.B(n_14652),
.Y(n_15444)
);

INVx1_ASAP7_75t_L g15445 ( 
.A(n_15101),
.Y(n_15445)
);

AND2x2_ASAP7_75t_L g15446 ( 
.A(n_14923),
.B(n_14653),
.Y(n_15446)
);

AND2x2_ASAP7_75t_L g15447 ( 
.A(n_14832),
.B(n_14675),
.Y(n_15447)
);

AND2x4_ASAP7_75t_SL g15448 ( 
.A(n_15238),
.B(n_15241),
.Y(n_15448)
);

INVx1_ASAP7_75t_L g15449 ( 
.A(n_15101),
.Y(n_15449)
);

HB1xp67_ASAP7_75t_L g15450 ( 
.A(n_14796),
.Y(n_15450)
);

AND2x2_ASAP7_75t_L g15451 ( 
.A(n_14783),
.B(n_14676),
.Y(n_15451)
);

OR2x2_ASAP7_75t_L g15452 ( 
.A(n_14855),
.B(n_14678),
.Y(n_15452)
);

AND2x2_ASAP7_75t_L g15453 ( 
.A(n_14910),
.B(n_14680),
.Y(n_15453)
);

CKINVDCx5p33_ASAP7_75t_R g15454 ( 
.A(n_14904),
.Y(n_15454)
);

AND2x4_ASAP7_75t_L g15455 ( 
.A(n_14853),
.B(n_14681),
.Y(n_15455)
);

INVx1_ASAP7_75t_L g15456 ( 
.A(n_14907),
.Y(n_15456)
);

INVx1_ASAP7_75t_L g15457 ( 
.A(n_14784),
.Y(n_15457)
);

AND2x2_ASAP7_75t_L g15458 ( 
.A(n_14980),
.B(n_14684),
.Y(n_15458)
);

INVx1_ASAP7_75t_L g15459 ( 
.A(n_14984),
.Y(n_15459)
);

AOI22xp5_ASAP7_75t_L g15460 ( 
.A1(n_14905),
.A2(n_14683),
.B1(n_14692),
.B2(n_14691),
.Y(n_15460)
);

INVx2_ASAP7_75t_L g15461 ( 
.A(n_15141),
.Y(n_15461)
);

OR2x2_ASAP7_75t_L g15462 ( 
.A(n_14892),
.B(n_14693),
.Y(n_15462)
);

AND2x2_ASAP7_75t_L g15463 ( 
.A(n_14823),
.B(n_14936),
.Y(n_15463)
);

AND2x2_ASAP7_75t_L g15464 ( 
.A(n_14972),
.B(n_14805),
.Y(n_15464)
);

INVx1_ASAP7_75t_L g15465 ( 
.A(n_14797),
.Y(n_15465)
);

AOI22xp33_ASAP7_75t_L g15466 ( 
.A1(n_15112),
.A2(n_14647),
.B1(n_14703),
.B2(n_14697),
.Y(n_15466)
);

INVx2_ASAP7_75t_L g15467 ( 
.A(n_14787),
.Y(n_15467)
);

NAND2x1_ASAP7_75t_L g15468 ( 
.A(n_14787),
.B(n_14696),
.Y(n_15468)
);

AND2x2_ASAP7_75t_L g15469 ( 
.A(n_14841),
.B(n_14709),
.Y(n_15469)
);

INVxp67_ASAP7_75t_SL g15470 ( 
.A(n_15138),
.Y(n_15470)
);

AND2x2_ASAP7_75t_L g15471 ( 
.A(n_14867),
.B(n_14729),
.Y(n_15471)
);

INVx1_ASAP7_75t_L g15472 ( 
.A(n_14797),
.Y(n_15472)
);

AND2x2_ASAP7_75t_L g15473 ( 
.A(n_14844),
.B(n_14731),
.Y(n_15473)
);

AND2x2_ASAP7_75t_L g15474 ( 
.A(n_14817),
.B(n_14733),
.Y(n_15474)
);

NAND2xp5_ASAP7_75t_L g15475 ( 
.A(n_14969),
.B(n_14735),
.Y(n_15475)
);

AND2x2_ASAP7_75t_L g15476 ( 
.A(n_14834),
.B(n_14737),
.Y(n_15476)
);

INVx1_ASAP7_75t_L g15477 ( 
.A(n_14785),
.Y(n_15477)
);

INVx2_ASAP7_75t_SL g15478 ( 
.A(n_14791),
.Y(n_15478)
);

INVx1_ASAP7_75t_L g15479 ( 
.A(n_14788),
.Y(n_15479)
);

NOR2xp33_ASAP7_75t_L g15480 ( 
.A(n_15187),
.B(n_14739),
.Y(n_15480)
);

INVxp33_ASAP7_75t_SL g15481 ( 
.A(n_15019),
.Y(n_15481)
);

INVx1_ASAP7_75t_L g15482 ( 
.A(n_14981),
.Y(n_15482)
);

AND2x2_ASAP7_75t_SL g15483 ( 
.A(n_14775),
.B(n_14747),
.Y(n_15483)
);

INVx1_ASAP7_75t_L g15484 ( 
.A(n_14793),
.Y(n_15484)
);

OR2x2_ASAP7_75t_L g15485 ( 
.A(n_15023),
.B(n_14752),
.Y(n_15485)
);

NAND2xp5_ASAP7_75t_L g15486 ( 
.A(n_15235),
.B(n_14753),
.Y(n_15486)
);

NAND4xp25_ASAP7_75t_SL g15487 ( 
.A(n_15133),
.B(n_14772),
.C(n_14700),
.D(n_9820),
.Y(n_15487)
);

NAND2xp5_ASAP7_75t_L g15488 ( 
.A(n_15258),
.B(n_10411),
.Y(n_15488)
);

INVx1_ASAP7_75t_L g15489 ( 
.A(n_14799),
.Y(n_15489)
);

HB1xp67_ASAP7_75t_L g15490 ( 
.A(n_14804),
.Y(n_15490)
);

NAND2xp5_ASAP7_75t_SL g15491 ( 
.A(n_15206),
.B(n_8175),
.Y(n_15491)
);

AND2x2_ASAP7_75t_L g15492 ( 
.A(n_14833),
.B(n_14780),
.Y(n_15492)
);

OR2x2_ASAP7_75t_L g15493 ( 
.A(n_14808),
.B(n_10412),
.Y(n_15493)
);

OR2x2_ASAP7_75t_L g15494 ( 
.A(n_15042),
.B(n_10412),
.Y(n_15494)
);

OR2x2_ASAP7_75t_L g15495 ( 
.A(n_14794),
.B(n_10421),
.Y(n_15495)
);

INVx1_ASAP7_75t_L g15496 ( 
.A(n_14819),
.Y(n_15496)
);

INVx1_ASAP7_75t_L g15497 ( 
.A(n_14806),
.Y(n_15497)
);

NAND2xp5_ASAP7_75t_L g15498 ( 
.A(n_15084),
.B(n_10421),
.Y(n_15498)
);

AND2x4_ASAP7_75t_L g15499 ( 
.A(n_14978),
.B(n_15022),
.Y(n_15499)
);

NAND2xp5_ASAP7_75t_L g15500 ( 
.A(n_14821),
.B(n_10423),
.Y(n_15500)
);

HB1xp67_ASAP7_75t_L g15501 ( 
.A(n_14839),
.Y(n_15501)
);

NAND2xp5_ASAP7_75t_L g15502 ( 
.A(n_14825),
.B(n_10423),
.Y(n_15502)
);

AND2x2_ASAP7_75t_L g15503 ( 
.A(n_14848),
.B(n_8952),
.Y(n_15503)
);

INVx1_ASAP7_75t_L g15504 ( 
.A(n_14816),
.Y(n_15504)
);

INVxp67_ASAP7_75t_L g15505 ( 
.A(n_15029),
.Y(n_15505)
);

NAND2xp5_ASAP7_75t_L g15506 ( 
.A(n_14842),
.B(n_10433),
.Y(n_15506)
);

AND2x4_ASAP7_75t_SL g15507 ( 
.A(n_15106),
.B(n_8861),
.Y(n_15507)
);

INVx1_ASAP7_75t_SL g15508 ( 
.A(n_14900),
.Y(n_15508)
);

INVx2_ASAP7_75t_L g15509 ( 
.A(n_14776),
.Y(n_15509)
);

AND2x2_ASAP7_75t_L g15510 ( 
.A(n_15083),
.B(n_10433),
.Y(n_15510)
);

NOR2xp33_ASAP7_75t_L g15511 ( 
.A(n_15048),
.B(n_10440),
.Y(n_15511)
);

OR2x2_ASAP7_75t_L g15512 ( 
.A(n_15231),
.B(n_10440),
.Y(n_15512)
);

INVx1_ASAP7_75t_L g15513 ( 
.A(n_14840),
.Y(n_15513)
);

INVx1_ASAP7_75t_L g15514 ( 
.A(n_14845),
.Y(n_15514)
);

NAND2xp5_ASAP7_75t_L g15515 ( 
.A(n_14871),
.B(n_10443),
.Y(n_15515)
);

NOR2xp33_ASAP7_75t_SL g15516 ( 
.A(n_15244),
.B(n_6772),
.Y(n_15516)
);

AND2x2_ASAP7_75t_L g15517 ( 
.A(n_15104),
.B(n_10443),
.Y(n_15517)
);

INVx1_ASAP7_75t_L g15518 ( 
.A(n_14851),
.Y(n_15518)
);

NAND2xp5_ASAP7_75t_L g15519 ( 
.A(n_14830),
.B(n_10449),
.Y(n_15519)
);

INVx1_ASAP7_75t_L g15520 ( 
.A(n_14864),
.Y(n_15520)
);

AND2x2_ASAP7_75t_L g15521 ( 
.A(n_14849),
.B(n_10449),
.Y(n_15521)
);

NAND2xp5_ASAP7_75t_L g15522 ( 
.A(n_14835),
.B(n_10461),
.Y(n_15522)
);

HB1xp67_ASAP7_75t_L g15523 ( 
.A(n_14870),
.Y(n_15523)
);

INVxp67_ASAP7_75t_SL g15524 ( 
.A(n_14922),
.Y(n_15524)
);

INVx2_ASAP7_75t_L g15525 ( 
.A(n_14776),
.Y(n_15525)
);

INVx2_ASAP7_75t_L g15526 ( 
.A(n_14778),
.Y(n_15526)
);

AND2x4_ASAP7_75t_L g15527 ( 
.A(n_15161),
.B(n_7767),
.Y(n_15527)
);

INVx1_ASAP7_75t_L g15528 ( 
.A(n_14973),
.Y(n_15528)
);

INVx1_ASAP7_75t_L g15529 ( 
.A(n_14843),
.Y(n_15529)
);

INVx4_ASAP7_75t_L g15530 ( 
.A(n_15162),
.Y(n_15530)
);

AND2x2_ASAP7_75t_L g15531 ( 
.A(n_14975),
.B(n_15251),
.Y(n_15531)
);

HB1xp67_ASAP7_75t_L g15532 ( 
.A(n_14882),
.Y(n_15532)
);

NAND2xp5_ASAP7_75t_L g15533 ( 
.A(n_15170),
.B(n_10461),
.Y(n_15533)
);

AND2x2_ASAP7_75t_L g15534 ( 
.A(n_14824),
.B(n_10479),
.Y(n_15534)
);

AND2x2_ASAP7_75t_L g15535 ( 
.A(n_14869),
.B(n_10479),
.Y(n_15535)
);

CKINVDCx16_ASAP7_75t_R g15536 ( 
.A(n_15189),
.Y(n_15536)
);

AND2x2_ASAP7_75t_L g15537 ( 
.A(n_14918),
.B(n_10491),
.Y(n_15537)
);

INVx1_ASAP7_75t_L g15538 ( 
.A(n_14828),
.Y(n_15538)
);

OR2x2_ASAP7_75t_L g15539 ( 
.A(n_15183),
.B(n_10491),
.Y(n_15539)
);

OR2x2_ASAP7_75t_L g15540 ( 
.A(n_14894),
.B(n_14897),
.Y(n_15540)
);

AND2x2_ASAP7_75t_L g15541 ( 
.A(n_14924),
.B(n_10492),
.Y(n_15541)
);

INVx2_ASAP7_75t_L g15542 ( 
.A(n_14786),
.Y(n_15542)
);

INVx2_ASAP7_75t_L g15543 ( 
.A(n_14886),
.Y(n_15543)
);

AND2x2_ASAP7_75t_L g15544 ( 
.A(n_14875),
.B(n_10492),
.Y(n_15544)
);

INVx1_ASAP7_75t_L g15545 ( 
.A(n_14829),
.Y(n_15545)
);

BUFx2_ASAP7_75t_L g15546 ( 
.A(n_15135),
.Y(n_15546)
);

AND2x2_ASAP7_75t_L g15547 ( 
.A(n_14856),
.B(n_10493),
.Y(n_15547)
);

NAND2xp5_ASAP7_75t_SL g15548 ( 
.A(n_14862),
.B(n_8207),
.Y(n_15548)
);

OR2x2_ASAP7_75t_L g15549 ( 
.A(n_14879),
.B(n_10493),
.Y(n_15549)
);

AND2x2_ASAP7_75t_L g15550 ( 
.A(n_15289),
.B(n_10500),
.Y(n_15550)
);

OR2x2_ASAP7_75t_L g15551 ( 
.A(n_14811),
.B(n_14789),
.Y(n_15551)
);

INVx1_ASAP7_75t_L g15552 ( 
.A(n_14790),
.Y(n_15552)
);

AND2x2_ASAP7_75t_L g15553 ( 
.A(n_14961),
.B(n_10500),
.Y(n_15553)
);

OR2x2_ASAP7_75t_L g15554 ( 
.A(n_15200),
.B(n_14837),
.Y(n_15554)
);

INVx1_ASAP7_75t_SL g15555 ( 
.A(n_15132),
.Y(n_15555)
);

INVx1_ASAP7_75t_L g15556 ( 
.A(n_14884),
.Y(n_15556)
);

INVx2_ASAP7_75t_L g15557 ( 
.A(n_14963),
.Y(n_15557)
);

INVx1_ASAP7_75t_L g15558 ( 
.A(n_15337),
.Y(n_15558)
);

INVx3_ASAP7_75t_L g15559 ( 
.A(n_14792),
.Y(n_15559)
);

AND2x2_ASAP7_75t_L g15560 ( 
.A(n_14899),
.B(n_10504),
.Y(n_15560)
);

NOR2xp33_ASAP7_75t_L g15561 ( 
.A(n_14802),
.B(n_10504),
.Y(n_15561)
);

NAND2xp5_ASAP7_75t_L g15562 ( 
.A(n_15194),
.B(n_10506),
.Y(n_15562)
);

AND2x2_ASAP7_75t_L g15563 ( 
.A(n_14854),
.B(n_10506),
.Y(n_15563)
);

AND2x2_ASAP7_75t_L g15564 ( 
.A(n_14927),
.B(n_10508),
.Y(n_15564)
);

AND2x2_ASAP7_75t_L g15565 ( 
.A(n_14926),
.B(n_15024),
.Y(n_15565)
);

AND2x2_ASAP7_75t_L g15566 ( 
.A(n_15031),
.B(n_10508),
.Y(n_15566)
);

NAND2xp5_ASAP7_75t_L g15567 ( 
.A(n_15197),
.B(n_10515),
.Y(n_15567)
);

AND2x2_ASAP7_75t_L g15568 ( 
.A(n_15034),
.B(n_10515),
.Y(n_15568)
);

OR2x2_ASAP7_75t_L g15569 ( 
.A(n_14795),
.B(n_10516),
.Y(n_15569)
);

OR2x2_ASAP7_75t_L g15570 ( 
.A(n_14917),
.B(n_10516),
.Y(n_15570)
);

OR2x2_ASAP7_75t_L g15571 ( 
.A(n_14919),
.B(n_14920),
.Y(n_15571)
);

INVx1_ASAP7_75t_SL g15572 ( 
.A(n_14942),
.Y(n_15572)
);

AND2x2_ASAP7_75t_L g15573 ( 
.A(n_15044),
.B(n_10532),
.Y(n_15573)
);

INVx3_ASAP7_75t_SL g15574 ( 
.A(n_14932),
.Y(n_15574)
);

INVx2_ASAP7_75t_SL g15575 ( 
.A(n_14826),
.Y(n_15575)
);

NAND2xp5_ASAP7_75t_L g15576 ( 
.A(n_14925),
.B(n_10532),
.Y(n_15576)
);

INVx1_ASAP7_75t_L g15577 ( 
.A(n_15367),
.Y(n_15577)
);

AND2x2_ASAP7_75t_L g15578 ( 
.A(n_14859),
.B(n_10557),
.Y(n_15578)
);

INVx2_ASAP7_75t_L g15579 ( 
.A(n_15010),
.Y(n_15579)
);

OR2x2_ASAP7_75t_L g15580 ( 
.A(n_14929),
.B(n_10557),
.Y(n_15580)
);

OR2x2_ASAP7_75t_L g15581 ( 
.A(n_14941),
.B(n_10563),
.Y(n_15581)
);

NAND2xp5_ASAP7_75t_L g15582 ( 
.A(n_14946),
.B(n_10563),
.Y(n_15582)
);

AND2x2_ASAP7_75t_L g15583 ( 
.A(n_14888),
.B(n_10568),
.Y(n_15583)
);

AND2x4_ASAP7_75t_L g15584 ( 
.A(n_15080),
.B(n_7845),
.Y(n_15584)
);

INVx2_ASAP7_75t_SL g15585 ( 
.A(n_14983),
.Y(n_15585)
);

NAND4xp25_ASAP7_75t_L g15586 ( 
.A(n_14846),
.B(n_8690),
.C(n_8634),
.D(n_6662),
.Y(n_15586)
);

OR2x2_ASAP7_75t_L g15587 ( 
.A(n_14949),
.B(n_10568),
.Y(n_15587)
);

INVx1_ASAP7_75t_L g15588 ( 
.A(n_14992),
.Y(n_15588)
);

NAND3xp33_ASAP7_75t_L g15589 ( 
.A(n_14947),
.B(n_10972),
.C(n_10668),
.Y(n_15589)
);

INVx1_ASAP7_75t_L g15590 ( 
.A(n_14893),
.Y(n_15590)
);

AND2x2_ASAP7_75t_L g15591 ( 
.A(n_14865),
.B(n_10579),
.Y(n_15591)
);

AND2x4_ASAP7_75t_L g15592 ( 
.A(n_14881),
.B(n_7845),
.Y(n_15592)
);

INVx1_ASAP7_75t_L g15593 ( 
.A(n_14885),
.Y(n_15593)
);

BUFx2_ASAP7_75t_L g15594 ( 
.A(n_15115),
.Y(n_15594)
);

AND2x2_ASAP7_75t_L g15595 ( 
.A(n_14911),
.B(n_10579),
.Y(n_15595)
);

OAI21xp5_ASAP7_75t_L g15596 ( 
.A1(n_14916),
.A2(n_11169),
.B(n_11134),
.Y(n_15596)
);

AND2x2_ASAP7_75t_L g15597 ( 
.A(n_14872),
.B(n_10588),
.Y(n_15597)
);

AND2x2_ASAP7_75t_L g15598 ( 
.A(n_14873),
.B(n_10588),
.Y(n_15598)
);

OR2x2_ASAP7_75t_L g15599 ( 
.A(n_15144),
.B(n_10591),
.Y(n_15599)
);

INVxp67_ASAP7_75t_L g15600 ( 
.A(n_15377),
.Y(n_15600)
);

AND2x2_ASAP7_75t_L g15601 ( 
.A(n_14954),
.B(n_10591),
.Y(n_15601)
);

INVx1_ASAP7_75t_L g15602 ( 
.A(n_14831),
.Y(n_15602)
);

AND2x2_ASAP7_75t_L g15603 ( 
.A(n_15292),
.B(n_10596),
.Y(n_15603)
);

AND2x2_ASAP7_75t_L g15604 ( 
.A(n_14887),
.B(n_10596),
.Y(n_15604)
);

AND2x2_ASAP7_75t_L g15605 ( 
.A(n_14891),
.B(n_10600),
.Y(n_15605)
);

AND2x4_ASAP7_75t_L g15606 ( 
.A(n_15180),
.B(n_7857),
.Y(n_15606)
);

NAND2x1p5_ASAP7_75t_L g15607 ( 
.A(n_14896),
.B(n_8057),
.Y(n_15607)
);

AND2x2_ASAP7_75t_L g15608 ( 
.A(n_14914),
.B(n_10600),
.Y(n_15608)
);

NAND2xp5_ASAP7_75t_L g15609 ( 
.A(n_14994),
.B(n_10615),
.Y(n_15609)
);

AND2x2_ASAP7_75t_L g15610 ( 
.A(n_14950),
.B(n_10615),
.Y(n_15610)
);

AND2x4_ASAP7_75t_L g15611 ( 
.A(n_15095),
.B(n_7857),
.Y(n_15611)
);

INVx1_ASAP7_75t_L g15612 ( 
.A(n_15000),
.Y(n_15612)
);

INVx1_ASAP7_75t_L g15613 ( 
.A(n_14838),
.Y(n_15613)
);

AND2x2_ASAP7_75t_L g15614 ( 
.A(n_15158),
.B(n_10625),
.Y(n_15614)
);

AND2x2_ASAP7_75t_L g15615 ( 
.A(n_14883),
.B(n_10625),
.Y(n_15615)
);

AND2x2_ASAP7_75t_L g15616 ( 
.A(n_14965),
.B(n_10635),
.Y(n_15616)
);

INVx2_ASAP7_75t_L g15617 ( 
.A(n_14876),
.Y(n_15617)
);

INVx1_ASAP7_75t_L g15618 ( 
.A(n_14877),
.Y(n_15618)
);

OR2x2_ASAP7_75t_L g15619 ( 
.A(n_14781),
.B(n_10635),
.Y(n_15619)
);

INVx1_ASAP7_75t_L g15620 ( 
.A(n_14815),
.Y(n_15620)
);

INVx1_ASAP7_75t_L g15621 ( 
.A(n_14866),
.Y(n_15621)
);

NOR2xp33_ASAP7_75t_L g15622 ( 
.A(n_15086),
.B(n_10640),
.Y(n_15622)
);

INVx2_ASAP7_75t_L g15623 ( 
.A(n_14939),
.Y(n_15623)
);

INVx1_ASAP7_75t_L g15624 ( 
.A(n_14976),
.Y(n_15624)
);

INVx1_ASAP7_75t_L g15625 ( 
.A(n_14861),
.Y(n_15625)
);

INVx1_ASAP7_75t_L g15626 ( 
.A(n_15164),
.Y(n_15626)
);

INVx1_ASAP7_75t_L g15627 ( 
.A(n_15172),
.Y(n_15627)
);

INVxp67_ASAP7_75t_L g15628 ( 
.A(n_15165),
.Y(n_15628)
);

AND2x2_ASAP7_75t_L g15629 ( 
.A(n_14959),
.B(n_10640),
.Y(n_15629)
);

AND2x2_ASAP7_75t_L g15630 ( 
.A(n_14960),
.B(n_10642),
.Y(n_15630)
);

AND2x2_ASAP7_75t_L g15631 ( 
.A(n_15303),
.B(n_10642),
.Y(n_15631)
);

NAND2xp5_ASAP7_75t_L g15632 ( 
.A(n_15310),
.B(n_10643),
.Y(n_15632)
);

AND2x2_ASAP7_75t_L g15633 ( 
.A(n_14977),
.B(n_10643),
.Y(n_15633)
);

AND2x2_ASAP7_75t_L g15634 ( 
.A(n_15052),
.B(n_10649),
.Y(n_15634)
);

AND2x2_ASAP7_75t_L g15635 ( 
.A(n_15281),
.B(n_10649),
.Y(n_15635)
);

INVx1_ASAP7_75t_L g15636 ( 
.A(n_15248),
.Y(n_15636)
);

INVx2_ASAP7_75t_SL g15637 ( 
.A(n_15089),
.Y(n_15637)
);

INVx1_ASAP7_75t_L g15638 ( 
.A(n_15263),
.Y(n_15638)
);

INVx1_ASAP7_75t_L g15639 ( 
.A(n_15193),
.Y(n_15639)
);

AND2x2_ASAP7_75t_L g15640 ( 
.A(n_14962),
.B(n_10651),
.Y(n_15640)
);

INVx4_ASAP7_75t_L g15641 ( 
.A(n_14895),
.Y(n_15641)
);

AND2x2_ASAP7_75t_L g15642 ( 
.A(n_15088),
.B(n_10651),
.Y(n_15642)
);

NAND2xp5_ASAP7_75t_L g15643 ( 
.A(n_15308),
.B(n_10654),
.Y(n_15643)
);

INVx6_ASAP7_75t_L g15644 ( 
.A(n_15265),
.Y(n_15644)
);

INVx1_ASAP7_75t_L g15645 ( 
.A(n_15198),
.Y(n_15645)
);

AND2x4_ASAP7_75t_L g15646 ( 
.A(n_15205),
.B(n_7857),
.Y(n_15646)
);

BUFx2_ASAP7_75t_L g15647 ( 
.A(n_14957),
.Y(n_15647)
);

AND2x2_ASAP7_75t_L g15648 ( 
.A(n_15105),
.B(n_10654),
.Y(n_15648)
);

INVx2_ASAP7_75t_L g15649 ( 
.A(n_15068),
.Y(n_15649)
);

INVx1_ASAP7_75t_L g15650 ( 
.A(n_15199),
.Y(n_15650)
);

AND2x2_ASAP7_75t_L g15651 ( 
.A(n_15316),
.B(n_10662),
.Y(n_15651)
);

INVx4_ASAP7_75t_L g15652 ( 
.A(n_15333),
.Y(n_15652)
);

AND2x2_ASAP7_75t_L g15653 ( 
.A(n_15299),
.B(n_10662),
.Y(n_15653)
);

OR2x2_ASAP7_75t_L g15654 ( 
.A(n_15335),
.B(n_10667),
.Y(n_15654)
);

INVx2_ASAP7_75t_SL g15655 ( 
.A(n_15219),
.Y(n_15655)
);

NAND2xp5_ASAP7_75t_L g15656 ( 
.A(n_15253),
.B(n_10667),
.Y(n_15656)
);

INVx2_ASAP7_75t_L g15657 ( 
.A(n_15077),
.Y(n_15657)
);

AND2x2_ASAP7_75t_L g15658 ( 
.A(n_14852),
.B(n_10678),
.Y(n_15658)
);

NAND2xp5_ASAP7_75t_L g15659 ( 
.A(n_15209),
.B(n_10678),
.Y(n_15659)
);

INVx2_ASAP7_75t_L g15660 ( 
.A(n_15219),
.Y(n_15660)
);

AND2x2_ASAP7_75t_L g15661 ( 
.A(n_15146),
.B(n_15074),
.Y(n_15661)
);

AND2x2_ASAP7_75t_L g15662 ( 
.A(n_15213),
.B(n_10682),
.Y(n_15662)
);

OR2x2_ASAP7_75t_L g15663 ( 
.A(n_14948),
.B(n_14801),
.Y(n_15663)
);

NOR2x1_ASAP7_75t_SL g15664 ( 
.A(n_14847),
.B(n_8207),
.Y(n_15664)
);

NAND2xp5_ASAP7_75t_L g15665 ( 
.A(n_15270),
.B(n_10682),
.Y(n_15665)
);

AND2x2_ASAP7_75t_L g15666 ( 
.A(n_14970),
.B(n_10695),
.Y(n_15666)
);

INVx4_ASAP7_75t_L g15667 ( 
.A(n_15207),
.Y(n_15667)
);

AND2x2_ASAP7_75t_L g15668 ( 
.A(n_15227),
.B(n_10695),
.Y(n_15668)
);

NAND2xp5_ASAP7_75t_L g15669 ( 
.A(n_15075),
.B(n_10697),
.Y(n_15669)
);

NAND2xp5_ASAP7_75t_L g15670 ( 
.A(n_15081),
.B(n_10697),
.Y(n_15670)
);

INVx1_ASAP7_75t_L g15671 ( 
.A(n_14836),
.Y(n_15671)
);

OR2x2_ASAP7_75t_L g15672 ( 
.A(n_14971),
.B(n_10698),
.Y(n_15672)
);

AND2x2_ASAP7_75t_L g15673 ( 
.A(n_15211),
.B(n_10698),
.Y(n_15673)
);

AND2x4_ASAP7_75t_L g15674 ( 
.A(n_15220),
.B(n_7918),
.Y(n_15674)
);

AND2x2_ASAP7_75t_L g15675 ( 
.A(n_15242),
.B(n_15246),
.Y(n_15675)
);

AND2x4_ASAP7_75t_SL g15676 ( 
.A(n_15225),
.B(n_8861),
.Y(n_15676)
);

AND2x2_ASAP7_75t_L g15677 ( 
.A(n_15278),
.B(n_10701),
.Y(n_15677)
);

INVx2_ASAP7_75t_L g15678 ( 
.A(n_15065),
.Y(n_15678)
);

NAND2xp5_ASAP7_75t_L g15679 ( 
.A(n_14901),
.B(n_10701),
.Y(n_15679)
);

AND2x2_ASAP7_75t_L g15680 ( 
.A(n_15342),
.B(n_10704),
.Y(n_15680)
);

NAND2xp5_ASAP7_75t_L g15681 ( 
.A(n_14909),
.B(n_10704),
.Y(n_15681)
);

AND2x2_ASAP7_75t_L g15682 ( 
.A(n_15365),
.B(n_10713),
.Y(n_15682)
);

NAND2xp5_ASAP7_75t_L g15683 ( 
.A(n_14912),
.B(n_10713),
.Y(n_15683)
);

INVx1_ASAP7_75t_L g15684 ( 
.A(n_14890),
.Y(n_15684)
);

INVx1_ASAP7_75t_L g15685 ( 
.A(n_14931),
.Y(n_15685)
);

HB1xp67_ASAP7_75t_L g15686 ( 
.A(n_15113),
.Y(n_15686)
);

INVx2_ASAP7_75t_L g15687 ( 
.A(n_15065),
.Y(n_15687)
);

AND2x2_ASAP7_75t_L g15688 ( 
.A(n_15323),
.B(n_10723),
.Y(n_15688)
);

INVx2_ASAP7_75t_L g15689 ( 
.A(n_15239),
.Y(n_15689)
);

INVx1_ASAP7_75t_L g15690 ( 
.A(n_14933),
.Y(n_15690)
);

AND2x2_ASAP7_75t_L g15691 ( 
.A(n_15329),
.B(n_10723),
.Y(n_15691)
);

INVx1_ASAP7_75t_L g15692 ( 
.A(n_14934),
.Y(n_15692)
);

AND2x2_ASAP7_75t_L g15693 ( 
.A(n_15334),
.B(n_10724),
.Y(n_15693)
);

AND2x2_ASAP7_75t_L g15694 ( 
.A(n_15336),
.B(n_10724),
.Y(n_15694)
);

NAND2xp5_ASAP7_75t_L g15695 ( 
.A(n_14913),
.B(n_10726),
.Y(n_15695)
);

HB1xp67_ASAP7_75t_L g15696 ( 
.A(n_15256),
.Y(n_15696)
);

OR2x2_ASAP7_75t_L g15697 ( 
.A(n_14777),
.B(n_10726),
.Y(n_15697)
);

NAND2xp5_ASAP7_75t_L g15698 ( 
.A(n_14898),
.B(n_10729),
.Y(n_15698)
);

NAND2xp5_ASAP7_75t_SL g15699 ( 
.A(n_14850),
.B(n_8207),
.Y(n_15699)
);

AND2x2_ASAP7_75t_L g15700 ( 
.A(n_15353),
.B(n_10729),
.Y(n_15700)
);

NAND2xp5_ASAP7_75t_L g15701 ( 
.A(n_15116),
.B(n_15122),
.Y(n_15701)
);

AND2x2_ASAP7_75t_L g15702 ( 
.A(n_15366),
.B(n_10730),
.Y(n_15702)
);

AND2x2_ASAP7_75t_L g15703 ( 
.A(n_15368),
.B(n_10730),
.Y(n_15703)
);

INVx2_ASAP7_75t_L g15704 ( 
.A(n_15262),
.Y(n_15704)
);

NAND2xp5_ASAP7_75t_L g15705 ( 
.A(n_15124),
.B(n_10731),
.Y(n_15705)
);

INVx1_ASAP7_75t_L g15706 ( 
.A(n_14935),
.Y(n_15706)
);

AND2x2_ASAP7_75t_L g15707 ( 
.A(n_15369),
.B(n_10731),
.Y(n_15707)
);

INVx1_ASAP7_75t_L g15708 ( 
.A(n_14822),
.Y(n_15708)
);

HB1xp67_ASAP7_75t_L g15709 ( 
.A(n_15119),
.Y(n_15709)
);

AND2x2_ASAP7_75t_L g15710 ( 
.A(n_15371),
.B(n_10732),
.Y(n_15710)
);

NOR2xp33_ASAP7_75t_L g15711 ( 
.A(n_15190),
.B(n_10732),
.Y(n_15711)
);

OR2x2_ASAP7_75t_L g15712 ( 
.A(n_14818),
.B(n_10736),
.Y(n_15712)
);

AND2x2_ASAP7_75t_L g15713 ( 
.A(n_15301),
.B(n_10736),
.Y(n_15713)
);

INVx1_ASAP7_75t_L g15714 ( 
.A(n_14940),
.Y(n_15714)
);

NAND2xp5_ASAP7_75t_L g15715 ( 
.A(n_15139),
.B(n_14930),
.Y(n_15715)
);

BUFx2_ASAP7_75t_L g15716 ( 
.A(n_15082),
.Y(n_15716)
);

INVx1_ASAP7_75t_L g15717 ( 
.A(n_14906),
.Y(n_15717)
);

NAND2xp5_ASAP7_75t_L g15718 ( 
.A(n_14979),
.B(n_10743),
.Y(n_15718)
);

AND2x2_ASAP7_75t_L g15719 ( 
.A(n_15378),
.B(n_15234),
.Y(n_15719)
);

INVx2_ASAP7_75t_SL g15720 ( 
.A(n_15117),
.Y(n_15720)
);

AND2x2_ASAP7_75t_L g15721 ( 
.A(n_14999),
.B(n_10743),
.Y(n_15721)
);

OAI211xp5_ASAP7_75t_L g15722 ( 
.A1(n_14807),
.A2(n_10972),
.B(n_10668),
.C(n_10599),
.Y(n_15722)
);

INVx3_ASAP7_75t_L g15723 ( 
.A(n_15020),
.Y(n_15723)
);

INVx2_ASAP7_75t_L g15724 ( 
.A(n_15240),
.Y(n_15724)
);

AND2x4_ASAP7_75t_L g15725 ( 
.A(n_15166),
.B(n_7918),
.Y(n_15725)
);

INVx1_ASAP7_75t_L g15726 ( 
.A(n_15027),
.Y(n_15726)
);

NAND2xp5_ASAP7_75t_L g15727 ( 
.A(n_14982),
.B(n_10746),
.Y(n_15727)
);

BUFx2_ASAP7_75t_L g15728 ( 
.A(n_15178),
.Y(n_15728)
);

INVx1_ASAP7_75t_L g15729 ( 
.A(n_14964),
.Y(n_15729)
);

INVx2_ASAP7_75t_L g15730 ( 
.A(n_15186),
.Y(n_15730)
);

AND2x2_ASAP7_75t_L g15731 ( 
.A(n_15305),
.B(n_10746),
.Y(n_15731)
);

INVx1_ASAP7_75t_L g15732 ( 
.A(n_14966),
.Y(n_15732)
);

AND2x2_ASAP7_75t_L g15733 ( 
.A(n_15306),
.B(n_10753),
.Y(n_15733)
);

NOR2xp33_ASAP7_75t_L g15734 ( 
.A(n_15040),
.B(n_10753),
.Y(n_15734)
);

AND2x4_ASAP7_75t_L g15735 ( 
.A(n_14987),
.B(n_7918),
.Y(n_15735)
);

AND2x2_ASAP7_75t_L g15736 ( 
.A(n_15307),
.B(n_10754),
.Y(n_15736)
);

INVx2_ASAP7_75t_L g15737 ( 
.A(n_15076),
.Y(n_15737)
);

INVxp67_ASAP7_75t_SL g15738 ( 
.A(n_15120),
.Y(n_15738)
);

AND2x4_ASAP7_75t_L g15739 ( 
.A(n_15015),
.B(n_7956),
.Y(n_15739)
);

AND2x2_ASAP7_75t_L g15740 ( 
.A(n_15070),
.B(n_10754),
.Y(n_15740)
);

AND2x2_ASAP7_75t_L g15741 ( 
.A(n_15130),
.B(n_10762),
.Y(n_15741)
);

AND2x2_ASAP7_75t_L g15742 ( 
.A(n_15311),
.B(n_10762),
.Y(n_15742)
);

AND2x4_ASAP7_75t_L g15743 ( 
.A(n_15053),
.B(n_7956),
.Y(n_15743)
);

INVx2_ASAP7_75t_L g15744 ( 
.A(n_15076),
.Y(n_15744)
);

INVx1_ASAP7_75t_L g15745 ( 
.A(n_14968),
.Y(n_15745)
);

INVx1_ASAP7_75t_L g15746 ( 
.A(n_14798),
.Y(n_15746)
);

INVx2_ASAP7_75t_L g15747 ( 
.A(n_15137),
.Y(n_15747)
);

INVx2_ASAP7_75t_L g15748 ( 
.A(n_15137),
.Y(n_15748)
);

INVx1_ASAP7_75t_L g15749 ( 
.A(n_15066),
.Y(n_15749)
);

INVx2_ASAP7_75t_L g15750 ( 
.A(n_14996),
.Y(n_15750)
);

INVxp67_ASAP7_75t_SL g15751 ( 
.A(n_15127),
.Y(n_15751)
);

INVx1_ASAP7_75t_L g15752 ( 
.A(n_15058),
.Y(n_15752)
);

INVx2_ASAP7_75t_L g15753 ( 
.A(n_15201),
.Y(n_15753)
);

AND2x2_ASAP7_75t_L g15754 ( 
.A(n_15045),
.B(n_10763),
.Y(n_15754)
);

NOR2xp67_ASAP7_75t_L g15755 ( 
.A(n_15297),
.B(n_10763),
.Y(n_15755)
);

BUFx2_ASAP7_75t_L g15756 ( 
.A(n_14991),
.Y(n_15756)
);

INVx1_ASAP7_75t_L g15757 ( 
.A(n_14952),
.Y(n_15757)
);

OR2x2_ASAP7_75t_L g15758 ( 
.A(n_15004),
.B(n_10764),
.Y(n_15758)
);

NAND2xp5_ASAP7_75t_L g15759 ( 
.A(n_14902),
.B(n_10764),
.Y(n_15759)
);

INVx1_ASAP7_75t_L g15760 ( 
.A(n_14958),
.Y(n_15760)
);

NAND3xp33_ASAP7_75t_L g15761 ( 
.A(n_14993),
.B(n_15001),
.C(n_14988),
.Y(n_15761)
);

INVx2_ASAP7_75t_L g15762 ( 
.A(n_15208),
.Y(n_15762)
);

AND2x2_ASAP7_75t_L g15763 ( 
.A(n_15142),
.B(n_10773),
.Y(n_15763)
);

INVx5_ASAP7_75t_L g15764 ( 
.A(n_15372),
.Y(n_15764)
);

INVx2_ASAP7_75t_L g15765 ( 
.A(n_15041),
.Y(n_15765)
);

INVxp67_ASAP7_75t_SL g15766 ( 
.A(n_14812),
.Y(n_15766)
);

OR2x2_ASAP7_75t_L g15767 ( 
.A(n_14974),
.B(n_10773),
.Y(n_15767)
);

INVx1_ASAP7_75t_L g15768 ( 
.A(n_15009),
.Y(n_15768)
);

OR2x2_ASAP7_75t_L g15769 ( 
.A(n_14951),
.B(n_14955),
.Y(n_15769)
);

INVx2_ASAP7_75t_L g15770 ( 
.A(n_15014),
.Y(n_15770)
);

HB1xp67_ASAP7_75t_L g15771 ( 
.A(n_15169),
.Y(n_15771)
);

NAND2xp5_ASAP7_75t_L g15772 ( 
.A(n_15011),
.B(n_10780),
.Y(n_15772)
);

INVx2_ASAP7_75t_L g15773 ( 
.A(n_15018),
.Y(n_15773)
);

INVx3_ASAP7_75t_L g15774 ( 
.A(n_15028),
.Y(n_15774)
);

HB1xp67_ASAP7_75t_L g15775 ( 
.A(n_15016),
.Y(n_15775)
);

OAI33xp33_ASAP7_75t_L g15776 ( 
.A1(n_15304),
.A2(n_10782),
.A3(n_10788),
.B1(n_10811),
.B2(n_10804),
.B3(n_10780),
.Y(n_15776)
);

INVx1_ASAP7_75t_L g15777 ( 
.A(n_15047),
.Y(n_15777)
);

OR2x2_ASAP7_75t_L g15778 ( 
.A(n_15163),
.B(n_10782),
.Y(n_15778)
);

INVx2_ASAP7_75t_SL g15779 ( 
.A(n_15087),
.Y(n_15779)
);

AND2x2_ASAP7_75t_L g15780 ( 
.A(n_15309),
.B(n_10788),
.Y(n_15780)
);

OR2x2_ASAP7_75t_L g15781 ( 
.A(n_15049),
.B(n_10804),
.Y(n_15781)
);

NAND2xp5_ASAP7_75t_L g15782 ( 
.A(n_15051),
.B(n_10811),
.Y(n_15782)
);

NAND2xp5_ASAP7_75t_L g15783 ( 
.A(n_15128),
.B(n_10814),
.Y(n_15783)
);

NAND2xp5_ASAP7_75t_L g15784 ( 
.A(n_15153),
.B(n_10814),
.Y(n_15784)
);

NOR2x1_ASAP7_75t_L g15785 ( 
.A(n_15160),
.B(n_10822),
.Y(n_15785)
);

NAND2xp5_ASAP7_75t_L g15786 ( 
.A(n_15035),
.B(n_10822),
.Y(n_15786)
);

OR2x2_ASAP7_75t_L g15787 ( 
.A(n_14945),
.B(n_10833),
.Y(n_15787)
);

INVx3_ASAP7_75t_L g15788 ( 
.A(n_15057),
.Y(n_15788)
);

HB1xp67_ASAP7_75t_L g15789 ( 
.A(n_15007),
.Y(n_15789)
);

AND2x2_ASAP7_75t_L g15790 ( 
.A(n_15147),
.B(n_10833),
.Y(n_15790)
);

BUFx2_ASAP7_75t_L g15791 ( 
.A(n_15375),
.Y(n_15791)
);

INVx1_ASAP7_75t_L g15792 ( 
.A(n_14937),
.Y(n_15792)
);

AND2x2_ASAP7_75t_L g15793 ( 
.A(n_15176),
.B(n_10837),
.Y(n_15793)
);

AND2x2_ASAP7_75t_L g15794 ( 
.A(n_14995),
.B(n_10837),
.Y(n_15794)
);

INVx1_ASAP7_75t_SL g15795 ( 
.A(n_15250),
.Y(n_15795)
);

OR2x2_ASAP7_75t_L g15796 ( 
.A(n_15294),
.B(n_10843),
.Y(n_15796)
);

AND2x2_ASAP7_75t_L g15797 ( 
.A(n_15043),
.B(n_10843),
.Y(n_15797)
);

AND2x2_ASAP7_75t_L g15798 ( 
.A(n_15056),
.B(n_15059),
.Y(n_15798)
);

AND2x2_ASAP7_75t_L g15799 ( 
.A(n_15182),
.B(n_10848),
.Y(n_15799)
);

INVx1_ASAP7_75t_L g15800 ( 
.A(n_14944),
.Y(n_15800)
);

INVx1_ASAP7_75t_L g15801 ( 
.A(n_15013),
.Y(n_15801)
);

INVx1_ASAP7_75t_SL g15802 ( 
.A(n_15103),
.Y(n_15802)
);

INVx1_ASAP7_75t_L g15803 ( 
.A(n_14956),
.Y(n_15803)
);

NAND2xp5_ASAP7_75t_L g15804 ( 
.A(n_15036),
.B(n_15214),
.Y(n_15804)
);

AND2x2_ASAP7_75t_L g15805 ( 
.A(n_15134),
.B(n_10848),
.Y(n_15805)
);

INVx1_ASAP7_75t_L g15806 ( 
.A(n_15006),
.Y(n_15806)
);

NAND4xp25_ASAP7_75t_L g15807 ( 
.A(n_15149),
.B(n_15062),
.C(n_15315),
.D(n_15218),
.Y(n_15807)
);

INVx2_ASAP7_75t_SL g15808 ( 
.A(n_15352),
.Y(n_15808)
);

INVx2_ASAP7_75t_L g15809 ( 
.A(n_15264),
.Y(n_15809)
);

AND2x2_ASAP7_75t_L g15810 ( 
.A(n_15266),
.B(n_10862),
.Y(n_15810)
);

INVx1_ASAP7_75t_L g15811 ( 
.A(n_15021),
.Y(n_15811)
);

OAI22xp5_ASAP7_75t_L g15812 ( 
.A1(n_15283),
.A2(n_15174),
.B1(n_15328),
.B2(n_15090),
.Y(n_15812)
);

NOR2xp33_ASAP7_75t_L g15813 ( 
.A(n_15217),
.B(n_15340),
.Y(n_15813)
);

INVx2_ASAP7_75t_L g15814 ( 
.A(n_15383),
.Y(n_15814)
);

NOR2x1_ASAP7_75t_SL g15815 ( 
.A(n_15129),
.B(n_8207),
.Y(n_15815)
);

INVx1_ASAP7_75t_L g15816 ( 
.A(n_15033),
.Y(n_15816)
);

AND2x2_ASAP7_75t_L g15817 ( 
.A(n_15267),
.B(n_10862),
.Y(n_15817)
);

AND2x2_ASAP7_75t_L g15818 ( 
.A(n_15271),
.B(n_10864),
.Y(n_15818)
);

INVx1_ASAP7_75t_L g15819 ( 
.A(n_15032),
.Y(n_15819)
);

AND2x4_ASAP7_75t_L g15820 ( 
.A(n_15230),
.B(n_7956),
.Y(n_15820)
);

INVx1_ASAP7_75t_L g15821 ( 
.A(n_15063),
.Y(n_15821)
);

AND2x2_ASAP7_75t_L g15822 ( 
.A(n_15275),
.B(n_10864),
.Y(n_15822)
);

NAND2xp5_ASAP7_75t_L g15823 ( 
.A(n_15233),
.B(n_10868),
.Y(n_15823)
);

HB1xp67_ASAP7_75t_L g15824 ( 
.A(n_15111),
.Y(n_15824)
);

OR2x2_ASAP7_75t_L g15825 ( 
.A(n_15005),
.B(n_15025),
.Y(n_15825)
);

INVx2_ASAP7_75t_L g15826 ( 
.A(n_15341),
.Y(n_15826)
);

INVx1_ASAP7_75t_L g15827 ( 
.A(n_15067),
.Y(n_15827)
);

BUFx2_ASAP7_75t_L g15828 ( 
.A(n_15243),
.Y(n_15828)
);

INVx1_ASAP7_75t_L g15829 ( 
.A(n_15072),
.Y(n_15829)
);

AND2x2_ASAP7_75t_L g15830 ( 
.A(n_15277),
.B(n_10868),
.Y(n_15830)
);

NOR2xp33_ASAP7_75t_L g15831 ( 
.A(n_15346),
.B(n_10874),
.Y(n_15831)
);

BUFx3_ASAP7_75t_L g15832 ( 
.A(n_15222),
.Y(n_15832)
);

INVx2_ASAP7_75t_L g15833 ( 
.A(n_15064),
.Y(n_15833)
);

INVx2_ASAP7_75t_L g15834 ( 
.A(n_15254),
.Y(n_15834)
);

NAND2xp5_ASAP7_75t_L g15835 ( 
.A(n_15295),
.B(n_15228),
.Y(n_15835)
);

INVx2_ASAP7_75t_SL g15836 ( 
.A(n_15114),
.Y(n_15836)
);

AND2x2_ASAP7_75t_L g15837 ( 
.A(n_14989),
.B(n_10874),
.Y(n_15837)
);

INVx2_ASAP7_75t_L g15838 ( 
.A(n_15046),
.Y(n_15838)
);

AND2x2_ASAP7_75t_L g15839 ( 
.A(n_15055),
.B(n_10882),
.Y(n_15839)
);

INVx2_ASAP7_75t_L g15840 ( 
.A(n_15345),
.Y(n_15840)
);

AOI22xp33_ASAP7_75t_L g15841 ( 
.A1(n_15268),
.A2(n_7823),
.B1(n_7800),
.B2(n_10668),
.Y(n_15841)
);

OR2x2_ASAP7_75t_L g15842 ( 
.A(n_14998),
.B(n_10882),
.Y(n_15842)
);

OR2x2_ASAP7_75t_L g15843 ( 
.A(n_15255),
.B(n_10894),
.Y(n_15843)
);

AND2x2_ASAP7_75t_L g15844 ( 
.A(n_15269),
.B(n_10894),
.Y(n_15844)
);

AND2x2_ASAP7_75t_L g15845 ( 
.A(n_15284),
.B(n_10915),
.Y(n_15845)
);

INVx1_ASAP7_75t_L g15846 ( 
.A(n_15054),
.Y(n_15846)
);

NAND2xp5_ASAP7_75t_L g15847 ( 
.A(n_15229),
.B(n_10915),
.Y(n_15847)
);

AND2x4_ASAP7_75t_L g15848 ( 
.A(n_15272),
.B(n_8023),
.Y(n_15848)
);

OR2x2_ASAP7_75t_L g15849 ( 
.A(n_15050),
.B(n_10920),
.Y(n_15849)
);

INVx2_ASAP7_75t_L g15850 ( 
.A(n_15349),
.Y(n_15850)
);

INVx1_ASAP7_75t_L g15851 ( 
.A(n_15060),
.Y(n_15851)
);

NAND2x1p5_ASAP7_75t_L g15852 ( 
.A(n_15097),
.B(n_8207),
.Y(n_15852)
);

INVx1_ASAP7_75t_L g15853 ( 
.A(n_15177),
.Y(n_15853)
);

AND2x2_ASAP7_75t_L g15854 ( 
.A(n_15291),
.B(n_15188),
.Y(n_15854)
);

AND2x2_ASAP7_75t_L g15855 ( 
.A(n_15192),
.B(n_10920),
.Y(n_15855)
);

INVx1_ASAP7_75t_L g15856 ( 
.A(n_15181),
.Y(n_15856)
);

INVx4_ASAP7_75t_L g15857 ( 
.A(n_15282),
.Y(n_15857)
);

AND2x2_ASAP7_75t_L g15858 ( 
.A(n_15093),
.B(n_15096),
.Y(n_15858)
);

INVx1_ASAP7_75t_L g15859 ( 
.A(n_14997),
.Y(n_15859)
);

HB1xp67_ASAP7_75t_L g15860 ( 
.A(n_15175),
.Y(n_15860)
);

INVx1_ASAP7_75t_L g15861 ( 
.A(n_15260),
.Y(n_15861)
);

OA21x2_ASAP7_75t_L g15862 ( 
.A1(n_15363),
.A2(n_10928),
.B(n_10924),
.Y(n_15862)
);

INVx1_ASAP7_75t_L g15863 ( 
.A(n_15276),
.Y(n_15863)
);

AND2x2_ASAP7_75t_L g15864 ( 
.A(n_15100),
.B(n_10924),
.Y(n_15864)
);

AND2x2_ASAP7_75t_L g15865 ( 
.A(n_15107),
.B(n_10928),
.Y(n_15865)
);

NOR2xp67_ASAP7_75t_L g15866 ( 
.A(n_15324),
.B(n_10930),
.Y(n_15866)
);

INVx1_ASAP7_75t_L g15867 ( 
.A(n_15168),
.Y(n_15867)
);

INVx1_ASAP7_75t_L g15868 ( 
.A(n_15259),
.Y(n_15868)
);

AND2x2_ASAP7_75t_L g15869 ( 
.A(n_15123),
.B(n_10930),
.Y(n_15869)
);

INVxp67_ASAP7_75t_SL g15870 ( 
.A(n_15150),
.Y(n_15870)
);

OR2x2_ASAP7_75t_L g15871 ( 
.A(n_15094),
.B(n_10936),
.Y(n_15871)
);

AND2x2_ASAP7_75t_L g15872 ( 
.A(n_15125),
.B(n_10936),
.Y(n_15872)
);

INVx1_ASAP7_75t_L g15873 ( 
.A(n_15079),
.Y(n_15873)
);

INVx1_ASAP7_75t_L g15874 ( 
.A(n_15285),
.Y(n_15874)
);

AND2x2_ASAP7_75t_L g15875 ( 
.A(n_15126),
.B(n_10938),
.Y(n_15875)
);

INVx2_ASAP7_75t_L g15876 ( 
.A(n_15356),
.Y(n_15876)
);

NAND2x1p5_ASAP7_75t_L g15877 ( 
.A(n_15237),
.B(n_8618),
.Y(n_15877)
);

AND2x2_ASAP7_75t_L g15878 ( 
.A(n_15136),
.B(n_15140),
.Y(n_15878)
);

OR2x2_ASAP7_75t_L g15879 ( 
.A(n_15202),
.B(n_10938),
.Y(n_15879)
);

NAND2xp5_ASAP7_75t_L g15880 ( 
.A(n_15287),
.B(n_10944),
.Y(n_15880)
);

INVx1_ASAP7_75t_L g15881 ( 
.A(n_15290),
.Y(n_15881)
);

NOR2x1_ASAP7_75t_SL g15882 ( 
.A(n_15286),
.B(n_8618),
.Y(n_15882)
);

AND2x2_ASAP7_75t_L g15883 ( 
.A(n_15143),
.B(n_10944),
.Y(n_15883)
);

OR2x2_ASAP7_75t_L g15884 ( 
.A(n_15203),
.B(n_10952),
.Y(n_15884)
);

INVx1_ASAP7_75t_L g15885 ( 
.A(n_15061),
.Y(n_15885)
);

AOI22xp33_ASAP7_75t_L g15886 ( 
.A1(n_15249),
.A2(n_10972),
.B1(n_10653),
.B2(n_10599),
.Y(n_15886)
);

INVx2_ASAP7_75t_L g15887 ( 
.A(n_15364),
.Y(n_15887)
);

INVx1_ASAP7_75t_L g15888 ( 
.A(n_15069),
.Y(n_15888)
);

AOI21xp5_ASAP7_75t_L g15889 ( 
.A1(n_15085),
.A2(n_10653),
.B(n_10647),
.Y(n_15889)
);

NOR3xp33_ASAP7_75t_SL g15890 ( 
.A(n_15204),
.B(n_8035),
.C(n_8033),
.Y(n_15890)
);

INVx2_ASAP7_75t_L g15891 ( 
.A(n_15151),
.Y(n_15891)
);

INVx2_ASAP7_75t_L g15892 ( 
.A(n_15152),
.Y(n_15892)
);

AND2x2_ASAP7_75t_L g15893 ( 
.A(n_15167),
.B(n_10952),
.Y(n_15893)
);

AND2x2_ASAP7_75t_L g15894 ( 
.A(n_15171),
.B(n_10953),
.Y(n_15894)
);

INVx1_ASAP7_75t_L g15895 ( 
.A(n_15091),
.Y(n_15895)
);

AND2x2_ASAP7_75t_L g15896 ( 
.A(n_15210),
.B(n_10953),
.Y(n_15896)
);

HB1xp67_ASAP7_75t_L g15897 ( 
.A(n_15280),
.Y(n_15897)
);

INVx2_ASAP7_75t_L g15898 ( 
.A(n_15156),
.Y(n_15898)
);

NAND5xp2_ASAP7_75t_L g15899 ( 
.A(n_15300),
.B(n_15321),
.C(n_15325),
.D(n_15318),
.E(n_15302),
.Y(n_15899)
);

OR2x2_ASAP7_75t_L g15900 ( 
.A(n_15212),
.B(n_10957),
.Y(n_15900)
);

AND2x2_ASAP7_75t_L g15901 ( 
.A(n_15179),
.B(n_10957),
.Y(n_15901)
);

AND2x2_ASAP7_75t_L g15902 ( 
.A(n_15216),
.B(n_10958),
.Y(n_15902)
);

AND2x2_ASAP7_75t_L g15903 ( 
.A(n_15026),
.B(n_10958),
.Y(n_15903)
);

INVx4_ASAP7_75t_L g15904 ( 
.A(n_15330),
.Y(n_15904)
);

INVx2_ASAP7_75t_L g15905 ( 
.A(n_15319),
.Y(n_15905)
);

NAND2xp5_ASAP7_75t_SL g15906 ( 
.A(n_15257),
.B(n_8618),
.Y(n_15906)
);

INVx1_ASAP7_75t_L g15907 ( 
.A(n_15131),
.Y(n_15907)
);

INVx1_ASAP7_75t_L g15908 ( 
.A(n_15073),
.Y(n_15908)
);

INVx1_ASAP7_75t_L g15909 ( 
.A(n_15261),
.Y(n_15909)
);

NAND2xp5_ASAP7_75t_L g15910 ( 
.A(n_15338),
.B(n_10959),
.Y(n_15910)
);

NOR2xp33_ASAP7_75t_SL g15911 ( 
.A(n_15092),
.B(n_6772),
.Y(n_15911)
);

INVx1_ASAP7_75t_L g15912 ( 
.A(n_15196),
.Y(n_15912)
);

AND2x2_ASAP7_75t_L g15913 ( 
.A(n_15039),
.B(n_10959),
.Y(n_15913)
);

NAND2xp5_ASAP7_75t_L g15914 ( 
.A(n_15343),
.B(n_10961),
.Y(n_15914)
);

INVx1_ASAP7_75t_L g15915 ( 
.A(n_15223),
.Y(n_15915)
);

INVx1_ASAP7_75t_L g15916 ( 
.A(n_15245),
.Y(n_15916)
);

AND2x2_ASAP7_75t_L g15917 ( 
.A(n_15312),
.B(n_10961),
.Y(n_15917)
);

NAND2xp5_ASAP7_75t_L g15918 ( 
.A(n_15396),
.B(n_15348),
.Y(n_15918)
);

INVx1_ASAP7_75t_L g15919 ( 
.A(n_15450),
.Y(n_15919)
);

OR2x2_ASAP7_75t_L g15920 ( 
.A(n_15536),
.B(n_15247),
.Y(n_15920)
);

INVx1_ASAP7_75t_L g15921 ( 
.A(n_15594),
.Y(n_15921)
);

AND2x4_ASAP7_75t_L g15922 ( 
.A(n_15400),
.B(n_15350),
.Y(n_15922)
);

INVx2_ASAP7_75t_L g15923 ( 
.A(n_15468),
.Y(n_15923)
);

AND2x2_ASAP7_75t_L g15924 ( 
.A(n_15574),
.B(n_15313),
.Y(n_15924)
);

AND2x2_ASAP7_75t_L g15925 ( 
.A(n_15448),
.B(n_15686),
.Y(n_15925)
);

AND2x2_ASAP7_75t_L g15926 ( 
.A(n_15531),
.B(n_15351),
.Y(n_15926)
);

NAND2x1p5_ASAP7_75t_L g15927 ( 
.A(n_15434),
.B(n_15357),
.Y(n_15927)
);

INVx1_ASAP7_75t_L g15928 ( 
.A(n_15594),
.Y(n_15928)
);

NAND2xp5_ASAP7_75t_L g15929 ( 
.A(n_15386),
.B(n_15358),
.Y(n_15929)
);

HB1xp67_ASAP7_75t_L g15930 ( 
.A(n_15442),
.Y(n_15930)
);

AND2x2_ASAP7_75t_L g15931 ( 
.A(n_15492),
.B(n_15359),
.Y(n_15931)
);

INVx1_ASAP7_75t_L g15932 ( 
.A(n_15470),
.Y(n_15932)
);

INVxp33_ASAP7_75t_L g15933 ( 
.A(n_15647),
.Y(n_15933)
);

INVx1_ASAP7_75t_L g15934 ( 
.A(n_15445),
.Y(n_15934)
);

AND2x2_ASAP7_75t_L g15935 ( 
.A(n_15559),
.B(n_15360),
.Y(n_15935)
);

INVx1_ASAP7_75t_L g15936 ( 
.A(n_15449),
.Y(n_15936)
);

AND2x2_ASAP7_75t_L g15937 ( 
.A(n_15641),
.B(n_15361),
.Y(n_15937)
);

OR2x2_ASAP7_75t_L g15938 ( 
.A(n_15467),
.B(n_15215),
.Y(n_15938)
);

AND2x4_ASAP7_75t_L g15939 ( 
.A(n_15478),
.B(n_15362),
.Y(n_15939)
);

AND2x2_ASAP7_75t_L g15940 ( 
.A(n_15565),
.B(n_15464),
.Y(n_15940)
);

AND2x2_ASAP7_75t_L g15941 ( 
.A(n_15463),
.B(n_15373),
.Y(n_15941)
);

INVx2_ASAP7_75t_L g15942 ( 
.A(n_15644),
.Y(n_15942)
);

AND2x2_ASAP7_75t_L g15943 ( 
.A(n_15403),
.B(n_15385),
.Y(n_15943)
);

INVxp67_ASAP7_75t_L g15944 ( 
.A(n_15647),
.Y(n_15944)
);

INVx2_ASAP7_75t_L g15945 ( 
.A(n_15644),
.Y(n_15945)
);

NAND2xp5_ASAP7_75t_L g15946 ( 
.A(n_15509),
.B(n_15274),
.Y(n_15946)
);

INVx1_ASAP7_75t_L g15947 ( 
.A(n_15696),
.Y(n_15947)
);

INVx1_ASAP7_75t_L g15948 ( 
.A(n_15490),
.Y(n_15948)
);

AND2x2_ASAP7_75t_L g15949 ( 
.A(n_15555),
.B(n_15332),
.Y(n_15949)
);

NOR2xp33_ASAP7_75t_L g15950 ( 
.A(n_15481),
.B(n_15296),
.Y(n_15950)
);

OR2x2_ASAP7_75t_L g15951 ( 
.A(n_15508),
.B(n_15288),
.Y(n_15951)
);

NOR3xp33_ASAP7_75t_L g15952 ( 
.A(n_15412),
.B(n_15226),
.C(n_15221),
.Y(n_15952)
);

INVx1_ASAP7_75t_L g15953 ( 
.A(n_15532),
.Y(n_15953)
);

NAND3xp33_ASAP7_75t_SL g15954 ( 
.A(n_15426),
.B(n_15191),
.C(n_15173),
.Y(n_15954)
);

INVx1_ASAP7_75t_L g15955 ( 
.A(n_15501),
.Y(n_15955)
);

INVx2_ASAP7_75t_L g15956 ( 
.A(n_15525),
.Y(n_15956)
);

AND2x2_ASAP7_75t_L g15957 ( 
.A(n_15441),
.B(n_15184),
.Y(n_15957)
);

OAI31xp33_ASAP7_75t_SL g15958 ( 
.A1(n_15524),
.A2(n_15008),
.A3(n_15102),
.B(n_15098),
.Y(n_15958)
);

AND2x2_ASAP7_75t_L g15959 ( 
.A(n_15397),
.B(n_15154),
.Y(n_15959)
);

INVx1_ASAP7_75t_SL g15960 ( 
.A(n_15483),
.Y(n_15960)
);

NAND2xp5_ASAP7_75t_L g15961 ( 
.A(n_15575),
.B(n_15195),
.Y(n_15961)
);

INVx1_ASAP7_75t_SL g15962 ( 
.A(n_15572),
.Y(n_15962)
);

NOR2x1_ASAP7_75t_L g15963 ( 
.A(n_15652),
.B(n_15232),
.Y(n_15963)
);

INVx1_ASAP7_75t_L g15964 ( 
.A(n_15523),
.Y(n_15964)
);

AND2x2_ASAP7_75t_L g15965 ( 
.A(n_15408),
.B(n_15314),
.Y(n_15965)
);

AND2x2_ASAP7_75t_L g15966 ( 
.A(n_15414),
.B(n_15370),
.Y(n_15966)
);

NAND2xp5_ASAP7_75t_L g15967 ( 
.A(n_15411),
.B(n_15252),
.Y(n_15967)
);

AND2x2_ASAP7_75t_L g15968 ( 
.A(n_15469),
.B(n_15279),
.Y(n_15968)
);

NOR2xp33_ASAP7_75t_L g15969 ( 
.A(n_15454),
.B(n_15530),
.Y(n_15969)
);

INVx1_ASAP7_75t_L g15970 ( 
.A(n_15419),
.Y(n_15970)
);

AND2x2_ASAP7_75t_L g15971 ( 
.A(n_15389),
.B(n_15236),
.Y(n_15971)
);

INVx1_ASAP7_75t_L g15972 ( 
.A(n_15465),
.Y(n_15972)
);

INVx2_ASAP7_75t_L g15973 ( 
.A(n_15637),
.Y(n_15973)
);

OR2x2_ASAP7_75t_L g15974 ( 
.A(n_15452),
.B(n_15293),
.Y(n_15974)
);

INVx1_ASAP7_75t_L g15975 ( 
.A(n_15472),
.Y(n_15975)
);

INVx1_ASAP7_75t_L g15976 ( 
.A(n_15459),
.Y(n_15976)
);

INVx1_ASAP7_75t_L g15977 ( 
.A(n_15416),
.Y(n_15977)
);

AND2x2_ASAP7_75t_L g15978 ( 
.A(n_15388),
.B(n_15317),
.Y(n_15978)
);

INVx2_ASAP7_75t_L g15979 ( 
.A(n_15391),
.Y(n_15979)
);

INVx1_ASAP7_75t_L g15980 ( 
.A(n_15462),
.Y(n_15980)
);

INVx1_ASAP7_75t_L g15981 ( 
.A(n_15390),
.Y(n_15981)
);

NAND2xp5_ASAP7_75t_L g15982 ( 
.A(n_15418),
.B(n_15320),
.Y(n_15982)
);

BUFx3_ASAP7_75t_L g15983 ( 
.A(n_15402),
.Y(n_15983)
);

INVx1_ASAP7_75t_L g15984 ( 
.A(n_15393),
.Y(n_15984)
);

AND2x4_ASAP7_75t_L g15985 ( 
.A(n_15557),
.B(n_15145),
.Y(n_15985)
);

INVx2_ASAP7_75t_SL g15986 ( 
.A(n_15461),
.Y(n_15986)
);

NAND2x1_ASAP7_75t_L g15987 ( 
.A(n_15395),
.B(n_15327),
.Y(n_15987)
);

NAND2xp5_ASAP7_75t_L g15988 ( 
.A(n_15420),
.B(n_15322),
.Y(n_15988)
);

HB1xp67_ASAP7_75t_L g15989 ( 
.A(n_15387),
.Y(n_15989)
);

AND2x2_ASAP7_75t_L g15990 ( 
.A(n_15471),
.B(n_15354),
.Y(n_15990)
);

NAND4xp25_ASAP7_75t_L g15991 ( 
.A(n_15466),
.B(n_15374),
.C(n_15381),
.D(n_15376),
.Y(n_15991)
);

INVx2_ASAP7_75t_L g15992 ( 
.A(n_15664),
.Y(n_15992)
);

NAND2xp5_ASAP7_75t_L g15993 ( 
.A(n_15457),
.B(n_15326),
.Y(n_15993)
);

INVx1_ASAP7_75t_L g15994 ( 
.A(n_15394),
.Y(n_15994)
);

AND2x2_ASAP7_75t_L g15995 ( 
.A(n_15661),
.B(n_15344),
.Y(n_15995)
);

INVx2_ASAP7_75t_L g15996 ( 
.A(n_15882),
.Y(n_15996)
);

NAND2xp5_ASAP7_75t_L g15997 ( 
.A(n_15456),
.B(n_15331),
.Y(n_15997)
);

AND2x2_ASAP7_75t_L g15998 ( 
.A(n_15431),
.B(n_15298),
.Y(n_15998)
);

NAND4xp25_ASAP7_75t_L g15999 ( 
.A(n_15480),
.B(n_15384),
.C(n_15382),
.D(n_15327),
.Y(n_15999)
);

INVx2_ASAP7_75t_L g16000 ( 
.A(n_15815),
.Y(n_16000)
);

INVx2_ASAP7_75t_L g16001 ( 
.A(n_15579),
.Y(n_16001)
);

NAND4xp25_ASAP7_75t_L g16002 ( 
.A(n_15734),
.B(n_15899),
.C(n_15715),
.D(n_15460),
.Y(n_16002)
);

AND2x2_ASAP7_75t_L g16003 ( 
.A(n_15719),
.B(n_15446),
.Y(n_16003)
);

NAND2xp5_ASAP7_75t_L g16004 ( 
.A(n_15499),
.B(n_15379),
.Y(n_16004)
);

OR2x2_ASAP7_75t_L g16005 ( 
.A(n_15551),
.B(n_15347),
.Y(n_16005)
);

NAND2xp5_ASAP7_75t_L g16006 ( 
.A(n_15482),
.B(n_15505),
.Y(n_16006)
);

AND2x4_ASAP7_75t_L g16007 ( 
.A(n_15623),
.B(n_15339),
.Y(n_16007)
);

AO211x2_ASAP7_75t_L g16008 ( 
.A1(n_15589),
.A2(n_15379),
.B(n_15380),
.C(n_15339),
.Y(n_16008)
);

INVx1_ASAP7_75t_L g16009 ( 
.A(n_15406),
.Y(n_16009)
);

INVx1_ASAP7_75t_L g16010 ( 
.A(n_15546),
.Y(n_16010)
);

OR2x2_ASAP7_75t_L g16011 ( 
.A(n_15554),
.B(n_15380),
.Y(n_16011)
);

INVx2_ASAP7_75t_L g16012 ( 
.A(n_15716),
.Y(n_16012)
);

INVx2_ASAP7_75t_L g16013 ( 
.A(n_15716),
.Y(n_16013)
);

AND2x2_ASAP7_75t_L g16014 ( 
.A(n_15451),
.B(n_10971),
.Y(n_16014)
);

INVx2_ASAP7_75t_L g16015 ( 
.A(n_15398),
.Y(n_16015)
);

INVx2_ASAP7_75t_SL g16016 ( 
.A(n_15405),
.Y(n_16016)
);

AND2x2_ASAP7_75t_L g16017 ( 
.A(n_15401),
.B(n_10971),
.Y(n_16017)
);

INVx1_ASAP7_75t_L g16018 ( 
.A(n_15546),
.Y(n_16018)
);

AND2x2_ASAP7_75t_L g16019 ( 
.A(n_15476),
.B(n_10981),
.Y(n_16019)
);

OR2x2_ASAP7_75t_L g16020 ( 
.A(n_15407),
.B(n_15443),
.Y(n_16020)
);

INVx1_ASAP7_75t_L g16021 ( 
.A(n_15789),
.Y(n_16021)
);

INVx1_ASAP7_75t_L g16022 ( 
.A(n_15413),
.Y(n_16022)
);

OAI33xp33_ASAP7_75t_L g16023 ( 
.A1(n_15475),
.A2(n_10982),
.A3(n_10985),
.B1(n_10998),
.B2(n_10986),
.B3(n_10981),
.Y(n_16023)
);

NAND2xp5_ASAP7_75t_SL g16024 ( 
.A(n_15516),
.B(n_8618),
.Y(n_16024)
);

INVx1_ASAP7_75t_L g16025 ( 
.A(n_15791),
.Y(n_16025)
);

NAND2xp5_ASAP7_75t_L g16026 ( 
.A(n_15756),
.B(n_10982),
.Y(n_16026)
);

NAND2xp5_ASAP7_75t_L g16027 ( 
.A(n_15756),
.B(n_10985),
.Y(n_16027)
);

INVx1_ASAP7_75t_L g16028 ( 
.A(n_15791),
.Y(n_16028)
);

NAND2xp5_ASAP7_75t_L g16029 ( 
.A(n_15526),
.B(n_10986),
.Y(n_16029)
);

INVx1_ASAP7_75t_L g16030 ( 
.A(n_15425),
.Y(n_16030)
);

INVx2_ASAP7_75t_L g16031 ( 
.A(n_15678),
.Y(n_16031)
);

NAND2xp5_ASAP7_75t_SL g16032 ( 
.A(n_15432),
.B(n_8618),
.Y(n_16032)
);

INVx2_ASAP7_75t_L g16033 ( 
.A(n_15687),
.Y(n_16033)
);

INVx1_ASAP7_75t_L g16034 ( 
.A(n_15428),
.Y(n_16034)
);

OR2x2_ASAP7_75t_L g16035 ( 
.A(n_15484),
.B(n_10998),
.Y(n_16035)
);

INVx1_ASAP7_75t_L g16036 ( 
.A(n_15410),
.Y(n_16036)
);

INVx1_ASAP7_75t_L g16037 ( 
.A(n_15473),
.Y(n_16037)
);

INVx1_ASAP7_75t_L g16038 ( 
.A(n_15435),
.Y(n_16038)
);

AND2x4_ASAP7_75t_L g16039 ( 
.A(n_15404),
.B(n_15489),
.Y(n_16039)
);

NAND2xp5_ASAP7_75t_L g16040 ( 
.A(n_15542),
.B(n_11004),
.Y(n_16040)
);

INVx1_ASAP7_75t_L g16041 ( 
.A(n_15828),
.Y(n_16041)
);

AND2x2_ASAP7_75t_L g16042 ( 
.A(n_15437),
.B(n_11004),
.Y(n_16042)
);

OAI31xp33_ASAP7_75t_SL g16043 ( 
.A1(n_15722),
.A2(n_11397),
.A3(n_11358),
.B(n_11373),
.Y(n_16043)
);

AND2x2_ASAP7_75t_L g16044 ( 
.A(n_15474),
.B(n_11007),
.Y(n_16044)
);

INVx2_ASAP7_75t_L g16045 ( 
.A(n_15737),
.Y(n_16045)
);

INVx2_ASAP7_75t_L g16046 ( 
.A(n_15744),
.Y(n_16046)
);

NAND2xp5_ASAP7_75t_SL g16047 ( 
.A(n_15429),
.B(n_8618),
.Y(n_16047)
);

BUFx2_ASAP7_75t_L g16048 ( 
.A(n_15709),
.Y(n_16048)
);

NAND2xp5_ASAP7_75t_L g16049 ( 
.A(n_15628),
.B(n_11007),
.Y(n_16049)
);

AND2x2_ASAP7_75t_L g16050 ( 
.A(n_15618),
.B(n_11012),
.Y(n_16050)
);

AND2x2_ASAP7_75t_L g16051 ( 
.A(n_15593),
.B(n_11012),
.Y(n_16051)
);

AND2x4_ASAP7_75t_L g16052 ( 
.A(n_15675),
.B(n_8023),
.Y(n_16052)
);

NAND2xp5_ASAP7_75t_L g16053 ( 
.A(n_15438),
.B(n_11016),
.Y(n_16053)
);

INVx1_ASAP7_75t_L g16054 ( 
.A(n_15828),
.Y(n_16054)
);

INVx1_ASAP7_75t_SL g16055 ( 
.A(n_15485),
.Y(n_16055)
);

BUFx2_ASAP7_75t_L g16056 ( 
.A(n_15738),
.Y(n_16056)
);

AOI21xp5_ASAP7_75t_L g16057 ( 
.A1(n_15766),
.A2(n_11018),
.B(n_11016),
.Y(n_16057)
);

AND2x2_ASAP7_75t_L g16058 ( 
.A(n_15590),
.B(n_15854),
.Y(n_16058)
);

INVx1_ASAP7_75t_L g16059 ( 
.A(n_15571),
.Y(n_16059)
);

NOR3xp33_ASAP7_75t_L g16060 ( 
.A(n_15761),
.B(n_15436),
.C(n_15813),
.Y(n_16060)
);

NAND2xp5_ASAP7_75t_L g16061 ( 
.A(n_15543),
.B(n_11018),
.Y(n_16061)
);

AND2x4_ASAP7_75t_L g16062 ( 
.A(n_15455),
.B(n_8023),
.Y(n_16062)
);

NOR2x1_ASAP7_75t_L g16063 ( 
.A(n_15667),
.B(n_11032),
.Y(n_16063)
);

AND2x4_ASAP7_75t_L g16064 ( 
.A(n_15458),
.B(n_8204),
.Y(n_16064)
);

AND2x2_ASAP7_75t_L g16065 ( 
.A(n_15798),
.B(n_11032),
.Y(n_16065)
);

AND2x2_ASAP7_75t_L g16066 ( 
.A(n_15858),
.B(n_11035),
.Y(n_16066)
);

INVxp67_ASAP7_75t_L g16067 ( 
.A(n_15771),
.Y(n_16067)
);

AND2x4_ASAP7_75t_L g16068 ( 
.A(n_15689),
.B(n_8204),
.Y(n_16068)
);

INVx1_ASAP7_75t_L g16069 ( 
.A(n_15540),
.Y(n_16069)
);

OAI211xp5_ASAP7_75t_SL g16070 ( 
.A1(n_15392),
.A2(n_15600),
.B(n_15663),
.C(n_15746),
.Y(n_16070)
);

INVx1_ASAP7_75t_L g16071 ( 
.A(n_15747),
.Y(n_16071)
);

AND2x4_ASAP7_75t_L g16072 ( 
.A(n_15836),
.B(n_15730),
.Y(n_16072)
);

AND2x2_ASAP7_75t_L g16073 ( 
.A(n_15878),
.B(n_11035),
.Y(n_16073)
);

AND2x2_ASAP7_75t_L g16074 ( 
.A(n_15826),
.B(n_11039),
.Y(n_16074)
);

HB1xp67_ASAP7_75t_L g16075 ( 
.A(n_15755),
.Y(n_16075)
);

OR2x2_ASAP7_75t_L g16076 ( 
.A(n_15617),
.B(n_11039),
.Y(n_16076)
);

AND2x2_ASAP7_75t_L g16077 ( 
.A(n_15840),
.B(n_11045),
.Y(n_16077)
);

OR2x2_ASAP7_75t_L g16078 ( 
.A(n_15409),
.B(n_11045),
.Y(n_16078)
);

INVx1_ASAP7_75t_L g16079 ( 
.A(n_15748),
.Y(n_16079)
);

NAND2xp5_ASAP7_75t_L g16080 ( 
.A(n_15558),
.B(n_11046),
.Y(n_16080)
);

NOR2xp33_ASAP7_75t_L g16081 ( 
.A(n_15655),
.B(n_11046),
.Y(n_16081)
);

AND2x2_ASAP7_75t_L g16082 ( 
.A(n_15850),
.B(n_15876),
.Y(n_16082)
);

INVx1_ASAP7_75t_L g16083 ( 
.A(n_15775),
.Y(n_16083)
);

AND2x4_ASAP7_75t_L g16084 ( 
.A(n_15887),
.B(n_8204),
.Y(n_16084)
);

INVx1_ASAP7_75t_L g16085 ( 
.A(n_15824),
.Y(n_16085)
);

AND2x2_ASAP7_75t_L g16086 ( 
.A(n_15453),
.B(n_11047),
.Y(n_16086)
);

INVx1_ASAP7_75t_L g16087 ( 
.A(n_15860),
.Y(n_16087)
);

NAND2xp5_ASAP7_75t_L g16088 ( 
.A(n_15577),
.B(n_11047),
.Y(n_16088)
);

INVx1_ASAP7_75t_L g16089 ( 
.A(n_15496),
.Y(n_16089)
);

AND2x2_ASAP7_75t_L g16090 ( 
.A(n_15704),
.B(n_11051),
.Y(n_16090)
);

AND2x2_ASAP7_75t_L g16091 ( 
.A(n_15724),
.B(n_11051),
.Y(n_16091)
);

AND2x2_ASAP7_75t_L g16092 ( 
.A(n_15905),
.B(n_11055),
.Y(n_16092)
);

OAI22xp5_ASAP7_75t_L g16093 ( 
.A1(n_15769),
.A2(n_8523),
.B1(n_8583),
.B2(n_8445),
.Y(n_16093)
);

OR2x2_ASAP7_75t_L g16094 ( 
.A(n_15486),
.B(n_11055),
.Y(n_16094)
);

INVx1_ASAP7_75t_SL g16095 ( 
.A(n_15512),
.Y(n_16095)
);

NAND2xp5_ASAP7_75t_L g16096 ( 
.A(n_15657),
.B(n_11063),
.Y(n_16096)
);

AND2x4_ASAP7_75t_SL g16097 ( 
.A(n_15897),
.B(n_5370),
.Y(n_16097)
);

AND2x2_ASAP7_75t_L g16098 ( 
.A(n_15750),
.B(n_11063),
.Y(n_16098)
);

NAND2xp5_ASAP7_75t_L g16099 ( 
.A(n_15477),
.B(n_11064),
.Y(n_16099)
);

OR2x2_ASAP7_75t_L g16100 ( 
.A(n_15701),
.B(n_11064),
.Y(n_16100)
);

AND2x2_ASAP7_75t_L g16101 ( 
.A(n_15765),
.B(n_11065),
.Y(n_16101)
);

NOR3xp33_ASAP7_75t_L g16102 ( 
.A(n_15807),
.B(n_8962),
.C(n_9019),
.Y(n_16102)
);

INVxp67_ASAP7_75t_L g16103 ( 
.A(n_15447),
.Y(n_16103)
);

BUFx3_ASAP7_75t_L g16104 ( 
.A(n_15723),
.Y(n_16104)
);

INVx2_ASAP7_75t_L g16105 ( 
.A(n_15649),
.Y(n_16105)
);

AND2x2_ASAP7_75t_L g16106 ( 
.A(n_15891),
.B(n_15892),
.Y(n_16106)
);

INVx2_ASAP7_75t_L g16107 ( 
.A(n_15503),
.Y(n_16107)
);

NAND2xp5_ASAP7_75t_L g16108 ( 
.A(n_15479),
.B(n_11065),
.Y(n_16108)
);

OR2x2_ASAP7_75t_L g16109 ( 
.A(n_15444),
.B(n_11067),
.Y(n_16109)
);

INVx1_ASAP7_75t_L g16110 ( 
.A(n_15417),
.Y(n_16110)
);

AND2x2_ASAP7_75t_L g16111 ( 
.A(n_15898),
.B(n_11067),
.Y(n_16111)
);

AND2x4_ASAP7_75t_L g16112 ( 
.A(n_15714),
.B(n_8445),
.Y(n_16112)
);

AND2x2_ASAP7_75t_L g16113 ( 
.A(n_15809),
.B(n_11078),
.Y(n_16113)
);

OR2x2_ASAP7_75t_L g16114 ( 
.A(n_15439),
.B(n_11078),
.Y(n_16114)
);

NAND2xp5_ASAP7_75t_L g16115 ( 
.A(n_15497),
.B(n_11080),
.Y(n_16115)
);

AND2x2_ASAP7_75t_L g16116 ( 
.A(n_15834),
.B(n_11080),
.Y(n_16116)
);

OR2x2_ASAP7_75t_L g16117 ( 
.A(n_15422),
.B(n_11089),
.Y(n_16117)
);

INVx1_ASAP7_75t_L g16118 ( 
.A(n_15399),
.Y(n_16118)
);

INVx1_ASAP7_75t_L g16119 ( 
.A(n_15504),
.Y(n_16119)
);

INVx2_ASAP7_75t_L g16120 ( 
.A(n_15862),
.Y(n_16120)
);

INVx1_ASAP7_75t_L g16121 ( 
.A(n_15614),
.Y(n_16121)
);

INVx2_ASAP7_75t_L g16122 ( 
.A(n_15862),
.Y(n_16122)
);

NAND2xp5_ASAP7_75t_L g16123 ( 
.A(n_15774),
.B(n_11089),
.Y(n_16123)
);

NOR3xp33_ASAP7_75t_L g16124 ( 
.A(n_15529),
.B(n_8962),
.C(n_11169),
.Y(n_16124)
);

AND2x2_ASAP7_75t_L g16125 ( 
.A(n_15773),
.B(n_11097),
.Y(n_16125)
);

AND2x2_ASAP7_75t_L g16126 ( 
.A(n_15833),
.B(n_11097),
.Y(n_16126)
);

INVx1_ASAP7_75t_L g16127 ( 
.A(n_15427),
.Y(n_16127)
);

INVx5_ASAP7_75t_L g16128 ( 
.A(n_15764),
.Y(n_16128)
);

HB1xp67_ASAP7_75t_L g16129 ( 
.A(n_15764),
.Y(n_16129)
);

INVx1_ASAP7_75t_L g16130 ( 
.A(n_15513),
.Y(n_16130)
);

AND2x2_ASAP7_75t_L g16131 ( 
.A(n_15838),
.B(n_15770),
.Y(n_16131)
);

AND2x2_ASAP7_75t_L g16132 ( 
.A(n_15433),
.B(n_11100),
.Y(n_16132)
);

INVx2_ASAP7_75t_L g16133 ( 
.A(n_15764),
.Y(n_16133)
);

XNOR2xp5_ASAP7_75t_L g16134 ( 
.A(n_15795),
.B(n_8236),
.Y(n_16134)
);

INVx1_ASAP7_75t_L g16135 ( 
.A(n_15514),
.Y(n_16135)
);

AND2x4_ASAP7_75t_L g16136 ( 
.A(n_15788),
.B(n_8445),
.Y(n_16136)
);

INVx1_ASAP7_75t_L g16137 ( 
.A(n_15518),
.Y(n_16137)
);

NAND2xp5_ASAP7_75t_SL g16138 ( 
.A(n_15728),
.B(n_8633),
.Y(n_16138)
);

NAND2xp5_ASAP7_75t_L g16139 ( 
.A(n_15520),
.B(n_15528),
.Y(n_16139)
);

NOR2xp33_ASAP7_75t_SL g16140 ( 
.A(n_15728),
.B(n_5370),
.Y(n_16140)
);

INVx1_ASAP7_75t_L g16141 ( 
.A(n_15423),
.Y(n_16141)
);

AND2x2_ASAP7_75t_L g16142 ( 
.A(n_15713),
.B(n_11100),
.Y(n_16142)
);

NAND3xp33_ASAP7_75t_SL g16143 ( 
.A(n_15802),
.B(n_8646),
.C(n_8417),
.Y(n_16143)
);

NAND2xp5_ASAP7_75t_L g16144 ( 
.A(n_15751),
.B(n_11106),
.Y(n_16144)
);

OR2x2_ASAP7_75t_L g16145 ( 
.A(n_15538),
.B(n_11106),
.Y(n_16145)
);

AND2x2_ASAP7_75t_L g16146 ( 
.A(n_15585),
.B(n_11108),
.Y(n_16146)
);

INVx1_ASAP7_75t_L g16147 ( 
.A(n_15424),
.Y(n_16147)
);

AND2x2_ASAP7_75t_L g16148 ( 
.A(n_15808),
.B(n_11108),
.Y(n_16148)
);

OR2x2_ASAP7_75t_L g16149 ( 
.A(n_15545),
.B(n_11110),
.Y(n_16149)
);

BUFx2_ASAP7_75t_L g16150 ( 
.A(n_15857),
.Y(n_16150)
);

INVx2_ASAP7_75t_L g16151 ( 
.A(n_15837),
.Y(n_16151)
);

NAND2xp5_ASAP7_75t_L g16152 ( 
.A(n_15556),
.B(n_11110),
.Y(n_16152)
);

INVx1_ASAP7_75t_L g16153 ( 
.A(n_15430),
.Y(n_16153)
);

INVx1_ASAP7_75t_L g16154 ( 
.A(n_15539),
.Y(n_16154)
);

INVx1_ASAP7_75t_SL g16155 ( 
.A(n_15654),
.Y(n_16155)
);

AOI22xp5_ASAP7_75t_L g16156 ( 
.A1(n_15911),
.A2(n_8642),
.B1(n_8644),
.B2(n_8633),
.Y(n_16156)
);

INVx1_ASAP7_75t_L g16157 ( 
.A(n_15421),
.Y(n_16157)
);

INVx1_ASAP7_75t_L g16158 ( 
.A(n_15608),
.Y(n_16158)
);

INVx1_ASAP7_75t_L g16159 ( 
.A(n_15550),
.Y(n_16159)
);

INVx1_ASAP7_75t_L g16160 ( 
.A(n_15488),
.Y(n_16160)
);

INVx1_ASAP7_75t_L g16161 ( 
.A(n_15493),
.Y(n_16161)
);

NAND2xp5_ASAP7_75t_L g16162 ( 
.A(n_15552),
.B(n_11117),
.Y(n_16162)
);

NOR2x1_ASAP7_75t_L g16163 ( 
.A(n_15904),
.B(n_11117),
.Y(n_16163)
);

NAND2xp5_ASAP7_75t_L g16164 ( 
.A(n_15640),
.B(n_11121),
.Y(n_16164)
);

AND2x2_ASAP7_75t_L g16165 ( 
.A(n_15660),
.B(n_11121),
.Y(n_16165)
);

INVx1_ASAP7_75t_L g16166 ( 
.A(n_15643),
.Y(n_16166)
);

AND2x4_ASAP7_75t_SL g16167 ( 
.A(n_15597),
.B(n_8861),
.Y(n_16167)
);

INVx2_ASAP7_75t_L g16168 ( 
.A(n_15611),
.Y(n_16168)
);

AND2x2_ASAP7_75t_L g16169 ( 
.A(n_15779),
.B(n_15598),
.Y(n_16169)
);

NAND2xp5_ASAP7_75t_L g16170 ( 
.A(n_15801),
.B(n_11124),
.Y(n_16170)
);

OAI21xp5_ASAP7_75t_L g16171 ( 
.A1(n_15812),
.A2(n_11191),
.B(n_11173),
.Y(n_16171)
);

INVx2_ASAP7_75t_L g16172 ( 
.A(n_15852),
.Y(n_16172)
);

OR2x2_ASAP7_75t_L g16173 ( 
.A(n_15636),
.B(n_11124),
.Y(n_16173)
);

INVx1_ASAP7_75t_L g16174 ( 
.A(n_15603),
.Y(n_16174)
);

AND2x2_ASAP7_75t_L g16175 ( 
.A(n_15720),
.B(n_11129),
.Y(n_16175)
);

NAND2xp5_ASAP7_75t_L g16176 ( 
.A(n_15819),
.B(n_11129),
.Y(n_16176)
);

INVx3_ASAP7_75t_L g16177 ( 
.A(n_15592),
.Y(n_16177)
);

AND2x2_ASAP7_75t_L g16178 ( 
.A(n_15753),
.B(n_11136),
.Y(n_16178)
);

INVxp67_ASAP7_75t_L g16179 ( 
.A(n_15511),
.Y(n_16179)
);

OR2x2_ASAP7_75t_L g16180 ( 
.A(n_15638),
.B(n_11136),
.Y(n_16180)
);

NAND2x1p5_ASAP7_75t_L g16181 ( 
.A(n_15832),
.B(n_8633),
.Y(n_16181)
);

INVx1_ASAP7_75t_L g16182 ( 
.A(n_15632),
.Y(n_16182)
);

INVx2_ASAP7_75t_L g16183 ( 
.A(n_15877),
.Y(n_16183)
);

OR2x2_ASAP7_75t_L g16184 ( 
.A(n_15639),
.B(n_11144),
.Y(n_16184)
);

AND2x2_ASAP7_75t_L g16185 ( 
.A(n_15762),
.B(n_11144),
.Y(n_16185)
);

OR2x2_ASAP7_75t_L g16186 ( 
.A(n_15624),
.B(n_11148),
.Y(n_16186)
);

NAND2xp5_ASAP7_75t_L g16187 ( 
.A(n_15588),
.B(n_11148),
.Y(n_16187)
);

NOR2xp33_ASAP7_75t_L g16188 ( 
.A(n_15440),
.B(n_11154),
.Y(n_16188)
);

INVxp33_ASAP7_75t_L g16189 ( 
.A(n_15586),
.Y(n_16189)
);

INVx1_ASAP7_75t_L g16190 ( 
.A(n_15544),
.Y(n_16190)
);

NAND2xp5_ASAP7_75t_L g16191 ( 
.A(n_15613),
.B(n_15861),
.Y(n_16191)
);

AND2x2_ASAP7_75t_L g16192 ( 
.A(n_15685),
.B(n_15690),
.Y(n_16192)
);

NAND2xp5_ASAP7_75t_L g16193 ( 
.A(n_15863),
.B(n_11154),
.Y(n_16193)
);

AND2x2_ASAP7_75t_L g16194 ( 
.A(n_15692),
.B(n_11155),
.Y(n_16194)
);

NOR2xp33_ASAP7_75t_L g16195 ( 
.A(n_15867),
.B(n_11155),
.Y(n_16195)
);

INVx1_ASAP7_75t_L g16196 ( 
.A(n_15547),
.Y(n_16196)
);

INVx2_ASAP7_75t_L g16197 ( 
.A(n_15553),
.Y(n_16197)
);

OR2x2_ASAP7_75t_L g16198 ( 
.A(n_15415),
.B(n_11158),
.Y(n_16198)
);

NAND2xp5_ASAP7_75t_L g16199 ( 
.A(n_15612),
.B(n_11158),
.Y(n_16199)
);

INVx1_ASAP7_75t_L g16200 ( 
.A(n_15631),
.Y(n_16200)
);

OR2x6_ASAP7_75t_L g16201 ( 
.A(n_15602),
.B(n_6162),
.Y(n_16201)
);

OA21x2_ASAP7_75t_L g16202 ( 
.A1(n_15814),
.A2(n_11166),
.B(n_11161),
.Y(n_16202)
);

AND2x2_ASAP7_75t_L g16203 ( 
.A(n_15621),
.B(n_15671),
.Y(n_16203)
);

AND2x2_ASAP7_75t_L g16204 ( 
.A(n_15708),
.B(n_11161),
.Y(n_16204)
);

AND2x2_ASAP7_75t_L g16205 ( 
.A(n_15666),
.B(n_11166),
.Y(n_16205)
);

AND2x2_ASAP7_75t_L g16206 ( 
.A(n_15620),
.B(n_11168),
.Y(n_16206)
);

HB1xp67_ASAP7_75t_L g16207 ( 
.A(n_15866),
.Y(n_16207)
);

INVx2_ASAP7_75t_L g16208 ( 
.A(n_15676),
.Y(n_16208)
);

AND2x2_ASAP7_75t_L g16209 ( 
.A(n_15706),
.B(n_11168),
.Y(n_16209)
);

INVx2_ASAP7_75t_L g16210 ( 
.A(n_15521),
.Y(n_16210)
);

AND2x2_ASAP7_75t_L g16211 ( 
.A(n_15684),
.B(n_11172),
.Y(n_16211)
);

NAND2xp5_ASAP7_75t_L g16212 ( 
.A(n_15626),
.B(n_15627),
.Y(n_16212)
);

INVx1_ASAP7_75t_L g16213 ( 
.A(n_15668),
.Y(n_16213)
);

HB1xp67_ASAP7_75t_L g16214 ( 
.A(n_15785),
.Y(n_16214)
);

AND2x2_ASAP7_75t_L g16215 ( 
.A(n_15615),
.B(n_11172),
.Y(n_16215)
);

INVx6_ASAP7_75t_L g16216 ( 
.A(n_15494),
.Y(n_16216)
);

NAND2xp5_ASAP7_75t_L g16217 ( 
.A(n_15645),
.B(n_11175),
.Y(n_16217)
);

NAND4xp25_ASAP7_75t_L g16218 ( 
.A(n_15561),
.B(n_6662),
.C(n_6718),
.D(n_6717),
.Y(n_16218)
);

INVx2_ASAP7_75t_L g16219 ( 
.A(n_15535),
.Y(n_16219)
);

INVx1_ASAP7_75t_L g16220 ( 
.A(n_15495),
.Y(n_16220)
);

INVx1_ASAP7_75t_L g16221 ( 
.A(n_15651),
.Y(n_16221)
);

AND2x4_ASAP7_75t_SL g16222 ( 
.A(n_15907),
.B(n_8896),
.Y(n_16222)
);

OR2x2_ASAP7_75t_L g16223 ( 
.A(n_15718),
.B(n_11175),
.Y(n_16223)
);

AND2x2_ASAP7_75t_L g16224 ( 
.A(n_15650),
.B(n_11181),
.Y(n_16224)
);

INVx2_ASAP7_75t_L g16225 ( 
.A(n_15578),
.Y(n_16225)
);

INVx2_ASAP7_75t_L g16226 ( 
.A(n_15583),
.Y(n_16226)
);

INVx1_ASAP7_75t_L g16227 ( 
.A(n_15563),
.Y(n_16227)
);

AND2x2_ASAP7_75t_L g16228 ( 
.A(n_15625),
.B(n_11181),
.Y(n_16228)
);

AND2x2_ASAP7_75t_L g16229 ( 
.A(n_15717),
.B(n_11185),
.Y(n_16229)
);

INVx2_ASAP7_75t_L g16230 ( 
.A(n_15591),
.Y(n_16230)
);

AND2x2_ASAP7_75t_L g16231 ( 
.A(n_15537),
.B(n_15541),
.Y(n_16231)
);

OR2x2_ASAP7_75t_L g16232 ( 
.A(n_15825),
.B(n_11185),
.Y(n_16232)
);

NOR2xp33_ASAP7_75t_SL g16233 ( 
.A(n_15870),
.B(n_6922),
.Y(n_16233)
);

OAI321xp33_ASAP7_75t_L g16234 ( 
.A1(n_15596),
.A2(n_8432),
.A3(n_8236),
.B1(n_8004),
.B2(n_8421),
.C(n_8633),
.Y(n_16234)
);

OR2x2_ASAP7_75t_L g16235 ( 
.A(n_15767),
.B(n_15498),
.Y(n_16235)
);

AND2x2_ASAP7_75t_L g16236 ( 
.A(n_15604),
.B(n_15605),
.Y(n_16236)
);

AOI22xp5_ASAP7_75t_L g16237 ( 
.A1(n_15487),
.A2(n_8642),
.B1(n_8644),
.B2(n_8633),
.Y(n_16237)
);

NAND2x1_ASAP7_75t_L g16238 ( 
.A(n_15606),
.B(n_11188),
.Y(n_16238)
);

INVx1_ASAP7_75t_L g16239 ( 
.A(n_15564),
.Y(n_16239)
);

AOI21xp5_ASAP7_75t_L g16240 ( 
.A1(n_15699),
.A2(n_11193),
.B(n_11188),
.Y(n_16240)
);

NAND2xp5_ASAP7_75t_L g16241 ( 
.A(n_15658),
.B(n_11193),
.Y(n_16241)
);

AND2x2_ASAP7_75t_L g16242 ( 
.A(n_15725),
.B(n_11198),
.Y(n_16242)
);

INVx2_ASAP7_75t_L g16243 ( 
.A(n_15534),
.Y(n_16243)
);

AND2x2_ASAP7_75t_L g16244 ( 
.A(n_15803),
.B(n_11198),
.Y(n_16244)
);

AO221x2_ASAP7_75t_L g16245 ( 
.A1(n_15792),
.A2(n_9820),
.B1(n_9818),
.B2(n_11206),
.C(n_11200),
.Y(n_16245)
);

NAND2xp5_ASAP7_75t_L g16246 ( 
.A(n_15853),
.B(n_15856),
.Y(n_16246)
);

NAND2xp5_ASAP7_75t_L g16247 ( 
.A(n_15885),
.B(n_11200),
.Y(n_16247)
);

OR2x2_ASAP7_75t_L g16248 ( 
.A(n_15726),
.B(n_11206),
.Y(n_16248)
);

NOR2x1p5_ASAP7_75t_L g16249 ( 
.A(n_15835),
.B(n_7882),
.Y(n_16249)
);

AOI22xp5_ASAP7_75t_L g16250 ( 
.A1(n_15507),
.A2(n_8642),
.B1(n_8644),
.B2(n_8633),
.Y(n_16250)
);

NAND2xp5_ASAP7_75t_L g16251 ( 
.A(n_15888),
.B(n_11209),
.Y(n_16251)
);

AND2x2_ASAP7_75t_SL g16252 ( 
.A(n_15796),
.B(n_7831),
.Y(n_16252)
);

INVx2_ASAP7_75t_L g16253 ( 
.A(n_15584),
.Y(n_16253)
);

INVx1_ASAP7_75t_L g16254 ( 
.A(n_15595),
.Y(n_16254)
);

INVx1_ASAP7_75t_L g16255 ( 
.A(n_15533),
.Y(n_16255)
);

OR2x2_ASAP7_75t_L g16256 ( 
.A(n_15752),
.B(n_11209),
.Y(n_16256)
);

NAND2xp5_ASAP7_75t_L g16257 ( 
.A(n_15912),
.B(n_11211),
.Y(n_16257)
);

OR2x2_ASAP7_75t_L g16258 ( 
.A(n_15895),
.B(n_11211),
.Y(n_16258)
);

INVx1_ASAP7_75t_L g16259 ( 
.A(n_15599),
.Y(n_16259)
);

INVxp67_ASAP7_75t_SL g16260 ( 
.A(n_15712),
.Y(n_16260)
);

OR2x2_ASAP7_75t_L g16261 ( 
.A(n_15506),
.B(n_11217),
.Y(n_16261)
);

BUFx2_ASAP7_75t_L g16262 ( 
.A(n_15560),
.Y(n_16262)
);

NAND2xp5_ASAP7_75t_L g16263 ( 
.A(n_15915),
.B(n_11217),
.Y(n_16263)
);

INVx2_ASAP7_75t_L g16264 ( 
.A(n_15610),
.Y(n_16264)
);

INVx1_ASAP7_75t_SL g16265 ( 
.A(n_15616),
.Y(n_16265)
);

AND2x2_ASAP7_75t_L g16266 ( 
.A(n_15642),
.B(n_11222),
.Y(n_16266)
);

BUFx4f_ASAP7_75t_SL g16267 ( 
.A(n_15800),
.Y(n_16267)
);

OAI21x1_ASAP7_75t_L g16268 ( 
.A1(n_15515),
.A2(n_11231),
.B(n_11222),
.Y(n_16268)
);

AND2x2_ASAP7_75t_L g16269 ( 
.A(n_15648),
.B(n_11231),
.Y(n_16269)
);

AND2x2_ASAP7_75t_L g16270 ( 
.A(n_15634),
.B(n_11244),
.Y(n_16270)
);

INVx1_ASAP7_75t_L g16271 ( 
.A(n_15549),
.Y(n_16271)
);

OAI33xp33_ASAP7_75t_L g16272 ( 
.A1(n_15729),
.A2(n_11247),
.A3(n_11250),
.B1(n_11264),
.B2(n_11258),
.B3(n_11244),
.Y(n_16272)
);

AND2x2_ASAP7_75t_SL g16273 ( 
.A(n_15868),
.B(n_7831),
.Y(n_16273)
);

NAND2xp5_ASAP7_75t_L g16274 ( 
.A(n_15732),
.B(n_11247),
.Y(n_16274)
);

OR2x2_ASAP7_75t_L g16275 ( 
.A(n_15697),
.B(n_11250),
.Y(n_16275)
);

INVx1_ASAP7_75t_L g16276 ( 
.A(n_15680),
.Y(n_16276)
);

AND2x4_ASAP7_75t_L g16277 ( 
.A(n_15745),
.B(n_8523),
.Y(n_16277)
);

NAND2xp5_ASAP7_75t_L g16278 ( 
.A(n_15510),
.B(n_11258),
.Y(n_16278)
);

INVxp67_ASAP7_75t_L g16279 ( 
.A(n_15622),
.Y(n_16279)
);

INVx1_ASAP7_75t_L g16280 ( 
.A(n_15682),
.Y(n_16280)
);

AND2x2_ASAP7_75t_L g16281 ( 
.A(n_15517),
.B(n_11264),
.Y(n_16281)
);

NAND2xp5_ASAP7_75t_L g16282 ( 
.A(n_15566),
.B(n_11277),
.Y(n_16282)
);

AND2x4_ASAP7_75t_SL g16283 ( 
.A(n_15601),
.B(n_15629),
.Y(n_16283)
);

AND2x2_ASAP7_75t_L g16284 ( 
.A(n_15568),
.B(n_11277),
.Y(n_16284)
);

NAND2xp5_ASAP7_75t_L g16285 ( 
.A(n_15573),
.B(n_15662),
.Y(n_16285)
);

INVx2_ASAP7_75t_L g16286 ( 
.A(n_15527),
.Y(n_16286)
);

INVx1_ASAP7_75t_L g16287 ( 
.A(n_15672),
.Y(n_16287)
);

INVx2_ASAP7_75t_SL g16288 ( 
.A(n_15646),
.Y(n_16288)
);

NOR3xp33_ASAP7_75t_L g16289 ( 
.A(n_15804),
.B(n_11191),
.C(n_11173),
.Y(n_16289)
);

NAND2x1_ASAP7_75t_SL g16290 ( 
.A(n_15633),
.B(n_9072),
.Y(n_16290)
);

AND2x2_ASAP7_75t_L g16291 ( 
.A(n_15630),
.B(n_11278),
.Y(n_16291)
);

OR2x2_ASAP7_75t_L g16292 ( 
.A(n_15619),
.B(n_11278),
.Y(n_16292)
);

OR2x2_ASAP7_75t_L g16293 ( 
.A(n_15759),
.B(n_11280),
.Y(n_16293)
);

HB1xp67_ASAP7_75t_L g16294 ( 
.A(n_15548),
.Y(n_16294)
);

INVxp67_ASAP7_75t_L g16295 ( 
.A(n_15711),
.Y(n_16295)
);

INVx1_ASAP7_75t_L g16296 ( 
.A(n_15570),
.Y(n_16296)
);

INVx2_ASAP7_75t_SL g16297 ( 
.A(n_15674),
.Y(n_16297)
);

AND2x2_ASAP7_75t_L g16298 ( 
.A(n_15757),
.B(n_11280),
.Y(n_16298)
);

INVx1_ASAP7_75t_L g16299 ( 
.A(n_15580),
.Y(n_16299)
);

OR2x2_ASAP7_75t_L g16300 ( 
.A(n_15519),
.B(n_11282),
.Y(n_16300)
);

INVx1_ASAP7_75t_L g16301 ( 
.A(n_15581),
.Y(n_16301)
);

AND2x2_ASAP7_75t_L g16302 ( 
.A(n_15760),
.B(n_11282),
.Y(n_16302)
);

AND2x2_ASAP7_75t_L g16303 ( 
.A(n_15768),
.B(n_11285),
.Y(n_16303)
);

INVxp33_ASAP7_75t_L g16304 ( 
.A(n_15831),
.Y(n_16304)
);

AND2x2_ASAP7_75t_L g16305 ( 
.A(n_15777),
.B(n_11285),
.Y(n_16305)
);

AND2x2_ASAP7_75t_L g16306 ( 
.A(n_15821),
.B(n_11286),
.Y(n_16306)
);

NAND2xp5_ASAP7_75t_L g16307 ( 
.A(n_15673),
.B(n_11286),
.Y(n_16307)
);

OR2x2_ASAP7_75t_L g16308 ( 
.A(n_15522),
.B(n_11287),
.Y(n_16308)
);

AND2x4_ASAP7_75t_L g16309 ( 
.A(n_15827),
.B(n_8523),
.Y(n_16309)
);

INVx2_ASAP7_75t_SL g16310 ( 
.A(n_15758),
.Y(n_16310)
);

NAND2xp5_ASAP7_75t_L g16311 ( 
.A(n_15677),
.B(n_11287),
.Y(n_16311)
);

NAND2xp5_ASAP7_75t_L g16312 ( 
.A(n_15741),
.B(n_9313),
.Y(n_16312)
);

HB1xp67_ASAP7_75t_L g16313 ( 
.A(n_15587),
.Y(n_16313)
);

NAND4xp25_ASAP7_75t_L g16314 ( 
.A(n_15576),
.B(n_15582),
.C(n_15500),
.D(n_15502),
.Y(n_16314)
);

AND2x2_ASAP7_75t_L g16315 ( 
.A(n_15754),
.B(n_11028),
.Y(n_16315)
);

OR2x2_ASAP7_75t_L g16316 ( 
.A(n_15569),
.B(n_9314),
.Y(n_16316)
);

INVx2_ASAP7_75t_L g16317 ( 
.A(n_15742),
.Y(n_16317)
);

AND2x2_ASAP7_75t_L g16318 ( 
.A(n_15805),
.B(n_11028),
.Y(n_16318)
);

AND2x2_ASAP7_75t_L g16319 ( 
.A(n_15635),
.B(n_11038),
.Y(n_16319)
);

AND2x2_ASAP7_75t_L g16320 ( 
.A(n_15653),
.B(n_11038),
.Y(n_16320)
);

OR2x2_ASAP7_75t_L g16321 ( 
.A(n_15656),
.B(n_9314),
.Y(n_16321)
);

INVx1_ASAP7_75t_L g16322 ( 
.A(n_15705),
.Y(n_16322)
);

NAND2xp5_ASAP7_75t_L g16323 ( 
.A(n_15790),
.B(n_9313),
.Y(n_16323)
);

INVxp67_ASAP7_75t_L g16324 ( 
.A(n_15688),
.Y(n_16324)
);

NAND2xp5_ASAP7_75t_L g16325 ( 
.A(n_15691),
.B(n_9329),
.Y(n_16325)
);

AND2x2_ASAP7_75t_L g16326 ( 
.A(n_15693),
.B(n_11091),
.Y(n_16326)
);

AND2x4_ASAP7_75t_L g16327 ( 
.A(n_15829),
.B(n_8583),
.Y(n_16327)
);

INVx1_ASAP7_75t_L g16328 ( 
.A(n_15781),
.Y(n_16328)
);

OR2x2_ASAP7_75t_L g16329 ( 
.A(n_15609),
.B(n_9314),
.Y(n_16329)
);

OR2x2_ASAP7_75t_L g16330 ( 
.A(n_15669),
.B(n_9314),
.Y(n_16330)
);

OR2x2_ASAP7_75t_L g16331 ( 
.A(n_15670),
.B(n_9317),
.Y(n_16331)
);

OR2x2_ASAP7_75t_L g16332 ( 
.A(n_15562),
.B(n_9317),
.Y(n_16332)
);

AOI21xp5_ASAP7_75t_L g16333 ( 
.A1(n_15491),
.A2(n_10653),
.B(n_10647),
.Y(n_16333)
);

HB1xp67_ASAP7_75t_L g16334 ( 
.A(n_15743),
.Y(n_16334)
);

OR2x2_ASAP7_75t_L g16335 ( 
.A(n_15567),
.B(n_9317),
.Y(n_16335)
);

AND2x4_ASAP7_75t_L g16336 ( 
.A(n_15859),
.B(n_8583),
.Y(n_16336)
);

AND2x2_ASAP7_75t_L g16337 ( 
.A(n_15694),
.B(n_11091),
.Y(n_16337)
);

AND2x2_ASAP7_75t_L g16338 ( 
.A(n_15700),
.B(n_11093),
.Y(n_16338)
);

NAND2xp5_ASAP7_75t_L g16339 ( 
.A(n_15702),
.B(n_9329),
.Y(n_16339)
);

NAND2xp5_ASAP7_75t_L g16340 ( 
.A(n_15703),
.B(n_9330),
.Y(n_16340)
);

OR2x2_ASAP7_75t_L g16341 ( 
.A(n_15659),
.B(n_9317),
.Y(n_16341)
);

OR2x2_ASAP7_75t_L g16342 ( 
.A(n_15665),
.B(n_8450),
.Y(n_16342)
);

INVx1_ASAP7_75t_L g16343 ( 
.A(n_15707),
.Y(n_16343)
);

HB1xp67_ASAP7_75t_L g16344 ( 
.A(n_15735),
.Y(n_16344)
);

AND2x2_ASAP7_75t_L g16345 ( 
.A(n_15710),
.B(n_11093),
.Y(n_16345)
);

INVx1_ASAP7_75t_L g16346 ( 
.A(n_15679),
.Y(n_16346)
);

INVx1_ASAP7_75t_L g16347 ( 
.A(n_15681),
.Y(n_16347)
);

NAND2xp5_ASAP7_75t_L g16348 ( 
.A(n_15873),
.B(n_9330),
.Y(n_16348)
);

INVx1_ASAP7_75t_SL g16349 ( 
.A(n_15787),
.Y(n_16349)
);

INVxp67_ASAP7_75t_SL g16350 ( 
.A(n_15683),
.Y(n_16350)
);

AND2x4_ASAP7_75t_L g16351 ( 
.A(n_15846),
.B(n_8827),
.Y(n_16351)
);

NAND2xp5_ASAP7_75t_L g16352 ( 
.A(n_15916),
.B(n_9335),
.Y(n_16352)
);

AND2x2_ASAP7_75t_L g16353 ( 
.A(n_15851),
.B(n_15874),
.Y(n_16353)
);

OR2x2_ASAP7_75t_L g16354 ( 
.A(n_15778),
.B(n_8458),
.Y(n_16354)
);

NAND2xp5_ASAP7_75t_SL g16355 ( 
.A(n_15890),
.B(n_8633),
.Y(n_16355)
);

OR2x2_ASAP7_75t_L g16356 ( 
.A(n_15695),
.B(n_8458),
.Y(n_16356)
);

AND2x2_ASAP7_75t_L g16357 ( 
.A(n_15881),
.B(n_10647),
.Y(n_16357)
);

NAND2xp5_ASAP7_75t_L g16358 ( 
.A(n_15908),
.B(n_9335),
.Y(n_16358)
);

NAND2xp5_ASAP7_75t_L g16359 ( 
.A(n_15909),
.B(n_15806),
.Y(n_16359)
);

NAND2xp5_ASAP7_75t_L g16360 ( 
.A(n_15811),
.B(n_9338),
.Y(n_16360)
);

NAND2xp5_ASAP7_75t_L g16361 ( 
.A(n_15816),
.B(n_9338),
.Y(n_16361)
);

INVx2_ASAP7_75t_L g16362 ( 
.A(n_15763),
.Y(n_16362)
);

AND2x2_ASAP7_75t_L g16363 ( 
.A(n_15739),
.B(n_10277),
.Y(n_16363)
);

INVx1_ASAP7_75t_SL g16364 ( 
.A(n_15843),
.Y(n_16364)
);

INVx2_ASAP7_75t_L g16365 ( 
.A(n_15793),
.Y(n_16365)
);

INVx1_ASAP7_75t_L g16366 ( 
.A(n_15698),
.Y(n_16366)
);

OR2x2_ASAP7_75t_L g16367 ( 
.A(n_15879),
.B(n_7626),
.Y(n_16367)
);

AND2x2_ASAP7_75t_L g16368 ( 
.A(n_15917),
.B(n_10277),
.Y(n_16368)
);

AND2x4_ASAP7_75t_SL g16369 ( 
.A(n_15820),
.B(n_8896),
.Y(n_16369)
);

AND2x2_ASAP7_75t_L g16370 ( 
.A(n_15749),
.B(n_10277),
.Y(n_16370)
);

NAND2xp5_ASAP7_75t_L g16371 ( 
.A(n_15848),
.B(n_9339),
.Y(n_16371)
);

OR2x2_ASAP7_75t_L g16372 ( 
.A(n_15884),
.B(n_7626),
.Y(n_16372)
);

AND2x2_ASAP7_75t_L g16373 ( 
.A(n_15731),
.B(n_7882),
.Y(n_16373)
);

INVx2_ASAP7_75t_L g16374 ( 
.A(n_15794),
.Y(n_16374)
);

NAND2xp5_ASAP7_75t_L g16375 ( 
.A(n_15721),
.B(n_9339),
.Y(n_16375)
);

AND2x2_ASAP7_75t_SL g16376 ( 
.A(n_15784),
.B(n_7831),
.Y(n_16376)
);

NAND2xp5_ASAP7_75t_L g16377 ( 
.A(n_15740),
.B(n_9342),
.Y(n_16377)
);

AND2x2_ASAP7_75t_L g16378 ( 
.A(n_15733),
.B(n_7882),
.Y(n_16378)
);

OR2x2_ASAP7_75t_L g16379 ( 
.A(n_15900),
.B(n_7626),
.Y(n_16379)
);

NAND2xp5_ASAP7_75t_L g16380 ( 
.A(n_15896),
.B(n_9342),
.Y(n_16380)
);

HB1xp67_ASAP7_75t_L g16381 ( 
.A(n_15849),
.Y(n_16381)
);

INVx1_ASAP7_75t_L g16382 ( 
.A(n_15727),
.Y(n_16382)
);

AND2x2_ASAP7_75t_L g16383 ( 
.A(n_15736),
.B(n_7882),
.Y(n_16383)
);

NAND2xp5_ASAP7_75t_L g16384 ( 
.A(n_15901),
.B(n_15799),
.Y(n_16384)
);

AOI221xp5_ASAP7_75t_L g16385 ( 
.A1(n_15776),
.A2(n_9820),
.B1(n_9818),
.B2(n_9146),
.C(n_9163),
.Y(n_16385)
);

NAND4xp25_ASAP7_75t_L g16386 ( 
.A(n_15772),
.B(n_6662),
.C(n_6718),
.D(n_6717),
.Y(n_16386)
);

INVx2_ASAP7_75t_L g16387 ( 
.A(n_15903),
.Y(n_16387)
);

BUFx2_ASAP7_75t_L g16388 ( 
.A(n_15842),
.Y(n_16388)
);

INVx1_ASAP7_75t_L g16389 ( 
.A(n_15782),
.Y(n_16389)
);

INVx1_ASAP7_75t_L g16390 ( 
.A(n_15783),
.Y(n_16390)
);

INVx2_ASAP7_75t_L g16391 ( 
.A(n_15913),
.Y(n_16391)
);

OAI21xp33_ASAP7_75t_L g16392 ( 
.A1(n_15810),
.A2(n_11358),
.B(n_11299),
.Y(n_16392)
);

NAND2xp5_ASAP7_75t_L g16393 ( 
.A(n_15786),
.B(n_9348),
.Y(n_16393)
);

INVx3_ASAP7_75t_L g16394 ( 
.A(n_15780),
.Y(n_16394)
);

INVx2_ASAP7_75t_L g16395 ( 
.A(n_15902),
.Y(n_16395)
);

AND2x2_ASAP7_75t_L g16396 ( 
.A(n_15817),
.B(n_7882),
.Y(n_16396)
);

OR2x2_ASAP7_75t_L g16397 ( 
.A(n_15871),
.B(n_15823),
.Y(n_16397)
);

NAND2xp33_ASAP7_75t_SL g16398 ( 
.A(n_15797),
.B(n_6922),
.Y(n_16398)
);

INVxp67_ASAP7_75t_SL g16399 ( 
.A(n_15847),
.Y(n_16399)
);

INVx1_ASAP7_75t_SL g16400 ( 
.A(n_15839),
.Y(n_16400)
);

INVx1_ASAP7_75t_L g16401 ( 
.A(n_15880),
.Y(n_16401)
);

AND2x2_ASAP7_75t_L g16402 ( 
.A(n_15818),
.B(n_7953),
.Y(n_16402)
);

INVx2_ASAP7_75t_L g16403 ( 
.A(n_15855),
.Y(n_16403)
);

INVxp67_ASAP7_75t_L g16404 ( 
.A(n_15910),
.Y(n_16404)
);

INVx2_ASAP7_75t_L g16405 ( 
.A(n_15864),
.Y(n_16405)
);

AND2x4_ASAP7_75t_L g16406 ( 
.A(n_15822),
.B(n_8827),
.Y(n_16406)
);

AND2x4_ASAP7_75t_L g16407 ( 
.A(n_15830),
.B(n_8827),
.Y(n_16407)
);

AND2x4_ASAP7_75t_L g16408 ( 
.A(n_15844),
.B(n_8876),
.Y(n_16408)
);

NAND2xp5_ASAP7_75t_L g16409 ( 
.A(n_15914),
.B(n_9348),
.Y(n_16409)
);

INVx2_ASAP7_75t_L g16410 ( 
.A(n_15865),
.Y(n_16410)
);

AND2x2_ASAP7_75t_L g16411 ( 
.A(n_15845),
.B(n_7953),
.Y(n_16411)
);

BUFx2_ASAP7_75t_L g16412 ( 
.A(n_15869),
.Y(n_16412)
);

INVx1_ASAP7_75t_L g16413 ( 
.A(n_15872),
.Y(n_16413)
);

INVx2_ASAP7_75t_L g16414 ( 
.A(n_15875),
.Y(n_16414)
);

AND2x2_ASAP7_75t_L g16415 ( 
.A(n_15883),
.B(n_7953),
.Y(n_16415)
);

INVx2_ASAP7_75t_L g16416 ( 
.A(n_16128),
.Y(n_16416)
);

AND2x2_ASAP7_75t_L g16417 ( 
.A(n_15925),
.B(n_15893),
.Y(n_16417)
);

NOR2xp67_ASAP7_75t_SL g16418 ( 
.A(n_15983),
.B(n_15894),
.Y(n_16418)
);

AND2x4_ASAP7_75t_L g16419 ( 
.A(n_15923),
.B(n_16128),
.Y(n_16419)
);

OA222x2_ASAP7_75t_L g16420 ( 
.A1(n_16120),
.A2(n_9818),
.B1(n_8977),
.B2(n_8957),
.C1(n_8980),
.C2(n_8964),
.Y(n_16420)
);

OR2x6_ASAP7_75t_L g16421 ( 
.A(n_15927),
.B(n_15607),
.Y(n_16421)
);

A2O1A1Ixp33_ASAP7_75t_L g16422 ( 
.A1(n_16060),
.A2(n_16188),
.B(n_15960),
.C(n_16043),
.Y(n_16422)
);

OR2x2_ASAP7_75t_L g16423 ( 
.A(n_15920),
.B(n_15906),
.Y(n_16423)
);

INVxp67_ASAP7_75t_SL g16424 ( 
.A(n_15989),
.Y(n_16424)
);

INVx1_ASAP7_75t_SL g16425 ( 
.A(n_15962),
.Y(n_16425)
);

INVx2_ASAP7_75t_SL g16426 ( 
.A(n_16128),
.Y(n_16426)
);

INVx2_ASAP7_75t_L g16427 ( 
.A(n_16129),
.Y(n_16427)
);

INVx1_ASAP7_75t_L g16428 ( 
.A(n_15930),
.Y(n_16428)
);

INVx1_ASAP7_75t_L g16429 ( 
.A(n_16214),
.Y(n_16429)
);

INVx1_ASAP7_75t_SL g16430 ( 
.A(n_16262),
.Y(n_16430)
);

O2A1O1Ixp5_ASAP7_75t_R g16431 ( 
.A1(n_16006),
.A2(n_15841),
.B(n_15889),
.C(n_15886),
.Y(n_16431)
);

AND2x2_ASAP7_75t_L g16432 ( 
.A(n_15924),
.B(n_10672),
.Y(n_16432)
);

OAI22xp33_ASAP7_75t_L g16433 ( 
.A1(n_16002),
.A2(n_8642),
.B1(n_8644),
.B2(n_8633),
.Y(n_16433)
);

AOI22xp33_ASAP7_75t_L g16434 ( 
.A1(n_16104),
.A2(n_11054),
.B1(n_8857),
.B2(n_9701),
.Y(n_16434)
);

INVx1_ASAP7_75t_L g16435 ( 
.A(n_16075),
.Y(n_16435)
);

O2A1O1Ixp5_ASAP7_75t_R g16436 ( 
.A1(n_15929),
.A2(n_15918),
.B(n_15961),
.C(n_16004),
.Y(n_16436)
);

NAND2xp5_ASAP7_75t_L g16437 ( 
.A(n_15940),
.B(n_9350),
.Y(n_16437)
);

NAND3xp33_ASAP7_75t_L g16438 ( 
.A(n_15958),
.B(n_8644),
.C(n_8642),
.Y(n_16438)
);

INVx2_ASAP7_75t_L g16439 ( 
.A(n_16133),
.Y(n_16439)
);

NAND2x1p5_ASAP7_75t_L g16440 ( 
.A(n_16150),
.B(n_8642),
.Y(n_16440)
);

AND2x2_ASAP7_75t_L g16441 ( 
.A(n_16003),
.B(n_10672),
.Y(n_16441)
);

AOI22xp5_ASAP7_75t_L g16442 ( 
.A1(n_15969),
.A2(n_8903),
.B1(n_8912),
.B2(n_8876),
.Y(n_16442)
);

INVx1_ASAP7_75t_L g16443 ( 
.A(n_16048),
.Y(n_16443)
);

INVx2_ASAP7_75t_L g16444 ( 
.A(n_15987),
.Y(n_16444)
);

NAND2xp5_ASAP7_75t_L g16445 ( 
.A(n_16025),
.B(n_9350),
.Y(n_16445)
);

OR2x2_ASAP7_75t_L g16446 ( 
.A(n_16012),
.B(n_9333),
.Y(n_16446)
);

AO22x1_ASAP7_75t_L g16447 ( 
.A1(n_15933),
.A2(n_6922),
.B1(n_9144),
.B2(n_9142),
.Y(n_16447)
);

O2A1O1Ixp33_ASAP7_75t_L g16448 ( 
.A1(n_15954),
.A2(n_9144),
.B(n_9146),
.C(n_9142),
.Y(n_16448)
);

AOI22xp5_ASAP7_75t_L g16449 ( 
.A1(n_16140),
.A2(n_8903),
.B1(n_8912),
.B2(n_8876),
.Y(n_16449)
);

INVx1_ASAP7_75t_L g16450 ( 
.A(n_16056),
.Y(n_16450)
);

INVx2_ASAP7_75t_L g16451 ( 
.A(n_16013),
.Y(n_16451)
);

AOI33xp33_ASAP7_75t_L g16452 ( 
.A1(n_15919),
.A2(n_8903),
.A3(n_8912),
.B1(n_9144),
.B2(n_9146),
.B3(n_9142),
.Y(n_16452)
);

O2A1O1Ixp5_ASAP7_75t_R g16453 ( 
.A1(n_16246),
.A2(n_15946),
.B(n_16384),
.C(n_15967),
.Y(n_16453)
);

AND2x2_ASAP7_75t_L g16454 ( 
.A(n_16169),
.B(n_10707),
.Y(n_16454)
);

INVx2_ASAP7_75t_L g16455 ( 
.A(n_16041),
.Y(n_16455)
);

INVx1_ASAP7_75t_L g16456 ( 
.A(n_16207),
.Y(n_16456)
);

AOI22xp33_ASAP7_75t_L g16457 ( 
.A1(n_15942),
.A2(n_11054),
.B1(n_8857),
.B2(n_9701),
.Y(n_16457)
);

INVx1_ASAP7_75t_L g16458 ( 
.A(n_16028),
.Y(n_16458)
);

NOR3x1_ASAP7_75t_L g16459 ( 
.A(n_15986),
.B(n_11246),
.C(n_11242),
.Y(n_16459)
);

INVx1_ASAP7_75t_SL g16460 ( 
.A(n_15974),
.Y(n_16460)
);

INVx1_ASAP7_75t_L g16461 ( 
.A(n_16054),
.Y(n_16461)
);

OAI32xp33_ASAP7_75t_L g16462 ( 
.A1(n_16010),
.A2(n_9192),
.A3(n_9203),
.B1(n_9176),
.B2(n_9163),
.Y(n_16462)
);

INVx1_ASAP7_75t_L g16463 ( 
.A(n_16122),
.Y(n_16463)
);

AND2x2_ASAP7_75t_L g16464 ( 
.A(n_16058),
.B(n_10707),
.Y(n_16464)
);

INVx2_ASAP7_75t_L g16465 ( 
.A(n_15973),
.Y(n_16465)
);

NOR2xp33_ASAP7_75t_L g16466 ( 
.A(n_16067),
.B(n_7510),
.Y(n_16466)
);

INVx1_ASAP7_75t_L g16467 ( 
.A(n_16018),
.Y(n_16467)
);

AND2x4_ASAP7_75t_L g16468 ( 
.A(n_15939),
.B(n_10755),
.Y(n_16468)
);

NAND2xp5_ASAP7_75t_L g16469 ( 
.A(n_15956),
.B(n_9360),
.Y(n_16469)
);

OR2x2_ASAP7_75t_L g16470 ( 
.A(n_15951),
.B(n_9333),
.Y(n_16470)
);

INVx1_ASAP7_75t_L g16471 ( 
.A(n_16412),
.Y(n_16471)
);

OAI322xp33_ASAP7_75t_L g16472 ( 
.A1(n_15955),
.A2(n_9203),
.A3(n_9176),
.B1(n_9221),
.B2(n_9232),
.C1(n_9192),
.C2(n_9163),
.Y(n_16472)
);

INVxp67_ASAP7_75t_L g16473 ( 
.A(n_16313),
.Y(n_16473)
);

AOI21x1_ASAP7_75t_L g16474 ( 
.A1(n_15921),
.A2(n_10760),
.B(n_10727),
.Y(n_16474)
);

INVx2_ASAP7_75t_L g16475 ( 
.A(n_15945),
.Y(n_16475)
);

INVx1_ASAP7_75t_L g16476 ( 
.A(n_15931),
.Y(n_16476)
);

O2A1O1Ixp33_ASAP7_75t_L g16477 ( 
.A1(n_15964),
.A2(n_16070),
.B(n_15928),
.C(n_15944),
.Y(n_16477)
);

INVx2_ASAP7_75t_L g16478 ( 
.A(n_16072),
.Y(n_16478)
);

AOI211xp5_ASAP7_75t_L g16479 ( 
.A1(n_16189),
.A2(n_7510),
.B(n_10401),
.C(n_10340),
.Y(n_16479)
);

INVx1_ASAP7_75t_L g16480 ( 
.A(n_15949),
.Y(n_16480)
);

INVx1_ASAP7_75t_L g16481 ( 
.A(n_15998),
.Y(n_16481)
);

INVx1_ASAP7_75t_L g16482 ( 
.A(n_15937),
.Y(n_16482)
);

OAI22xp33_ASAP7_75t_L g16483 ( 
.A1(n_16233),
.A2(n_8644),
.B1(n_8748),
.B2(n_8642),
.Y(n_16483)
);

OR2x2_ASAP7_75t_L g16484 ( 
.A(n_15970),
.B(n_9333),
.Y(n_16484)
);

INVx1_ASAP7_75t_L g16485 ( 
.A(n_15926),
.Y(n_16485)
);

INVx3_ASAP7_75t_L g16486 ( 
.A(n_15922),
.Y(n_16486)
);

INVx1_ASAP7_75t_L g16487 ( 
.A(n_15941),
.Y(n_16487)
);

OR2x2_ASAP7_75t_L g16488 ( 
.A(n_15979),
.B(n_9333),
.Y(n_16488)
);

XOR2x2_ASAP7_75t_L g16489 ( 
.A(n_15950),
.B(n_7510),
.Y(n_16489)
);

INVx1_ASAP7_75t_L g16490 ( 
.A(n_15932),
.Y(n_16490)
);

INVx1_ASAP7_75t_L g16491 ( 
.A(n_15935),
.Y(n_16491)
);

INVxp67_ASAP7_75t_SL g16492 ( 
.A(n_16163),
.Y(n_16492)
);

INVx1_ASAP7_75t_L g16493 ( 
.A(n_16020),
.Y(n_16493)
);

INVx1_ASAP7_75t_L g16494 ( 
.A(n_15953),
.Y(n_16494)
);

INVx1_ASAP7_75t_L g16495 ( 
.A(n_16082),
.Y(n_16495)
);

INVx1_ASAP7_75t_L g16496 ( 
.A(n_16131),
.Y(n_16496)
);

OAI211xp5_ASAP7_75t_L g16497 ( 
.A1(n_15948),
.A2(n_11054),
.B(n_11373),
.C(n_11299),
.Y(n_16497)
);

AND2x4_ASAP7_75t_L g16498 ( 
.A(n_16021),
.B(n_10755),
.Y(n_16498)
);

INVx1_ASAP7_75t_L g16499 ( 
.A(n_16106),
.Y(n_16499)
);

HB1xp67_ASAP7_75t_L g16500 ( 
.A(n_15992),
.Y(n_16500)
);

INVx1_ASAP7_75t_SL g16501 ( 
.A(n_16216),
.Y(n_16501)
);

INVx1_ASAP7_75t_L g16502 ( 
.A(n_15943),
.Y(n_16502)
);

AOI22xp5_ASAP7_75t_L g16503 ( 
.A1(n_16055),
.A2(n_8644),
.B1(n_8748),
.B2(n_8642),
.Y(n_16503)
);

INVx2_ASAP7_75t_L g16504 ( 
.A(n_16216),
.Y(n_16504)
);

OAI22xp33_ASAP7_75t_L g16505 ( 
.A1(n_16267),
.A2(n_8748),
.B1(n_8947),
.B2(n_8644),
.Y(n_16505)
);

BUFx3_ASAP7_75t_L g16506 ( 
.A(n_16039),
.Y(n_16506)
);

NAND2xp67_ASAP7_75t_SL g16507 ( 
.A(n_15995),
.B(n_7782),
.Y(n_16507)
);

INVx1_ASAP7_75t_L g16508 ( 
.A(n_16083),
.Y(n_16508)
);

OAI31xp33_ASAP7_75t_L g16509 ( 
.A1(n_16398),
.A2(n_9192),
.A3(n_9203),
.B(n_9176),
.Y(n_16509)
);

OAI22xp5_ASAP7_75t_L g16510 ( 
.A1(n_16103),
.A2(n_8947),
.B1(n_8748),
.B2(n_7953),
.Y(n_16510)
);

NAND2xp5_ASAP7_75t_L g16511 ( 
.A(n_16085),
.B(n_9360),
.Y(n_16511)
);

NOR2xp33_ASAP7_75t_L g16512 ( 
.A(n_16265),
.B(n_7510),
.Y(n_16512)
);

INVxp33_ASAP7_75t_L g16513 ( 
.A(n_15959),
.Y(n_16513)
);

AND2x2_ASAP7_75t_L g16514 ( 
.A(n_15965),
.B(n_10340),
.Y(n_16514)
);

INVx1_ASAP7_75t_L g16515 ( 
.A(n_16087),
.Y(n_16515)
);

AOI22xp5_ASAP7_75t_L g16516 ( 
.A1(n_16143),
.A2(n_8947),
.B1(n_8748),
.B2(n_7953),
.Y(n_16516)
);

OR2x2_ASAP7_75t_L g16517 ( 
.A(n_16400),
.B(n_9349),
.Y(n_16517)
);

NAND2x2_ASAP7_75t_L g16518 ( 
.A(n_16016),
.B(n_16288),
.Y(n_16518)
);

INVx1_ASAP7_75t_L g16519 ( 
.A(n_16036),
.Y(n_16519)
);

NAND4xp75_ASAP7_75t_L g16520 ( 
.A(n_15963),
.B(n_9872),
.C(n_9870),
.D(n_9653),
.Y(n_16520)
);

INVx1_ASAP7_75t_L g16521 ( 
.A(n_16031),
.Y(n_16521)
);

INVx1_ASAP7_75t_SL g16522 ( 
.A(n_16005),
.Y(n_16522)
);

INVx1_ASAP7_75t_L g16523 ( 
.A(n_16033),
.Y(n_16523)
);

AND2x4_ASAP7_75t_L g16524 ( 
.A(n_16260),
.B(n_10401),
.Y(n_16524)
);

INVx1_ASAP7_75t_L g16525 ( 
.A(n_16381),
.Y(n_16525)
);

INVxp67_ASAP7_75t_L g16526 ( 
.A(n_16388),
.Y(n_16526)
);

AND2x2_ASAP7_75t_L g16527 ( 
.A(n_15957),
.B(n_7972),
.Y(n_16527)
);

INVx1_ASAP7_75t_L g16528 ( 
.A(n_16022),
.Y(n_16528)
);

AND2x4_ASAP7_75t_L g16529 ( 
.A(n_16283),
.B(n_11242),
.Y(n_16529)
);

NAND4xp75_ASAP7_75t_SL g16530 ( 
.A(n_15966),
.B(n_8432),
.C(n_8421),
.D(n_9870),
.Y(n_16530)
);

AO22x1_ASAP7_75t_L g16531 ( 
.A1(n_15980),
.A2(n_9232),
.B1(n_9234),
.B2(n_9221),
.Y(n_16531)
);

OAI22xp33_ASAP7_75t_L g16532 ( 
.A1(n_16095),
.A2(n_8947),
.B1(n_8748),
.B2(n_9221),
.Y(n_16532)
);

XNOR2xp5_ASAP7_75t_L g16533 ( 
.A(n_16134),
.B(n_8236),
.Y(n_16533)
);

HB1xp67_ASAP7_75t_L g16534 ( 
.A(n_16063),
.Y(n_16534)
);

OR2x2_ASAP7_75t_L g16535 ( 
.A(n_16394),
.B(n_9349),
.Y(n_16535)
);

NAND5xp2_ASAP7_75t_L g16536 ( 
.A(n_15952),
.B(n_8432),
.C(n_7942),
.D(n_7949),
.E(n_7881),
.Y(n_16536)
);

NAND2xp67_ASAP7_75t_SL g16537 ( 
.A(n_16231),
.B(n_7782),
.Y(n_16537)
);

O2A1O1Ixp33_ASAP7_75t_L g16538 ( 
.A1(n_16138),
.A2(n_9234),
.B(n_9237),
.C(n_9232),
.Y(n_16538)
);

INVx2_ASAP7_75t_L g16539 ( 
.A(n_16011),
.Y(n_16539)
);

NOR2xp67_ASAP7_75t_SL g16540 ( 
.A(n_16059),
.B(n_16069),
.Y(n_16540)
);

O2A1O1Ixp5_ASAP7_75t_R g16541 ( 
.A1(n_16191),
.A2(n_8035),
.B(n_8046),
.C(n_8033),
.Y(n_16541)
);

INVx1_ASAP7_75t_L g16542 ( 
.A(n_16038),
.Y(n_16542)
);

OAI211xp5_ASAP7_75t_L g16543 ( 
.A1(n_15991),
.A2(n_9673),
.B(n_9694),
.C(n_9653),
.Y(n_16543)
);

INVx1_ASAP7_75t_L g16544 ( 
.A(n_16105),
.Y(n_16544)
);

AND2x2_ASAP7_75t_L g16545 ( 
.A(n_16030),
.B(n_16034),
.Y(n_16545)
);

OR2x2_ASAP7_75t_L g16546 ( 
.A(n_16151),
.B(n_16045),
.Y(n_16546)
);

INVx1_ASAP7_75t_L g16547 ( 
.A(n_16121),
.Y(n_16547)
);

NAND2xp5_ASAP7_75t_L g16548 ( 
.A(n_16007),
.B(n_9361),
.Y(n_16548)
);

AOI21xp5_ASAP7_75t_L g16549 ( 
.A1(n_16008),
.A2(n_11260),
.B(n_11246),
.Y(n_16549)
);

NAND2xp5_ASAP7_75t_L g16550 ( 
.A(n_16037),
.B(n_15947),
.Y(n_16550)
);

OAI22xp33_ASAP7_75t_L g16551 ( 
.A1(n_16155),
.A2(n_8947),
.B1(n_8748),
.B2(n_9234),
.Y(n_16551)
);

INVx1_ASAP7_75t_L g16552 ( 
.A(n_16236),
.Y(n_16552)
);

HB1xp67_ASAP7_75t_L g16553 ( 
.A(n_15996),
.Y(n_16553)
);

AND4x1_ASAP7_75t_L g16554 ( 
.A(n_16071),
.B(n_7380),
.C(n_7358),
.D(n_8046),
.Y(n_16554)
);

XNOR2xp5_ASAP7_75t_L g16555 ( 
.A(n_16134),
.B(n_6662),
.Y(n_16555)
);

AOI211xp5_ASAP7_75t_L g16556 ( 
.A1(n_15999),
.A2(n_7510),
.B(n_11260),
.C(n_9236),
.Y(n_16556)
);

AND2x2_ASAP7_75t_L g16557 ( 
.A(n_15971),
.B(n_7972),
.Y(n_16557)
);

INVxp67_ASAP7_75t_SL g16558 ( 
.A(n_16026),
.Y(n_16558)
);

INVx1_ASAP7_75t_L g16559 ( 
.A(n_15938),
.Y(n_16559)
);

OAI22x1_ASAP7_75t_L g16560 ( 
.A1(n_16197),
.A2(n_9168),
.B1(n_9072),
.B2(n_8139),
.Y(n_16560)
);

INVx1_ASAP7_75t_L g16561 ( 
.A(n_16046),
.Y(n_16561)
);

NAND4xp75_ASAP7_75t_SL g16562 ( 
.A(n_15978),
.B(n_8421),
.C(n_9872),
.D(n_9870),
.Y(n_16562)
);

INVx1_ASAP7_75t_L g16563 ( 
.A(n_16213),
.Y(n_16563)
);

INVx1_ASAP7_75t_L g16564 ( 
.A(n_16285),
.Y(n_16564)
);

AND2x2_ASAP7_75t_L g16565 ( 
.A(n_16107),
.B(n_7972),
.Y(n_16565)
);

AND2x4_ASAP7_75t_L g16566 ( 
.A(n_16310),
.B(n_11411),
.Y(n_16566)
);

INVx2_ASAP7_75t_SL g16567 ( 
.A(n_16097),
.Y(n_16567)
);

OR2x2_ASAP7_75t_L g16568 ( 
.A(n_16243),
.B(n_9349),
.Y(n_16568)
);

NAND2xp5_ASAP7_75t_L g16569 ( 
.A(n_15934),
.B(n_9361),
.Y(n_16569)
);

INVx4_ASAP7_75t_L g16570 ( 
.A(n_16015),
.Y(n_16570)
);

NAND2xp5_ASAP7_75t_L g16571 ( 
.A(n_15936),
.B(n_9366),
.Y(n_16571)
);

NAND2xp5_ASAP7_75t_SL g16572 ( 
.A(n_16273),
.B(n_8748),
.Y(n_16572)
);

NAND2xp5_ASAP7_75t_L g16573 ( 
.A(n_16079),
.B(n_9366),
.Y(n_16573)
);

OA222x2_ASAP7_75t_L g16574 ( 
.A1(n_16027),
.A2(n_15984),
.B1(n_15994),
.B2(n_16009),
.C1(n_15981),
.C2(n_16139),
.Y(n_16574)
);

OR2x2_ASAP7_75t_L g16575 ( 
.A(n_16264),
.B(n_9349),
.Y(n_16575)
);

AOI22xp5_ASAP7_75t_L g16576 ( 
.A1(n_16218),
.A2(n_8947),
.B1(n_7972),
.B2(n_8158),
.Y(n_16576)
);

INVx1_ASAP7_75t_L g16577 ( 
.A(n_15968),
.Y(n_16577)
);

INVx2_ASAP7_75t_L g16578 ( 
.A(n_16000),
.Y(n_16578)
);

INVx2_ASAP7_75t_L g16579 ( 
.A(n_16001),
.Y(n_16579)
);

A2O1A1Ixp33_ASAP7_75t_L g16580 ( 
.A1(n_16290),
.A2(n_16171),
.B(n_16081),
.C(n_15976),
.Y(n_16580)
);

OR2x2_ASAP7_75t_L g16581 ( 
.A(n_16210),
.B(n_16219),
.Y(n_16581)
);

INVx1_ASAP7_75t_L g16582 ( 
.A(n_16174),
.Y(n_16582)
);

OAI322xp33_ASAP7_75t_L g16583 ( 
.A1(n_15972),
.A2(n_9246),
.A3(n_9240),
.B1(n_9256),
.B2(n_9258),
.C1(n_9244),
.C2(n_9237),
.Y(n_16583)
);

O2A1O1Ixp33_ASAP7_75t_L g16584 ( 
.A1(n_16344),
.A2(n_9240),
.B(n_9244),
.C(n_9237),
.Y(n_16584)
);

NOR2xp33_ASAP7_75t_L g16585 ( 
.A(n_16158),
.B(n_8947),
.Y(n_16585)
);

AND2x4_ASAP7_75t_L g16586 ( 
.A(n_16225),
.B(n_11411),
.Y(n_16586)
);

INVx1_ASAP7_75t_L g16587 ( 
.A(n_15990),
.Y(n_16587)
);

AOI211xp5_ASAP7_75t_L g16588 ( 
.A1(n_16304),
.A2(n_9236),
.B(n_8947),
.C(n_8690),
.Y(n_16588)
);

OAI33xp33_ASAP7_75t_L g16589 ( 
.A1(n_15975),
.A2(n_9256),
.A3(n_9244),
.B1(n_9258),
.B2(n_9246),
.B3(n_9240),
.Y(n_16589)
);

AOI22xp5_ASAP7_75t_L g16590 ( 
.A1(n_16386),
.A2(n_7972),
.B1(n_8158),
.B2(n_8139),
.Y(n_16590)
);

OR2x2_ASAP7_75t_L g16591 ( 
.A(n_16226),
.B(n_7736),
.Y(n_16591)
);

AOI22xp5_ASAP7_75t_L g16592 ( 
.A1(n_16208),
.A2(n_8158),
.B1(n_8254),
.B2(n_8139),
.Y(n_16592)
);

AO221x1_ASAP7_75t_L g16593 ( 
.A1(n_16177),
.A2(n_8254),
.B1(n_8269),
.B2(n_8158),
.C(n_8139),
.Y(n_16593)
);

INVx1_ASAP7_75t_L g16594 ( 
.A(n_16334),
.Y(n_16594)
);

INVx1_ASAP7_75t_L g16595 ( 
.A(n_16190),
.Y(n_16595)
);

INVx1_ASAP7_75t_L g16596 ( 
.A(n_16196),
.Y(n_16596)
);

NAND3xp33_ASAP7_75t_L g16597 ( 
.A(n_15977),
.B(n_9168),
.C(n_9072),
.Y(n_16597)
);

INVx1_ASAP7_75t_L g16598 ( 
.A(n_16227),
.Y(n_16598)
);

INVx1_ASAP7_75t_L g16599 ( 
.A(n_16239),
.Y(n_16599)
);

INVx1_ASAP7_75t_L g16600 ( 
.A(n_16254),
.Y(n_16600)
);

AOI221xp5_ASAP7_75t_L g16601 ( 
.A1(n_16179),
.A2(n_9258),
.B1(n_9259),
.B2(n_9256),
.C(n_9246),
.Y(n_16601)
);

AOI32xp33_ASAP7_75t_L g16602 ( 
.A1(n_16127),
.A2(n_10564),
.A3(n_10545),
.B1(n_10460),
.B2(n_10727),
.Y(n_16602)
);

BUFx2_ASAP7_75t_L g16603 ( 
.A(n_16220),
.Y(n_16603)
);

NOR2xp33_ASAP7_75t_L g16604 ( 
.A(n_16200),
.B(n_8139),
.Y(n_16604)
);

OR2x2_ASAP7_75t_L g16605 ( 
.A(n_16230),
.B(n_7736),
.Y(n_16605)
);

INVx2_ASAP7_75t_L g16606 ( 
.A(n_16317),
.Y(n_16606)
);

INVx1_ASAP7_75t_L g16607 ( 
.A(n_16276),
.Y(n_16607)
);

INVxp67_ASAP7_75t_SL g16608 ( 
.A(n_16181),
.Y(n_16608)
);

INVx1_ASAP7_75t_SL g16609 ( 
.A(n_16364),
.Y(n_16609)
);

AOI22xp5_ASAP7_75t_L g16610 ( 
.A1(n_16110),
.A2(n_8254),
.B1(n_8269),
.B2(n_8158),
.Y(n_16610)
);

INVx1_ASAP7_75t_L g16611 ( 
.A(n_16280),
.Y(n_16611)
);

CKINVDCx16_ASAP7_75t_R g16612 ( 
.A(n_16192),
.Y(n_16612)
);

INVx2_ASAP7_75t_L g16613 ( 
.A(n_16362),
.Y(n_16613)
);

HB1xp67_ASAP7_75t_L g16614 ( 
.A(n_16201),
.Y(n_16614)
);

INVx1_ASAP7_75t_L g16615 ( 
.A(n_16148),
.Y(n_16615)
);

INVx1_ASAP7_75t_SL g16616 ( 
.A(n_16235),
.Y(n_16616)
);

INVx1_ASAP7_75t_L g16617 ( 
.A(n_16413),
.Y(n_16617)
);

INVx2_ASAP7_75t_L g16618 ( 
.A(n_16365),
.Y(n_16618)
);

INVx1_ASAP7_75t_L g16619 ( 
.A(n_16146),
.Y(n_16619)
);

AOI21xp5_ASAP7_75t_L g16620 ( 
.A1(n_16024),
.A2(n_10760),
.B(n_11087),
.Y(n_16620)
);

OR2x2_ASAP7_75t_L g16621 ( 
.A(n_16374),
.B(n_7736),
.Y(n_16621)
);

O2A1O1Ixp33_ASAP7_75t_L g16622 ( 
.A1(n_16294),
.A2(n_16212),
.B(n_16119),
.C(n_16130),
.Y(n_16622)
);

INVx1_ASAP7_75t_L g16623 ( 
.A(n_16387),
.Y(n_16623)
);

HB1xp67_ASAP7_75t_L g16624 ( 
.A(n_16201),
.Y(n_16624)
);

OR2x2_ASAP7_75t_L g16625 ( 
.A(n_16391),
.B(n_7849),
.Y(n_16625)
);

INVx1_ASAP7_75t_L g16626 ( 
.A(n_16395),
.Y(n_16626)
);

NAND2xp5_ASAP7_75t_SL g16627 ( 
.A(n_16252),
.B(n_8254),
.Y(n_16627)
);

AND2x2_ASAP7_75t_L g16628 ( 
.A(n_16403),
.B(n_8254),
.Y(n_16628)
);

OAI322xp33_ASAP7_75t_L g16629 ( 
.A1(n_16089),
.A2(n_16135),
.A3(n_16137),
.B1(n_16114),
.B2(n_16324),
.C1(n_16049),
.C2(n_16295),
.Y(n_16629)
);

INVxp67_ASAP7_75t_SL g16630 ( 
.A(n_16144),
.Y(n_16630)
);

OR2x2_ASAP7_75t_L g16631 ( 
.A(n_16405),
.B(n_7849),
.Y(n_16631)
);

AOI22xp5_ASAP7_75t_L g16632 ( 
.A1(n_15985),
.A2(n_8269),
.B1(n_8518),
.B2(n_8433),
.Y(n_16632)
);

INVx2_ASAP7_75t_SL g16633 ( 
.A(n_16222),
.Y(n_16633)
);

OAI31xp33_ASAP7_75t_L g16634 ( 
.A1(n_16349),
.A2(n_9266),
.A3(n_9276),
.B(n_9259),
.Y(n_16634)
);

BUFx2_ASAP7_75t_L g16635 ( 
.A(n_16271),
.Y(n_16635)
);

INVx1_ASAP7_75t_L g16636 ( 
.A(n_16410),
.Y(n_16636)
);

INVx1_ASAP7_75t_L g16637 ( 
.A(n_16414),
.Y(n_16637)
);

INVx1_ASAP7_75t_L g16638 ( 
.A(n_16044),
.Y(n_16638)
);

INVx1_ASAP7_75t_L g16639 ( 
.A(n_16042),
.Y(n_16639)
);

OR2x2_ASAP7_75t_L g16640 ( 
.A(n_16159),
.B(n_7849),
.Y(n_16640)
);

AOI22xp5_ASAP7_75t_L g16641 ( 
.A1(n_16136),
.A2(n_8269),
.B1(n_8518),
.B2(n_8433),
.Y(n_16641)
);

OAI22xp5_ASAP7_75t_L g16642 ( 
.A1(n_16279),
.A2(n_8269),
.B1(n_8518),
.B2(n_8433),
.Y(n_16642)
);

NAND2xp5_ASAP7_75t_L g16643 ( 
.A(n_16297),
.B(n_9368),
.Y(n_16643)
);

INVx1_ASAP7_75t_L g16644 ( 
.A(n_16221),
.Y(n_16644)
);

INVx2_ASAP7_75t_SL g16645 ( 
.A(n_16249),
.Y(n_16645)
);

NAND2xp5_ASAP7_75t_L g16646 ( 
.A(n_16154),
.B(n_9368),
.Y(n_16646)
);

AOI32xp33_ASAP7_75t_L g16647 ( 
.A1(n_16203),
.A2(n_10564),
.A3(n_10545),
.B1(n_10460),
.B2(n_9276),
.Y(n_16647)
);

OAI31xp67_ASAP7_75t_L g16648 ( 
.A1(n_16168),
.A2(n_9266),
.A3(n_9276),
.B(n_9259),
.Y(n_16648)
);

OAI22xp33_ASAP7_75t_L g16649 ( 
.A1(n_16237),
.A2(n_16253),
.B1(n_15982),
.B2(n_16286),
.Y(n_16649)
);

AND2x2_ASAP7_75t_L g16650 ( 
.A(n_16175),
.B(n_8433),
.Y(n_16650)
);

INVx1_ASAP7_75t_L g16651 ( 
.A(n_16014),
.Y(n_16651)
);

O2A1O1Ixp33_ASAP7_75t_L g16652 ( 
.A1(n_15988),
.A2(n_16287),
.B(n_16299),
.C(n_16296),
.Y(n_16652)
);

O2A1O1Ixp5_ASAP7_75t_L g16653 ( 
.A1(n_16032),
.A2(n_9284),
.B(n_9285),
.C(n_9266),
.Y(n_16653)
);

OR2x2_ASAP7_75t_L g16654 ( 
.A(n_16343),
.B(n_7868),
.Y(n_16654)
);

NOR2xp33_ASAP7_75t_L g16655 ( 
.A(n_16314),
.B(n_8433),
.Y(n_16655)
);

BUFx2_ASAP7_75t_L g16656 ( 
.A(n_16301),
.Y(n_16656)
);

INVx2_ASAP7_75t_L g16657 ( 
.A(n_16202),
.Y(n_16657)
);

INVx1_ASAP7_75t_L g16658 ( 
.A(n_16017),
.Y(n_16658)
);

INVx1_ASAP7_75t_L g16659 ( 
.A(n_16019),
.Y(n_16659)
);

AND2x2_ASAP7_75t_L g16660 ( 
.A(n_16376),
.B(n_8518),
.Y(n_16660)
);

NAND2xp5_ASAP7_75t_L g16661 ( 
.A(n_16161),
.B(n_16086),
.Y(n_16661)
);

OA222x2_ASAP7_75t_L g16662 ( 
.A1(n_16141),
.A2(n_8977),
.B1(n_8957),
.B2(n_8980),
.C1(n_8964),
.C2(n_8953),
.Y(n_16662)
);

INVxp67_ASAP7_75t_SL g16663 ( 
.A(n_16123),
.Y(n_16663)
);

INVx1_ASAP7_75t_L g16664 ( 
.A(n_16132),
.Y(n_16664)
);

INVx2_ASAP7_75t_L g16665 ( 
.A(n_16202),
.Y(n_16665)
);

AOI22xp33_ASAP7_75t_L g16666 ( 
.A1(n_16102),
.A2(n_8857),
.B1(n_9701),
.B2(n_8225),
.Y(n_16666)
);

INVx1_ASAP7_75t_L g16667 ( 
.A(n_16076),
.Y(n_16667)
);

INVx1_ASAP7_75t_L g16668 ( 
.A(n_16178),
.Y(n_16668)
);

INVx2_ASAP7_75t_L g16669 ( 
.A(n_16065),
.Y(n_16669)
);

OR2x2_ASAP7_75t_L g16670 ( 
.A(n_15997),
.B(n_7868),
.Y(n_16670)
);

BUFx3_ASAP7_75t_L g16671 ( 
.A(n_16328),
.Y(n_16671)
);

INVx1_ASAP7_75t_L g16672 ( 
.A(n_16185),
.Y(n_16672)
);

AOI21xp33_ASAP7_75t_L g16673 ( 
.A1(n_16118),
.A2(n_11142),
.B(n_11087),
.Y(n_16673)
);

NAND3xp33_ASAP7_75t_L g16674 ( 
.A(n_16259),
.B(n_9168),
.C(n_9701),
.Y(n_16674)
);

OR2x2_ASAP7_75t_L g16675 ( 
.A(n_15993),
.B(n_7868),
.Y(n_16675)
);

NAND4xp25_ASAP7_75t_L g16676 ( 
.A(n_16195),
.B(n_6718),
.C(n_6740),
.D(n_6717),
.Y(n_16676)
);

INVx2_ASAP7_75t_L g16677 ( 
.A(n_16066),
.Y(n_16677)
);

INVx1_ASAP7_75t_L g16678 ( 
.A(n_16090),
.Y(n_16678)
);

INVx1_ASAP7_75t_L g16679 ( 
.A(n_16091),
.Y(n_16679)
);

INVx1_ASAP7_75t_L g16680 ( 
.A(n_16092),
.Y(n_16680)
);

AND2x2_ASAP7_75t_L g16681 ( 
.A(n_16166),
.B(n_8518),
.Y(n_16681)
);

XNOR2xp5_ASAP7_75t_L g16682 ( 
.A(n_16073),
.B(n_6717),
.Y(n_16682)
);

AND2x2_ASAP7_75t_L g16683 ( 
.A(n_16165),
.B(n_8528),
.Y(n_16683)
);

AND2x4_ASAP7_75t_L g16684 ( 
.A(n_16160),
.B(n_10775),
.Y(n_16684)
);

NOR3x1_ASAP7_75t_L g16685 ( 
.A(n_16350),
.B(n_9732),
.C(n_9724),
.Y(n_16685)
);

INVx2_ASAP7_75t_L g16686 ( 
.A(n_16062),
.Y(n_16686)
);

INVx2_ASAP7_75t_SL g16687 ( 
.A(n_16369),
.Y(n_16687)
);

INVx2_ASAP7_75t_SL g16688 ( 
.A(n_16167),
.Y(n_16688)
);

OR2x6_ASAP7_75t_L g16689 ( 
.A(n_16353),
.B(n_16359),
.Y(n_16689)
);

INVx1_ASAP7_75t_L g16690 ( 
.A(n_16035),
.Y(n_16690)
);

INVx1_ASAP7_75t_L g16691 ( 
.A(n_16050),
.Y(n_16691)
);

INVx1_ASAP7_75t_L g16692 ( 
.A(n_16051),
.Y(n_16692)
);

XNOR2xp5_ASAP7_75t_L g16693 ( 
.A(n_16074),
.B(n_6718),
.Y(n_16693)
);

NAND2xp5_ASAP7_75t_L g16694 ( 
.A(n_16077),
.B(n_9369),
.Y(n_16694)
);

OR2x2_ASAP7_75t_L g16695 ( 
.A(n_16397),
.B(n_8382),
.Y(n_16695)
);

NAND2xp33_ASAP7_75t_L g16696 ( 
.A(n_16183),
.B(n_8785),
.Y(n_16696)
);

NAND2xp5_ASAP7_75t_L g16697 ( 
.A(n_16098),
.B(n_9369),
.Y(n_16697)
);

AND2x2_ASAP7_75t_L g16698 ( 
.A(n_16113),
.B(n_8528),
.Y(n_16698)
);

A2O1A1Ixp33_ASAP7_75t_L g16699 ( 
.A1(n_16057),
.A2(n_10787),
.B(n_10812),
.C(n_10775),
.Y(n_16699)
);

INVx1_ASAP7_75t_L g16700 ( 
.A(n_16029),
.Y(n_16700)
);

NAND2xp5_ASAP7_75t_L g16701 ( 
.A(n_16101),
.B(n_9381),
.Y(n_16701)
);

INVx1_ASAP7_75t_L g16702 ( 
.A(n_16040),
.Y(n_16702)
);

AOI22xp5_ASAP7_75t_L g16703 ( 
.A1(n_16068),
.A2(n_8544),
.B1(n_8589),
.B2(n_8528),
.Y(n_16703)
);

INVx1_ASAP7_75t_L g16704 ( 
.A(n_16061),
.Y(n_16704)
);

OR2x2_ASAP7_75t_L g16705 ( 
.A(n_16053),
.B(n_8382),
.Y(n_16705)
);

A2O1A1Ixp33_ASAP7_75t_L g16706 ( 
.A1(n_16172),
.A2(n_10812),
.B(n_10841),
.C(n_10787),
.Y(n_16706)
);

NAND2xp5_ASAP7_75t_L g16707 ( 
.A(n_16111),
.B(n_9381),
.Y(n_16707)
);

NAND2xp5_ASAP7_75t_L g16708 ( 
.A(n_16125),
.B(n_9382),
.Y(n_16708)
);

OA222x2_ASAP7_75t_L g16709 ( 
.A1(n_16147),
.A2(n_8977),
.B1(n_8957),
.B2(n_8980),
.C1(n_8964),
.C2(n_8953),
.Y(n_16709)
);

INVx1_ASAP7_75t_L g16710 ( 
.A(n_16126),
.Y(n_16710)
);

INVx1_ASAP7_75t_L g16711 ( 
.A(n_16116),
.Y(n_16711)
);

OR2x2_ASAP7_75t_L g16712 ( 
.A(n_16354),
.B(n_8393),
.Y(n_16712)
);

INVx1_ASAP7_75t_L g16713 ( 
.A(n_16096),
.Y(n_16713)
);

INVx1_ASAP7_75t_SL g16714 ( 
.A(n_16142),
.Y(n_16714)
);

INVx2_ASAP7_75t_L g16715 ( 
.A(n_16064),
.Y(n_16715)
);

INVx1_ASAP7_75t_L g16716 ( 
.A(n_16258),
.Y(n_16716)
);

INVx2_ASAP7_75t_SL g16717 ( 
.A(n_16232),
.Y(n_16717)
);

AND2x4_ASAP7_75t_L g16718 ( 
.A(n_16399),
.B(n_10841),
.Y(n_16718)
);

INVx2_ASAP7_75t_L g16719 ( 
.A(n_16205),
.Y(n_16719)
);

AND2x2_ASAP7_75t_L g16720 ( 
.A(n_16182),
.B(n_8528),
.Y(n_16720)
);

INVx1_ASAP7_75t_L g16721 ( 
.A(n_16224),
.Y(n_16721)
);

INVx1_ASAP7_75t_L g16722 ( 
.A(n_16173),
.Y(n_16722)
);

INVx1_ASAP7_75t_L g16723 ( 
.A(n_16180),
.Y(n_16723)
);

OAI322xp33_ASAP7_75t_L g16724 ( 
.A1(n_16094),
.A2(n_9334),
.A3(n_9285),
.B1(n_9336),
.B2(n_9340),
.C1(n_9322),
.C2(n_9284),
.Y(n_16724)
);

NOR2xp33_ASAP7_75t_L g16725 ( 
.A(n_16404),
.B(n_8528),
.Y(n_16725)
);

AND2x4_ASAP7_75t_L g16726 ( 
.A(n_16255),
.B(n_10853),
.Y(n_16726)
);

AOI211xp5_ASAP7_75t_L g16727 ( 
.A1(n_16047),
.A2(n_8634),
.B(n_9787),
.C(n_11239),
.Y(n_16727)
);

INVx1_ASAP7_75t_L g16728 ( 
.A(n_16184),
.Y(n_16728)
);

OR2x2_ASAP7_75t_L g16729 ( 
.A(n_16164),
.B(n_8393),
.Y(n_16729)
);

OR2x2_ASAP7_75t_L g16730 ( 
.A(n_16109),
.B(n_8550),
.Y(n_16730)
);

INVx1_ASAP7_75t_L g16731 ( 
.A(n_16186),
.Y(n_16731)
);

HB1xp67_ASAP7_75t_L g16732 ( 
.A(n_16238),
.Y(n_16732)
);

INVx1_ASAP7_75t_L g16733 ( 
.A(n_16145),
.Y(n_16733)
);

AOI22xp5_ASAP7_75t_L g16734 ( 
.A1(n_16084),
.A2(n_8589),
.B1(n_8652),
.B2(n_8544),
.Y(n_16734)
);

BUFx3_ASAP7_75t_L g16735 ( 
.A(n_16322),
.Y(n_16735)
);

INVx1_ASAP7_75t_L g16736 ( 
.A(n_16149),
.Y(n_16736)
);

OAI211xp5_ASAP7_75t_L g16737 ( 
.A1(n_16080),
.A2(n_9653),
.B(n_9694),
.C(n_9673),
.Y(n_16737)
);

AND2x4_ASAP7_75t_L g16738 ( 
.A(n_16153),
.B(n_10853),
.Y(n_16738)
);

A2O1A1Ixp33_ASAP7_75t_L g16739 ( 
.A1(n_16157),
.A2(n_10857),
.B(n_10865),
.C(n_10855),
.Y(n_16739)
);

INVx2_ASAP7_75t_L g16740 ( 
.A(n_16215),
.Y(n_16740)
);

AND2x2_ASAP7_75t_L g16741 ( 
.A(n_16204),
.B(n_8544),
.Y(n_16741)
);

NAND3xp33_ASAP7_75t_L g16742 ( 
.A(n_16088),
.B(n_9872),
.C(n_9870),
.Y(n_16742)
);

INVx1_ASAP7_75t_L g16743 ( 
.A(n_16170),
.Y(n_16743)
);

INVx1_ASAP7_75t_L g16744 ( 
.A(n_16193),
.Y(n_16744)
);

INVx1_ASAP7_75t_L g16745 ( 
.A(n_16247),
.Y(n_16745)
);

INVx1_ASAP7_75t_L g16746 ( 
.A(n_16251),
.Y(n_16746)
);

INVx2_ASAP7_75t_L g16747 ( 
.A(n_16291),
.Y(n_16747)
);

OR2x2_ASAP7_75t_L g16748 ( 
.A(n_16117),
.B(n_8550),
.Y(n_16748)
);

OAI32xp33_ASAP7_75t_L g16749 ( 
.A1(n_16078),
.A2(n_9322),
.A3(n_9334),
.B1(n_9285),
.B2(n_9284),
.Y(n_16749)
);

INVxp33_ASAP7_75t_L g16750 ( 
.A(n_16257),
.Y(n_16750)
);

AND2x2_ASAP7_75t_L g16751 ( 
.A(n_16206),
.B(n_8544),
.Y(n_16751)
);

AND2x2_ASAP7_75t_L g16752 ( 
.A(n_16209),
.B(n_8544),
.Y(n_16752)
);

INVx1_ASAP7_75t_L g16753 ( 
.A(n_16263),
.Y(n_16753)
);

INVx1_ASAP7_75t_L g16754 ( 
.A(n_16176),
.Y(n_16754)
);

AOI22xp5_ASAP7_75t_L g16755 ( 
.A1(n_16052),
.A2(n_8652),
.B1(n_8666),
.B2(n_8589),
.Y(n_16755)
);

OAI33xp33_ASAP7_75t_L g16756 ( 
.A1(n_16099),
.A2(n_9340),
.A3(n_9334),
.B1(n_9355),
.B2(n_9336),
.B3(n_9322),
.Y(n_16756)
);

HB1xp67_ASAP7_75t_L g16757 ( 
.A(n_16266),
.Y(n_16757)
);

INVx1_ASAP7_75t_L g16758 ( 
.A(n_16298),
.Y(n_16758)
);

INVx1_ASAP7_75t_L g16759 ( 
.A(n_16302),
.Y(n_16759)
);

AOI22xp5_ASAP7_75t_L g16760 ( 
.A1(n_16112),
.A2(n_8652),
.B1(n_8666),
.B2(n_8589),
.Y(n_16760)
);

INVx1_ASAP7_75t_L g16761 ( 
.A(n_16303),
.Y(n_16761)
);

INVx1_ASAP7_75t_L g16762 ( 
.A(n_16305),
.Y(n_16762)
);

NAND2xp5_ASAP7_75t_L g16763 ( 
.A(n_16194),
.B(n_9382),
.Y(n_16763)
);

INVx2_ASAP7_75t_L g16764 ( 
.A(n_16269),
.Y(n_16764)
);

NAND2xp5_ASAP7_75t_L g16765 ( 
.A(n_16211),
.B(n_9396),
.Y(n_16765)
);

AOI322xp5_ASAP7_75t_L g16766 ( 
.A1(n_16346),
.A2(n_9356),
.A3(n_9340),
.B1(n_9362),
.B2(n_9363),
.C1(n_9355),
.C2(n_9336),
.Y(n_16766)
);

INVx2_ASAP7_75t_SL g16767 ( 
.A(n_16270),
.Y(n_16767)
);

AOI22xp5_ASAP7_75t_L g16768 ( 
.A1(n_16406),
.A2(n_8652),
.B1(n_8666),
.B2(n_8589),
.Y(n_16768)
);

INVx1_ASAP7_75t_L g16769 ( 
.A(n_16306),
.Y(n_16769)
);

INVx1_ASAP7_75t_L g16770 ( 
.A(n_16248),
.Y(n_16770)
);

OAI32xp33_ASAP7_75t_L g16771 ( 
.A1(n_16198),
.A2(n_9362),
.A3(n_9363),
.B1(n_9356),
.B2(n_9355),
.Y(n_16771)
);

INVxp67_ASAP7_75t_L g16772 ( 
.A(n_16228),
.Y(n_16772)
);

INVx1_ASAP7_75t_L g16773 ( 
.A(n_16256),
.Y(n_16773)
);

NAND2xp5_ASAP7_75t_L g16774 ( 
.A(n_16244),
.B(n_9396),
.Y(n_16774)
);

OA222x2_ASAP7_75t_L g16775 ( 
.A1(n_16108),
.A2(n_8994),
.B1(n_8987),
.B2(n_8996),
.C1(n_8993),
.C2(n_8953),
.Y(n_16775)
);

OAI32xp33_ASAP7_75t_L g16776 ( 
.A1(n_16115),
.A2(n_9363),
.A3(n_9367),
.B1(n_9362),
.B2(n_9356),
.Y(n_16776)
);

INVx1_ASAP7_75t_L g16777 ( 
.A(n_16217),
.Y(n_16777)
);

INVxp67_ASAP7_75t_L g16778 ( 
.A(n_16229),
.Y(n_16778)
);

AND2x2_ASAP7_75t_L g16779 ( 
.A(n_16347),
.B(n_8652),
.Y(n_16779)
);

AND3x1_ASAP7_75t_L g16780 ( 
.A(n_16366),
.B(n_8822),
.C(n_8666),
.Y(n_16780)
);

OAI22xp5_ASAP7_75t_L g16781 ( 
.A1(n_16367),
.A2(n_8822),
.B1(n_8866),
.B2(n_8666),
.Y(n_16781)
);

INVx1_ASAP7_75t_L g16782 ( 
.A(n_16152),
.Y(n_16782)
);

OAI22xp33_ASAP7_75t_L g16783 ( 
.A1(n_16156),
.A2(n_9367),
.B1(n_8993),
.B2(n_8994),
.Y(n_16783)
);

NOR2xp33_ASAP7_75t_L g16784 ( 
.A(n_16382),
.B(n_8822),
.Y(n_16784)
);

INVx1_ASAP7_75t_L g16785 ( 
.A(n_16162),
.Y(n_16785)
);

INVx1_ASAP7_75t_L g16786 ( 
.A(n_16187),
.Y(n_16786)
);

AND2x2_ASAP7_75t_L g16787 ( 
.A(n_16389),
.B(n_8822),
.Y(n_16787)
);

AOI32xp33_ASAP7_75t_L g16788 ( 
.A1(n_16277),
.A2(n_9367),
.A3(n_10857),
.B1(n_10865),
.B2(n_10855),
.Y(n_16788)
);

NAND2xp5_ASAP7_75t_L g16789 ( 
.A(n_16390),
.B(n_9398),
.Y(n_16789)
);

AOI33xp33_ASAP7_75t_L g16790 ( 
.A1(n_16401),
.A2(n_8915),
.A3(n_8933),
.B1(n_8646),
.B2(n_8993),
.B3(n_8987),
.Y(n_16790)
);

NAND2x2_ASAP7_75t_L g16791 ( 
.A(n_16100),
.B(n_6740),
.Y(n_16791)
);

NOR2xp33_ASAP7_75t_SL g16792 ( 
.A(n_16309),
.B(n_16327),
.Y(n_16792)
);

NAND2xp5_ASAP7_75t_L g16793 ( 
.A(n_16336),
.B(n_9398),
.Y(n_16793)
);

HB1xp67_ASAP7_75t_L g16794 ( 
.A(n_16281),
.Y(n_16794)
);

NAND3xp33_ASAP7_75t_L g16795 ( 
.A(n_16199),
.B(n_9872),
.C(n_9673),
.Y(n_16795)
);

AOI22xp5_ASAP7_75t_L g16796 ( 
.A1(n_16407),
.A2(n_8866),
.B1(n_8822),
.B2(n_8416),
.Y(n_16796)
);

AND2x2_ASAP7_75t_L g16797 ( 
.A(n_16242),
.B(n_8866),
.Y(n_16797)
);

O2A1O1Ixp5_ASAP7_75t_R g16798 ( 
.A1(n_16274),
.A2(n_8065),
.B(n_6913),
.C(n_6932),
.Y(n_16798)
);

INVx1_ASAP7_75t_L g16799 ( 
.A(n_16293),
.Y(n_16799)
);

INVx2_ASAP7_75t_L g16800 ( 
.A(n_16284),
.Y(n_16800)
);

AOI22xp33_ASAP7_75t_L g16801 ( 
.A1(n_16289),
.A2(n_8857),
.B1(n_9673),
.B2(n_9653),
.Y(n_16801)
);

NAND4xp75_ASAP7_75t_L g16802 ( 
.A(n_16278),
.B(n_9694),
.C(n_9635),
.D(n_10077),
.Y(n_16802)
);

OR2x2_ASAP7_75t_L g16803 ( 
.A(n_16342),
.B(n_10077),
.Y(n_16803)
);

NAND4xp25_ASAP7_75t_L g16804 ( 
.A(n_16348),
.B(n_6750),
.C(n_6759),
.D(n_6740),
.Y(n_16804)
);

INVx1_ASAP7_75t_L g16805 ( 
.A(n_16223),
.Y(n_16805)
);

AND2x2_ASAP7_75t_L g16806 ( 
.A(n_16351),
.B(n_8866),
.Y(n_16806)
);

AND2x4_ASAP7_75t_L g16807 ( 
.A(n_16360),
.B(n_10867),
.Y(n_16807)
);

INVx1_ASAP7_75t_SL g16808 ( 
.A(n_16275),
.Y(n_16808)
);

OAI22xp5_ASAP7_75t_L g16809 ( 
.A1(n_16372),
.A2(n_8866),
.B1(n_8994),
.B2(n_8987),
.Y(n_16809)
);

INVx2_ASAP7_75t_L g16810 ( 
.A(n_16292),
.Y(n_16810)
);

AOI22xp5_ASAP7_75t_L g16811 ( 
.A1(n_16408),
.A2(n_8416),
.B1(n_8420),
.B2(n_8247),
.Y(n_16811)
);

AND2x2_ASAP7_75t_L g16812 ( 
.A(n_16356),
.B(n_8416),
.Y(n_16812)
);

AND2x2_ASAP7_75t_L g16813 ( 
.A(n_16373),
.B(n_8416),
.Y(n_16813)
);

NAND2xp5_ASAP7_75t_L g16814 ( 
.A(n_16282),
.B(n_9406),
.Y(n_16814)
);

AND2x2_ASAP7_75t_L g16815 ( 
.A(n_16378),
.B(n_8416),
.Y(n_16815)
);

INVx1_ASAP7_75t_L g16816 ( 
.A(n_16300),
.Y(n_16816)
);

INVx1_ASAP7_75t_L g16817 ( 
.A(n_16308),
.Y(n_16817)
);

OAI22xp33_ASAP7_75t_L g16818 ( 
.A1(n_16379),
.A2(n_8996),
.B1(n_9005),
.B2(n_9004),
.Y(n_16818)
);

NAND2xp5_ASAP7_75t_L g16819 ( 
.A(n_16307),
.B(n_9406),
.Y(n_16819)
);

NAND2xp5_ASAP7_75t_SL g16820 ( 
.A(n_16612),
.B(n_16370),
.Y(n_16820)
);

OR2x2_ASAP7_75t_L g16821 ( 
.A(n_16430),
.B(n_16241),
.Y(n_16821)
);

AND2x2_ASAP7_75t_L g16822 ( 
.A(n_16417),
.B(n_16383),
.Y(n_16822)
);

INVx1_ASAP7_75t_SL g16823 ( 
.A(n_16501),
.Y(n_16823)
);

AND2x2_ASAP7_75t_L g16824 ( 
.A(n_16486),
.B(n_16396),
.Y(n_16824)
);

OR2x2_ASAP7_75t_L g16825 ( 
.A(n_16460),
.B(n_16311),
.Y(n_16825)
);

AND4x1_ASAP7_75t_L g16826 ( 
.A(n_16418),
.B(n_16361),
.C(n_16352),
.D(n_16358),
.Y(n_16826)
);

AND2x2_ASAP7_75t_L g16827 ( 
.A(n_16594),
.B(n_16402),
.Y(n_16827)
);

AND2x2_ASAP7_75t_L g16828 ( 
.A(n_16539),
.B(n_16506),
.Y(n_16828)
);

INVx1_ASAP7_75t_L g16829 ( 
.A(n_16426),
.Y(n_16829)
);

HB1xp67_ASAP7_75t_L g16830 ( 
.A(n_16534),
.Y(n_16830)
);

INVx1_ASAP7_75t_L g16831 ( 
.A(n_16732),
.Y(n_16831)
);

NOR2xp33_ASAP7_75t_L g16832 ( 
.A(n_16513),
.B(n_16261),
.Y(n_16832)
);

INVx1_ASAP7_75t_L g16833 ( 
.A(n_16657),
.Y(n_16833)
);

NAND2xp5_ASAP7_75t_SL g16834 ( 
.A(n_16425),
.B(n_16093),
.Y(n_16834)
);

INVx1_ASAP7_75t_L g16835 ( 
.A(n_16665),
.Y(n_16835)
);

OR2x2_ASAP7_75t_L g16836 ( 
.A(n_16481),
.B(n_16375),
.Y(n_16836)
);

AND2x4_ASAP7_75t_L g16837 ( 
.A(n_16478),
.B(n_16411),
.Y(n_16837)
);

OAI33xp33_ASAP7_75t_L g16838 ( 
.A1(n_16433),
.A2(n_16409),
.A3(n_16393),
.B1(n_16339),
.B2(n_16340),
.B3(n_16325),
.Y(n_16838)
);

INVx1_ASAP7_75t_L g16839 ( 
.A(n_16424),
.Y(n_16839)
);

INVx1_ASAP7_75t_L g16840 ( 
.A(n_16500),
.Y(n_16840)
);

AND2x2_ASAP7_75t_L g16841 ( 
.A(n_16480),
.B(n_16415),
.Y(n_16841)
);

NAND2xp5_ASAP7_75t_L g16842 ( 
.A(n_16444),
.B(n_16312),
.Y(n_16842)
);

NAND2xp5_ASAP7_75t_L g16843 ( 
.A(n_16427),
.B(n_16323),
.Y(n_16843)
);

OR2x2_ASAP7_75t_L g16844 ( 
.A(n_16546),
.B(n_16377),
.Y(n_16844)
);

OR2x2_ASAP7_75t_L g16845 ( 
.A(n_16609),
.B(n_16380),
.Y(n_16845)
);

AND2x2_ASAP7_75t_L g16846 ( 
.A(n_16504),
.B(n_16451),
.Y(n_16846)
);

NAND4xp25_ASAP7_75t_L g16847 ( 
.A(n_16477),
.B(n_16371),
.C(n_16357),
.D(n_16240),
.Y(n_16847)
);

AOI211x1_ASAP7_75t_SL g16848 ( 
.A1(n_16422),
.A2(n_16355),
.B(n_16333),
.C(n_16023),
.Y(n_16848)
);

AND2x4_ASAP7_75t_L g16849 ( 
.A(n_16471),
.B(n_16319),
.Y(n_16849)
);

INVx1_ASAP7_75t_L g16850 ( 
.A(n_16553),
.Y(n_16850)
);

OAI22xp5_ASAP7_75t_L g16851 ( 
.A1(n_16518),
.A2(n_16250),
.B1(n_16330),
.B2(n_16329),
.Y(n_16851)
);

OAI31xp33_ASAP7_75t_L g16852 ( 
.A1(n_16431),
.A2(n_16574),
.A3(n_16580),
.B(n_16616),
.Y(n_16852)
);

NOR2x1_ASAP7_75t_L g16853 ( 
.A(n_16689),
.B(n_16315),
.Y(n_16853)
);

AND2x2_ASAP7_75t_L g16854 ( 
.A(n_16545),
.B(n_16318),
.Y(n_16854)
);

AND2x2_ASAP7_75t_L g16855 ( 
.A(n_16476),
.B(n_16320),
.Y(n_16855)
);

AND2x2_ASAP7_75t_L g16856 ( 
.A(n_16485),
.B(n_16326),
.Y(n_16856)
);

INVx1_ASAP7_75t_L g16857 ( 
.A(n_16416),
.Y(n_16857)
);

AND2x2_ASAP7_75t_L g16858 ( 
.A(n_16465),
.B(n_16337),
.Y(n_16858)
);

INVx2_ASAP7_75t_L g16859 ( 
.A(n_16419),
.Y(n_16859)
);

NAND2xp5_ASAP7_75t_L g16860 ( 
.A(n_16443),
.B(n_16338),
.Y(n_16860)
);

AND2x2_ASAP7_75t_L g16861 ( 
.A(n_16491),
.B(n_16345),
.Y(n_16861)
);

OAI33xp33_ASAP7_75t_L g16862 ( 
.A1(n_16649),
.A2(n_16331),
.A3(n_16341),
.B1(n_16335),
.B2(n_16332),
.B3(n_16321),
.Y(n_16862)
);

NOR2xp33_ASAP7_75t_L g16863 ( 
.A(n_16570),
.B(n_16272),
.Y(n_16863)
);

NAND2xp5_ASAP7_75t_SL g16864 ( 
.A(n_16526),
.B(n_16234),
.Y(n_16864)
);

INVxp67_ASAP7_75t_L g16865 ( 
.A(n_16540),
.Y(n_16865)
);

INVx1_ASAP7_75t_L g16866 ( 
.A(n_16419),
.Y(n_16866)
);

NAND2xp5_ASAP7_75t_L g16867 ( 
.A(n_16428),
.B(n_16363),
.Y(n_16867)
);

INVx1_ASAP7_75t_L g16868 ( 
.A(n_16492),
.Y(n_16868)
);

AOI221xp5_ASAP7_75t_L g16869 ( 
.A1(n_16622),
.A2(n_16392),
.B1(n_16124),
.B2(n_16385),
.C(n_16368),
.Y(n_16869)
);

OAI211xp5_ASAP7_75t_SL g16870 ( 
.A1(n_16436),
.A2(n_16316),
.B(n_16268),
.C(n_16245),
.Y(n_16870)
);

INVx1_ASAP7_75t_L g16871 ( 
.A(n_16757),
.Y(n_16871)
);

AND2x4_ASAP7_75t_L g16872 ( 
.A(n_16671),
.B(n_8196),
.Y(n_16872)
);

AND2x2_ASAP7_75t_L g16873 ( 
.A(n_16475),
.B(n_16245),
.Y(n_16873)
);

INVx1_ASAP7_75t_L g16874 ( 
.A(n_16794),
.Y(n_16874)
);

INVx2_ASAP7_75t_L g16875 ( 
.A(n_16421),
.Y(n_16875)
);

HB1xp67_ASAP7_75t_L g16876 ( 
.A(n_16421),
.Y(n_16876)
);

OR2x2_ASAP7_75t_L g16877 ( 
.A(n_16581),
.B(n_10077),
.Y(n_16877)
);

HB1xp67_ASAP7_75t_L g16878 ( 
.A(n_16603),
.Y(n_16878)
);

INVx2_ASAP7_75t_L g16879 ( 
.A(n_16439),
.Y(n_16879)
);

INVx1_ASAP7_75t_L g16880 ( 
.A(n_16635),
.Y(n_16880)
);

OR2x6_ASAP7_75t_L g16881 ( 
.A(n_16689),
.B(n_6740),
.Y(n_16881)
);

INVx1_ASAP7_75t_L g16882 ( 
.A(n_16656),
.Y(n_16882)
);

HB1xp67_ASAP7_75t_L g16883 ( 
.A(n_16525),
.Y(n_16883)
);

CKINVDCx6p67_ASAP7_75t_R g16884 ( 
.A(n_16735),
.Y(n_16884)
);

NOR4xp25_ASAP7_75t_SL g16885 ( 
.A(n_16453),
.B(n_9411),
.C(n_9415),
.D(n_9409),
.Y(n_16885)
);

NOR2xp33_ASAP7_75t_R g16886 ( 
.A(n_16493),
.B(n_8896),
.Y(n_16886)
);

OAI21xp5_ASAP7_75t_L g16887 ( 
.A1(n_16473),
.A2(n_11239),
.B(n_10907),
.Y(n_16887)
);

AOI22xp5_ASAP7_75t_L g16888 ( 
.A1(n_16522),
.A2(n_10169),
.B1(n_10226),
.B2(n_10077),
.Y(n_16888)
);

INVx1_ASAP7_75t_L g16889 ( 
.A(n_16463),
.Y(n_16889)
);

OR2x2_ASAP7_75t_L g16890 ( 
.A(n_16450),
.B(n_10169),
.Y(n_16890)
);

CKINVDCx16_ASAP7_75t_R g16891 ( 
.A(n_16423),
.Y(n_16891)
);

INVx1_ASAP7_75t_L g16892 ( 
.A(n_16482),
.Y(n_16892)
);

NAND2xp5_ASAP7_75t_L g16893 ( 
.A(n_16767),
.B(n_9409),
.Y(n_16893)
);

INVx1_ASAP7_75t_L g16894 ( 
.A(n_16552),
.Y(n_16894)
);

AND2x2_ASAP7_75t_L g16895 ( 
.A(n_16487),
.B(n_10169),
.Y(n_16895)
);

NAND2xp5_ASAP7_75t_L g16896 ( 
.A(n_16714),
.B(n_9411),
.Y(n_16896)
);

INVx1_ASAP7_75t_L g16897 ( 
.A(n_16502),
.Y(n_16897)
);

NAND3xp33_ASAP7_75t_L g16898 ( 
.A(n_16429),
.B(n_9694),
.C(n_9635),
.Y(n_16898)
);

NAND2xp5_ASAP7_75t_L g16899 ( 
.A(n_16578),
.B(n_9415),
.Y(n_16899)
);

OAI31xp33_ASAP7_75t_L g16900 ( 
.A1(n_16438),
.A2(n_9004),
.A3(n_9005),
.B(n_8996),
.Y(n_16900)
);

INVx1_ASAP7_75t_L g16901 ( 
.A(n_16495),
.Y(n_16901)
);

NOR2xp33_ASAP7_75t_R g16902 ( 
.A(n_16559),
.B(n_8896),
.Y(n_16902)
);

NOR2xp33_ASAP7_75t_L g16903 ( 
.A(n_16496),
.B(n_8915),
.Y(n_16903)
);

INVx1_ASAP7_75t_L g16904 ( 
.A(n_16499),
.Y(n_16904)
);

INVx1_ASAP7_75t_SL g16905 ( 
.A(n_16808),
.Y(n_16905)
);

INVx1_ASAP7_75t_L g16906 ( 
.A(n_16455),
.Y(n_16906)
);

INVx1_ASAP7_75t_SL g16907 ( 
.A(n_16661),
.Y(n_16907)
);

NAND3xp33_ASAP7_75t_SL g16908 ( 
.A(n_16652),
.B(n_8933),
.C(n_8066),
.Y(n_16908)
);

HB1xp67_ASAP7_75t_L g16909 ( 
.A(n_16440),
.Y(n_16909)
);

AND2x4_ASAP7_75t_L g16910 ( 
.A(n_16606),
.B(n_8196),
.Y(n_16910)
);

CKINVDCx16_ASAP7_75t_R g16911 ( 
.A(n_16567),
.Y(n_16911)
);

AND2x2_ASAP7_75t_L g16912 ( 
.A(n_16613),
.B(n_10169),
.Y(n_16912)
);

NOR3xp33_ASAP7_75t_L g16913 ( 
.A(n_16550),
.B(n_9787),
.C(n_10867),
.Y(n_16913)
);

AOI21xp5_ASAP7_75t_L g16914 ( 
.A1(n_16696),
.A2(n_11142),
.B(n_11087),
.Y(n_16914)
);

NOR2x1_ASAP7_75t_L g16915 ( 
.A(n_16716),
.B(n_9004),
.Y(n_16915)
);

NOR2xp33_ASAP7_75t_L g16916 ( 
.A(n_16615),
.B(n_8065),
.Y(n_16916)
);

INVx1_ASAP7_75t_L g16917 ( 
.A(n_16619),
.Y(n_16917)
);

OR2x2_ASAP7_75t_L g16918 ( 
.A(n_16669),
.B(n_16677),
.Y(n_16918)
);

OR2x2_ASAP7_75t_L g16919 ( 
.A(n_16618),
.B(n_10226),
.Y(n_16919)
);

INVx1_ASAP7_75t_L g16920 ( 
.A(n_16458),
.Y(n_16920)
);

INVx1_ASAP7_75t_L g16921 ( 
.A(n_16461),
.Y(n_16921)
);

NOR2xp33_ASAP7_75t_L g16922 ( 
.A(n_16639),
.B(n_8201),
.Y(n_16922)
);

NAND2x1p5_ASAP7_75t_L g16923 ( 
.A(n_16717),
.B(n_6750),
.Y(n_16923)
);

NAND3xp33_ASAP7_75t_L g16924 ( 
.A(n_16435),
.B(n_9635),
.C(n_10226),
.Y(n_16924)
);

NAND2xp5_ASAP7_75t_L g16925 ( 
.A(n_16456),
.B(n_9417),
.Y(n_16925)
);

AND2x2_ASAP7_75t_L g16926 ( 
.A(n_16623),
.B(n_16626),
.Y(n_16926)
);

NAND2xp5_ASAP7_75t_L g16927 ( 
.A(n_16467),
.B(n_9417),
.Y(n_16927)
);

INVx1_ASAP7_75t_L g16928 ( 
.A(n_16638),
.Y(n_16928)
);

OR2x2_ASAP7_75t_L g16929 ( 
.A(n_16651),
.B(n_10226),
.Y(n_16929)
);

AND2x4_ASAP7_75t_L g16930 ( 
.A(n_16636),
.B(n_16637),
.Y(n_16930)
);

AND2x2_ASAP7_75t_L g16931 ( 
.A(n_16577),
.B(n_16587),
.Y(n_16931)
);

NOR2x1_ASAP7_75t_L g16932 ( 
.A(n_16629),
.B(n_16690),
.Y(n_16932)
);

AND2x2_ASAP7_75t_L g16933 ( 
.A(n_16579),
.B(n_10234),
.Y(n_16933)
);

NAND2xp5_ASAP7_75t_L g16934 ( 
.A(n_16658),
.B(n_9419),
.Y(n_16934)
);

NOR3xp33_ASAP7_75t_L g16935 ( 
.A(n_16564),
.B(n_9787),
.C(n_10906),
.Y(n_16935)
);

AND2x2_ASAP7_75t_L g16936 ( 
.A(n_16715),
.B(n_10234),
.Y(n_16936)
);

INVx2_ASAP7_75t_L g16937 ( 
.A(n_16719),
.Y(n_16937)
);

HB1xp67_ASAP7_75t_L g16938 ( 
.A(n_16614),
.Y(n_16938)
);

NAND2xp5_ASAP7_75t_L g16939 ( 
.A(n_16659),
.B(n_9419),
.Y(n_16939)
);

NAND2xp33_ASAP7_75t_L g16940 ( 
.A(n_16624),
.B(n_9420),
.Y(n_16940)
);

NAND4xp25_ASAP7_75t_L g16941 ( 
.A(n_16512),
.B(n_6759),
.C(n_6811),
.D(n_6750),
.Y(n_16941)
);

NAND2xp5_ASAP7_75t_L g16942 ( 
.A(n_16664),
.B(n_9420),
.Y(n_16942)
);

INVx1_ASAP7_75t_L g16943 ( 
.A(n_16740),
.Y(n_16943)
);

OR2x2_ASAP7_75t_L g16944 ( 
.A(n_16747),
.B(n_10234),
.Y(n_16944)
);

AND2x2_ASAP7_75t_L g16945 ( 
.A(n_16764),
.B(n_10234),
.Y(n_16945)
);

INVx1_ASAP7_75t_L g16946 ( 
.A(n_16691),
.Y(n_16946)
);

BUFx3_ASAP7_75t_L g16947 ( 
.A(n_16521),
.Y(n_16947)
);

NAND2x1p5_ASAP7_75t_L g16948 ( 
.A(n_16490),
.B(n_6750),
.Y(n_16948)
);

NAND2xp33_ASAP7_75t_SL g16949 ( 
.A(n_16750),
.B(n_16722),
.Y(n_16949)
);

INVx1_ASAP7_75t_L g16950 ( 
.A(n_16692),
.Y(n_16950)
);

AND2x2_ASAP7_75t_L g16951 ( 
.A(n_16686),
.B(n_10254),
.Y(n_16951)
);

INVxp67_ASAP7_75t_SL g16952 ( 
.A(n_16608),
.Y(n_16952)
);

OAI33xp33_ASAP7_75t_L g16953 ( 
.A1(n_16508),
.A2(n_9016),
.A3(n_9006),
.B1(n_9018),
.B2(n_9010),
.B3(n_9005),
.Y(n_16953)
);

OR2x2_ASAP7_75t_L g16954 ( 
.A(n_16800),
.B(n_10254),
.Y(n_16954)
);

NAND5xp2_ASAP7_75t_SL g16955 ( 
.A(n_16527),
.B(n_7892),
.C(n_7900),
.D(n_7875),
.E(n_7782),
.Y(n_16955)
);

NOR2xp33_ASAP7_75t_L g16956 ( 
.A(n_16772),
.B(n_8201),
.Y(n_16956)
);

NAND2xp5_ASAP7_75t_L g16957 ( 
.A(n_16523),
.B(n_9421),
.Y(n_16957)
);

AND2x2_ASAP7_75t_L g16958 ( 
.A(n_16561),
.B(n_10254),
.Y(n_16958)
);

NAND2xp33_ASAP7_75t_SL g16959 ( 
.A(n_16723),
.B(n_8441),
.Y(n_16959)
);

NOR2x1_ASAP7_75t_L g16960 ( 
.A(n_16728),
.B(n_9006),
.Y(n_16960)
);

NOR2xp33_ASAP7_75t_L g16961 ( 
.A(n_16778),
.B(n_8209),
.Y(n_16961)
);

INVx1_ASAP7_75t_L g16962 ( 
.A(n_16544),
.Y(n_16962)
);

AND2x2_ASAP7_75t_SL g16963 ( 
.A(n_16792),
.B(n_7831),
.Y(n_16963)
);

AND2x2_ASAP7_75t_L g16964 ( 
.A(n_16633),
.B(n_10254),
.Y(n_16964)
);

OR2x2_ASAP7_75t_L g16965 ( 
.A(n_16582),
.B(n_10271),
.Y(n_16965)
);

INVx1_ASAP7_75t_L g16966 ( 
.A(n_16595),
.Y(n_16966)
);

INVx2_ASAP7_75t_L g16967 ( 
.A(n_16517),
.Y(n_16967)
);

INVx1_ASAP7_75t_L g16968 ( 
.A(n_16596),
.Y(n_16968)
);

INVxp67_ASAP7_75t_L g16969 ( 
.A(n_16466),
.Y(n_16969)
);

INVx2_ASAP7_75t_L g16970 ( 
.A(n_16489),
.Y(n_16970)
);

OR2x2_ASAP7_75t_L g16971 ( 
.A(n_16598),
.B(n_10271),
.Y(n_16971)
);

NAND2xp5_ASAP7_75t_L g16972 ( 
.A(n_16599),
.B(n_9421),
.Y(n_16972)
);

INVx1_ASAP7_75t_L g16973 ( 
.A(n_16600),
.Y(n_16973)
);

AND2x2_ASAP7_75t_L g16974 ( 
.A(n_16519),
.B(n_10271),
.Y(n_16974)
);

NOR2x2_ASAP7_75t_L g16975 ( 
.A(n_16810),
.B(n_7769),
.Y(n_16975)
);

AND2x2_ASAP7_75t_L g16976 ( 
.A(n_16542),
.B(n_10271),
.Y(n_16976)
);

INVx1_ASAP7_75t_L g16977 ( 
.A(n_16617),
.Y(n_16977)
);

NAND4xp25_ASAP7_75t_L g16978 ( 
.A(n_16655),
.B(n_16804),
.C(n_16676),
.D(n_16515),
.Y(n_16978)
);

INVx1_ASAP7_75t_L g16979 ( 
.A(n_16528),
.Y(n_16979)
);

OR2x2_ASAP7_75t_L g16980 ( 
.A(n_16721),
.B(n_9006),
.Y(n_16980)
);

INVx2_ASAP7_75t_L g16981 ( 
.A(n_16484),
.Y(n_16981)
);

AND2x2_ASAP7_75t_L g16982 ( 
.A(n_16687),
.B(n_8420),
.Y(n_16982)
);

AND2x2_ASAP7_75t_L g16983 ( 
.A(n_16607),
.B(n_8420),
.Y(n_16983)
);

NOR3xp33_ASAP7_75t_SL g16984 ( 
.A(n_16494),
.B(n_6826),
.C(n_7024),
.Y(n_16984)
);

AND2x2_ASAP7_75t_L g16985 ( 
.A(n_16611),
.B(n_8420),
.Y(n_16985)
);

OR2x2_ASAP7_75t_L g16986 ( 
.A(n_16758),
.B(n_9010),
.Y(n_16986)
);

AND2x2_ASAP7_75t_L g16987 ( 
.A(n_16688),
.B(n_8420),
.Y(n_16987)
);

INVx1_ASAP7_75t_L g16988 ( 
.A(n_16759),
.Y(n_16988)
);

INVx2_ASAP7_75t_L g16989 ( 
.A(n_16591),
.Y(n_16989)
);

NOR2xp67_ASAP7_75t_SL g16990 ( 
.A(n_16547),
.B(n_6759),
.Y(n_16990)
);

INVx1_ASAP7_75t_L g16991 ( 
.A(n_16761),
.Y(n_16991)
);

NAND2xp5_ASAP7_75t_L g16992 ( 
.A(n_16762),
.B(n_9422),
.Y(n_16992)
);

AND2x2_ASAP7_75t_L g16993 ( 
.A(n_16563),
.B(n_16668),
.Y(n_16993)
);

INVx3_ASAP7_75t_SL g16994 ( 
.A(n_16644),
.Y(n_16994)
);

NOR2xp33_ASAP7_75t_L g16995 ( 
.A(n_16769),
.B(n_8209),
.Y(n_16995)
);

AND2x2_ASAP7_75t_L g16996 ( 
.A(n_16672),
.B(n_8420),
.Y(n_16996)
);

NOR2xp33_ASAP7_75t_L g16997 ( 
.A(n_16678),
.B(n_16679),
.Y(n_16997)
);

INVxp67_ASAP7_75t_SL g16998 ( 
.A(n_16731),
.Y(n_16998)
);

AND2x2_ASAP7_75t_L g16999 ( 
.A(n_16680),
.B(n_7875),
.Y(n_16999)
);

INVx1_ASAP7_75t_L g17000 ( 
.A(n_16710),
.Y(n_17000)
);

NOR2xp33_ASAP7_75t_R g17001 ( 
.A(n_16711),
.B(n_8896),
.Y(n_17001)
);

AND2x2_ASAP7_75t_L g17002 ( 
.A(n_16630),
.B(n_7875),
.Y(n_17002)
);

A2O1A1Ixp33_ASAP7_75t_L g17003 ( 
.A1(n_16549),
.A2(n_10907),
.B(n_10927),
.C(n_10906),
.Y(n_17003)
);

AND2x2_ASAP7_75t_L g17004 ( 
.A(n_16663),
.B(n_7892),
.Y(n_17004)
);

AND2x4_ASAP7_75t_L g17005 ( 
.A(n_16558),
.B(n_8211),
.Y(n_17005)
);

AND2x4_ASAP7_75t_L g17006 ( 
.A(n_16733),
.B(n_8211),
.Y(n_17006)
);

NOR2xp33_ASAP7_75t_L g17007 ( 
.A(n_16736),
.B(n_8216),
.Y(n_17007)
);

AOI21xp5_ASAP7_75t_L g17008 ( 
.A1(n_16770),
.A2(n_11142),
.B(n_9016),
.Y(n_17008)
);

INVx1_ASAP7_75t_L g17009 ( 
.A(n_16773),
.Y(n_17009)
);

NAND2xp5_ASAP7_75t_L g17010 ( 
.A(n_16667),
.B(n_9422),
.Y(n_17010)
);

AOI31xp33_ASAP7_75t_SL g17011 ( 
.A1(n_16693),
.A2(n_9010),
.A3(n_9018),
.B(n_9016),
.Y(n_17011)
);

INVx1_ASAP7_75t_L g17012 ( 
.A(n_16548),
.Y(n_17012)
);

INVx2_ASAP7_75t_L g17013 ( 
.A(n_16605),
.Y(n_17013)
);

NOR3xp33_ASAP7_75t_SL g17014 ( 
.A(n_16799),
.B(n_7024),
.C(n_7866),
.Y(n_17014)
);

OR2x2_ASAP7_75t_L g17015 ( 
.A(n_16640),
.B(n_9018),
.Y(n_17015)
);

OAI21xp33_ASAP7_75t_L g17016 ( 
.A1(n_16555),
.A2(n_9526),
.B(n_9525),
.Y(n_17016)
);

AOI22xp5_ASAP7_75t_L g17017 ( 
.A1(n_16682),
.A2(n_9635),
.B1(n_8247),
.B2(n_9375),
.Y(n_17017)
);

NOR2xp33_ASAP7_75t_L g17018 ( 
.A(n_16805),
.B(n_16816),
.Y(n_17018)
);

OR2x2_ASAP7_75t_L g17019 ( 
.A(n_16654),
.B(n_9023),
.Y(n_17019)
);

OR2x2_ASAP7_75t_L g17020 ( 
.A(n_16621),
.B(n_9023),
.Y(n_17020)
);

NAND2xp5_ASAP7_75t_L g17021 ( 
.A(n_16645),
.B(n_9423),
.Y(n_17021)
);

OR2x2_ASAP7_75t_L g17022 ( 
.A(n_16625),
.B(n_9023),
.Y(n_17022)
);

AND2x2_ASAP7_75t_SL g17023 ( 
.A(n_16817),
.B(n_8862),
.Y(n_17023)
);

INVx2_ASAP7_75t_L g17024 ( 
.A(n_16631),
.Y(n_17024)
);

INVx4_ASAP7_75t_L g17025 ( 
.A(n_16700),
.Y(n_17025)
);

INVx1_ASAP7_75t_L g17026 ( 
.A(n_16437),
.Y(n_17026)
);

OR2x2_ASAP7_75t_L g17027 ( 
.A(n_16670),
.B(n_9051),
.Y(n_17027)
);

AND2x2_ASAP7_75t_L g17028 ( 
.A(n_16557),
.B(n_7892),
.Y(n_17028)
);

NOR2xp33_ASAP7_75t_L g17029 ( 
.A(n_16743),
.B(n_8216),
.Y(n_17029)
);

OR2x2_ASAP7_75t_L g17030 ( 
.A(n_16675),
.B(n_9051),
.Y(n_17030)
);

INVx1_ASAP7_75t_SL g17031 ( 
.A(n_16628),
.Y(n_17031)
);

CKINVDCx16_ASAP7_75t_R g17032 ( 
.A(n_16744),
.Y(n_17032)
);

AND2x2_ASAP7_75t_SL g17033 ( 
.A(n_16745),
.B(n_8862),
.Y(n_17033)
);

NAND2xp33_ASAP7_75t_R g17034 ( 
.A(n_16746),
.B(n_16753),
.Y(n_17034)
);

NAND2xp5_ASAP7_75t_L g17035 ( 
.A(n_16702),
.B(n_9423),
.Y(n_17035)
);

INVx2_ASAP7_75t_L g17036 ( 
.A(n_16446),
.Y(n_17036)
);

INVx4_ASAP7_75t_L g17037 ( 
.A(n_16704),
.Y(n_17037)
);

AND2x2_ASAP7_75t_L g17038 ( 
.A(n_16754),
.B(n_7900),
.Y(n_17038)
);

NAND2xp5_ASAP7_75t_L g17039 ( 
.A(n_16713),
.B(n_9424),
.Y(n_17039)
);

OR2x2_ASAP7_75t_L g17040 ( 
.A(n_16695),
.B(n_9051),
.Y(n_17040)
);

INVx1_ASAP7_75t_L g17041 ( 
.A(n_16643),
.Y(n_17041)
);

INVx1_ASAP7_75t_L g17042 ( 
.A(n_16445),
.Y(n_17042)
);

AND2x2_ASAP7_75t_L g17043 ( 
.A(n_16565),
.B(n_7900),
.Y(n_17043)
);

AOI21xp33_ASAP7_75t_L g17044 ( 
.A1(n_16556),
.A2(n_9526),
.B(n_9525),
.Y(n_17044)
);

OR2x6_ASAP7_75t_L g17045 ( 
.A(n_16777),
.B(n_6759),
.Y(n_17045)
);

AND2x4_ASAP7_75t_L g17046 ( 
.A(n_16782),
.B(n_16785),
.Y(n_17046)
);

OAI33xp33_ASAP7_75t_L g17047 ( 
.A1(n_16507),
.A2(n_9077),
.A3(n_9063),
.B1(n_9084),
.B2(n_9071),
.B3(n_9062),
.Y(n_17047)
);

OR2x2_ASAP7_75t_L g17048 ( 
.A(n_16730),
.B(n_9062),
.Y(n_17048)
);

OAI33xp33_ASAP7_75t_L g17049 ( 
.A1(n_16537),
.A2(n_9077),
.A3(n_9063),
.B1(n_9084),
.B2(n_9071),
.B3(n_9062),
.Y(n_17049)
);

CKINVDCx16_ASAP7_75t_R g17050 ( 
.A(n_16786),
.Y(n_17050)
);

NOR2xp33_ASAP7_75t_L g17051 ( 
.A(n_16646),
.B(n_8218),
.Y(n_17051)
);

NAND2xp5_ASAP7_75t_L g17052 ( 
.A(n_16585),
.B(n_9424),
.Y(n_17052)
);

AOI21xp33_ASAP7_75t_SL g17053 ( 
.A1(n_16572),
.A2(n_10956),
.B(n_10927),
.Y(n_17053)
);

INVx1_ASAP7_75t_SL g17054 ( 
.A(n_16720),
.Y(n_17054)
);

CKINVDCx20_ASAP7_75t_R g17055 ( 
.A(n_16511),
.Y(n_17055)
);

NAND2xp5_ASAP7_75t_L g17056 ( 
.A(n_16604),
.B(n_16681),
.Y(n_17056)
);

INVx2_ASAP7_75t_L g17057 ( 
.A(n_16474),
.Y(n_17057)
);

NOR2xp33_ASAP7_75t_L g17058 ( 
.A(n_16469),
.B(n_8218),
.Y(n_17058)
);

NAND2xp33_ASAP7_75t_SL g17059 ( 
.A(n_16454),
.B(n_16432),
.Y(n_17059)
);

AND2x2_ASAP7_75t_L g17060 ( 
.A(n_16660),
.B(n_7911),
.Y(n_17060)
);

NOR2xp33_ASAP7_75t_L g17061 ( 
.A(n_16573),
.B(n_16554),
.Y(n_17061)
);

AND2x2_ASAP7_75t_L g17062 ( 
.A(n_16514),
.B(n_7911),
.Y(n_17062)
);

INVx1_ASAP7_75t_SL g17063 ( 
.A(n_16779),
.Y(n_17063)
);

OR2x2_ASAP7_75t_L g17064 ( 
.A(n_16748),
.B(n_9063),
.Y(n_17064)
);

INVx2_ASAP7_75t_L g17065 ( 
.A(n_16470),
.Y(n_17065)
);

NAND2xp5_ASAP7_75t_L g17066 ( 
.A(n_16787),
.B(n_9425),
.Y(n_17066)
);

NOR2xp33_ASAP7_75t_L g17067 ( 
.A(n_16569),
.B(n_16571),
.Y(n_17067)
);

AND2x4_ASAP7_75t_L g17068 ( 
.A(n_16441),
.B(n_8224),
.Y(n_17068)
);

NOR2xp67_ASAP7_75t_L g17069 ( 
.A(n_16464),
.B(n_9425),
.Y(n_17069)
);

OR2x2_ASAP7_75t_L g17070 ( 
.A(n_16705),
.B(n_9071),
.Y(n_17070)
);

NAND2xp5_ASAP7_75t_L g17071 ( 
.A(n_16725),
.B(n_9427),
.Y(n_17071)
);

AND2x2_ASAP7_75t_L g17072 ( 
.A(n_16650),
.B(n_7911),
.Y(n_17072)
);

INVx2_ASAP7_75t_L g17073 ( 
.A(n_16488),
.Y(n_17073)
);

INVx3_ASAP7_75t_SL g17074 ( 
.A(n_16627),
.Y(n_17074)
);

HB1xp67_ASAP7_75t_L g17075 ( 
.A(n_16791),
.Y(n_17075)
);

INVxp67_ASAP7_75t_L g17076 ( 
.A(n_16784),
.Y(n_17076)
);

INVx1_ASAP7_75t_L g17077 ( 
.A(n_16789),
.Y(n_17077)
);

NOR2xp33_ASAP7_75t_R g17078 ( 
.A(n_16541),
.B(n_6811),
.Y(n_17078)
);

NAND2xp5_ASAP7_75t_L g17079 ( 
.A(n_16814),
.B(n_9427),
.Y(n_17079)
);

INVx2_ASAP7_75t_L g17080 ( 
.A(n_16529),
.Y(n_17080)
);

NAND2xp33_ASAP7_75t_SL g17081 ( 
.A(n_16683),
.B(n_8441),
.Y(n_17081)
);

NOR2xp33_ASAP7_75t_SL g17082 ( 
.A(n_16448),
.B(n_8656),
.Y(n_17082)
);

INVx1_ASAP7_75t_L g17083 ( 
.A(n_16763),
.Y(n_17083)
);

INVx1_ASAP7_75t_SL g17084 ( 
.A(n_16741),
.Y(n_17084)
);

NOR3xp33_ASAP7_75t_SL g17085 ( 
.A(n_16483),
.B(n_7921),
.C(n_7866),
.Y(n_17085)
);

INVx1_ASAP7_75t_L g17086 ( 
.A(n_16765),
.Y(n_17086)
);

INVx2_ASAP7_75t_L g17087 ( 
.A(n_16529),
.Y(n_17087)
);

INVx1_ASAP7_75t_L g17088 ( 
.A(n_16774),
.Y(n_17088)
);

NAND2xp33_ASAP7_75t_R g17089 ( 
.A(n_16718),
.B(n_16751),
.Y(n_17089)
);

INVx1_ASAP7_75t_L g17090 ( 
.A(n_16694),
.Y(n_17090)
);

AND2x2_ASAP7_75t_L g17091 ( 
.A(n_16797),
.B(n_7940),
.Y(n_17091)
);

INVx2_ASAP7_75t_L g17092 ( 
.A(n_16568),
.Y(n_17092)
);

INVx1_ASAP7_75t_L g17093 ( 
.A(n_16697),
.Y(n_17093)
);

OR2x2_ASAP7_75t_L g17094 ( 
.A(n_16712),
.B(n_9077),
.Y(n_17094)
);

INVx2_ASAP7_75t_L g17095 ( 
.A(n_16575),
.Y(n_17095)
);

OR2x2_ASAP7_75t_L g17096 ( 
.A(n_16729),
.B(n_9084),
.Y(n_17096)
);

NAND2xp33_ASAP7_75t_SL g17097 ( 
.A(n_16701),
.B(n_8441),
.Y(n_17097)
);

AOI22xp33_ASAP7_75t_L g17098 ( 
.A1(n_16597),
.A2(n_7963),
.B1(n_7979),
.B2(n_8386),
.Y(n_17098)
);

CKINVDCx16_ASAP7_75t_R g17099 ( 
.A(n_16798),
.Y(n_17099)
);

CKINVDCx16_ASAP7_75t_R g17100 ( 
.A(n_16533),
.Y(n_17100)
);

AND2x2_ASAP7_75t_L g17101 ( 
.A(n_16752),
.B(n_7940),
.Y(n_17101)
);

INVx1_ASAP7_75t_L g17102 ( 
.A(n_16707),
.Y(n_17102)
);

AND2x2_ASAP7_75t_L g17103 ( 
.A(n_16698),
.B(n_7940),
.Y(n_17103)
);

NAND2xp5_ASAP7_75t_L g17104 ( 
.A(n_16819),
.B(n_9434),
.Y(n_17104)
);

AND2x2_ASAP7_75t_L g17105 ( 
.A(n_16806),
.B(n_7959),
.Y(n_17105)
);

INVx1_ASAP7_75t_SL g17106 ( 
.A(n_16708),
.Y(n_17106)
);

CKINVDCx5p33_ASAP7_75t_R g17107 ( 
.A(n_16442),
.Y(n_17107)
);

OR2x2_ASAP7_75t_L g17108 ( 
.A(n_16793),
.B(n_9085),
.Y(n_17108)
);

INVx1_ASAP7_75t_L g17109 ( 
.A(n_16790),
.Y(n_17109)
);

INVx1_ASAP7_75t_L g17110 ( 
.A(n_16780),
.Y(n_17110)
);

INVx1_ASAP7_75t_L g17111 ( 
.A(n_16452),
.Y(n_17111)
);

INVx1_ASAP7_75t_L g17112 ( 
.A(n_16459),
.Y(n_17112)
);

NAND2xp5_ASAP7_75t_L g17113 ( 
.A(n_16503),
.B(n_9434),
.Y(n_17113)
);

OR2x2_ASAP7_75t_L g17114 ( 
.A(n_16536),
.B(n_9085),
.Y(n_17114)
);

NAND2xp5_ASAP7_75t_L g17115 ( 
.A(n_16449),
.B(n_9437),
.Y(n_17115)
);

NAND2xp5_ASAP7_75t_L g17116 ( 
.A(n_16516),
.B(n_9437),
.Y(n_17116)
);

INVx1_ASAP7_75t_L g17117 ( 
.A(n_16807),
.Y(n_17117)
);

INVxp67_ASAP7_75t_L g17118 ( 
.A(n_16718),
.Y(n_17118)
);

NAND2xp5_ASAP7_75t_L g17119 ( 
.A(n_16468),
.B(n_16666),
.Y(n_17119)
);

NAND3xp33_ASAP7_75t_SL g17120 ( 
.A(n_16479),
.B(n_8066),
.C(n_8043),
.Y(n_17120)
);

NAND2x1_ASAP7_75t_SL g17121 ( 
.A(n_16468),
.B(n_9085),
.Y(n_17121)
);

OR2x2_ASAP7_75t_L g17122 ( 
.A(n_16803),
.B(n_9089),
.Y(n_17122)
);

AND2x2_ASAP7_75t_L g17123 ( 
.A(n_16592),
.B(n_7959),
.Y(n_17123)
);

INVx1_ASAP7_75t_L g17124 ( 
.A(n_16807),
.Y(n_17124)
);

OAI31xp33_ASAP7_75t_L g17125 ( 
.A1(n_16505),
.A2(n_9098),
.A3(n_9113),
.B(n_9089),
.Y(n_17125)
);

OR2x2_ASAP7_75t_L g17126 ( 
.A(n_16535),
.B(n_9089),
.Y(n_17126)
);

NOR2xp33_ASAP7_75t_L g17127 ( 
.A(n_16576),
.B(n_16510),
.Y(n_17127)
);

INVx1_ASAP7_75t_L g17128 ( 
.A(n_16566),
.Y(n_17128)
);

AND2x2_ASAP7_75t_L g17129 ( 
.A(n_16812),
.B(n_7959),
.Y(n_17129)
);

NOR2xp33_ASAP7_75t_L g17130 ( 
.A(n_16632),
.B(n_8224),
.Y(n_17130)
);

INVx2_ASAP7_75t_L g17131 ( 
.A(n_16566),
.Y(n_17131)
);

NAND2xp5_ASAP7_75t_L g17132 ( 
.A(n_16509),
.B(n_9439),
.Y(n_17132)
);

INVx1_ASAP7_75t_L g17133 ( 
.A(n_16531),
.Y(n_17133)
);

NAND2xp5_ASAP7_75t_L g17134 ( 
.A(n_16498),
.B(n_9439),
.Y(n_17134)
);

NOR2xp33_ASAP7_75t_L g17135 ( 
.A(n_16610),
.B(n_16642),
.Y(n_17135)
);

INVxp33_ASAP7_75t_L g17136 ( 
.A(n_16524),
.Y(n_17136)
);

INVxp67_ASAP7_75t_SL g17137 ( 
.A(n_16532),
.Y(n_17137)
);

NAND2xp5_ASAP7_75t_L g17138 ( 
.A(n_16498),
.B(n_9444),
.Y(n_17138)
);

AND2x2_ASAP7_75t_L g17139 ( 
.A(n_16590),
.B(n_7978),
.Y(n_17139)
);

AND2x2_ASAP7_75t_L g17140 ( 
.A(n_16685),
.B(n_7978),
.Y(n_17140)
);

INVx2_ASAP7_75t_L g17141 ( 
.A(n_16738),
.Y(n_17141)
);

INVx3_ASAP7_75t_L g17142 ( 
.A(n_16738),
.Y(n_17142)
);

AND2x2_ASAP7_75t_L g17143 ( 
.A(n_16813),
.B(n_7978),
.Y(n_17143)
);

XNOR2x1_ASAP7_75t_L g17144 ( 
.A(n_16447),
.B(n_6811),
.Y(n_17144)
);

OAI33xp33_ASAP7_75t_L g17145 ( 
.A1(n_16551),
.A2(n_9126),
.A3(n_9113),
.B1(n_9130),
.B2(n_9121),
.B3(n_9098),
.Y(n_17145)
);

NAND2xp5_ASAP7_75t_SL g17146 ( 
.A(n_16524),
.B(n_10156),
.Y(n_17146)
);

AND2x2_ASAP7_75t_L g17147 ( 
.A(n_16815),
.B(n_7988),
.Y(n_17147)
);

INVx1_ASAP7_75t_L g17148 ( 
.A(n_16653),
.Y(n_17148)
);

NAND2xp33_ASAP7_75t_SL g17149 ( 
.A(n_16560),
.B(n_8653),
.Y(n_17149)
);

NAND2xp5_ASAP7_75t_L g17150 ( 
.A(n_16602),
.B(n_9444),
.Y(n_17150)
);

AND2x2_ASAP7_75t_SL g17151 ( 
.A(n_16684),
.B(n_8862),
.Y(n_17151)
);

OR2x2_ASAP7_75t_L g17152 ( 
.A(n_16674),
.B(n_9098),
.Y(n_17152)
);

NAND2xp5_ASAP7_75t_L g17153 ( 
.A(n_16788),
.B(n_9447),
.Y(n_17153)
);

INVx2_ASAP7_75t_SL g17154 ( 
.A(n_16593),
.Y(n_17154)
);

AND2x2_ASAP7_75t_L g17155 ( 
.A(n_16684),
.B(n_7988),
.Y(n_17155)
);

AOI21xp33_ASAP7_75t_L g17156 ( 
.A1(n_16497),
.A2(n_9526),
.B(n_9525),
.Y(n_17156)
);

AOI211xp5_ASAP7_75t_L g17157 ( 
.A1(n_16673),
.A2(n_16699),
.B(n_16739),
.C(n_16706),
.Y(n_17157)
);

NOR2xp33_ASAP7_75t_R g17158 ( 
.A(n_16726),
.B(n_6811),
.Y(n_17158)
);

INVx1_ASAP7_75t_SL g17159 ( 
.A(n_16726),
.Y(n_17159)
);

NAND2xp5_ASAP7_75t_L g17160 ( 
.A(n_16647),
.B(n_9447),
.Y(n_17160)
);

INVxp67_ASAP7_75t_L g17161 ( 
.A(n_16586),
.Y(n_17161)
);

NOR3xp33_ASAP7_75t_L g17162 ( 
.A(n_16588),
.B(n_10973),
.C(n_10956),
.Y(n_17162)
);

CKINVDCx8_ASAP7_75t_R g17163 ( 
.A(n_16586),
.Y(n_17163)
);

AND2x2_ASAP7_75t_L g17164 ( 
.A(n_16641),
.B(n_16760),
.Y(n_17164)
);

NAND2xp5_ASAP7_75t_L g17165 ( 
.A(n_16634),
.B(n_9448),
.Y(n_17165)
);

OR2x2_ASAP7_75t_L g17166 ( 
.A(n_16781),
.B(n_9113),
.Y(n_17166)
);

AND2x2_ASAP7_75t_L g17167 ( 
.A(n_16755),
.B(n_16768),
.Y(n_17167)
);

INVx1_ASAP7_75t_L g17168 ( 
.A(n_16462),
.Y(n_17168)
);

INVx2_ASAP7_75t_L g17169 ( 
.A(n_16520),
.Y(n_17169)
);

NAND3xp33_ASAP7_75t_SL g17170 ( 
.A(n_16727),
.B(n_8066),
.C(n_8043),
.Y(n_17170)
);

NOR2xp33_ASAP7_75t_L g17171 ( 
.A(n_16543),
.B(n_8227),
.Y(n_17171)
);

NOR3xp33_ASAP7_75t_L g17172 ( 
.A(n_16783),
.B(n_10973),
.C(n_9732),
.Y(n_17172)
);

OR2x2_ASAP7_75t_L g17173 ( 
.A(n_16742),
.B(n_9121),
.Y(n_17173)
);

OAI21xp5_ASAP7_75t_L g17174 ( 
.A1(n_16620),
.A2(n_16801),
.B(n_16795),
.Y(n_17174)
);

INVx1_ASAP7_75t_L g17175 ( 
.A(n_16584),
.Y(n_17175)
);

INVx1_ASAP7_75t_L g17176 ( 
.A(n_16776),
.Y(n_17176)
);

NAND2xp5_ASAP7_75t_L g17177 ( 
.A(n_16703),
.B(n_9448),
.Y(n_17177)
);

INVx1_ASAP7_75t_L g17178 ( 
.A(n_16538),
.Y(n_17178)
);

INVx1_ASAP7_75t_L g17179 ( 
.A(n_16749),
.Y(n_17179)
);

INVx1_ASAP7_75t_L g17180 ( 
.A(n_16771),
.Y(n_17180)
);

NAND2xp33_ASAP7_75t_R g17181 ( 
.A(n_16648),
.B(n_16530),
.Y(n_17181)
);

INVx1_ASAP7_75t_L g17182 ( 
.A(n_16809),
.Y(n_17182)
);

OR2x4_ASAP7_75t_L g17183 ( 
.A(n_16562),
.B(n_7320),
.Y(n_17183)
);

INVx1_ASAP7_75t_L g17184 ( 
.A(n_16818),
.Y(n_17184)
);

NOR2xp33_ASAP7_75t_L g17185 ( 
.A(n_16734),
.B(n_8227),
.Y(n_17185)
);

NAND2xp5_ASAP7_75t_L g17186 ( 
.A(n_16796),
.B(n_9450),
.Y(n_17186)
);

NAND2xp5_ASAP7_75t_L g17187 ( 
.A(n_16457),
.B(n_9450),
.Y(n_17187)
);

NAND3xp33_ASAP7_75t_SL g17188 ( 
.A(n_16434),
.B(n_8066),
.C(n_8043),
.Y(n_17188)
);

AND2x2_ASAP7_75t_L g17189 ( 
.A(n_16420),
.B(n_7988),
.Y(n_17189)
);

INVx1_ASAP7_75t_L g17190 ( 
.A(n_16802),
.Y(n_17190)
);

AND2x2_ASAP7_75t_L g17191 ( 
.A(n_16811),
.B(n_16775),
.Y(n_17191)
);

NAND2xp5_ASAP7_75t_L g17192 ( 
.A(n_16737),
.B(n_9454),
.Y(n_17192)
);

CKINVDCx16_ASAP7_75t_R g17193 ( 
.A(n_16662),
.Y(n_17193)
);

INVx2_ASAP7_75t_L g17194 ( 
.A(n_16709),
.Y(n_17194)
);

CKINVDCx20_ASAP7_75t_L g17195 ( 
.A(n_16589),
.Y(n_17195)
);

NAND2xp5_ASAP7_75t_L g17196 ( 
.A(n_16601),
.B(n_9454),
.Y(n_17196)
);

OR2x2_ASAP7_75t_L g17197 ( 
.A(n_16756),
.B(n_9121),
.Y(n_17197)
);

INVx1_ASAP7_75t_L g17198 ( 
.A(n_16472),
.Y(n_17198)
);

INVx1_ASAP7_75t_SL g17199 ( 
.A(n_16583),
.Y(n_17199)
);

INVx2_ASAP7_75t_L g17200 ( 
.A(n_16724),
.Y(n_17200)
);

NAND2xp5_ASAP7_75t_L g17201 ( 
.A(n_16766),
.B(n_9456),
.Y(n_17201)
);

NAND2xp5_ASAP7_75t_L g17202 ( 
.A(n_16417),
.B(n_9456),
.Y(n_17202)
);

AND2x2_ASAP7_75t_L g17203 ( 
.A(n_16417),
.B(n_8070),
.Y(n_17203)
);

AND2x2_ASAP7_75t_L g17204 ( 
.A(n_16417),
.B(n_8070),
.Y(n_17204)
);

INVx1_ASAP7_75t_L g17205 ( 
.A(n_16426),
.Y(n_17205)
);

AND2x2_ASAP7_75t_L g17206 ( 
.A(n_16417),
.B(n_8070),
.Y(n_17206)
);

NAND2xp5_ASAP7_75t_L g17207 ( 
.A(n_16911),
.B(n_9457),
.Y(n_17207)
);

OAI21x1_ASAP7_75t_L g17208 ( 
.A1(n_16853),
.A2(n_17194),
.B(n_17142),
.Y(n_17208)
);

OAI21xp33_ASAP7_75t_L g17209 ( 
.A1(n_16823),
.A2(n_9533),
.B(n_9531),
.Y(n_17209)
);

HB1xp67_ASAP7_75t_L g17210 ( 
.A(n_17193),
.Y(n_17210)
);

INVx2_ASAP7_75t_L g17211 ( 
.A(n_17121),
.Y(n_17211)
);

NAND2xp5_ASAP7_75t_L g17212 ( 
.A(n_16891),
.B(n_9457),
.Y(n_17212)
);

INVxp67_ASAP7_75t_L g17213 ( 
.A(n_16878),
.Y(n_17213)
);

NOR2xp33_ASAP7_75t_L g17214 ( 
.A(n_16865),
.B(n_8318),
.Y(n_17214)
);

INVx1_ASAP7_75t_SL g17215 ( 
.A(n_16884),
.Y(n_17215)
);

NAND2xp5_ASAP7_75t_SL g17216 ( 
.A(n_16852),
.B(n_10156),
.Y(n_17216)
);

INVx4_ASAP7_75t_L g17217 ( 
.A(n_16994),
.Y(n_17217)
);

OR2x2_ASAP7_75t_L g17218 ( 
.A(n_16859),
.B(n_9126),
.Y(n_17218)
);

AOI221xp5_ASAP7_75t_L g17219 ( 
.A1(n_16869),
.A2(n_9130),
.B1(n_9135),
.B2(n_9126),
.C(n_8656),
.Y(n_17219)
);

OR2x2_ASAP7_75t_L g17220 ( 
.A(n_16866),
.B(n_9130),
.Y(n_17220)
);

AOI22xp33_ASAP7_75t_L g17221 ( 
.A1(n_16932),
.A2(n_7963),
.B1(n_7979),
.B2(n_8386),
.Y(n_17221)
);

INVx2_ASAP7_75t_L g17222 ( 
.A(n_16828),
.Y(n_17222)
);

NOR2xp33_ASAP7_75t_L g17223 ( 
.A(n_16938),
.B(n_8318),
.Y(n_17223)
);

INVx1_ASAP7_75t_L g17224 ( 
.A(n_16883),
.Y(n_17224)
);

OR2x2_ASAP7_75t_L g17225 ( 
.A(n_16918),
.B(n_9135),
.Y(n_17225)
);

NOR2xp33_ASAP7_75t_L g17226 ( 
.A(n_16905),
.B(n_8326),
.Y(n_17226)
);

AND2x2_ASAP7_75t_L g17227 ( 
.A(n_16822),
.B(n_9274),
.Y(n_17227)
);

INVx1_ASAP7_75t_L g17228 ( 
.A(n_16876),
.Y(n_17228)
);

INVx1_ASAP7_75t_L g17229 ( 
.A(n_16952),
.Y(n_17229)
);

INVx3_ASAP7_75t_L g17230 ( 
.A(n_16881),
.Y(n_17230)
);

AND2x2_ASAP7_75t_L g17231 ( 
.A(n_16824),
.B(n_9278),
.Y(n_17231)
);

AND2x2_ASAP7_75t_L g17232 ( 
.A(n_16846),
.B(n_9287),
.Y(n_17232)
);

INVx1_ASAP7_75t_L g17233 ( 
.A(n_16854),
.Y(n_17233)
);

NOR2xp33_ASAP7_75t_L g17234 ( 
.A(n_16829),
.B(n_8326),
.Y(n_17234)
);

NOR2xp33_ASAP7_75t_L g17235 ( 
.A(n_17205),
.B(n_16880),
.Y(n_17235)
);

INVx1_ASAP7_75t_SL g17236 ( 
.A(n_16949),
.Y(n_17236)
);

AND2x4_ASAP7_75t_L g17237 ( 
.A(n_16882),
.B(n_8328),
.Y(n_17237)
);

INVx1_ASAP7_75t_L g17238 ( 
.A(n_16830),
.Y(n_17238)
);

OAI21x1_ASAP7_75t_L g17239 ( 
.A1(n_16820),
.A2(n_9303),
.B(n_9287),
.Y(n_17239)
);

CKINVDCx16_ASAP7_75t_R g17240 ( 
.A(n_17032),
.Y(n_17240)
);

INVxp67_ASAP7_75t_L g17241 ( 
.A(n_16990),
.Y(n_17241)
);

AND2x2_ASAP7_75t_L g17242 ( 
.A(n_16931),
.B(n_9287),
.Y(n_17242)
);

INVx1_ASAP7_75t_L g17243 ( 
.A(n_16839),
.Y(n_17243)
);

INVx1_ASAP7_75t_SL g17244 ( 
.A(n_16959),
.Y(n_17244)
);

INVx1_ASAP7_75t_L g17245 ( 
.A(n_17128),
.Y(n_17245)
);

INVx1_ASAP7_75t_L g17246 ( 
.A(n_16871),
.Y(n_17246)
);

AND2x2_ASAP7_75t_L g17247 ( 
.A(n_16937),
.B(n_9303),
.Y(n_17247)
);

INVx1_ASAP7_75t_L g17248 ( 
.A(n_16874),
.Y(n_17248)
);

NAND2xp5_ASAP7_75t_L g17249 ( 
.A(n_16831),
.B(n_9459),
.Y(n_17249)
);

BUFx3_ASAP7_75t_L g17250 ( 
.A(n_16881),
.Y(n_17250)
);

INVx1_ASAP7_75t_L g17251 ( 
.A(n_16840),
.Y(n_17251)
);

INVx1_ASAP7_75t_SL g17252 ( 
.A(n_16825),
.Y(n_17252)
);

INVx1_ASAP7_75t_L g17253 ( 
.A(n_16850),
.Y(n_17253)
);

INVx1_ASAP7_75t_L g17254 ( 
.A(n_16998),
.Y(n_17254)
);

INVx2_ASAP7_75t_L g17255 ( 
.A(n_17203),
.Y(n_17255)
);

BUFx2_ASAP7_75t_L g17256 ( 
.A(n_17158),
.Y(n_17256)
);

INVx1_ASAP7_75t_L g17257 ( 
.A(n_17131),
.Y(n_17257)
);

INVx1_ASAP7_75t_L g17258 ( 
.A(n_16833),
.Y(n_17258)
);

INVx1_ASAP7_75t_SL g17259 ( 
.A(n_17074),
.Y(n_17259)
);

OR2x2_ASAP7_75t_L g17260 ( 
.A(n_16879),
.B(n_9135),
.Y(n_17260)
);

INVx2_ASAP7_75t_L g17261 ( 
.A(n_17204),
.Y(n_17261)
);

INVx1_ASAP7_75t_L g17262 ( 
.A(n_16835),
.Y(n_17262)
);

INVx2_ASAP7_75t_L g17263 ( 
.A(n_17206),
.Y(n_17263)
);

NAND2xp5_ASAP7_75t_L g17264 ( 
.A(n_16857),
.B(n_9459),
.Y(n_17264)
);

INVx1_ASAP7_75t_SL g17265 ( 
.A(n_16923),
.Y(n_17265)
);

INVx1_ASAP7_75t_L g17266 ( 
.A(n_16861),
.Y(n_17266)
);

INVx2_ASAP7_75t_L g17267 ( 
.A(n_17189),
.Y(n_17267)
);

OR2x2_ASAP7_75t_L g17268 ( 
.A(n_16847),
.B(n_10156),
.Y(n_17268)
);

AO21x2_ASAP7_75t_L g17269 ( 
.A1(n_16868),
.A2(n_9732),
.B(n_9724),
.Y(n_17269)
);

HB1xp67_ASAP7_75t_L g17270 ( 
.A(n_17133),
.Y(n_17270)
);

INVx1_ASAP7_75t_L g17271 ( 
.A(n_17080),
.Y(n_17271)
);

NOR2xp33_ASAP7_75t_L g17272 ( 
.A(n_16907),
.B(n_16943),
.Y(n_17272)
);

AOI22xp33_ASAP7_75t_L g17273 ( 
.A1(n_16875),
.A2(n_7963),
.B1(n_7979),
.B2(n_7968),
.Y(n_17273)
);

INVx1_ASAP7_75t_L g17274 ( 
.A(n_17087),
.Y(n_17274)
);

AOI22xp33_ASAP7_75t_L g17275 ( 
.A1(n_16947),
.A2(n_7963),
.B1(n_7968),
.B2(n_7951),
.Y(n_17275)
);

OR2x2_ASAP7_75t_L g17276 ( 
.A(n_16821),
.B(n_10171),
.Y(n_17276)
);

INVx1_ASAP7_75t_L g17277 ( 
.A(n_17141),
.Y(n_17277)
);

NAND4xp75_ASAP7_75t_L g17278 ( 
.A(n_16926),
.B(n_9393),
.C(n_8247),
.D(n_7980),
.Y(n_17278)
);

INVx1_ASAP7_75t_L g17279 ( 
.A(n_16855),
.Y(n_17279)
);

INVx1_ASAP7_75t_L g17280 ( 
.A(n_16856),
.Y(n_17280)
);

INVx1_ASAP7_75t_L g17281 ( 
.A(n_17057),
.Y(n_17281)
);

INVx1_ASAP7_75t_SL g17282 ( 
.A(n_17059),
.Y(n_17282)
);

INVx1_ASAP7_75t_L g17283 ( 
.A(n_16858),
.Y(n_17283)
);

INVx1_ASAP7_75t_L g17284 ( 
.A(n_16993),
.Y(n_17284)
);

NOR3xp33_ASAP7_75t_L g17285 ( 
.A(n_17050),
.B(n_9748),
.C(n_9724),
.Y(n_17285)
);

NAND2xp5_ASAP7_75t_L g17286 ( 
.A(n_16849),
.B(n_9462),
.Y(n_17286)
);

AND2x2_ASAP7_75t_L g17287 ( 
.A(n_16963),
.B(n_9303),
.Y(n_17287)
);

OR2x2_ASAP7_75t_L g17288 ( 
.A(n_16894),
.B(n_10171),
.Y(n_17288)
);

HB1xp67_ASAP7_75t_L g17289 ( 
.A(n_16948),
.Y(n_17289)
);

INVx1_ASAP7_75t_SL g17290 ( 
.A(n_16975),
.Y(n_17290)
);

HB1xp67_ASAP7_75t_L g17291 ( 
.A(n_16909),
.Y(n_17291)
);

INVx1_ASAP7_75t_SL g17292 ( 
.A(n_16845),
.Y(n_17292)
);

INVx1_ASAP7_75t_L g17293 ( 
.A(n_16873),
.Y(n_17293)
);

INVx1_ASAP7_75t_SL g17294 ( 
.A(n_17159),
.Y(n_17294)
);

AO21x2_ASAP7_75t_L g17295 ( 
.A1(n_17009),
.A2(n_9748),
.B(n_9323),
.Y(n_17295)
);

NOR2x1_ASAP7_75t_L g17296 ( 
.A(n_17025),
.B(n_9462),
.Y(n_17296)
);

AOI22xp33_ASAP7_75t_L g17297 ( 
.A1(n_17109),
.A2(n_7980),
.B1(n_7987),
.B2(n_7951),
.Y(n_17297)
);

AND2x2_ASAP7_75t_L g17298 ( 
.A(n_16841),
.B(n_9323),
.Y(n_17298)
);

INVx1_ASAP7_75t_SL g17299 ( 
.A(n_16844),
.Y(n_17299)
);

NAND2xp5_ASAP7_75t_L g17300 ( 
.A(n_16837),
.B(n_9468),
.Y(n_17300)
);

NAND2xp5_ASAP7_75t_L g17301 ( 
.A(n_16930),
.B(n_9468),
.Y(n_17301)
);

INVx1_ASAP7_75t_L g17302 ( 
.A(n_16827),
.Y(n_17302)
);

INVx2_ASAP7_75t_L g17303 ( 
.A(n_17004),
.Y(n_17303)
);

INVx2_ASAP7_75t_L g17304 ( 
.A(n_17002),
.Y(n_17304)
);

INVx2_ASAP7_75t_L g17305 ( 
.A(n_16999),
.Y(n_17305)
);

OR2x6_ASAP7_75t_L g17306 ( 
.A(n_17037),
.B(n_6905),
.Y(n_17306)
);

INVx2_ASAP7_75t_L g17307 ( 
.A(n_17062),
.Y(n_17307)
);

NOR2x1_ASAP7_75t_L g17308 ( 
.A(n_17055),
.B(n_9474),
.Y(n_17308)
);

BUFx3_ASAP7_75t_L g17309 ( 
.A(n_16928),
.Y(n_17309)
);

HB1xp67_ASAP7_75t_L g17310 ( 
.A(n_17089),
.Y(n_17310)
);

OR2x2_ASAP7_75t_L g17311 ( 
.A(n_16860),
.B(n_10171),
.Y(n_17311)
);

INVx2_ASAP7_75t_L g17312 ( 
.A(n_17155),
.Y(n_17312)
);

INVx3_ASAP7_75t_L g17313 ( 
.A(n_17163),
.Y(n_17313)
);

NOR2x1_ASAP7_75t_L g17314 ( 
.A(n_16906),
.B(n_9474),
.Y(n_17314)
);

NAND3xp33_ASAP7_75t_L g17315 ( 
.A(n_16826),
.B(n_16863),
.C(n_17112),
.Y(n_17315)
);

CKINVDCx16_ASAP7_75t_R g17316 ( 
.A(n_17100),
.Y(n_17316)
);

AND2x4_ASAP7_75t_L g17317 ( 
.A(n_16989),
.B(n_8328),
.Y(n_17317)
);

INVx1_ASAP7_75t_L g17318 ( 
.A(n_16867),
.Y(n_17318)
);

INVx2_ASAP7_75t_L g17319 ( 
.A(n_17140),
.Y(n_17319)
);

CKINVDCx16_ASAP7_75t_R g17320 ( 
.A(n_17034),
.Y(n_17320)
);

INVx3_ASAP7_75t_SL g17321 ( 
.A(n_17046),
.Y(n_17321)
);

AND2x2_ASAP7_75t_L g17322 ( 
.A(n_17013),
.B(n_9323),
.Y(n_17322)
);

INVx1_ASAP7_75t_L g17323 ( 
.A(n_16892),
.Y(n_17323)
);

AND2x2_ASAP7_75t_L g17324 ( 
.A(n_17024),
.B(n_8072),
.Y(n_17324)
);

NOR2x1_ASAP7_75t_L g17325 ( 
.A(n_16920),
.B(n_9480),
.Y(n_17325)
);

OR2x2_ASAP7_75t_L g17326 ( 
.A(n_17099),
.B(n_10173),
.Y(n_17326)
);

CKINVDCx20_ASAP7_75t_R g17327 ( 
.A(n_16834),
.Y(n_17327)
);

AND2x2_ASAP7_75t_L g17328 ( 
.A(n_17075),
.B(n_8072),
.Y(n_17328)
);

OR2x2_ASAP7_75t_L g17329 ( 
.A(n_17199),
.B(n_10173),
.Y(n_17329)
);

AND2x2_ASAP7_75t_L g17330 ( 
.A(n_16897),
.B(n_8072),
.Y(n_17330)
);

AND2x2_ASAP7_75t_L g17331 ( 
.A(n_16901),
.B(n_16904),
.Y(n_17331)
);

OAI221xp5_ASAP7_75t_SL g17332 ( 
.A1(n_17198),
.A2(n_8653),
.B1(n_8519),
.B2(n_8353),
.C(n_9373),
.Y(n_17332)
);

HB1xp67_ASAP7_75t_L g17333 ( 
.A(n_17045),
.Y(n_17333)
);

INVx1_ASAP7_75t_L g17334 ( 
.A(n_16917),
.Y(n_17334)
);

NOR2x1_ASAP7_75t_L g17335 ( 
.A(n_16921),
.B(n_9480),
.Y(n_17335)
);

INVx6_ASAP7_75t_L g17336 ( 
.A(n_16836),
.Y(n_17336)
);

INVx3_ASAP7_75t_L g17337 ( 
.A(n_16872),
.Y(n_17337)
);

INVx4_ASAP7_75t_L g17338 ( 
.A(n_16946),
.Y(n_17338)
);

AND2x2_ASAP7_75t_L g17339 ( 
.A(n_16832),
.B(n_8094),
.Y(n_17339)
);

INVx1_ASAP7_75t_SL g17340 ( 
.A(n_17054),
.Y(n_17340)
);

OR2x6_ASAP7_75t_L g17341 ( 
.A(n_16843),
.B(n_6905),
.Y(n_17341)
);

INVx1_ASAP7_75t_L g17342 ( 
.A(n_16842),
.Y(n_17342)
);

INVx1_ASAP7_75t_L g17343 ( 
.A(n_16889),
.Y(n_17343)
);

OR2x2_ASAP7_75t_L g17344 ( 
.A(n_17084),
.B(n_10173),
.Y(n_17344)
);

INVx1_ASAP7_75t_L g17345 ( 
.A(n_16950),
.Y(n_17345)
);

OR2x2_ASAP7_75t_L g17346 ( 
.A(n_16988),
.B(n_10179),
.Y(n_17346)
);

INVx1_ASAP7_75t_L g17347 ( 
.A(n_16991),
.Y(n_17347)
);

INVx1_ASAP7_75t_L g17348 ( 
.A(n_17117),
.Y(n_17348)
);

AND3x2_ASAP7_75t_L g17349 ( 
.A(n_17118),
.B(n_9488),
.C(n_9483),
.Y(n_17349)
);

INVx1_ASAP7_75t_L g17350 ( 
.A(n_17124),
.Y(n_17350)
);

AND2x2_ASAP7_75t_L g17351 ( 
.A(n_17038),
.B(n_8094),
.Y(n_17351)
);

INVx2_ASAP7_75t_L g17352 ( 
.A(n_16982),
.Y(n_17352)
);

INVx1_ASAP7_75t_SL g17353 ( 
.A(n_17063),
.Y(n_17353)
);

INVx1_ASAP7_75t_L g17354 ( 
.A(n_17000),
.Y(n_17354)
);

NOR2xp33_ASAP7_75t_L g17355 ( 
.A(n_17136),
.B(n_6905),
.Y(n_17355)
);

OR2x2_ASAP7_75t_L g17356 ( 
.A(n_17031),
.B(n_10179),
.Y(n_17356)
);

AND2x2_ASAP7_75t_L g17357 ( 
.A(n_16997),
.B(n_8094),
.Y(n_17357)
);

INVx1_ASAP7_75t_L g17358 ( 
.A(n_17065),
.Y(n_17358)
);

OR2x2_ASAP7_75t_L g17359 ( 
.A(n_17200),
.B(n_10179),
.Y(n_17359)
);

NAND2xp5_ASAP7_75t_L g17360 ( 
.A(n_17168),
.B(n_9483),
.Y(n_17360)
);

CKINVDCx16_ASAP7_75t_R g17361 ( 
.A(n_17018),
.Y(n_17361)
);

INVx1_ASAP7_75t_L g17362 ( 
.A(n_17202),
.Y(n_17362)
);

INVx2_ASAP7_75t_L g17363 ( 
.A(n_16987),
.Y(n_17363)
);

OR2x2_ASAP7_75t_L g17364 ( 
.A(n_16978),
.B(n_10182),
.Y(n_17364)
);

OR2x2_ASAP7_75t_L g17365 ( 
.A(n_16962),
.B(n_10182),
.Y(n_17365)
);

AND2x2_ASAP7_75t_L g17366 ( 
.A(n_17045),
.B(n_8098),
.Y(n_17366)
);

INVx2_ASAP7_75t_L g17367 ( 
.A(n_17144),
.Y(n_17367)
);

OR2x2_ASAP7_75t_L g17368 ( 
.A(n_16966),
.B(n_10182),
.Y(n_17368)
);

INVx3_ASAP7_75t_L g17369 ( 
.A(n_16910),
.Y(n_17369)
);

INVx1_ASAP7_75t_L g17370 ( 
.A(n_17110),
.Y(n_17370)
);

AND2x2_ASAP7_75t_L g17371 ( 
.A(n_16903),
.B(n_8098),
.Y(n_17371)
);

INVx2_ASAP7_75t_L g17372 ( 
.A(n_17151),
.Y(n_17372)
);

INVx3_ASAP7_75t_L g17373 ( 
.A(n_17005),
.Y(n_17373)
);

INVx1_ASAP7_75t_SL g17374 ( 
.A(n_16886),
.Y(n_17374)
);

HB1xp67_ASAP7_75t_L g17375 ( 
.A(n_17069),
.Y(n_17375)
);

INVx1_ASAP7_75t_SL g17376 ( 
.A(n_16902),
.Y(n_17376)
);

CKINVDCx16_ASAP7_75t_R g17377 ( 
.A(n_16885),
.Y(n_17377)
);

OR2x2_ASAP7_75t_L g17378 ( 
.A(n_16968),
.B(n_10187),
.Y(n_17378)
);

INVx1_ASAP7_75t_L g17379 ( 
.A(n_16940),
.Y(n_17379)
);

INVx1_ASAP7_75t_L g17380 ( 
.A(n_16981),
.Y(n_17380)
);

INVx1_ASAP7_75t_L g17381 ( 
.A(n_17161),
.Y(n_17381)
);

AND2x2_ASAP7_75t_L g17382 ( 
.A(n_17023),
.B(n_8098),
.Y(n_17382)
);

INVx1_ASAP7_75t_L g17383 ( 
.A(n_17179),
.Y(n_17383)
);

HB1xp67_ASAP7_75t_L g17384 ( 
.A(n_17148),
.Y(n_17384)
);

AOI22xp33_ASAP7_75t_L g17385 ( 
.A1(n_16864),
.A2(n_7987),
.B1(n_7322),
.B2(n_7350),
.Y(n_17385)
);

NOR2x1_ASAP7_75t_L g17386 ( 
.A(n_16870),
.B(n_9488),
.Y(n_17386)
);

OR2x2_ASAP7_75t_L g17387 ( 
.A(n_16973),
.B(n_16977),
.Y(n_17387)
);

INVx1_ASAP7_75t_SL g17388 ( 
.A(n_17191),
.Y(n_17388)
);

NOR2xp33_ASAP7_75t_L g17389 ( 
.A(n_16941),
.B(n_6905),
.Y(n_17389)
);

AND2x4_ASAP7_75t_L g17390 ( 
.A(n_16979),
.B(n_16970),
.Y(n_17390)
);

INVxp67_ASAP7_75t_L g17391 ( 
.A(n_17061),
.Y(n_17391)
);

NOR2xp67_ASAP7_75t_L g17392 ( 
.A(n_16908),
.B(n_9506),
.Y(n_17392)
);

AND2x2_ASAP7_75t_L g17393 ( 
.A(n_16916),
.B(n_8118),
.Y(n_17393)
);

INVx2_ASAP7_75t_L g17394 ( 
.A(n_16983),
.Y(n_17394)
);

BUFx2_ASAP7_75t_L g17395 ( 
.A(n_17149),
.Y(n_17395)
);

AO21x1_ASAP7_75t_L g17396 ( 
.A1(n_17190),
.A2(n_9748),
.B(n_9533),
.Y(n_17396)
);

INVx3_ASAP7_75t_L g17397 ( 
.A(n_17006),
.Y(n_17397)
);

AND2x2_ASAP7_75t_L g17398 ( 
.A(n_17033),
.B(n_17014),
.Y(n_17398)
);

INVx1_ASAP7_75t_L g17399 ( 
.A(n_17180),
.Y(n_17399)
);

INVx1_ASAP7_75t_L g17400 ( 
.A(n_17176),
.Y(n_17400)
);

INVx1_ASAP7_75t_L g17401 ( 
.A(n_17137),
.Y(n_17401)
);

NAND2xp5_ASAP7_75t_SL g17402 ( 
.A(n_17078),
.B(n_10187),
.Y(n_17402)
);

NAND2xp5_ASAP7_75t_L g17403 ( 
.A(n_16848),
.B(n_9506),
.Y(n_17403)
);

OAI21xp5_ASAP7_75t_SL g17404 ( 
.A1(n_17111),
.A2(n_7881),
.B(n_7825),
.Y(n_17404)
);

OR2x2_ASAP7_75t_L g17405 ( 
.A(n_17184),
.B(n_10187),
.Y(n_17405)
);

AND2x2_ASAP7_75t_L g17406 ( 
.A(n_17106),
.B(n_8118),
.Y(n_17406)
);

NOR2xp33_ASAP7_75t_L g17407 ( 
.A(n_16838),
.B(n_16862),
.Y(n_17407)
);

INVx1_ASAP7_75t_L g17408 ( 
.A(n_16896),
.Y(n_17408)
);

INVx2_ASAP7_75t_L g17409 ( 
.A(n_16985),
.Y(n_17409)
);

OR2x2_ASAP7_75t_L g17410 ( 
.A(n_17154),
.B(n_17056),
.Y(n_17410)
);

HB1xp67_ASAP7_75t_L g17411 ( 
.A(n_16915),
.Y(n_17411)
);

AO21x2_ASAP7_75t_L g17412 ( 
.A1(n_17036),
.A2(n_9253),
.B(n_8656),
.Y(n_17412)
);

INVxp67_ASAP7_75t_SL g17413 ( 
.A(n_16967),
.Y(n_17413)
);

AND2x2_ASAP7_75t_L g17414 ( 
.A(n_16969),
.B(n_8118),
.Y(n_17414)
);

INVx1_ASAP7_75t_L g17415 ( 
.A(n_17175),
.Y(n_17415)
);

OR2x2_ASAP7_75t_L g17416 ( 
.A(n_16851),
.B(n_10198),
.Y(n_17416)
);

AND2x2_ASAP7_75t_L g17417 ( 
.A(n_16984),
.B(n_8138),
.Y(n_17417)
);

INVx1_ASAP7_75t_L g17418 ( 
.A(n_17169),
.Y(n_17418)
);

AND2x2_ASAP7_75t_L g17419 ( 
.A(n_17107),
.B(n_8138),
.Y(n_17419)
);

OR2x2_ASAP7_75t_L g17420 ( 
.A(n_17178),
.B(n_16893),
.Y(n_17420)
);

INVxp67_ASAP7_75t_L g17421 ( 
.A(n_17127),
.Y(n_17421)
);

INVx1_ASAP7_75t_L g17422 ( 
.A(n_17092),
.Y(n_17422)
);

INVx1_ASAP7_75t_L g17423 ( 
.A(n_17095),
.Y(n_17423)
);

HB1xp67_ASAP7_75t_L g17424 ( 
.A(n_16960),
.Y(n_17424)
);

AND2x2_ASAP7_75t_L g17425 ( 
.A(n_17076),
.B(n_8138),
.Y(n_17425)
);

INVx1_ASAP7_75t_SL g17426 ( 
.A(n_17001),
.Y(n_17426)
);

INVx4_ASAP7_75t_L g17427 ( 
.A(n_17042),
.Y(n_17427)
);

INVx1_ASAP7_75t_SL g17428 ( 
.A(n_17167),
.Y(n_17428)
);

INVx1_ASAP7_75t_L g17429 ( 
.A(n_16899),
.Y(n_17429)
);

NAND2xp5_ASAP7_75t_L g17430 ( 
.A(n_16922),
.B(n_9521),
.Y(n_17430)
);

INVx1_ASAP7_75t_SL g17431 ( 
.A(n_17164),
.Y(n_17431)
);

OAI221xp5_ASAP7_75t_L g17432 ( 
.A1(n_17174),
.A2(n_8217),
.B1(n_8396),
.B2(n_8140),
.C(n_8043),
.Y(n_17432)
);

BUFx2_ASAP7_75t_L g17433 ( 
.A(n_17183),
.Y(n_17433)
);

OR2x2_ASAP7_75t_L g17434 ( 
.A(n_17182),
.B(n_10198),
.Y(n_17434)
);

NAND2x1p5_ASAP7_75t_L g17435 ( 
.A(n_17041),
.B(n_6906),
.Y(n_17435)
);

AND2x2_ASAP7_75t_L g17436 ( 
.A(n_17060),
.B(n_8152),
.Y(n_17436)
);

INVx1_ASAP7_75t_L g17437 ( 
.A(n_17073),
.Y(n_17437)
);

INVx1_ASAP7_75t_SL g17438 ( 
.A(n_17081),
.Y(n_17438)
);

INVx1_ASAP7_75t_L g17439 ( 
.A(n_16925),
.Y(n_17439)
);

AND2x2_ASAP7_75t_L g17440 ( 
.A(n_16956),
.B(n_8152),
.Y(n_17440)
);

NAND2xp5_ASAP7_75t_L g17441 ( 
.A(n_17007),
.B(n_9521),
.Y(n_17441)
);

OR2x2_ASAP7_75t_L g17442 ( 
.A(n_17201),
.B(n_10198),
.Y(n_17442)
);

OR2x2_ASAP7_75t_L g17443 ( 
.A(n_17114),
.B(n_10207),
.Y(n_17443)
);

BUFx3_ASAP7_75t_L g17444 ( 
.A(n_17083),
.Y(n_17444)
);

INVx2_ASAP7_75t_L g17445 ( 
.A(n_16929),
.Y(n_17445)
);

OR2x2_ASAP7_75t_L g17446 ( 
.A(n_17097),
.B(n_10207),
.Y(n_17446)
);

INVx1_ASAP7_75t_SL g17447 ( 
.A(n_17119),
.Y(n_17447)
);

AND2x4_ASAP7_75t_L g17448 ( 
.A(n_17026),
.B(n_9530),
.Y(n_17448)
);

INVx2_ASAP7_75t_L g17449 ( 
.A(n_17043),
.Y(n_17449)
);

OAI21x1_ASAP7_75t_L g17450 ( 
.A1(n_16890),
.A2(n_9445),
.B(n_9435),
.Y(n_17450)
);

NOR2xp33_ASAP7_75t_L g17451 ( 
.A(n_16961),
.B(n_6906),
.Y(n_17451)
);

AND2x4_ASAP7_75t_L g17452 ( 
.A(n_17086),
.B(n_9530),
.Y(n_17452)
);

INVxp67_ASAP7_75t_L g17453 ( 
.A(n_17067),
.Y(n_17453)
);

BUFx3_ASAP7_75t_L g17454 ( 
.A(n_17088),
.Y(n_17454)
);

AND2x2_ASAP7_75t_L g17455 ( 
.A(n_16995),
.B(n_8152),
.Y(n_17455)
);

HB1xp67_ASAP7_75t_L g17456 ( 
.A(n_17181),
.Y(n_17456)
);

AND2x2_ASAP7_75t_L g17457 ( 
.A(n_17090),
.B(n_8162),
.Y(n_17457)
);

BUFx3_ASAP7_75t_L g17458 ( 
.A(n_17093),
.Y(n_17458)
);

AND2x2_ASAP7_75t_L g17459 ( 
.A(n_17102),
.B(n_8162),
.Y(n_17459)
);

INVx1_ASAP7_75t_L g17460 ( 
.A(n_16934),
.Y(n_17460)
);

INVx1_ASAP7_75t_SL g17461 ( 
.A(n_17010),
.Y(n_17461)
);

HB1xp67_ASAP7_75t_L g17462 ( 
.A(n_16927),
.Y(n_17462)
);

INVx1_ASAP7_75t_L g17463 ( 
.A(n_16939),
.Y(n_17463)
);

AND2x2_ASAP7_75t_L g17464 ( 
.A(n_17012),
.B(n_8162),
.Y(n_17464)
);

INVxp67_ASAP7_75t_L g17465 ( 
.A(n_17135),
.Y(n_17465)
);

NAND2xp5_ASAP7_75t_L g17466 ( 
.A(n_17157),
.B(n_17029),
.Y(n_17466)
);

AOI22xp33_ASAP7_75t_L g17467 ( 
.A1(n_16955),
.A2(n_7987),
.B1(n_7322),
.B2(n_7350),
.Y(n_17467)
);

INVx1_ASAP7_75t_SL g17468 ( 
.A(n_17021),
.Y(n_17468)
);

INVx1_ASAP7_75t_L g17469 ( 
.A(n_16942),
.Y(n_17469)
);

INVx1_ASAP7_75t_L g17470 ( 
.A(n_16992),
.Y(n_17470)
);

INVx1_ASAP7_75t_L g17471 ( 
.A(n_16972),
.Y(n_17471)
);

INVx1_ASAP7_75t_L g17472 ( 
.A(n_16957),
.Y(n_17472)
);

OR2x2_ASAP7_75t_L g17473 ( 
.A(n_17160),
.B(n_17153),
.Y(n_17473)
);

AOI22xp33_ASAP7_75t_L g17474 ( 
.A1(n_17195),
.A2(n_7987),
.B1(n_7322),
.B2(n_7350),
.Y(n_17474)
);

OR2x2_ASAP7_75t_L g17475 ( 
.A(n_17150),
.B(n_10207),
.Y(n_17475)
);

AOI22xp33_ASAP7_75t_L g17476 ( 
.A1(n_17139),
.A2(n_7987),
.B1(n_7322),
.B2(n_7350),
.Y(n_17476)
);

INVx1_ASAP7_75t_SL g17477 ( 
.A(n_16964),
.Y(n_17477)
);

AOI22xp33_ASAP7_75t_L g17478 ( 
.A1(n_17123),
.A2(n_7987),
.B1(n_7322),
.B2(n_7350),
.Y(n_17478)
);

NAND2xp5_ASAP7_75t_L g17479 ( 
.A(n_17077),
.B(n_9535),
.Y(n_17479)
);

INVx1_ASAP7_75t_SL g17480 ( 
.A(n_17035),
.Y(n_17480)
);

AND2x2_ASAP7_75t_L g17481 ( 
.A(n_17105),
.B(n_8280),
.Y(n_17481)
);

INVx1_ASAP7_75t_SL g17482 ( 
.A(n_17039),
.Y(n_17482)
);

BUFx3_ASAP7_75t_L g17483 ( 
.A(n_17051),
.Y(n_17483)
);

INVx2_ASAP7_75t_L g17484 ( 
.A(n_16996),
.Y(n_17484)
);

NAND2xp5_ASAP7_75t_L g17485 ( 
.A(n_17058),
.B(n_9535),
.Y(n_17485)
);

OR2x2_ASAP7_75t_L g17486 ( 
.A(n_17115),
.B(n_10208),
.Y(n_17486)
);

AND2x2_ASAP7_75t_L g17487 ( 
.A(n_17028),
.B(n_8280),
.Y(n_17487)
);

OR2x2_ASAP7_75t_L g17488 ( 
.A(n_16980),
.B(n_10208),
.Y(n_17488)
);

NOR2xp33_ASAP7_75t_L g17489 ( 
.A(n_17079),
.B(n_6906),
.Y(n_17489)
);

INVx1_ASAP7_75t_L g17490 ( 
.A(n_17104),
.Y(n_17490)
);

AND2x2_ASAP7_75t_L g17491 ( 
.A(n_17103),
.B(n_17101),
.Y(n_17491)
);

OR2x2_ASAP7_75t_L g17492 ( 
.A(n_16986),
.B(n_10208),
.Y(n_17492)
);

INVx2_ASAP7_75t_SL g17493 ( 
.A(n_16936),
.Y(n_17493)
);

AOI21xp5_ASAP7_75t_SL g17494 ( 
.A1(n_17003),
.A2(n_9393),
.B(n_6906),
.Y(n_17494)
);

BUFx3_ASAP7_75t_L g17495 ( 
.A(n_17071),
.Y(n_17495)
);

INVx1_ASAP7_75t_L g17496 ( 
.A(n_17134),
.Y(n_17496)
);

OR2x2_ASAP7_75t_L g17497 ( 
.A(n_17165),
.B(n_10212),
.Y(n_17497)
);

INVx1_ASAP7_75t_L g17498 ( 
.A(n_17138),
.Y(n_17498)
);

CKINVDCx14_ASAP7_75t_R g17499 ( 
.A(n_17120),
.Y(n_17499)
);

AND2x2_ASAP7_75t_L g17500 ( 
.A(n_17072),
.B(n_9253),
.Y(n_17500)
);

INVx1_ASAP7_75t_L g17501 ( 
.A(n_17066),
.Y(n_17501)
);

INVx3_ASAP7_75t_L g17502 ( 
.A(n_17068),
.Y(n_17502)
);

INVx2_ASAP7_75t_L g17503 ( 
.A(n_16877),
.Y(n_17503)
);

INVx1_ASAP7_75t_L g17504 ( 
.A(n_17052),
.Y(n_17504)
);

AND2x4_ASAP7_75t_L g17505 ( 
.A(n_17091),
.B(n_9539),
.Y(n_17505)
);

NAND2xp5_ASAP7_75t_L g17506 ( 
.A(n_17171),
.B(n_9539),
.Y(n_17506)
);

AND2x2_ASAP7_75t_L g17507 ( 
.A(n_17085),
.B(n_17129),
.Y(n_17507)
);

NAND2xp5_ASAP7_75t_L g17508 ( 
.A(n_16951),
.B(n_16895),
.Y(n_17508)
);

AND2x2_ASAP7_75t_L g17509 ( 
.A(n_17143),
.B(n_9253),
.Y(n_17509)
);

NAND2xp5_ASAP7_75t_L g17510 ( 
.A(n_16974),
.B(n_16976),
.Y(n_17510)
);

INVx1_ASAP7_75t_L g17511 ( 
.A(n_17197),
.Y(n_17511)
);

INVx2_ASAP7_75t_L g17512 ( 
.A(n_16965),
.Y(n_17512)
);

INVx2_ASAP7_75t_L g17513 ( 
.A(n_16971),
.Y(n_17513)
);

OR2x2_ASAP7_75t_L g17514 ( 
.A(n_17132),
.B(n_10212),
.Y(n_17514)
);

INVx2_ASAP7_75t_L g17515 ( 
.A(n_17152),
.Y(n_17515)
);

NAND2xp5_ASAP7_75t_L g17516 ( 
.A(n_16912),
.B(n_9540),
.Y(n_17516)
);

INVx1_ASAP7_75t_SL g17517 ( 
.A(n_16958),
.Y(n_17517)
);

AOI22xp33_ASAP7_75t_L g17518 ( 
.A1(n_17170),
.A2(n_17188),
.B1(n_17162),
.B2(n_17172),
.Y(n_17518)
);

AND2x2_ASAP7_75t_L g17519 ( 
.A(n_17147),
.B(n_8247),
.Y(n_17519)
);

AND2x2_ASAP7_75t_L g17520 ( 
.A(n_16945),
.B(n_10212),
.Y(n_17520)
);

NOR2xp33_ASAP7_75t_L g17521 ( 
.A(n_17016),
.B(n_9540),
.Y(n_17521)
);

NAND2xp5_ASAP7_75t_L g17522 ( 
.A(n_17185),
.B(n_9546),
.Y(n_17522)
);

OR2x2_ASAP7_75t_L g17523 ( 
.A(n_17196),
.B(n_10227),
.Y(n_17523)
);

OR2x2_ASAP7_75t_L g17524 ( 
.A(n_17177),
.B(n_10227),
.Y(n_17524)
);

INVx1_ASAP7_75t_SL g17525 ( 
.A(n_16933),
.Y(n_17525)
);

CKINVDCx16_ASAP7_75t_R g17526 ( 
.A(n_17082),
.Y(n_17526)
);

NOR2xp33_ASAP7_75t_L g17527 ( 
.A(n_17130),
.B(n_9546),
.Y(n_17527)
);

AND2x2_ASAP7_75t_L g17528 ( 
.A(n_17321),
.B(n_16887),
.Y(n_17528)
);

OAI21xp5_ASAP7_75t_L g17529 ( 
.A1(n_17210),
.A2(n_17192),
.B(n_17187),
.Y(n_17529)
);

INVx2_ASAP7_75t_L g17530 ( 
.A(n_17240),
.Y(n_17530)
);

AOI21xp33_ASAP7_75t_SL g17531 ( 
.A1(n_17320),
.A2(n_16919),
.B(n_17113),
.Y(n_17531)
);

AOI211xp5_ASAP7_75t_L g17532 ( 
.A1(n_17332),
.A2(n_17011),
.B(n_17053),
.C(n_17044),
.Y(n_17532)
);

INVx1_ASAP7_75t_L g17533 ( 
.A(n_17411),
.Y(n_17533)
);

AOI21xp33_ASAP7_75t_SL g17534 ( 
.A1(n_17377),
.A2(n_17116),
.B(n_16954),
.Y(n_17534)
);

INVx1_ASAP7_75t_L g17535 ( 
.A(n_17424),
.Y(n_17535)
);

AOI22x1_ASAP7_75t_L g17536 ( 
.A1(n_17395),
.A2(n_16944),
.B1(n_17108),
.B2(n_17173),
.Y(n_17536)
);

BUFx2_ASAP7_75t_L g17537 ( 
.A(n_17310),
.Y(n_17537)
);

AOI211xp5_ASAP7_75t_L g17538 ( 
.A1(n_17216),
.A2(n_17146),
.B(n_17156),
.C(n_17186),
.Y(n_17538)
);

AND2x2_ASAP7_75t_L g17539 ( 
.A(n_17316),
.B(n_17040),
.Y(n_17539)
);

AOI21xp5_ASAP7_75t_L g17540 ( 
.A1(n_17236),
.A2(n_16914),
.B(n_17008),
.Y(n_17540)
);

NAND2xp5_ASAP7_75t_L g17541 ( 
.A(n_17401),
.B(n_16900),
.Y(n_17541)
);

INVxp67_ASAP7_75t_SL g17542 ( 
.A(n_17291),
.Y(n_17542)
);

NAND4xp25_ASAP7_75t_SL g17543 ( 
.A(n_17244),
.B(n_16913),
.C(n_16935),
.D(n_17125),
.Y(n_17543)
);

AND2x2_ASAP7_75t_L g17544 ( 
.A(n_17419),
.B(n_17096),
.Y(n_17544)
);

NAND2xp5_ASAP7_75t_L g17545 ( 
.A(n_17215),
.B(n_17070),
.Y(n_17545)
);

AND2x2_ASAP7_75t_L g17546 ( 
.A(n_17357),
.B(n_17027),
.Y(n_17546)
);

HB1xp67_ASAP7_75t_L g17547 ( 
.A(n_17306),
.Y(n_17547)
);

OAI22xp33_ASAP7_75t_SL g17548 ( 
.A1(n_17336),
.A2(n_17122),
.B1(n_17126),
.B2(n_17022),
.Y(n_17548)
);

NOR2xp33_ASAP7_75t_SL g17549 ( 
.A(n_17217),
.B(n_17047),
.Y(n_17549)
);

OR2x2_ASAP7_75t_L g17550 ( 
.A(n_17361),
.B(n_17030),
.Y(n_17550)
);

INVx1_ASAP7_75t_L g17551 ( 
.A(n_17267),
.Y(n_17551)
);

OAI22xp5_ASAP7_75t_L g17552 ( 
.A1(n_17327),
.A2(n_16924),
.B1(n_17020),
.B2(n_17048),
.Y(n_17552)
);

INVx1_ASAP7_75t_L g17553 ( 
.A(n_17228),
.Y(n_17553)
);

NAND2xp5_ASAP7_75t_L g17554 ( 
.A(n_17282),
.B(n_17064),
.Y(n_17554)
);

AOI31xp33_ASAP7_75t_L g17555 ( 
.A1(n_17213),
.A2(n_17019),
.A3(n_17015),
.B(n_17094),
.Y(n_17555)
);

INVx1_ASAP7_75t_SL g17556 ( 
.A(n_17336),
.Y(n_17556)
);

NAND2xp5_ASAP7_75t_L g17557 ( 
.A(n_17388),
.B(n_17098),
.Y(n_17557)
);

AND2x2_ASAP7_75t_L g17558 ( 
.A(n_17330),
.B(n_17017),
.Y(n_17558)
);

OAI32xp33_ASAP7_75t_L g17559 ( 
.A1(n_17407),
.A2(n_17166),
.A3(n_16898),
.B1(n_17049),
.B2(n_17145),
.Y(n_17559)
);

OR2x2_ASAP7_75t_L g17560 ( 
.A(n_17294),
.B(n_16888),
.Y(n_17560)
);

AND2x2_ASAP7_75t_L g17561 ( 
.A(n_17233),
.B(n_10227),
.Y(n_17561)
);

INVx2_ASAP7_75t_L g17562 ( 
.A(n_17208),
.Y(n_17562)
);

INVx1_ASAP7_75t_L g17563 ( 
.A(n_17433),
.Y(n_17563)
);

NAND3xp33_ASAP7_75t_L g17564 ( 
.A(n_17315),
.B(n_16953),
.C(n_9393),
.Y(n_17564)
);

AND2x4_ASAP7_75t_SL g17565 ( 
.A(n_17222),
.B(n_6940),
.Y(n_17565)
);

AOI21xp5_ASAP7_75t_L g17566 ( 
.A1(n_17413),
.A2(n_9533),
.B(n_9531),
.Y(n_17566)
);

AOI22xp5_ASAP7_75t_L g17567 ( 
.A1(n_17235),
.A2(n_9534),
.B1(n_9553),
.B2(n_9531),
.Y(n_17567)
);

INVx1_ASAP7_75t_L g17568 ( 
.A(n_17456),
.Y(n_17568)
);

OAI322xp33_ASAP7_75t_L g17569 ( 
.A1(n_17499),
.A2(n_9376),
.A3(n_9375),
.B1(n_9392),
.B2(n_9395),
.C1(n_9391),
.C2(n_9373),
.Y(n_17569)
);

NAND2xp5_ASAP7_75t_L g17570 ( 
.A(n_17302),
.B(n_9547),
.Y(n_17570)
);

INVx1_ASAP7_75t_L g17571 ( 
.A(n_17375),
.Y(n_17571)
);

INVx1_ASAP7_75t_L g17572 ( 
.A(n_17229),
.Y(n_17572)
);

NAND2xp5_ASAP7_75t_L g17573 ( 
.A(n_17438),
.B(n_9547),
.Y(n_17573)
);

INVx2_ASAP7_75t_L g17574 ( 
.A(n_17328),
.Y(n_17574)
);

NAND2xp5_ASAP7_75t_L g17575 ( 
.A(n_17266),
.B(n_9550),
.Y(n_17575)
);

OAI321xp33_ASAP7_75t_L g17576 ( 
.A1(n_17383),
.A2(n_7942),
.A3(n_7825),
.B1(n_8030),
.B2(n_7949),
.C(n_7881),
.Y(n_17576)
);

NOR2xp33_ASAP7_75t_L g17577 ( 
.A(n_17338),
.B(n_9550),
.Y(n_17577)
);

OAI21xp5_ASAP7_75t_SL g17578 ( 
.A1(n_17428),
.A2(n_8217),
.B(n_8140),
.Y(n_17578)
);

NOR2xp33_ASAP7_75t_L g17579 ( 
.A(n_17279),
.B(n_9555),
.Y(n_17579)
);

AOI222xp33_ASAP7_75t_L g17580 ( 
.A1(n_17386),
.A2(n_9575),
.B1(n_9553),
.B2(n_9584),
.C1(n_9559),
.C2(n_9534),
.Y(n_17580)
);

OR2x2_ASAP7_75t_L g17581 ( 
.A(n_17303),
.B(n_17304),
.Y(n_17581)
);

INVx1_ASAP7_75t_SL g17582 ( 
.A(n_17252),
.Y(n_17582)
);

INVx1_ASAP7_75t_L g17583 ( 
.A(n_17333),
.Y(n_17583)
);

NOR2x1_ASAP7_75t_L g17584 ( 
.A(n_17224),
.B(n_9555),
.Y(n_17584)
);

NAND2xp5_ASAP7_75t_L g17585 ( 
.A(n_17280),
.B(n_9568),
.Y(n_17585)
);

NAND3xp33_ASAP7_75t_L g17586 ( 
.A(n_17399),
.B(n_9393),
.C(n_9534),
.Y(n_17586)
);

INVx1_ASAP7_75t_SL g17587 ( 
.A(n_17265),
.Y(n_17587)
);

OAI21xp5_ASAP7_75t_SL g17588 ( 
.A1(n_17431),
.A2(n_8217),
.B(n_8140),
.Y(n_17588)
);

INVx1_ASAP7_75t_L g17589 ( 
.A(n_17319),
.Y(n_17589)
);

NOR2xp33_ASAP7_75t_L g17590 ( 
.A(n_17340),
.B(n_9568),
.Y(n_17590)
);

NOR3xp33_ASAP7_75t_SL g17591 ( 
.A(n_17526),
.B(n_6913),
.C(n_6911),
.Y(n_17591)
);

AOI22xp33_ASAP7_75t_L g17592 ( 
.A1(n_17400),
.A2(n_9559),
.B1(n_9575),
.B2(n_9553),
.Y(n_17592)
);

BUFx2_ASAP7_75t_L g17593 ( 
.A(n_17306),
.Y(n_17593)
);

OAI21xp33_ASAP7_75t_SL g17594 ( 
.A1(n_17392),
.A2(n_9445),
.B(n_9435),
.Y(n_17594)
);

AOI21xp33_ASAP7_75t_SL g17595 ( 
.A1(n_17238),
.A2(n_9445),
.B(n_9435),
.Y(n_17595)
);

AOI21xp5_ASAP7_75t_L g17596 ( 
.A1(n_17292),
.A2(n_17299),
.B(n_17259),
.Y(n_17596)
);

INVx1_ASAP7_75t_L g17597 ( 
.A(n_17270),
.Y(n_17597)
);

AND2x2_ASAP7_75t_L g17598 ( 
.A(n_17491),
.B(n_10249),
.Y(n_17598)
);

A2O1A1Ixp33_ASAP7_75t_L g17599 ( 
.A1(n_17272),
.A2(n_9528),
.B(n_9577),
.C(n_9461),
.Y(n_17599)
);

HB1xp67_ASAP7_75t_L g17600 ( 
.A(n_17289),
.Y(n_17600)
);

AOI21xp33_ASAP7_75t_L g17601 ( 
.A1(n_17410),
.A2(n_9575),
.B(n_9559),
.Y(n_17601)
);

INVx1_ASAP7_75t_L g17602 ( 
.A(n_17254),
.Y(n_17602)
);

INVx1_ASAP7_75t_L g17603 ( 
.A(n_17384),
.Y(n_17603)
);

NAND2xp5_ASAP7_75t_L g17604 ( 
.A(n_17373),
.B(n_9573),
.Y(n_17604)
);

OAI32xp33_ASAP7_75t_L g17605 ( 
.A1(n_17447),
.A2(n_9589),
.A3(n_9591),
.B1(n_9587),
.B2(n_9584),
.Y(n_17605)
);

INVx1_ASAP7_75t_L g17606 ( 
.A(n_17284),
.Y(n_17606)
);

INVx1_ASAP7_75t_L g17607 ( 
.A(n_17207),
.Y(n_17607)
);

INVx1_ASAP7_75t_L g17608 ( 
.A(n_17331),
.Y(n_17608)
);

NOR3xp33_ASAP7_75t_L g17609 ( 
.A(n_17313),
.B(n_5652),
.C(n_5627),
.Y(n_17609)
);

AND2x2_ASAP7_75t_L g17610 ( 
.A(n_17255),
.B(n_10249),
.Y(n_17610)
);

INVx1_ASAP7_75t_L g17611 ( 
.A(n_17277),
.Y(n_17611)
);

INVx1_ASAP7_75t_L g17612 ( 
.A(n_17271),
.Y(n_17612)
);

OAI21xp5_ASAP7_75t_L g17613 ( 
.A1(n_17421),
.A2(n_17241),
.B(n_17465),
.Y(n_17613)
);

INVx1_ASAP7_75t_L g17614 ( 
.A(n_17274),
.Y(n_17614)
);

AOI21xp33_ASAP7_75t_L g17615 ( 
.A1(n_17353),
.A2(n_9587),
.B(n_9584),
.Y(n_17615)
);

INVx1_ASAP7_75t_L g17616 ( 
.A(n_17283),
.Y(n_17616)
);

AOI21xp33_ASAP7_75t_L g17617 ( 
.A1(n_17355),
.A2(n_9589),
.B(n_9587),
.Y(n_17617)
);

AOI21xp33_ASAP7_75t_L g17618 ( 
.A1(n_17511),
.A2(n_17358),
.B(n_17370),
.Y(n_17618)
);

AOI221xp5_ASAP7_75t_L g17619 ( 
.A1(n_17223),
.A2(n_9600),
.B1(n_9620),
.B2(n_9591),
.C(n_9589),
.Y(n_17619)
);

O2A1O1Ixp33_ASAP7_75t_SL g17620 ( 
.A1(n_17212),
.A2(n_17379),
.B(n_17403),
.C(n_17211),
.Y(n_17620)
);

INVx1_ASAP7_75t_L g17621 ( 
.A(n_17337),
.Y(n_17621)
);

NOR2xp67_ASAP7_75t_SL g17622 ( 
.A(n_17309),
.B(n_7077),
.Y(n_17622)
);

OAI21xp5_ASAP7_75t_L g17623 ( 
.A1(n_17391),
.A2(n_10222),
.B(n_10192),
.Y(n_17623)
);

AND2x2_ASAP7_75t_L g17624 ( 
.A(n_17261),
.B(n_10249),
.Y(n_17624)
);

OAI21xp33_ASAP7_75t_SL g17625 ( 
.A1(n_17474),
.A2(n_9528),
.B(n_9461),
.Y(n_17625)
);

AOI22xp33_ASAP7_75t_L g17626 ( 
.A1(n_17418),
.A2(n_9600),
.B1(n_9620),
.B2(n_9591),
.Y(n_17626)
);

INVx1_ASAP7_75t_L g17627 ( 
.A(n_17263),
.Y(n_17627)
);

NOR2xp33_ASAP7_75t_L g17628 ( 
.A(n_17397),
.B(n_9573),
.Y(n_17628)
);

AND2x2_ASAP7_75t_L g17629 ( 
.A(n_17414),
.B(n_10261),
.Y(n_17629)
);

NAND2xp5_ASAP7_75t_L g17630 ( 
.A(n_17324),
.B(n_9574),
.Y(n_17630)
);

OAI31xp33_ASAP7_75t_L g17631 ( 
.A1(n_17290),
.A2(n_8217),
.A3(n_8396),
.B(n_8140),
.Y(n_17631)
);

INVx1_ASAP7_75t_L g17632 ( 
.A(n_17257),
.Y(n_17632)
);

AND4x1_ASAP7_75t_L g17633 ( 
.A(n_17381),
.B(n_7380),
.C(n_7358),
.D(n_7419),
.Y(n_17633)
);

AOI21xp33_ASAP7_75t_SL g17634 ( 
.A1(n_17435),
.A2(n_9528),
.B(n_9461),
.Y(n_17634)
);

AOI222xp33_ASAP7_75t_L g17635 ( 
.A1(n_17415),
.A2(n_9628),
.B1(n_9620),
.B2(n_9641),
.C1(n_9622),
.C2(n_9600),
.Y(n_17635)
);

INVxp67_ASAP7_75t_L g17636 ( 
.A(n_17256),
.Y(n_17636)
);

OR2x2_ASAP7_75t_L g17637 ( 
.A(n_17307),
.B(n_10261),
.Y(n_17637)
);

INVx2_ASAP7_75t_L g17638 ( 
.A(n_17349),
.Y(n_17638)
);

NAND2xp5_ASAP7_75t_L g17639 ( 
.A(n_17369),
.B(n_9574),
.Y(n_17639)
);

AOI22xp33_ASAP7_75t_SL g17640 ( 
.A1(n_17250),
.A2(n_7322),
.B1(n_7350),
.B2(n_7320),
.Y(n_17640)
);

INVx2_ASAP7_75t_L g17641 ( 
.A(n_17366),
.Y(n_17641)
);

NAND2xp5_ASAP7_75t_L g17642 ( 
.A(n_17339),
.B(n_9579),
.Y(n_17642)
);

NOR2xp33_ASAP7_75t_L g17643 ( 
.A(n_17230),
.B(n_9579),
.Y(n_17643)
);

INVx1_ASAP7_75t_L g17644 ( 
.A(n_17245),
.Y(n_17644)
);

NAND2xp5_ASAP7_75t_L g17645 ( 
.A(n_17502),
.B(n_9580),
.Y(n_17645)
);

INVx1_ASAP7_75t_SL g17646 ( 
.A(n_17387),
.Y(n_17646)
);

INVx1_ASAP7_75t_L g17647 ( 
.A(n_17251),
.Y(n_17647)
);

INVx1_ASAP7_75t_L g17648 ( 
.A(n_17253),
.Y(n_17648)
);

INVx1_ASAP7_75t_L g17649 ( 
.A(n_17246),
.Y(n_17649)
);

INVxp67_ASAP7_75t_L g17650 ( 
.A(n_17341),
.Y(n_17650)
);

AOI21xp5_ASAP7_75t_L g17651 ( 
.A1(n_17510),
.A2(n_9628),
.B(n_9622),
.Y(n_17651)
);

AND2x2_ASAP7_75t_L g17652 ( 
.A(n_17449),
.B(n_10261),
.Y(n_17652)
);

INVxp67_ASAP7_75t_SL g17653 ( 
.A(n_17296),
.Y(n_17653)
);

AOI21xp33_ASAP7_75t_SL g17654 ( 
.A1(n_17380),
.A2(n_9590),
.B(n_9577),
.Y(n_17654)
);

NOR2xp33_ASAP7_75t_R g17655 ( 
.A(n_17422),
.B(n_6729),
.Y(n_17655)
);

OAI221xp5_ASAP7_75t_L g17656 ( 
.A1(n_17518),
.A2(n_8549),
.B1(n_8608),
.B2(n_8429),
.C(n_8396),
.Y(n_17656)
);

OR2x2_ASAP7_75t_L g17657 ( 
.A(n_17305),
.B(n_10268),
.Y(n_17657)
);

INVx2_ASAP7_75t_L g17658 ( 
.A(n_17406),
.Y(n_17658)
);

OR2x2_ASAP7_75t_L g17659 ( 
.A(n_17312),
.B(n_10268),
.Y(n_17659)
);

INVx1_ASAP7_75t_L g17660 ( 
.A(n_17248),
.Y(n_17660)
);

INVx1_ASAP7_75t_L g17661 ( 
.A(n_17507),
.Y(n_17661)
);

INVxp33_ASAP7_75t_L g17662 ( 
.A(n_17226),
.Y(n_17662)
);

AND2x2_ASAP7_75t_L g17663 ( 
.A(n_17425),
.B(n_10268),
.Y(n_17663)
);

O2A1O1Ixp33_ASAP7_75t_L g17664 ( 
.A1(n_17466),
.A2(n_9628),
.B(n_9641),
.C(n_9622),
.Y(n_17664)
);

OAI22xp5_ASAP7_75t_L g17665 ( 
.A1(n_17326),
.A2(n_9373),
.B1(n_9376),
.B2(n_9375),
.Y(n_17665)
);

INVxp67_ASAP7_75t_SL g17666 ( 
.A(n_17508),
.Y(n_17666)
);

OR2x2_ASAP7_75t_L g17667 ( 
.A(n_17477),
.B(n_10272),
.Y(n_17667)
);

NAND2xp5_ASAP7_75t_L g17668 ( 
.A(n_17348),
.B(n_9580),
.Y(n_17668)
);

INVx1_ASAP7_75t_L g17669 ( 
.A(n_17350),
.Y(n_17669)
);

OR2x2_ASAP7_75t_L g17670 ( 
.A(n_17341),
.B(n_10272),
.Y(n_17670)
);

INVx1_ASAP7_75t_L g17671 ( 
.A(n_17243),
.Y(n_17671)
);

OR2x2_ASAP7_75t_L g17672 ( 
.A(n_17423),
.B(n_10272),
.Y(n_17672)
);

AND2x2_ASAP7_75t_L g17673 ( 
.A(n_17457),
.B(n_10279),
.Y(n_17673)
);

AOI21xp5_ASAP7_75t_L g17674 ( 
.A1(n_17437),
.A2(n_9647),
.B(n_9641),
.Y(n_17674)
);

INVx1_ASAP7_75t_L g17675 ( 
.A(n_17258),
.Y(n_17675)
);

INVx1_ASAP7_75t_L g17676 ( 
.A(n_17262),
.Y(n_17676)
);

NAND2xp67_ASAP7_75t_L g17677 ( 
.A(n_17367),
.B(n_10279),
.Y(n_17677)
);

INVx1_ASAP7_75t_SL g17678 ( 
.A(n_17517),
.Y(n_17678)
);

INVx3_ASAP7_75t_L g17679 ( 
.A(n_17317),
.Y(n_17679)
);

NOR2x1_ASAP7_75t_L g17680 ( 
.A(n_17427),
.B(n_9581),
.Y(n_17680)
);

AOI221xp5_ASAP7_75t_L g17681 ( 
.A1(n_17389),
.A2(n_9647),
.B1(n_10280),
.B2(n_10282),
.C(n_10279),
.Y(n_17681)
);

AOI22xp5_ASAP7_75t_L g17682 ( 
.A1(n_17390),
.A2(n_9647),
.B1(n_10150),
.B2(n_10135),
.Y(n_17682)
);

INVx1_ASAP7_75t_L g17683 ( 
.A(n_17308),
.Y(n_17683)
);

AO221x1_ASAP7_75t_L g17684 ( 
.A1(n_17293),
.A2(n_8284),
.B1(n_9391),
.B2(n_9392),
.C(n_9376),
.Y(n_17684)
);

A2O1A1Ixp33_ASAP7_75t_L g17685 ( 
.A1(n_17214),
.A2(n_9590),
.B(n_9615),
.C(n_9577),
.Y(n_17685)
);

NAND2xp5_ASAP7_75t_L g17686 ( 
.A(n_17459),
.B(n_9581),
.Y(n_17686)
);

OAI22xp5_ASAP7_75t_L g17687 ( 
.A1(n_17385),
.A2(n_9391),
.B1(n_9395),
.B2(n_9392),
.Y(n_17687)
);

INVx1_ASAP7_75t_L g17688 ( 
.A(n_17398),
.Y(n_17688)
);

INVx1_ASAP7_75t_L g17689 ( 
.A(n_17394),
.Y(n_17689)
);

INVx2_ASAP7_75t_L g17690 ( 
.A(n_17382),
.Y(n_17690)
);

NOR3xp33_ASAP7_75t_L g17691 ( 
.A(n_17318),
.B(n_5652),
.C(n_5627),
.Y(n_17691)
);

INVx1_ASAP7_75t_L g17692 ( 
.A(n_17409),
.Y(n_17692)
);

NAND2x1p5_ASAP7_75t_L g17693 ( 
.A(n_17444),
.B(n_17454),
.Y(n_17693)
);

NAND2xp5_ASAP7_75t_L g17694 ( 
.A(n_17493),
.B(n_9582),
.Y(n_17694)
);

A2O1A1Ixp33_ASAP7_75t_L g17695 ( 
.A1(n_17234),
.A2(n_9615),
.B(n_9590),
.C(n_9792),
.Y(n_17695)
);

OR2x2_ASAP7_75t_L g17696 ( 
.A(n_17352),
.B(n_10280),
.Y(n_17696)
);

OAI22xp5_ASAP7_75t_L g17697 ( 
.A1(n_17329),
.A2(n_9395),
.B1(n_9402),
.B2(n_9397),
.Y(n_17697)
);

AOI22x1_ASAP7_75t_SL g17698 ( 
.A1(n_17342),
.A2(n_9402),
.B1(n_9405),
.B2(n_9397),
.Y(n_17698)
);

INVx2_ASAP7_75t_L g17699 ( 
.A(n_17371),
.Y(n_17699)
);

AND2x2_ASAP7_75t_L g17700 ( 
.A(n_17464),
.B(n_10280),
.Y(n_17700)
);

INVx1_ASAP7_75t_L g17701 ( 
.A(n_17484),
.Y(n_17701)
);

AND2x2_ASAP7_75t_L g17702 ( 
.A(n_17372),
.B(n_10282),
.Y(n_17702)
);

AND2x2_ASAP7_75t_L g17703 ( 
.A(n_17451),
.B(n_10282),
.Y(n_17703)
);

OAI22xp5_ASAP7_75t_L g17704 ( 
.A1(n_17359),
.A2(n_9397),
.B1(n_9405),
.B2(n_9402),
.Y(n_17704)
);

INVx2_ASAP7_75t_L g17705 ( 
.A(n_17220),
.Y(n_17705)
);

NAND2xp5_ASAP7_75t_L g17706 ( 
.A(n_17525),
.B(n_9582),
.Y(n_17706)
);

OAI32xp33_ASAP7_75t_L g17707 ( 
.A1(n_17360),
.A2(n_9704),
.A3(n_9677),
.B1(n_9655),
.B2(n_10135),
.Y(n_17707)
);

AOI21xp33_ASAP7_75t_L g17708 ( 
.A1(n_17473),
.A2(n_9677),
.B(n_9655),
.Y(n_17708)
);

OAI21xp5_ASAP7_75t_L g17709 ( 
.A1(n_17453),
.A2(n_10222),
.B(n_10192),
.Y(n_17709)
);

INVx1_ASAP7_75t_L g17710 ( 
.A(n_17363),
.Y(n_17710)
);

OAI21xp5_ASAP7_75t_SL g17711 ( 
.A1(n_17374),
.A2(n_8429),
.B(n_8396),
.Y(n_17711)
);

OAI21xp5_ASAP7_75t_L g17712 ( 
.A1(n_17323),
.A2(n_10222),
.B(n_10192),
.Y(n_17712)
);

O2A1O1Ixp33_ASAP7_75t_L g17713 ( 
.A1(n_17515),
.A2(n_9677),
.B(n_9704),
.C(n_9655),
.Y(n_17713)
);

NAND2xp5_ASAP7_75t_L g17714 ( 
.A(n_17334),
.B(n_17345),
.Y(n_17714)
);

AND2x2_ASAP7_75t_L g17715 ( 
.A(n_17417),
.B(n_10283),
.Y(n_17715)
);

NOR2xp67_ASAP7_75t_L g17716 ( 
.A(n_17347),
.B(n_9585),
.Y(n_17716)
);

HB1xp67_ASAP7_75t_L g17717 ( 
.A(n_17314),
.Y(n_17717)
);

AND2x2_ASAP7_75t_L g17718 ( 
.A(n_17483),
.B(n_10283),
.Y(n_17718)
);

INVx1_ASAP7_75t_L g17719 ( 
.A(n_17300),
.Y(n_17719)
);

AOI21xp33_ASAP7_75t_SL g17720 ( 
.A1(n_17354),
.A2(n_9615),
.B(n_8549),
.Y(n_17720)
);

OAI322xp33_ASAP7_75t_L g17721 ( 
.A1(n_17416),
.A2(n_9426),
.A3(n_9413),
.B1(n_9430),
.B2(n_9432),
.C1(n_9429),
.C2(n_9405),
.Y(n_17721)
);

AOI221xp5_ASAP7_75t_L g17722 ( 
.A1(n_17343),
.A2(n_10290),
.B1(n_10285),
.B2(n_10283),
.C(n_10155),
.Y(n_17722)
);

NOR2xp33_ASAP7_75t_L g17723 ( 
.A(n_17468),
.B(n_9585),
.Y(n_17723)
);

OAI22xp5_ASAP7_75t_L g17724 ( 
.A1(n_17432),
.A2(n_9413),
.B1(n_9429),
.B2(n_9426),
.Y(n_17724)
);

NOR2x1_ASAP7_75t_L g17725 ( 
.A(n_17458),
.B(n_17420),
.Y(n_17725)
);

OAI21xp5_ASAP7_75t_L g17726 ( 
.A1(n_17489),
.A2(n_10235),
.B(n_10232),
.Y(n_17726)
);

AOI221xp5_ASAP7_75t_L g17727 ( 
.A1(n_17402),
.A2(n_17376),
.B1(n_17426),
.B2(n_17281),
.C(n_17237),
.Y(n_17727)
);

OAI21xp33_ASAP7_75t_SL g17728 ( 
.A1(n_17325),
.A2(n_9817),
.B(n_9792),
.Y(n_17728)
);

INVx2_ASAP7_75t_L g17729 ( 
.A(n_17218),
.Y(n_17729)
);

INVx1_ASAP7_75t_L g17730 ( 
.A(n_17286),
.Y(n_17730)
);

NOR2xp33_ASAP7_75t_L g17731 ( 
.A(n_17461),
.B(n_9594),
.Y(n_17731)
);

NAND2xp5_ASAP7_75t_L g17732 ( 
.A(n_17480),
.B(n_9594),
.Y(n_17732)
);

AOI221xp5_ASAP7_75t_L g17733 ( 
.A1(n_17408),
.A2(n_10290),
.B1(n_10285),
.B2(n_10155),
.C(n_10150),
.Y(n_17733)
);

XOR2x2_ASAP7_75t_L g17734 ( 
.A(n_17482),
.B(n_7825),
.Y(n_17734)
);

INVx1_ASAP7_75t_L g17735 ( 
.A(n_17503),
.Y(n_17735)
);

INVx1_ASAP7_75t_SL g17736 ( 
.A(n_17405),
.Y(n_17736)
);

AOI332xp33_ASAP7_75t_L g17737 ( 
.A1(n_17439),
.A2(n_9413),
.A3(n_9432),
.B1(n_9429),
.B2(n_9426),
.B3(n_9441),
.C1(n_9440),
.C2(n_9430),
.Y(n_17737)
);

BUFx2_ASAP7_75t_L g17738 ( 
.A(n_17335),
.Y(n_17738)
);

AOI32xp33_ASAP7_75t_L g17739 ( 
.A1(n_17495),
.A2(n_9850),
.A3(n_9817),
.B1(n_9792),
.B2(n_9440),
.Y(n_17739)
);

INVx1_ASAP7_75t_L g17740 ( 
.A(n_17301),
.Y(n_17740)
);

INVxp67_ASAP7_75t_L g17741 ( 
.A(n_17462),
.Y(n_17741)
);

INVx1_ASAP7_75t_L g17742 ( 
.A(n_17445),
.Y(n_17742)
);

AND2x2_ASAP7_75t_L g17743 ( 
.A(n_17440),
.B(n_10285),
.Y(n_17743)
);

NOR2xp33_ASAP7_75t_L g17744 ( 
.A(n_17362),
.B(n_9598),
.Y(n_17744)
);

NOR2x1p5_ASAP7_75t_L g17745 ( 
.A(n_17364),
.B(n_6932),
.Y(n_17745)
);

OAI21xp33_ASAP7_75t_L g17746 ( 
.A1(n_17404),
.A2(n_10150),
.B(n_10135),
.Y(n_17746)
);

HB1xp67_ASAP7_75t_L g17747 ( 
.A(n_17512),
.Y(n_17747)
);

INVx1_ASAP7_75t_L g17748 ( 
.A(n_17513),
.Y(n_17748)
);

OAI21xp5_ASAP7_75t_L g17749 ( 
.A1(n_17268),
.A2(n_10235),
.B(n_10232),
.Y(n_17749)
);

OAI21xp5_ASAP7_75t_L g17750 ( 
.A1(n_17249),
.A2(n_10235),
.B(n_10232),
.Y(n_17750)
);

INVx1_ASAP7_75t_L g17751 ( 
.A(n_17264),
.Y(n_17751)
);

HB1xp67_ASAP7_75t_L g17752 ( 
.A(n_17225),
.Y(n_17752)
);

OAI22xp33_ASAP7_75t_SL g17753 ( 
.A1(n_17443),
.A2(n_10290),
.B1(n_10155),
.B2(n_9704),
.Y(n_17753)
);

OAI21xp33_ASAP7_75t_L g17754 ( 
.A1(n_17351),
.A2(n_9432),
.B(n_9430),
.Y(n_17754)
);

INVxp67_ASAP7_75t_L g17755 ( 
.A(n_17434),
.Y(n_17755)
);

AND2x2_ASAP7_75t_L g17756 ( 
.A(n_17455),
.B(n_17393),
.Y(n_17756)
);

INVx1_ASAP7_75t_SL g17757 ( 
.A(n_17356),
.Y(n_17757)
);

NAND2xp5_ASAP7_75t_L g17758 ( 
.A(n_17448),
.B(n_9598),
.Y(n_17758)
);

NAND2xp5_ASAP7_75t_L g17759 ( 
.A(n_17452),
.B(n_9601),
.Y(n_17759)
);

A2O1A1Ixp33_ASAP7_75t_L g17760 ( 
.A1(n_17521),
.A2(n_9850),
.B(n_9817),
.C(n_9441),
.Y(n_17760)
);

AOI221xp5_ASAP7_75t_L g17761 ( 
.A1(n_17494),
.A2(n_9441),
.B1(n_9465),
.B2(n_9451),
.C(n_9440),
.Y(n_17761)
);

INVx1_ASAP7_75t_SL g17762 ( 
.A(n_17344),
.Y(n_17762)
);

INVx1_ASAP7_75t_L g17763 ( 
.A(n_17479),
.Y(n_17763)
);

INVx1_ASAP7_75t_SL g17764 ( 
.A(n_17276),
.Y(n_17764)
);

INVx1_ASAP7_75t_L g17765 ( 
.A(n_17441),
.Y(n_17765)
);

INVx1_ASAP7_75t_L g17766 ( 
.A(n_17430),
.Y(n_17766)
);

NAND3xp33_ASAP7_75t_SL g17767 ( 
.A(n_17460),
.B(n_8549),
.C(n_8429),
.Y(n_17767)
);

INVx1_ASAP7_75t_L g17768 ( 
.A(n_17496),
.Y(n_17768)
);

AND2x2_ASAP7_75t_L g17769 ( 
.A(n_17436),
.B(n_9601),
.Y(n_17769)
);

NAND2xp5_ASAP7_75t_L g17770 ( 
.A(n_17429),
.B(n_9607),
.Y(n_17770)
);

OAI21xp33_ASAP7_75t_L g17771 ( 
.A1(n_17209),
.A2(n_9465),
.B(n_9451),
.Y(n_17771)
);

AOI21xp33_ASAP7_75t_SL g17772 ( 
.A1(n_17463),
.A2(n_17470),
.B(n_17469),
.Y(n_17772)
);

OAI221xp5_ASAP7_75t_L g17773 ( 
.A1(n_17442),
.A2(n_8608),
.B1(n_8687),
.B2(n_8549),
.C(n_8429),
.Y(n_17773)
);

AND2x2_ASAP7_75t_L g17774 ( 
.A(n_17504),
.B(n_9607),
.Y(n_17774)
);

OAI221xp5_ASAP7_75t_L g17775 ( 
.A1(n_17506),
.A2(n_8740),
.B1(n_8754),
.B2(n_8687),
.C(n_8608),
.Y(n_17775)
);

NAND2xp5_ASAP7_75t_L g17776 ( 
.A(n_17501),
.B(n_9610),
.Y(n_17776)
);

INVx1_ASAP7_75t_L g17777 ( 
.A(n_17498),
.Y(n_17777)
);

INVxp33_ASAP7_75t_L g17778 ( 
.A(n_17311),
.Y(n_17778)
);

NAND2xp5_ASAP7_75t_L g17779 ( 
.A(n_17472),
.B(n_9610),
.Y(n_17779)
);

OAI21xp5_ASAP7_75t_L g17780 ( 
.A1(n_17490),
.A2(n_10252),
.B(n_7955),
.Y(n_17780)
);

INVx2_ASAP7_75t_L g17781 ( 
.A(n_17488),
.Y(n_17781)
);

INVx1_ASAP7_75t_L g17782 ( 
.A(n_17288),
.Y(n_17782)
);

OAI21xp5_ASAP7_75t_L g17783 ( 
.A1(n_17471),
.A2(n_17322),
.B(n_17475),
.Y(n_17783)
);

NAND2xp5_ASAP7_75t_L g17784 ( 
.A(n_17527),
.B(n_9612),
.Y(n_17784)
);

AND2x2_ASAP7_75t_L g17785 ( 
.A(n_17505),
.B(n_9612),
.Y(n_17785)
);

AOI22xp33_ASAP7_75t_L g17786 ( 
.A1(n_17219),
.A2(n_17231),
.B1(n_17285),
.B2(n_17519),
.Y(n_17786)
);

NAND2xp33_ASAP7_75t_SL g17787 ( 
.A(n_17260),
.B(n_8653),
.Y(n_17787)
);

INVxp67_ASAP7_75t_L g17788 ( 
.A(n_17365),
.Y(n_17788)
);

OAI22xp5_ASAP7_75t_L g17789 ( 
.A1(n_17221),
.A2(n_9451),
.B1(n_9476),
.B2(n_9465),
.Y(n_17789)
);

OR2x2_ASAP7_75t_L g17790 ( 
.A(n_17522),
.B(n_9476),
.Y(n_17790)
);

INVx1_ASAP7_75t_L g17791 ( 
.A(n_17346),
.Y(n_17791)
);

NOR2xp33_ASAP7_75t_L g17792 ( 
.A(n_17485),
.B(n_9613),
.Y(n_17792)
);

INVx1_ASAP7_75t_SL g17793 ( 
.A(n_17368),
.Y(n_17793)
);

NAND2xp5_ASAP7_75t_L g17794 ( 
.A(n_17378),
.B(n_9613),
.Y(n_17794)
);

AOI22xp5_ASAP7_75t_L g17795 ( 
.A1(n_17232),
.A2(n_9477),
.B1(n_9478),
.B2(n_9476),
.Y(n_17795)
);

INVx1_ASAP7_75t_L g17796 ( 
.A(n_17516),
.Y(n_17796)
);

OR2x2_ASAP7_75t_L g17797 ( 
.A(n_17556),
.B(n_17497),
.Y(n_17797)
);

NOR2xp33_ASAP7_75t_L g17798 ( 
.A(n_17530),
.B(n_17514),
.Y(n_17798)
);

INVx1_ASAP7_75t_L g17799 ( 
.A(n_17542),
.Y(n_17799)
);

NAND2xp5_ASAP7_75t_L g17800 ( 
.A(n_17562),
.B(n_17242),
.Y(n_17800)
);

INVx1_ASAP7_75t_L g17801 ( 
.A(n_17600),
.Y(n_17801)
);

AOI221xp5_ASAP7_75t_L g17802 ( 
.A1(n_17559),
.A2(n_17247),
.B1(n_17298),
.B2(n_17287),
.C(n_17523),
.Y(n_17802)
);

INVx2_ASAP7_75t_L g17803 ( 
.A(n_17693),
.Y(n_17803)
);

AOI22xp5_ASAP7_75t_L g17804 ( 
.A1(n_17582),
.A2(n_17396),
.B1(n_17227),
.B2(n_17520),
.Y(n_17804)
);

NAND2xp5_ASAP7_75t_L g17805 ( 
.A(n_17574),
.B(n_17486),
.Y(n_17805)
);

HB1xp67_ASAP7_75t_L g17806 ( 
.A(n_17717),
.Y(n_17806)
);

INVx1_ASAP7_75t_L g17807 ( 
.A(n_17738),
.Y(n_17807)
);

AOI222xp33_ASAP7_75t_L g17808 ( 
.A1(n_17564),
.A2(n_17500),
.B1(n_17509),
.B2(n_17481),
.C1(n_17487),
.C2(n_17297),
.Y(n_17808)
);

OAI222xp33_ASAP7_75t_L g17809 ( 
.A1(n_17622),
.A2(n_17446),
.B1(n_17524),
.B2(n_17492),
.C1(n_17476),
.C2(n_17478),
.Y(n_17809)
);

INVx1_ASAP7_75t_L g17810 ( 
.A(n_17537),
.Y(n_17810)
);

INVxp33_ASAP7_75t_L g17811 ( 
.A(n_17725),
.Y(n_17811)
);

INVx2_ASAP7_75t_L g17812 ( 
.A(n_17581),
.Y(n_17812)
);

INVxp67_ASAP7_75t_L g17813 ( 
.A(n_17539),
.Y(n_17813)
);

OR2x2_ASAP7_75t_L g17814 ( 
.A(n_17551),
.B(n_17467),
.Y(n_17814)
);

INVx1_ASAP7_75t_L g17815 ( 
.A(n_17747),
.Y(n_17815)
);

OAI22xp5_ASAP7_75t_L g17816 ( 
.A1(n_17587),
.A2(n_17273),
.B1(n_17278),
.B2(n_17275),
.Y(n_17816)
);

NOR2xp33_ASAP7_75t_L g17817 ( 
.A(n_17646),
.B(n_17412),
.Y(n_17817)
);

INVx1_ASAP7_75t_L g17818 ( 
.A(n_17550),
.Y(n_17818)
);

AND2x2_ASAP7_75t_L g17819 ( 
.A(n_17756),
.B(n_17269),
.Y(n_17819)
);

INVx1_ASAP7_75t_L g17820 ( 
.A(n_17653),
.Y(n_17820)
);

NAND2xp5_ASAP7_75t_L g17821 ( 
.A(n_17679),
.B(n_17239),
.Y(n_17821)
);

NAND2xp5_ASAP7_75t_L g17822 ( 
.A(n_17679),
.B(n_17295),
.Y(n_17822)
);

INVx1_ASAP7_75t_L g17823 ( 
.A(n_17544),
.Y(n_17823)
);

INVx1_ASAP7_75t_L g17824 ( 
.A(n_17547),
.Y(n_17824)
);

AND2x2_ASAP7_75t_L g17825 ( 
.A(n_17583),
.B(n_17450),
.Y(n_17825)
);

AOI311xp33_ASAP7_75t_L g17826 ( 
.A1(n_17538),
.A2(n_17532),
.A3(n_17618),
.B(n_17548),
.C(n_17552),
.Y(n_17826)
);

NAND2xp5_ASAP7_75t_L g17827 ( 
.A(n_17568),
.B(n_9626),
.Y(n_17827)
);

O2A1O1Ixp33_ASAP7_75t_L g17828 ( 
.A1(n_17534),
.A2(n_9478),
.B(n_9479),
.C(n_9477),
.Y(n_17828)
);

INVx1_ASAP7_75t_L g17829 ( 
.A(n_17752),
.Y(n_17829)
);

NAND2xp5_ASAP7_75t_L g17830 ( 
.A(n_17627),
.B(n_9626),
.Y(n_17830)
);

AND2x2_ASAP7_75t_L g17831 ( 
.A(n_17699),
.B(n_9630),
.Y(n_17831)
);

AOI21xp33_ASAP7_75t_L g17832 ( 
.A1(n_17778),
.A2(n_17662),
.B(n_17678),
.Y(n_17832)
);

O2A1O1Ixp5_ASAP7_75t_SL g17833 ( 
.A1(n_17563),
.A2(n_9631),
.B(n_9633),
.C(n_9630),
.Y(n_17833)
);

INVx1_ASAP7_75t_SL g17834 ( 
.A(n_17593),
.Y(n_17834)
);

INVx1_ASAP7_75t_L g17835 ( 
.A(n_17546),
.Y(n_17835)
);

NAND2x1p5_ASAP7_75t_L g17836 ( 
.A(n_17597),
.B(n_8593),
.Y(n_17836)
);

A2O1A1Ixp33_ASAP7_75t_L g17837 ( 
.A1(n_17596),
.A2(n_9850),
.B(n_9478),
.C(n_9479),
.Y(n_17837)
);

INVx1_ASAP7_75t_L g17838 ( 
.A(n_17545),
.Y(n_17838)
);

NAND2xp5_ASAP7_75t_L g17839 ( 
.A(n_17736),
.B(n_9631),
.Y(n_17839)
);

NAND2xp5_ASAP7_75t_L g17840 ( 
.A(n_17621),
.B(n_9633),
.Y(n_17840)
);

INVxp67_ASAP7_75t_SL g17841 ( 
.A(n_17683),
.Y(n_17841)
);

NAND2xp5_ASAP7_75t_L g17842 ( 
.A(n_17553),
.B(n_9640),
.Y(n_17842)
);

AOI21xp33_ASAP7_75t_SL g17843 ( 
.A1(n_17555),
.A2(n_8687),
.B(n_8608),
.Y(n_17843)
);

OR2x2_ASAP7_75t_L g17844 ( 
.A(n_17554),
.B(n_9477),
.Y(n_17844)
);

OAI21xp5_ASAP7_75t_SL g17845 ( 
.A1(n_17636),
.A2(n_8740),
.B(n_8687),
.Y(n_17845)
);

OR4x1_ASAP7_75t_L g17846 ( 
.A(n_17543),
.B(n_9644),
.C(n_9645),
.D(n_9640),
.Y(n_17846)
);

INVx2_ASAP7_75t_L g17847 ( 
.A(n_17536),
.Y(n_17847)
);

INVx2_ASAP7_75t_L g17848 ( 
.A(n_17658),
.Y(n_17848)
);

NAND2xp5_ASAP7_75t_L g17849 ( 
.A(n_17589),
.B(n_9644),
.Y(n_17849)
);

INVx1_ASAP7_75t_L g17850 ( 
.A(n_17608),
.Y(n_17850)
);

NAND2xp5_ASAP7_75t_L g17851 ( 
.A(n_17603),
.B(n_17690),
.Y(n_17851)
);

OAI22xp5_ASAP7_75t_L g17852 ( 
.A1(n_17735),
.A2(n_9479),
.B1(n_9503),
.B2(n_9502),
.Y(n_17852)
);

OAI322xp33_ASAP7_75t_L g17853 ( 
.A1(n_17549),
.A2(n_9505),
.A3(n_9502),
.B1(n_9508),
.B2(n_9514),
.C1(n_9512),
.C2(n_9503),
.Y(n_17853)
);

AOI21xp5_ASAP7_75t_L g17854 ( 
.A1(n_17540),
.A2(n_17620),
.B(n_17529),
.Y(n_17854)
);

A2O1A1Ixp33_ASAP7_75t_L g17855 ( 
.A1(n_17643),
.A2(n_9503),
.B(n_9505),
.C(n_9502),
.Y(n_17855)
);

INVx1_ASAP7_75t_L g17856 ( 
.A(n_17677),
.Y(n_17856)
);

INVx2_ASAP7_75t_L g17857 ( 
.A(n_17638),
.Y(n_17857)
);

OAI32xp33_ASAP7_75t_L g17858 ( 
.A1(n_17560),
.A2(n_9508),
.A3(n_9514),
.B1(n_9512),
.B2(n_9505),
.Y(n_17858)
);

NOR2x1_ASAP7_75t_L g17859 ( 
.A(n_17533),
.B(n_9645),
.Y(n_17859)
);

OR2x2_ASAP7_75t_L g17860 ( 
.A(n_17641),
.B(n_9508),
.Y(n_17860)
);

OAI22xp33_ASAP7_75t_L g17861 ( 
.A1(n_17541),
.A2(n_9512),
.B1(n_9518),
.B2(n_9514),
.Y(n_17861)
);

OR2x2_ASAP7_75t_L g17862 ( 
.A(n_17611),
.B(n_9518),
.Y(n_17862)
);

OR2x2_ASAP7_75t_L g17863 ( 
.A(n_17612),
.B(n_9518),
.Y(n_17863)
);

AND2x2_ASAP7_75t_L g17864 ( 
.A(n_17528),
.B(n_17616),
.Y(n_17864)
);

NAND2xp5_ASAP7_75t_L g17865 ( 
.A(n_17614),
.B(n_17632),
.Y(n_17865)
);

AND2x2_ASAP7_75t_L g17866 ( 
.A(n_17710),
.B(n_9650),
.Y(n_17866)
);

NAND3xp33_ASAP7_75t_L g17867 ( 
.A(n_17727),
.B(n_17531),
.C(n_17535),
.Y(n_17867)
);

INVx1_ASAP7_75t_L g17868 ( 
.A(n_17680),
.Y(n_17868)
);

OAI221xp5_ASAP7_75t_L g17869 ( 
.A1(n_17786),
.A2(n_9522),
.B1(n_8925),
.B2(n_8754),
.C(n_8740),
.Y(n_17869)
);

INVx1_ASAP7_75t_SL g17870 ( 
.A(n_17757),
.Y(n_17870)
);

INVx1_ASAP7_75t_L g17871 ( 
.A(n_17644),
.Y(n_17871)
);

OAI221xp5_ASAP7_75t_L g17872 ( 
.A1(n_17613),
.A2(n_9522),
.B1(n_8925),
.B2(n_8754),
.C(n_8740),
.Y(n_17872)
);

AO221x1_ASAP7_75t_L g17873 ( 
.A1(n_17772),
.A2(n_9522),
.B1(n_8284),
.B2(n_7196),
.C(n_7199),
.Y(n_17873)
);

NAND2xp5_ASAP7_75t_L g17874 ( 
.A(n_17669),
.B(n_9650),
.Y(n_17874)
);

AND2x2_ASAP7_75t_L g17875 ( 
.A(n_17661),
.B(n_17689),
.Y(n_17875)
);

NAND2xp5_ASAP7_75t_L g17876 ( 
.A(n_17606),
.B(n_9658),
.Y(n_17876)
);

NAND2xp5_ASAP7_75t_L g17877 ( 
.A(n_17762),
.B(n_9658),
.Y(n_17877)
);

NOR2xp33_ASAP7_75t_L g17878 ( 
.A(n_17650),
.B(n_17692),
.Y(n_17878)
);

INVx2_ASAP7_75t_L g17879 ( 
.A(n_17705),
.Y(n_17879)
);

AOI22xp5_ASAP7_75t_L g17880 ( 
.A1(n_17688),
.A2(n_9660),
.B1(n_9669),
.B2(n_9666),
.Y(n_17880)
);

OAI21xp33_ASAP7_75t_L g17881 ( 
.A1(n_17655),
.A2(n_8353),
.B(n_7950),
.Y(n_17881)
);

NOR2xp33_ASAP7_75t_L g17882 ( 
.A(n_17701),
.B(n_9660),
.Y(n_17882)
);

INVx1_ASAP7_75t_L g17883 ( 
.A(n_17571),
.Y(n_17883)
);

OAI211xp5_ASAP7_75t_L g17884 ( 
.A1(n_17557),
.A2(n_9669),
.B(n_9670),
.C(n_9666),
.Y(n_17884)
);

AOI21xp33_ASAP7_75t_L g17885 ( 
.A1(n_17742),
.A2(n_8012),
.B(n_10252),
.Y(n_17885)
);

INVx1_ASAP7_75t_L g17886 ( 
.A(n_17748),
.Y(n_17886)
);

INVx1_ASAP7_75t_L g17887 ( 
.A(n_17573),
.Y(n_17887)
);

AOI211xp5_ASAP7_75t_L g17888 ( 
.A1(n_17647),
.A2(n_7955),
.B(n_7971),
.C(n_7932),
.Y(n_17888)
);

AOI21xp5_ASAP7_75t_L g17889 ( 
.A1(n_17666),
.A2(n_9672),
.B(n_9670),
.Y(n_17889)
);

AND2x2_ASAP7_75t_L g17890 ( 
.A(n_17591),
.B(n_9672),
.Y(n_17890)
);

NAND2xp5_ASAP7_75t_SL g17891 ( 
.A(n_17648),
.B(n_9675),
.Y(n_17891)
);

OAI21xp5_ASAP7_75t_L g17892 ( 
.A1(n_17741),
.A2(n_10252),
.B(n_7955),
.Y(n_17892)
);

INVx1_ASAP7_75t_L g17893 ( 
.A(n_17649),
.Y(n_17893)
);

OAI21xp5_ASAP7_75t_SL g17894 ( 
.A1(n_17572),
.A2(n_8925),
.B(n_8754),
.Y(n_17894)
);

NAND2xp5_ASAP7_75t_L g17895 ( 
.A(n_17793),
.B(n_9675),
.Y(n_17895)
);

INVx1_ASAP7_75t_L g17896 ( 
.A(n_17660),
.Y(n_17896)
);

OAI22xp33_ASAP7_75t_SL g17897 ( 
.A1(n_17696),
.A2(n_9686),
.B1(n_9688),
.B2(n_9684),
.Y(n_17897)
);

INVx1_ASAP7_75t_SL g17898 ( 
.A(n_17764),
.Y(n_17898)
);

NAND2xp5_ASAP7_75t_L g17899 ( 
.A(n_17755),
.B(n_9684),
.Y(n_17899)
);

NAND2xp5_ASAP7_75t_L g17900 ( 
.A(n_17602),
.B(n_9686),
.Y(n_17900)
);

INVx1_ASAP7_75t_L g17901 ( 
.A(n_17714),
.Y(n_17901)
);

INVxp67_ASAP7_75t_L g17902 ( 
.A(n_17590),
.Y(n_17902)
);

OAI22xp5_ASAP7_75t_L g17903 ( 
.A1(n_17656),
.A2(n_9688),
.B1(n_9699),
.B2(n_9696),
.Y(n_17903)
);

INVx1_ASAP7_75t_L g17904 ( 
.A(n_17671),
.Y(n_17904)
);

BUFx2_ASAP7_75t_L g17905 ( 
.A(n_17584),
.Y(n_17905)
);

INVx1_ASAP7_75t_L g17906 ( 
.A(n_17729),
.Y(n_17906)
);

INVx1_ASAP7_75t_L g17907 ( 
.A(n_17675),
.Y(n_17907)
);

NAND2xp5_ASAP7_75t_L g17908 ( 
.A(n_17782),
.B(n_9696),
.Y(n_17908)
);

INVx1_ASAP7_75t_L g17909 ( 
.A(n_17676),
.Y(n_17909)
);

INVx1_ASAP7_75t_L g17910 ( 
.A(n_17791),
.Y(n_17910)
);

A2O1A1Ixp33_ASAP7_75t_L g17911 ( 
.A1(n_17628),
.A2(n_10275),
.B(n_9709),
.C(n_9710),
.Y(n_17911)
);

INVx1_ASAP7_75t_L g17912 ( 
.A(n_17604),
.Y(n_17912)
);

AOI221x1_ASAP7_75t_SL g17913 ( 
.A1(n_17768),
.A2(n_9710),
.B1(n_9713),
.B2(n_9709),
.C(n_9699),
.Y(n_17913)
);

INVx1_ASAP7_75t_L g17914 ( 
.A(n_17645),
.Y(n_17914)
);

OR2x6_ASAP7_75t_L g17915 ( 
.A(n_17777),
.B(n_7077),
.Y(n_17915)
);

NOR2xp33_ASAP7_75t_L g17916 ( 
.A(n_17788),
.B(n_9713),
.Y(n_17916)
);

AOI22xp5_ASAP7_75t_L g17917 ( 
.A1(n_17787),
.A2(n_9715),
.B1(n_9721),
.B2(n_9720),
.Y(n_17917)
);

INVx1_ASAP7_75t_L g17918 ( 
.A(n_17558),
.Y(n_17918)
);

INVx1_ASAP7_75t_L g17919 ( 
.A(n_17706),
.Y(n_17919)
);

NAND2xp5_ASAP7_75t_L g17920 ( 
.A(n_17781),
.B(n_9715),
.Y(n_17920)
);

O2A1O1Ixp33_ASAP7_75t_SL g17921 ( 
.A1(n_17668),
.A2(n_9720),
.B(n_9723),
.C(n_9721),
.Y(n_17921)
);

NAND2xp5_ASAP7_75t_L g17922 ( 
.A(n_17579),
.B(n_9723),
.Y(n_17922)
);

AOI221xp5_ASAP7_75t_L g17923 ( 
.A1(n_17601),
.A2(n_8284),
.B1(n_9745),
.B2(n_9746),
.C(n_9731),
.Y(n_17923)
);

O2A1O1Ixp33_ASAP7_75t_SL g17924 ( 
.A1(n_17732),
.A2(n_9731),
.B(n_9746),
.C(n_9745),
.Y(n_17924)
);

INVx1_ASAP7_75t_L g17925 ( 
.A(n_17639),
.Y(n_17925)
);

INVx1_ASAP7_75t_L g17926 ( 
.A(n_17694),
.Y(n_17926)
);

OAI22xp5_ASAP7_75t_L g17927 ( 
.A1(n_17640),
.A2(n_9749),
.B1(n_9753),
.B2(n_9751),
.Y(n_17927)
);

OAI21xp5_ASAP7_75t_L g17928 ( 
.A1(n_17783),
.A2(n_7971),
.B(n_7932),
.Y(n_17928)
);

NOR2xp33_ASAP7_75t_L g17929 ( 
.A(n_17607),
.B(n_17740),
.Y(n_17929)
);

NOR2x1_ASAP7_75t_L g17930 ( 
.A(n_17751),
.B(n_9749),
.Y(n_17930)
);

INVx1_ASAP7_75t_L g17931 ( 
.A(n_17716),
.Y(n_17931)
);

INVx1_ASAP7_75t_L g17932 ( 
.A(n_17570),
.Y(n_17932)
);

INVx1_ASAP7_75t_L g17933 ( 
.A(n_17575),
.Y(n_17933)
);

OAI211xp5_ASAP7_75t_L g17934 ( 
.A1(n_17730),
.A2(n_9753),
.B(n_9754),
.C(n_9751),
.Y(n_17934)
);

NAND2x1p5_ASAP7_75t_L g17935 ( 
.A(n_17763),
.B(n_8593),
.Y(n_17935)
);

OAI21xp5_ASAP7_75t_SL g17936 ( 
.A1(n_17565),
.A2(n_8925),
.B(n_7881),
.Y(n_17936)
);

NAND2x1_ASAP7_75t_L g17937 ( 
.A(n_17577),
.B(n_9754),
.Y(n_17937)
);

AOI22xp33_ASAP7_75t_L g17938 ( 
.A1(n_17609),
.A2(n_7322),
.B1(n_7350),
.B2(n_7320),
.Y(n_17938)
);

NOR2xp33_ASAP7_75t_L g17939 ( 
.A(n_17719),
.B(n_9757),
.Y(n_17939)
);

AND2x2_ASAP7_75t_L g17940 ( 
.A(n_17745),
.B(n_9757),
.Y(n_17940)
);

INVx1_ASAP7_75t_L g17941 ( 
.A(n_17585),
.Y(n_17941)
);

AOI21xp5_ASAP7_75t_L g17942 ( 
.A1(n_17796),
.A2(n_9763),
.B(n_9762),
.Y(n_17942)
);

NAND2xp5_ASAP7_75t_L g17943 ( 
.A(n_17561),
.B(n_9762),
.Y(n_17943)
);

OR2x2_ASAP7_75t_L g17944 ( 
.A(n_17642),
.B(n_9763),
.Y(n_17944)
);

INVx3_ASAP7_75t_L g17945 ( 
.A(n_17734),
.Y(n_17945)
);

INVx1_ASAP7_75t_L g17946 ( 
.A(n_17774),
.Y(n_17946)
);

INVx2_ASAP7_75t_L g17947 ( 
.A(n_17769),
.Y(n_17947)
);

OAI21xp33_ASAP7_75t_SL g17948 ( 
.A1(n_17631),
.A2(n_10275),
.B(n_10026),
.Y(n_17948)
);

OAI22xp5_ASAP7_75t_L g17949 ( 
.A1(n_17578),
.A2(n_9773),
.B1(n_9781),
.B2(n_9776),
.Y(n_17949)
);

NAND2xp5_ASAP7_75t_L g17950 ( 
.A(n_17723),
.B(n_9773),
.Y(n_17950)
);

INVx1_ASAP7_75t_L g17951 ( 
.A(n_17731),
.Y(n_17951)
);

NOR2xp33_ASAP7_75t_L g17952 ( 
.A(n_17765),
.B(n_17766),
.Y(n_17952)
);

AOI22xp5_ASAP7_75t_L g17953 ( 
.A1(n_17715),
.A2(n_9776),
.B1(n_9801),
.B2(n_9781),
.Y(n_17953)
);

INVx2_ASAP7_75t_L g17954 ( 
.A(n_17785),
.Y(n_17954)
);

NAND2xp5_ASAP7_75t_L g17955 ( 
.A(n_17744),
.B(n_9801),
.Y(n_17955)
);

INVx2_ASAP7_75t_L g17956 ( 
.A(n_17670),
.Y(n_17956)
);

OAI22xp5_ASAP7_75t_L g17957 ( 
.A1(n_17588),
.A2(n_9806),
.B1(n_9813),
.B2(n_9809),
.Y(n_17957)
);

NAND2xp5_ASAP7_75t_L g17958 ( 
.A(n_17792),
.B(n_17702),
.Y(n_17958)
);

AND2x2_ASAP7_75t_L g17959 ( 
.A(n_17633),
.B(n_17610),
.Y(n_17959)
);

OAI221xp5_ASAP7_75t_L g17960 ( 
.A1(n_17691),
.A2(n_7942),
.B1(n_8030),
.B2(n_7949),
.C(n_7825),
.Y(n_17960)
);

AOI21xp33_ASAP7_75t_L g17961 ( 
.A1(n_17667),
.A2(n_8012),
.B(n_9806),
.Y(n_17961)
);

OAI21xp5_ASAP7_75t_L g17962 ( 
.A1(n_17624),
.A2(n_7971),
.B(n_7932),
.Y(n_17962)
);

INVx1_ASAP7_75t_L g17963 ( 
.A(n_17776),
.Y(n_17963)
);

INVx1_ASAP7_75t_L g17964 ( 
.A(n_17770),
.Y(n_17964)
);

NAND2xp5_ASAP7_75t_L g17965 ( 
.A(n_17652),
.B(n_9809),
.Y(n_17965)
);

INVx1_ASAP7_75t_L g17966 ( 
.A(n_17779),
.Y(n_17966)
);

INVx1_ASAP7_75t_L g17967 ( 
.A(n_17758),
.Y(n_17967)
);

O2A1O1Ixp33_ASAP7_75t_SL g17968 ( 
.A1(n_17672),
.A2(n_9813),
.B(n_8353),
.C(n_8519),
.Y(n_17968)
);

AOI32xp33_ASAP7_75t_L g17969 ( 
.A1(n_17718),
.A2(n_17598),
.A3(n_17703),
.B1(n_17637),
.B2(n_17659),
.Y(n_17969)
);

NAND2xp5_ASAP7_75t_L g17970 ( 
.A(n_17686),
.B(n_8012),
.Y(n_17970)
);

INVxp67_ASAP7_75t_SL g17971 ( 
.A(n_17657),
.Y(n_17971)
);

INVxp67_ASAP7_75t_L g17972 ( 
.A(n_17630),
.Y(n_17972)
);

INVx1_ASAP7_75t_L g17973 ( 
.A(n_17759),
.Y(n_17973)
);

OR2x2_ASAP7_75t_L g17974 ( 
.A(n_17794),
.B(n_8519),
.Y(n_17974)
);

NAND2xp5_ASAP7_75t_L g17975 ( 
.A(n_17784),
.B(n_8012),
.Y(n_17975)
);

AOI211x1_ASAP7_75t_SL g17976 ( 
.A1(n_17615),
.A2(n_7921),
.B(n_8016),
.C(n_7950),
.Y(n_17976)
);

NAND2xp5_ASAP7_75t_SL g17977 ( 
.A(n_17594),
.B(n_7320),
.Y(n_17977)
);

AOI221x1_ASAP7_75t_L g17978 ( 
.A1(n_17566),
.A2(n_8940),
.B1(n_8916),
.B2(n_8908),
.C(n_8727),
.Y(n_17978)
);

NAND3xp33_ASAP7_75t_L g17979 ( 
.A(n_17586),
.B(n_8016),
.C(n_7322),
.Y(n_17979)
);

INVx1_ASAP7_75t_L g17980 ( 
.A(n_17629),
.Y(n_17980)
);

NOR2xp33_ASAP7_75t_L g17981 ( 
.A(n_17790),
.B(n_8692),
.Y(n_17981)
);

INVx2_ASAP7_75t_L g17982 ( 
.A(n_17673),
.Y(n_17982)
);

INVx1_ASAP7_75t_L g17983 ( 
.A(n_17663),
.Y(n_17983)
);

OR2x2_ASAP7_75t_L g17984 ( 
.A(n_17700),
.B(n_8692),
.Y(n_17984)
);

AOI211xp5_ASAP7_75t_L g17985 ( 
.A1(n_17708),
.A2(n_8231),
.B(n_8593),
.C(n_10275),
.Y(n_17985)
);

INVx1_ASAP7_75t_L g17986 ( 
.A(n_17698),
.Y(n_17986)
);

AOI221xp5_ASAP7_75t_L g17987 ( 
.A1(n_17674),
.A2(n_8401),
.B1(n_8400),
.B2(n_8727),
.C(n_8908),
.Y(n_17987)
);

NAND2xp5_ASAP7_75t_L g17988 ( 
.A(n_17743),
.B(n_8012),
.Y(n_17988)
);

AOI221xp5_ASAP7_75t_L g17989 ( 
.A1(n_17746),
.A2(n_8401),
.B1(n_8400),
.B2(n_8940),
.C(n_8916),
.Y(n_17989)
);

INVx3_ASAP7_75t_L g17990 ( 
.A(n_17711),
.Y(n_17990)
);

OAI22xp5_ASAP7_75t_L g17991 ( 
.A1(n_17592),
.A2(n_7998),
.B1(n_8029),
.B2(n_7966),
.Y(n_17991)
);

INVx2_ASAP7_75t_L g17992 ( 
.A(n_17684),
.Y(n_17992)
);

OAI21xp5_ASAP7_75t_L g17993 ( 
.A1(n_17625),
.A2(n_7730),
.B(n_8231),
.Y(n_17993)
);

INVx1_ASAP7_75t_L g17994 ( 
.A(n_17664),
.Y(n_17994)
);

AOI221xp5_ASAP7_75t_L g17995 ( 
.A1(n_17617),
.A2(n_8401),
.B1(n_8400),
.B2(n_8626),
.C(n_8597),
.Y(n_17995)
);

INVx2_ASAP7_75t_L g17996 ( 
.A(n_17682),
.Y(n_17996)
);

INVxp67_ASAP7_75t_L g17997 ( 
.A(n_17767),
.Y(n_17997)
);

INVx1_ASAP7_75t_L g17998 ( 
.A(n_17753),
.Y(n_17998)
);

AND2x4_ASAP7_75t_L g17999 ( 
.A(n_17651),
.B(n_17749),
.Y(n_17999)
);

INVx1_ASAP7_75t_L g18000 ( 
.A(n_17728),
.Y(n_18000)
);

INVx1_ASAP7_75t_L g18001 ( 
.A(n_17605),
.Y(n_18001)
);

INVx1_ASAP7_75t_L g18002 ( 
.A(n_17771),
.Y(n_18002)
);

INVx1_ASAP7_75t_L g18003 ( 
.A(n_17567),
.Y(n_18003)
);

INVx1_ASAP7_75t_L g18004 ( 
.A(n_17724),
.Y(n_18004)
);

INVx2_ASAP7_75t_SL g18005 ( 
.A(n_17697),
.Y(n_18005)
);

AOI22xp5_ASAP7_75t_SL g18006 ( 
.A1(n_17789),
.A2(n_7384),
.B1(n_8307),
.B2(n_8179),
.Y(n_18006)
);

AOI221xp5_ASAP7_75t_L g18007 ( 
.A1(n_17720),
.A2(n_8651),
.B1(n_8679),
.B2(n_8626),
.C(n_8597),
.Y(n_18007)
);

AOI221xp5_ASAP7_75t_SL g18008 ( 
.A1(n_17626),
.A2(n_7350),
.B1(n_7364),
.B2(n_7322),
.C(n_7320),
.Y(n_18008)
);

NOR2xp33_ASAP7_75t_SL g18009 ( 
.A(n_17773),
.B(n_17775),
.Y(n_18009)
);

AOI22xp33_ASAP7_75t_L g18010 ( 
.A1(n_17754),
.A2(n_7350),
.B1(n_7364),
.B2(n_7320),
.Y(n_18010)
);

INVx1_ASAP7_75t_L g18011 ( 
.A(n_17713),
.Y(n_18011)
);

HB1xp67_ASAP7_75t_L g18012 ( 
.A(n_17623),
.Y(n_18012)
);

AOI211xp5_ASAP7_75t_L g18013 ( 
.A1(n_17634),
.A2(n_8231),
.B(n_7179),
.C(n_7274),
.Y(n_18013)
);

AND2x2_ASAP7_75t_L g18014 ( 
.A(n_17726),
.B(n_8480),
.Y(n_18014)
);

INVx3_ASAP7_75t_SL g18015 ( 
.A(n_17576),
.Y(n_18015)
);

AND2x2_ASAP7_75t_L g18016 ( 
.A(n_17712),
.B(n_8480),
.Y(n_18016)
);

INVx1_ASAP7_75t_L g18017 ( 
.A(n_17707),
.Y(n_18017)
);

INVx1_ASAP7_75t_L g18018 ( 
.A(n_17704),
.Y(n_18018)
);

AOI32xp33_ASAP7_75t_L g18019 ( 
.A1(n_17665),
.A2(n_17681),
.A3(n_17722),
.B1(n_17733),
.B2(n_17687),
.Y(n_18019)
);

INVx1_ASAP7_75t_L g18020 ( 
.A(n_17709),
.Y(n_18020)
);

O2A1O1Ixp33_ASAP7_75t_SL g18021 ( 
.A1(n_17760),
.A2(n_7440),
.B(n_7443),
.C(n_7428),
.Y(n_18021)
);

OR2x2_ASAP7_75t_L g18022 ( 
.A(n_17750),
.B(n_8651),
.Y(n_18022)
);

NAND2xp5_ASAP7_75t_L g18023 ( 
.A(n_17739),
.B(n_8129),
.Y(n_18023)
);

AOI22xp5_ASAP7_75t_L g18024 ( 
.A1(n_17795),
.A2(n_17761),
.B1(n_17635),
.B2(n_17580),
.Y(n_18024)
);

AOI22xp5_ASAP7_75t_L g18025 ( 
.A1(n_17619),
.A2(n_8179),
.B1(n_7440),
.B2(n_7443),
.Y(n_18025)
);

INVx2_ASAP7_75t_SL g18026 ( 
.A(n_17737),
.Y(n_18026)
);

OAI21xp33_ASAP7_75t_L g18027 ( 
.A1(n_17654),
.A2(n_8679),
.B(n_7998),
.Y(n_18027)
);

AOI21xp5_ASAP7_75t_L g18028 ( 
.A1(n_17780),
.A2(n_8453),
.B(n_7730),
.Y(n_18028)
);

O2A1O1Ixp33_ASAP7_75t_L g18029 ( 
.A1(n_17595),
.A2(n_7949),
.B(n_8030),
.C(n_7942),
.Y(n_18029)
);

OR2x2_ASAP7_75t_L g18030 ( 
.A(n_17685),
.B(n_17599),
.Y(n_18030)
);

NAND2xp5_ASAP7_75t_L g18031 ( 
.A(n_17695),
.B(n_8129),
.Y(n_18031)
);

INVx2_ASAP7_75t_L g18032 ( 
.A(n_17569),
.Y(n_18032)
);

HB1xp67_ASAP7_75t_L g18033 ( 
.A(n_17721),
.Y(n_18033)
);

INVx1_ASAP7_75t_L g18034 ( 
.A(n_17542),
.Y(n_18034)
);

AND2x2_ASAP7_75t_L g18035 ( 
.A(n_17530),
.B(n_8480),
.Y(n_18035)
);

NAND2xp5_ASAP7_75t_SL g18036 ( 
.A(n_17556),
.B(n_7320),
.Y(n_18036)
);

INVx1_ASAP7_75t_L g18037 ( 
.A(n_17542),
.Y(n_18037)
);

OAI32xp33_ASAP7_75t_L g18038 ( 
.A1(n_17562),
.A2(n_8030),
.A3(n_7886),
.B1(n_7998),
.B2(n_8029),
.Y(n_18038)
);

INVx1_ASAP7_75t_L g18039 ( 
.A(n_17542),
.Y(n_18039)
);

AND2x2_ASAP7_75t_L g18040 ( 
.A(n_17835),
.B(n_8480),
.Y(n_18040)
);

NAND2x1_ASAP7_75t_SL g18041 ( 
.A(n_17819),
.B(n_7721),
.Y(n_18041)
);

INVx1_ASAP7_75t_L g18042 ( 
.A(n_17905),
.Y(n_18042)
);

NAND2xp5_ASAP7_75t_L g18043 ( 
.A(n_17834),
.B(n_8129),
.Y(n_18043)
);

AOI22xp33_ASAP7_75t_L g18044 ( 
.A1(n_17801),
.A2(n_7364),
.B1(n_7385),
.B2(n_7320),
.Y(n_18044)
);

NAND2xp5_ASAP7_75t_L g18045 ( 
.A(n_17823),
.B(n_8129),
.Y(n_18045)
);

NAND2xp5_ASAP7_75t_L g18046 ( 
.A(n_17799),
.B(n_8129),
.Y(n_18046)
);

INVx2_ASAP7_75t_L g18047 ( 
.A(n_17812),
.Y(n_18047)
);

NOR2xp33_ASAP7_75t_L g18048 ( 
.A(n_17811),
.B(n_7077),
.Y(n_18048)
);

INVx3_ASAP7_75t_SL g18049 ( 
.A(n_17898),
.Y(n_18049)
);

NAND2xp5_ASAP7_75t_L g18050 ( 
.A(n_18034),
.B(n_8149),
.Y(n_18050)
);

INVx1_ASAP7_75t_L g18051 ( 
.A(n_18037),
.Y(n_18051)
);

NAND2xp5_ASAP7_75t_L g18052 ( 
.A(n_18039),
.B(n_8149),
.Y(n_18052)
);

INVx1_ASAP7_75t_L g18053 ( 
.A(n_17806),
.Y(n_18053)
);

INVx2_ASAP7_75t_L g18054 ( 
.A(n_17915),
.Y(n_18054)
);

NOR2xp33_ASAP7_75t_L g18055 ( 
.A(n_17813),
.B(n_17810),
.Y(n_18055)
);

NAND2xp5_ASAP7_75t_L g18056 ( 
.A(n_17829),
.B(n_8149),
.Y(n_18056)
);

NAND2xp5_ASAP7_75t_L g18057 ( 
.A(n_17824),
.B(n_17815),
.Y(n_18057)
);

AND2x2_ASAP7_75t_L g18058 ( 
.A(n_17875),
.B(n_8480),
.Y(n_18058)
);

NAND2x1p5_ASAP7_75t_L g18059 ( 
.A(n_17870),
.B(n_5993),
.Y(n_18059)
);

INVx6_ASAP7_75t_L g18060 ( 
.A(n_17797),
.Y(n_18060)
);

AOI22xp33_ASAP7_75t_L g18061 ( 
.A1(n_17818),
.A2(n_7364),
.B1(n_7385),
.B2(n_7320),
.Y(n_18061)
);

NOR2xp33_ASAP7_75t_L g18062 ( 
.A(n_17918),
.B(n_17848),
.Y(n_18062)
);

NAND2xp5_ASAP7_75t_L g18063 ( 
.A(n_17841),
.B(n_8149),
.Y(n_18063)
);

INVx1_ASAP7_75t_L g18064 ( 
.A(n_17851),
.Y(n_18064)
);

NAND2xp5_ASAP7_75t_L g18065 ( 
.A(n_17883),
.B(n_8149),
.Y(n_18065)
);

AOI222xp33_ASAP7_75t_L g18066 ( 
.A1(n_18000),
.A2(n_7723),
.B1(n_7712),
.B2(n_7818),
.C1(n_7827),
.C2(n_7817),
.Y(n_18066)
);

INVx1_ASAP7_75t_L g18067 ( 
.A(n_17856),
.Y(n_18067)
);

NAND2xp5_ASAP7_75t_L g18068 ( 
.A(n_17879),
.B(n_8453),
.Y(n_18068)
);

INVx1_ASAP7_75t_L g18069 ( 
.A(n_17864),
.Y(n_18069)
);

OR2x2_ASAP7_75t_L g18070 ( 
.A(n_17982),
.B(n_7657),
.Y(n_18070)
);

NAND2xp5_ASAP7_75t_L g18071 ( 
.A(n_17850),
.B(n_8453),
.Y(n_18071)
);

NAND2xp5_ASAP7_75t_L g18072 ( 
.A(n_17980),
.B(n_8453),
.Y(n_18072)
);

OR2x2_ASAP7_75t_L g18073 ( 
.A(n_17906),
.B(n_7657),
.Y(n_18073)
);

INVx1_ASAP7_75t_L g18074 ( 
.A(n_17822),
.Y(n_18074)
);

AND2x2_ASAP7_75t_L g18075 ( 
.A(n_17915),
.B(n_8480),
.Y(n_18075)
);

INVx1_ASAP7_75t_L g18076 ( 
.A(n_17825),
.Y(n_18076)
);

NOR2xp33_ASAP7_75t_L g18077 ( 
.A(n_17867),
.B(n_7077),
.Y(n_18077)
);

INVx1_ASAP7_75t_L g18078 ( 
.A(n_17959),
.Y(n_18078)
);

HB1xp67_ASAP7_75t_L g18079 ( 
.A(n_17868),
.Y(n_18079)
);

NAND2xp33_ASAP7_75t_L g18080 ( 
.A(n_17826),
.B(n_7127),
.Y(n_18080)
);

NAND2xp5_ASAP7_75t_L g18081 ( 
.A(n_17983),
.B(n_8453),
.Y(n_18081)
);

INVxp67_ASAP7_75t_SL g18082 ( 
.A(n_17804),
.Y(n_18082)
);

NOR2xp33_ASAP7_75t_L g18083 ( 
.A(n_17886),
.B(n_7436),
.Y(n_18083)
);

NAND2xp5_ASAP7_75t_L g18084 ( 
.A(n_17971),
.B(n_8240),
.Y(n_18084)
);

INVx1_ASAP7_75t_L g18085 ( 
.A(n_17910),
.Y(n_18085)
);

AND2x2_ASAP7_75t_SL g18086 ( 
.A(n_17803),
.B(n_8862),
.Y(n_18086)
);

AND2x2_ASAP7_75t_L g18087 ( 
.A(n_17838),
.B(n_18035),
.Y(n_18087)
);

BUFx2_ASAP7_75t_L g18088 ( 
.A(n_17859),
.Y(n_18088)
);

OR2x2_ASAP7_75t_L g18089 ( 
.A(n_17814),
.B(n_17805),
.Y(n_18089)
);

OR2x2_ASAP7_75t_L g18090 ( 
.A(n_17974),
.B(n_7657),
.Y(n_18090)
);

OAI22xp5_ASAP7_75t_L g18091 ( 
.A1(n_17938),
.A2(n_17807),
.B1(n_17847),
.B2(n_17857),
.Y(n_18091)
);

AND2x2_ASAP7_75t_L g18092 ( 
.A(n_18015),
.B(n_8480),
.Y(n_18092)
);

NOR2xp33_ASAP7_75t_SL g18093 ( 
.A(n_17832),
.B(n_5676),
.Y(n_18093)
);

OAI21xp5_ASAP7_75t_L g18094 ( 
.A1(n_17854),
.A2(n_7723),
.B(n_7817),
.Y(n_18094)
);

AND2x2_ASAP7_75t_L g18095 ( 
.A(n_17947),
.B(n_8480),
.Y(n_18095)
);

NOR2xp33_ASAP7_75t_SL g18096 ( 
.A(n_17878),
.B(n_5676),
.Y(n_18096)
);

INVx1_ASAP7_75t_L g18097 ( 
.A(n_17800),
.Y(n_18097)
);

OR2x2_ASAP7_75t_L g18098 ( 
.A(n_17865),
.B(n_7657),
.Y(n_18098)
);

NAND2xp5_ASAP7_75t_L g18099 ( 
.A(n_17969),
.B(n_8240),
.Y(n_18099)
);

OR2x2_ASAP7_75t_L g18100 ( 
.A(n_18026),
.B(n_7657),
.Y(n_18100)
);

NAND2x1_ASAP7_75t_SL g18101 ( 
.A(n_17931),
.B(n_7721),
.Y(n_18101)
);

AND2x2_ASAP7_75t_L g18102 ( 
.A(n_17798),
.B(n_8500),
.Y(n_18102)
);

NAND2xp5_ASAP7_75t_L g18103 ( 
.A(n_17820),
.B(n_17871),
.Y(n_18103)
);

INVx1_ASAP7_75t_L g18104 ( 
.A(n_17821),
.Y(n_18104)
);

NAND2xp5_ASAP7_75t_L g18105 ( 
.A(n_17893),
.B(n_8240),
.Y(n_18105)
);

NAND2xp5_ASAP7_75t_L g18106 ( 
.A(n_17896),
.B(n_8240),
.Y(n_18106)
);

NAND2xp5_ASAP7_75t_L g18107 ( 
.A(n_17904),
.B(n_8240),
.Y(n_18107)
);

OA21x2_ASAP7_75t_L g18108 ( 
.A1(n_17817),
.A2(n_10026),
.B(n_10022),
.Y(n_18108)
);

INVx2_ASAP7_75t_L g18109 ( 
.A(n_17846),
.Y(n_18109)
);

INVx1_ASAP7_75t_L g18110 ( 
.A(n_17831),
.Y(n_18110)
);

NAND2xp5_ASAP7_75t_L g18111 ( 
.A(n_17907),
.B(n_8249),
.Y(n_18111)
);

AND2x2_ASAP7_75t_L g18112 ( 
.A(n_17954),
.B(n_8500),
.Y(n_18112)
);

OR2x2_ASAP7_75t_L g18113 ( 
.A(n_17909),
.B(n_7657),
.Y(n_18113)
);

INVx2_ASAP7_75t_SL g18114 ( 
.A(n_18036),
.Y(n_18114)
);

NAND2xp5_ASAP7_75t_L g18115 ( 
.A(n_18033),
.B(n_17986),
.Y(n_18115)
);

HB1xp67_ASAP7_75t_L g18116 ( 
.A(n_17930),
.Y(n_18116)
);

NOR2xp33_ASAP7_75t_L g18117 ( 
.A(n_17946),
.B(n_7436),
.Y(n_18117)
);

INVx1_ASAP7_75t_L g18118 ( 
.A(n_17866),
.Y(n_18118)
);

OAI21xp5_ASAP7_75t_L g18119 ( 
.A1(n_17997),
.A2(n_7723),
.B(n_7817),
.Y(n_18119)
);

INVx1_ASAP7_75t_L g18120 ( 
.A(n_17839),
.Y(n_18120)
);

NOR2x1_ASAP7_75t_L g18121 ( 
.A(n_17956),
.B(n_8249),
.Y(n_18121)
);

INVx1_ASAP7_75t_L g18122 ( 
.A(n_17895),
.Y(n_18122)
);

NOR3xp33_ASAP7_75t_L g18123 ( 
.A(n_17901),
.B(n_5676),
.C(n_6558),
.Y(n_18123)
);

INVx1_ASAP7_75t_SL g18124 ( 
.A(n_17958),
.Y(n_18124)
);

AND2x2_ASAP7_75t_L g18125 ( 
.A(n_17945),
.B(n_17990),
.Y(n_18125)
);

INVxp67_ASAP7_75t_L g18126 ( 
.A(n_17929),
.Y(n_18126)
);

INVx2_ASAP7_75t_L g18127 ( 
.A(n_17940),
.Y(n_18127)
);

INVx1_ASAP7_75t_L g18128 ( 
.A(n_17877),
.Y(n_18128)
);

OR2x2_ASAP7_75t_L g18129 ( 
.A(n_18032),
.B(n_7657),
.Y(n_18129)
);

HB1xp67_ASAP7_75t_L g18130 ( 
.A(n_18001),
.Y(n_18130)
);

NAND2xp5_ASAP7_75t_L g18131 ( 
.A(n_17802),
.B(n_8249),
.Y(n_18131)
);

OR2x2_ASAP7_75t_L g18132 ( 
.A(n_17984),
.B(n_7657),
.Y(n_18132)
);

NAND2xp5_ASAP7_75t_L g18133 ( 
.A(n_18017),
.B(n_8249),
.Y(n_18133)
);

OR2x2_ASAP7_75t_L g18134 ( 
.A(n_17992),
.B(n_8895),
.Y(n_18134)
);

INVx1_ASAP7_75t_L g18135 ( 
.A(n_17920),
.Y(n_18135)
);

NOR2xp33_ASAP7_75t_L g18136 ( 
.A(n_17902),
.B(n_7436),
.Y(n_18136)
);

NAND2xp5_ASAP7_75t_L g18137 ( 
.A(n_17890),
.B(n_8249),
.Y(n_18137)
);

AOI21xp5_ASAP7_75t_L g18138 ( 
.A1(n_17816),
.A2(n_10026),
.B(n_10022),
.Y(n_18138)
);

OAI211xp5_ASAP7_75t_L g18139 ( 
.A1(n_18004),
.A2(n_7721),
.B(n_7991),
.C(n_10022),
.Y(n_18139)
);

NAND2xp5_ASAP7_75t_L g18140 ( 
.A(n_17998),
.B(n_18005),
.Y(n_18140)
);

INVx1_ASAP7_75t_L g18141 ( 
.A(n_17830),
.Y(n_18141)
);

INVx1_ASAP7_75t_L g18142 ( 
.A(n_17849),
.Y(n_18142)
);

NOR2xp33_ASAP7_75t_L g18143 ( 
.A(n_17990),
.B(n_7436),
.Y(n_18143)
);

NOR2xp33_ASAP7_75t_L g18144 ( 
.A(n_17945),
.B(n_7436),
.Y(n_18144)
);

INVx1_ASAP7_75t_L g18145 ( 
.A(n_17827),
.Y(n_18145)
);

NOR2x1_ASAP7_75t_L g18146 ( 
.A(n_17887),
.B(n_17919),
.Y(n_18146)
);

NAND2xp5_ASAP7_75t_SL g18147 ( 
.A(n_17808),
.B(n_7364),
.Y(n_18147)
);

NOR2xp33_ASAP7_75t_L g18148 ( 
.A(n_17951),
.B(n_7436),
.Y(n_18148)
);

NAND2xp5_ASAP7_75t_L g18149 ( 
.A(n_17882),
.B(n_8252),
.Y(n_18149)
);

INVx1_ASAP7_75t_L g18150 ( 
.A(n_17908),
.Y(n_18150)
);

HB1xp67_ASAP7_75t_L g18151 ( 
.A(n_18011),
.Y(n_18151)
);

HB1xp67_ASAP7_75t_L g18152 ( 
.A(n_18012),
.Y(n_18152)
);

NOR2xp33_ASAP7_75t_L g18153 ( 
.A(n_18002),
.B(n_7436),
.Y(n_18153)
);

AOI22xp33_ASAP7_75t_L g18154 ( 
.A1(n_17869),
.A2(n_7385),
.B1(n_7421),
.B2(n_7364),
.Y(n_18154)
);

INVx1_ASAP7_75t_L g18155 ( 
.A(n_17842),
.Y(n_18155)
);

AND2x2_ASAP7_75t_L g18156 ( 
.A(n_17952),
.B(n_17972),
.Y(n_18156)
);

AND2x2_ASAP7_75t_L g18157 ( 
.A(n_17996),
.B(n_8500),
.Y(n_18157)
);

AOI22xp5_ASAP7_75t_L g18158 ( 
.A1(n_18009),
.A2(n_8179),
.B1(n_7440),
.B2(n_7443),
.Y(n_18158)
);

HB1xp67_ASAP7_75t_L g18159 ( 
.A(n_17891),
.Y(n_18159)
);

NAND2xp5_ASAP7_75t_L g18160 ( 
.A(n_17916),
.B(n_8252),
.Y(n_18160)
);

INVx1_ASAP7_75t_SL g18161 ( 
.A(n_17844),
.Y(n_18161)
);

NOR2xp33_ASAP7_75t_L g18162 ( 
.A(n_17912),
.B(n_7497),
.Y(n_18162)
);

OR2x2_ASAP7_75t_L g18163 ( 
.A(n_17840),
.B(n_8895),
.Y(n_18163)
);

AND2x2_ASAP7_75t_L g18164 ( 
.A(n_17914),
.B(n_8500),
.Y(n_18164)
);

NAND2xp5_ASAP7_75t_L g18165 ( 
.A(n_18018),
.B(n_8252),
.Y(n_18165)
);

INVx1_ASAP7_75t_L g18166 ( 
.A(n_17876),
.Y(n_18166)
);

NAND2xp5_ASAP7_75t_L g18167 ( 
.A(n_17994),
.B(n_8252),
.Y(n_18167)
);

INVx1_ASAP7_75t_L g18168 ( 
.A(n_17900),
.Y(n_18168)
);

INVx2_ASAP7_75t_L g18169 ( 
.A(n_17944),
.Y(n_18169)
);

NAND2xp5_ASAP7_75t_L g18170 ( 
.A(n_18024),
.B(n_8252),
.Y(n_18170)
);

AND2x2_ASAP7_75t_L g18171 ( 
.A(n_17925),
.B(n_8500),
.Y(n_18171)
);

INVx2_ASAP7_75t_L g18172 ( 
.A(n_17860),
.Y(n_18172)
);

INVx2_ASAP7_75t_L g18173 ( 
.A(n_17862),
.Y(n_18173)
);

INVx1_ASAP7_75t_L g18174 ( 
.A(n_17899),
.Y(n_18174)
);

INVx2_ASAP7_75t_SL g18175 ( 
.A(n_17863),
.Y(n_18175)
);

AOI22xp5_ASAP7_75t_L g18176 ( 
.A1(n_17881),
.A2(n_8179),
.B1(n_7440),
.B2(n_7469),
.Y(n_18176)
);

NOR2xp33_ASAP7_75t_L g18177 ( 
.A(n_17809),
.B(n_7497),
.Y(n_18177)
);

HB1xp67_ASAP7_75t_L g18178 ( 
.A(n_17999),
.Y(n_18178)
);

OR2x2_ASAP7_75t_L g18179 ( 
.A(n_18003),
.B(n_8895),
.Y(n_18179)
);

INVx2_ASAP7_75t_L g18180 ( 
.A(n_18030),
.Y(n_18180)
);

INVx1_ASAP7_75t_L g18181 ( 
.A(n_17874),
.Y(n_18181)
);

INVx1_ASAP7_75t_L g18182 ( 
.A(n_17937),
.Y(n_18182)
);

NAND2xp5_ASAP7_75t_L g18183 ( 
.A(n_17976),
.B(n_8469),
.Y(n_18183)
);

OAI22xp5_ASAP7_75t_L g18184 ( 
.A1(n_17979),
.A2(n_8029),
.B1(n_7966),
.B2(n_7886),
.Y(n_18184)
);

INVx2_ASAP7_75t_L g18185 ( 
.A(n_18022),
.Y(n_18185)
);

AND2x2_ASAP7_75t_L g18186 ( 
.A(n_17926),
.B(n_8500),
.Y(n_18186)
);

NAND2xp5_ASAP7_75t_L g18187 ( 
.A(n_18020),
.B(n_8469),
.Y(n_18187)
);

INVx1_ASAP7_75t_L g18188 ( 
.A(n_17950),
.Y(n_18188)
);

INVx1_ASAP7_75t_L g18189 ( 
.A(n_17999),
.Y(n_18189)
);

NOR3xp33_ASAP7_75t_L g18190 ( 
.A(n_17967),
.B(n_5676),
.C(n_6558),
.Y(n_18190)
);

INVxp33_ASAP7_75t_L g18191 ( 
.A(n_17939),
.Y(n_18191)
);

NAND2xp5_ASAP7_75t_L g18192 ( 
.A(n_17932),
.B(n_8469),
.Y(n_18192)
);

AOI22xp33_ASAP7_75t_L g18193 ( 
.A1(n_17873),
.A2(n_7385),
.B1(n_7421),
.B2(n_7364),
.Y(n_18193)
);

OR2x2_ASAP7_75t_L g18194 ( 
.A(n_17943),
.B(n_8895),
.Y(n_18194)
);

NOR2x1_ASAP7_75t_L g18195 ( 
.A(n_17933),
.B(n_8469),
.Y(n_18195)
);

AND2x2_ASAP7_75t_L g18196 ( 
.A(n_17973),
.B(n_8500),
.Y(n_18196)
);

NAND2x1_ASAP7_75t_SL g18197 ( 
.A(n_17941),
.B(n_17963),
.Y(n_18197)
);

INVx1_ASAP7_75t_L g18198 ( 
.A(n_17955),
.Y(n_18198)
);

INVx1_ASAP7_75t_L g18199 ( 
.A(n_17922),
.Y(n_18199)
);

INVx1_ASAP7_75t_L g18200 ( 
.A(n_17964),
.Y(n_18200)
);

NAND2xp5_ASAP7_75t_L g18201 ( 
.A(n_17966),
.B(n_8469),
.Y(n_18201)
);

INVx1_ASAP7_75t_L g18202 ( 
.A(n_17965),
.Y(n_18202)
);

AND2x2_ASAP7_75t_L g18203 ( 
.A(n_17981),
.B(n_8500),
.Y(n_18203)
);

OR2x2_ASAP7_75t_L g18204 ( 
.A(n_17903),
.B(n_8895),
.Y(n_18204)
);

NAND2x1_ASAP7_75t_L g18205 ( 
.A(n_17917),
.B(n_7497),
.Y(n_18205)
);

NAND2xp5_ASAP7_75t_L g18206 ( 
.A(n_18019),
.B(n_8485),
.Y(n_18206)
);

AND2x2_ASAP7_75t_L g18207 ( 
.A(n_18016),
.B(n_8836),
.Y(n_18207)
);

NAND2xp5_ASAP7_75t_L g18208 ( 
.A(n_17889),
.B(n_8485),
.Y(n_18208)
);

NOR2xp33_ASAP7_75t_L g18209 ( 
.A(n_17977),
.B(n_7497),
.Y(n_18209)
);

NOR2xp33_ASAP7_75t_L g18210 ( 
.A(n_17843),
.B(n_7497),
.Y(n_18210)
);

AND2x4_ASAP7_75t_L g18211 ( 
.A(n_17942),
.B(n_7912),
.Y(n_18211)
);

INVx1_ASAP7_75t_SL g18212 ( 
.A(n_17975),
.Y(n_18212)
);

NAND2xp5_ASAP7_75t_L g18213 ( 
.A(n_17913),
.B(n_8485),
.Y(n_18213)
);

INVx1_ASAP7_75t_L g18214 ( 
.A(n_17924),
.Y(n_18214)
);

NOR2xp33_ASAP7_75t_L g18215 ( 
.A(n_17884),
.B(n_7497),
.Y(n_18215)
);

INVx1_ASAP7_75t_L g18216 ( 
.A(n_17921),
.Y(n_18216)
);

AND2x2_ASAP7_75t_L g18217 ( 
.A(n_18014),
.B(n_8836),
.Y(n_18217)
);

AND2x2_ASAP7_75t_L g18218 ( 
.A(n_18008),
.B(n_8836),
.Y(n_18218)
);

NAND2xp5_ASAP7_75t_L g18219 ( 
.A(n_18027),
.B(n_8485),
.Y(n_18219)
);

INVx1_ASAP7_75t_L g18220 ( 
.A(n_17968),
.Y(n_18220)
);

NOR2xp33_ASAP7_75t_L g18221 ( 
.A(n_17948),
.B(n_7497),
.Y(n_18221)
);

NAND2xp5_ASAP7_75t_L g18222 ( 
.A(n_17978),
.B(n_8485),
.Y(n_18222)
);

INVx2_ASAP7_75t_L g18223 ( 
.A(n_17970),
.Y(n_18223)
);

INVx1_ASAP7_75t_L g18224 ( 
.A(n_17897),
.Y(n_18224)
);

AND2x2_ASAP7_75t_L g18225 ( 
.A(n_18010),
.B(n_8836),
.Y(n_18225)
);

INVx1_ASAP7_75t_L g18226 ( 
.A(n_18021),
.Y(n_18226)
);

AND2x2_ASAP7_75t_L g18227 ( 
.A(n_17880),
.B(n_8836),
.Y(n_18227)
);

INVx1_ASAP7_75t_L g18228 ( 
.A(n_18023),
.Y(n_18228)
);

INVx1_ASAP7_75t_L g18229 ( 
.A(n_17988),
.Y(n_18229)
);

INVx1_ASAP7_75t_L g18230 ( 
.A(n_17837),
.Y(n_18230)
);

INVx1_ASAP7_75t_L g18231 ( 
.A(n_18031),
.Y(n_18231)
);

NAND2xp5_ASAP7_75t_L g18232 ( 
.A(n_17949),
.B(n_8537),
.Y(n_18232)
);

INVx1_ASAP7_75t_L g18233 ( 
.A(n_17934),
.Y(n_18233)
);

INVx1_ASAP7_75t_L g18234 ( 
.A(n_17828),
.Y(n_18234)
);

NOR2xp33_ASAP7_75t_L g18235 ( 
.A(n_17936),
.B(n_7364),
.Y(n_18235)
);

INVxp33_ASAP7_75t_L g18236 ( 
.A(n_17957),
.Y(n_18236)
);

INVx1_ASAP7_75t_L g18237 ( 
.A(n_17953),
.Y(n_18237)
);

NAND2xp5_ASAP7_75t_L g18238 ( 
.A(n_17833),
.B(n_8537),
.Y(n_18238)
);

INVx1_ASAP7_75t_SL g18239 ( 
.A(n_17961),
.Y(n_18239)
);

INVx2_ASAP7_75t_L g18240 ( 
.A(n_17836),
.Y(n_18240)
);

NAND2xp33_ASAP7_75t_L g18241 ( 
.A(n_17935),
.B(n_7127),
.Y(n_18241)
);

INVx1_ASAP7_75t_L g18242 ( 
.A(n_17927),
.Y(n_18242)
);

INVx1_ASAP7_75t_L g18243 ( 
.A(n_17861),
.Y(n_18243)
);

OR2x2_ASAP7_75t_L g18244 ( 
.A(n_17845),
.B(n_8895),
.Y(n_18244)
);

INVx2_ASAP7_75t_L g18245 ( 
.A(n_17960),
.Y(n_18245)
);

AND2x2_ASAP7_75t_L g18246 ( 
.A(n_17894),
.B(n_8836),
.Y(n_18246)
);

NOR2xp33_ASAP7_75t_L g18247 ( 
.A(n_17872),
.B(n_18038),
.Y(n_18247)
);

NOR2xp33_ASAP7_75t_L g18248 ( 
.A(n_18029),
.B(n_17885),
.Y(n_18248)
);

NAND2x1_ASAP7_75t_SL g18249 ( 
.A(n_18025),
.B(n_18013),
.Y(n_18249)
);

NAND2xp5_ASAP7_75t_L g18250 ( 
.A(n_17923),
.B(n_17985),
.Y(n_18250)
);

OR2x2_ASAP7_75t_L g18251 ( 
.A(n_17991),
.B(n_8895),
.Y(n_18251)
);

OR2x2_ASAP7_75t_L g18252 ( 
.A(n_17993),
.B(n_8895),
.Y(n_18252)
);

NOR2xp33_ASAP7_75t_L g18253 ( 
.A(n_17852),
.B(n_7364),
.Y(n_18253)
);

AOI221xp5_ASAP7_75t_L g18254 ( 
.A1(n_17858),
.A2(n_7422),
.B1(n_7450),
.B2(n_7421),
.C(n_7385),
.Y(n_18254)
);

NAND2x1_ASAP7_75t_SL g18255 ( 
.A(n_18006),
.B(n_7140),
.Y(n_18255)
);

AND2x2_ASAP7_75t_L g18256 ( 
.A(n_18007),
.B(n_8836),
.Y(n_18256)
);

INVx1_ASAP7_75t_L g18257 ( 
.A(n_17911),
.Y(n_18257)
);

NAND2xp5_ASAP7_75t_L g18258 ( 
.A(n_17995),
.B(n_8537),
.Y(n_18258)
);

AND2x2_ASAP7_75t_L g18259 ( 
.A(n_17989),
.B(n_8836),
.Y(n_18259)
);

INVx1_ASAP7_75t_L g18260 ( 
.A(n_18028),
.Y(n_18260)
);

INVx1_ASAP7_75t_L g18261 ( 
.A(n_17855),
.Y(n_18261)
);

NOR2xp33_ASAP7_75t_L g18262 ( 
.A(n_17853),
.B(n_7385),
.Y(n_18262)
);

INVx1_ASAP7_75t_L g18263 ( 
.A(n_17987),
.Y(n_18263)
);

INVx1_ASAP7_75t_L g18264 ( 
.A(n_17892),
.Y(n_18264)
);

INVx1_ASAP7_75t_SL g18265 ( 
.A(n_17928),
.Y(n_18265)
);

NAND2xp5_ASAP7_75t_L g18266 ( 
.A(n_17888),
.B(n_8537),
.Y(n_18266)
);

NOR2xp33_ASAP7_75t_L g18267 ( 
.A(n_17962),
.B(n_7385),
.Y(n_18267)
);

INVx1_ASAP7_75t_L g18268 ( 
.A(n_17835),
.Y(n_18268)
);

INVx1_ASAP7_75t_L g18269 ( 
.A(n_17835),
.Y(n_18269)
);

INVx1_ASAP7_75t_SL g18270 ( 
.A(n_17898),
.Y(n_18270)
);

AND2x2_ASAP7_75t_L g18271 ( 
.A(n_17835),
.B(n_8609),
.Y(n_18271)
);

NOR2xp33_ASAP7_75t_L g18272 ( 
.A(n_17811),
.B(n_7385),
.Y(n_18272)
);

NAND2xp5_ASAP7_75t_L g18273 ( 
.A(n_17835),
.B(n_8537),
.Y(n_18273)
);

NAND2xp5_ASAP7_75t_L g18274 ( 
.A(n_17835),
.B(n_8572),
.Y(n_18274)
);

INVx1_ASAP7_75t_L g18275 ( 
.A(n_17835),
.Y(n_18275)
);

OR2x2_ASAP7_75t_L g18276 ( 
.A(n_17835),
.B(n_7658),
.Y(n_18276)
);

INVx1_ASAP7_75t_L g18277 ( 
.A(n_17835),
.Y(n_18277)
);

NAND2xp5_ASAP7_75t_L g18278 ( 
.A(n_17835),
.B(n_8572),
.Y(n_18278)
);

AND2x2_ASAP7_75t_L g18279 ( 
.A(n_17835),
.B(n_8609),
.Y(n_18279)
);

INVx1_ASAP7_75t_L g18280 ( 
.A(n_17835),
.Y(n_18280)
);

OAI221xp5_ASAP7_75t_L g18281 ( 
.A1(n_17813),
.A2(n_7469),
.B1(n_7428),
.B2(n_7179),
.C(n_7274),
.Y(n_18281)
);

INVxp67_ASAP7_75t_L g18282 ( 
.A(n_17835),
.Y(n_18282)
);

AND2x4_ASAP7_75t_L g18283 ( 
.A(n_17835),
.B(n_7912),
.Y(n_18283)
);

NAND2xp5_ASAP7_75t_L g18284 ( 
.A(n_17835),
.B(n_8572),
.Y(n_18284)
);

NAND2xp5_ASAP7_75t_L g18285 ( 
.A(n_17835),
.B(n_8572),
.Y(n_18285)
);

NAND3x1_ASAP7_75t_L g18286 ( 
.A(n_18146),
.B(n_7588),
.C(n_7587),
.Y(n_18286)
);

CKINVDCx5p33_ASAP7_75t_R g18287 ( 
.A(n_18049),
.Y(n_18287)
);

NAND2xp5_ASAP7_75t_SL g18288 ( 
.A(n_18053),
.B(n_7385),
.Y(n_18288)
);

NAND2xp5_ASAP7_75t_L g18289 ( 
.A(n_18177),
.B(n_8572),
.Y(n_18289)
);

NOR2x1_ASAP7_75t_L g18290 ( 
.A(n_18088),
.B(n_8580),
.Y(n_18290)
);

XNOR2x2_ASAP7_75t_L g18291 ( 
.A(n_18270),
.B(n_7912),
.Y(n_18291)
);

NOR2xp33_ASAP7_75t_L g18292 ( 
.A(n_18060),
.B(n_7421),
.Y(n_18292)
);

INVx1_ASAP7_75t_L g18293 ( 
.A(n_18060),
.Y(n_18293)
);

NAND2xp5_ASAP7_75t_L g18294 ( 
.A(n_18130),
.B(n_8580),
.Y(n_18294)
);

INVx8_ASAP7_75t_L g18295 ( 
.A(n_18156),
.Y(n_18295)
);

AND2x2_ASAP7_75t_L g18296 ( 
.A(n_18047),
.B(n_18069),
.Y(n_18296)
);

INVx1_ASAP7_75t_L g18297 ( 
.A(n_18116),
.Y(n_18297)
);

NAND2xp5_ASAP7_75t_L g18298 ( 
.A(n_18077),
.B(n_8580),
.Y(n_18298)
);

INVx2_ASAP7_75t_L g18299 ( 
.A(n_18059),
.Y(n_18299)
);

AOI22xp5_ASAP7_75t_L g18300 ( 
.A1(n_18055),
.A2(n_8179),
.B1(n_7469),
.B2(n_7428),
.Y(n_18300)
);

INVx2_ASAP7_75t_L g18301 ( 
.A(n_18086),
.Y(n_18301)
);

NAND2xp5_ASAP7_75t_L g18302 ( 
.A(n_18082),
.B(n_18268),
.Y(n_18302)
);

OAI221xp5_ASAP7_75t_L g18303 ( 
.A1(n_18080),
.A2(n_7469),
.B1(n_7179),
.B2(n_7274),
.C(n_7140),
.Y(n_18303)
);

OR2x2_ASAP7_75t_L g18304 ( 
.A(n_18057),
.B(n_7967),
.Y(n_18304)
);

INVx1_ASAP7_75t_L g18305 ( 
.A(n_18079),
.Y(n_18305)
);

NOR2x1_ASAP7_75t_L g18306 ( 
.A(n_18182),
.B(n_8580),
.Y(n_18306)
);

CKINVDCx20_ASAP7_75t_L g18307 ( 
.A(n_18197),
.Y(n_18307)
);

INVx1_ASAP7_75t_L g18308 ( 
.A(n_18178),
.Y(n_18308)
);

INVx1_ASAP7_75t_L g18309 ( 
.A(n_18269),
.Y(n_18309)
);

INVx1_ASAP7_75t_L g18310 ( 
.A(n_18275),
.Y(n_18310)
);

INVx2_ASAP7_75t_L g18311 ( 
.A(n_18277),
.Y(n_18311)
);

HB1xp67_ASAP7_75t_L g18312 ( 
.A(n_18220),
.Y(n_18312)
);

INVx1_ASAP7_75t_L g18313 ( 
.A(n_18280),
.Y(n_18313)
);

NOR3x1_ASAP7_75t_L g18314 ( 
.A(n_18115),
.B(n_7920),
.C(n_7827),
.Y(n_18314)
);

NAND2xp5_ASAP7_75t_L g18315 ( 
.A(n_18215),
.B(n_18083),
.Y(n_18315)
);

NAND2xp5_ASAP7_75t_L g18316 ( 
.A(n_18048),
.B(n_8580),
.Y(n_18316)
);

NAND2xp5_ASAP7_75t_L g18317 ( 
.A(n_18282),
.B(n_7933),
.Y(n_18317)
);

INVx1_ASAP7_75t_L g18318 ( 
.A(n_18151),
.Y(n_18318)
);

INVx1_ASAP7_75t_L g18319 ( 
.A(n_18152),
.Y(n_18319)
);

INVx1_ASAP7_75t_L g18320 ( 
.A(n_18076),
.Y(n_18320)
);

AOI22xp5_ASAP7_75t_L g18321 ( 
.A1(n_18062),
.A2(n_8179),
.B1(n_7561),
.B2(n_7568),
.Y(n_18321)
);

INVx1_ASAP7_75t_L g18322 ( 
.A(n_18103),
.Y(n_18322)
);

INVx1_ASAP7_75t_L g18323 ( 
.A(n_18085),
.Y(n_18323)
);

NAND2xp5_ASAP7_75t_L g18324 ( 
.A(n_18117),
.B(n_7933),
.Y(n_18324)
);

INVxp67_ASAP7_75t_L g18325 ( 
.A(n_18144),
.Y(n_18325)
);

INVx1_ASAP7_75t_L g18326 ( 
.A(n_18078),
.Y(n_18326)
);

INVx1_ASAP7_75t_L g18327 ( 
.A(n_18051),
.Y(n_18327)
);

NAND2xp5_ASAP7_75t_L g18328 ( 
.A(n_18042),
.B(n_7933),
.Y(n_18328)
);

INVx1_ASAP7_75t_L g18329 ( 
.A(n_18089),
.Y(n_18329)
);

AND2x2_ASAP7_75t_L g18330 ( 
.A(n_18153),
.B(n_8609),
.Y(n_18330)
);

AOI21xp5_ASAP7_75t_L g18331 ( 
.A1(n_18140),
.A2(n_6935),
.B(n_6933),
.Y(n_18331)
);

INVxp67_ASAP7_75t_L g18332 ( 
.A(n_18159),
.Y(n_18332)
);

AOI21xp5_ASAP7_75t_L g18333 ( 
.A1(n_18147),
.A2(n_6935),
.B(n_6933),
.Y(n_18333)
);

AND2x2_ASAP7_75t_L g18334 ( 
.A(n_18125),
.B(n_8609),
.Y(n_18334)
);

INVx1_ASAP7_75t_L g18335 ( 
.A(n_18272),
.Y(n_18335)
);

NAND2xp5_ASAP7_75t_SL g18336 ( 
.A(n_18180),
.B(n_7421),
.Y(n_18336)
);

NAND2xp33_ASAP7_75t_SL g18337 ( 
.A(n_18191),
.B(n_7140),
.Y(n_18337)
);

NAND2xp5_ASAP7_75t_L g18338 ( 
.A(n_18175),
.B(n_18143),
.Y(n_18338)
);

AND2x2_ASAP7_75t_L g18339 ( 
.A(n_18148),
.B(n_8609),
.Y(n_18339)
);

NOR4xp25_ASAP7_75t_SL g18340 ( 
.A(n_18216),
.B(n_7560),
.C(n_7582),
.D(n_7539),
.Y(n_18340)
);

INVx1_ASAP7_75t_L g18341 ( 
.A(n_18129),
.Y(n_18341)
);

NAND2x1_ASAP7_75t_L g18342 ( 
.A(n_18214),
.B(n_8069),
.Y(n_18342)
);

INVxp67_ASAP7_75t_L g18343 ( 
.A(n_18093),
.Y(n_18343)
);

INVx1_ASAP7_75t_L g18344 ( 
.A(n_18189),
.Y(n_18344)
);

NOR3xp33_ASAP7_75t_SL g18345 ( 
.A(n_18091),
.B(n_18104),
.C(n_18064),
.Y(n_18345)
);

XOR2x2_ASAP7_75t_L g18346 ( 
.A(n_18136),
.B(n_5993),
.Y(n_18346)
);

NOR3xp33_ASAP7_75t_L g18347 ( 
.A(n_18097),
.B(n_5676),
.C(n_6558),
.Y(n_18347)
);

INVx1_ASAP7_75t_L g18348 ( 
.A(n_18173),
.Y(n_18348)
);

NAND2xp5_ASAP7_75t_L g18349 ( 
.A(n_18209),
.B(n_7933),
.Y(n_18349)
);

NAND2x1_ASAP7_75t_L g18350 ( 
.A(n_18226),
.B(n_8069),
.Y(n_18350)
);

NOR4xp25_ASAP7_75t_SL g18351 ( 
.A(n_18224),
.B(n_7560),
.C(n_7582),
.D(n_7539),
.Y(n_18351)
);

BUFx2_ASAP7_75t_L g18352 ( 
.A(n_18114),
.Y(n_18352)
);

AOI22xp33_ASAP7_75t_SL g18353 ( 
.A1(n_18092),
.A2(n_7384),
.B1(n_7190),
.B2(n_7196),
.Y(n_18353)
);

NAND2xp5_ASAP7_75t_L g18354 ( 
.A(n_18162),
.B(n_7945),
.Y(n_18354)
);

INVx1_ASAP7_75t_L g18355 ( 
.A(n_18100),
.Y(n_18355)
);

NAND3xp33_ASAP7_75t_L g18356 ( 
.A(n_18126),
.B(n_7422),
.C(n_7421),
.Y(n_18356)
);

INVx1_ASAP7_75t_L g18357 ( 
.A(n_18118),
.Y(n_18357)
);

OR2x2_ASAP7_75t_L g18358 ( 
.A(n_18134),
.B(n_7967),
.Y(n_18358)
);

INVx1_ASAP7_75t_SL g18359 ( 
.A(n_18161),
.Y(n_18359)
);

OR2x2_ASAP7_75t_L g18360 ( 
.A(n_18179),
.B(n_7967),
.Y(n_18360)
);

NOR2xp67_ASAP7_75t_SL g18361 ( 
.A(n_18110),
.B(n_18200),
.Y(n_18361)
);

AND2x2_ASAP7_75t_L g18362 ( 
.A(n_18124),
.B(n_8609),
.Y(n_18362)
);

INVx1_ASAP7_75t_L g18363 ( 
.A(n_18109),
.Y(n_18363)
);

INVx1_ASAP7_75t_L g18364 ( 
.A(n_18113),
.Y(n_18364)
);

AOI21xp33_ASAP7_75t_L g18365 ( 
.A1(n_18236),
.A2(n_6806),
.B(n_6729),
.Y(n_18365)
);

AOI22xp5_ASAP7_75t_L g18366 ( 
.A1(n_18210),
.A2(n_18221),
.B1(n_18247),
.B2(n_18262),
.Y(n_18366)
);

INVx2_ASAP7_75t_L g18367 ( 
.A(n_18058),
.Y(n_18367)
);

INVx1_ASAP7_75t_L g18368 ( 
.A(n_18172),
.Y(n_18368)
);

INVx1_ASAP7_75t_L g18369 ( 
.A(n_18067),
.Y(n_18369)
);

INVx1_ASAP7_75t_L g18370 ( 
.A(n_18087),
.Y(n_18370)
);

NAND2xp5_ASAP7_75t_L g18371 ( 
.A(n_18234),
.B(n_7945),
.Y(n_18371)
);

NOR2xp33_ASAP7_75t_L g18372 ( 
.A(n_18127),
.B(n_7421),
.Y(n_18372)
);

NAND2xp5_ASAP7_75t_L g18373 ( 
.A(n_18233),
.B(n_7945),
.Y(n_18373)
);

XOR2x2_ASAP7_75t_L g18374 ( 
.A(n_18249),
.B(n_5993),
.Y(n_18374)
);

INVx1_ASAP7_75t_L g18375 ( 
.A(n_18073),
.Y(n_18375)
);

INVxp67_ASAP7_75t_SL g18376 ( 
.A(n_18240),
.Y(n_18376)
);

INVx1_ASAP7_75t_L g18377 ( 
.A(n_18098),
.Y(n_18377)
);

INVx1_ASAP7_75t_L g18378 ( 
.A(n_18054),
.Y(n_18378)
);

NOR5xp2_ASAP7_75t_L g18379 ( 
.A(n_18074),
.B(n_6342),
.C(n_8006),
.D(n_8109),
.E(n_7967),
.Y(n_18379)
);

XNOR2xp5_ASAP7_75t_L g18380 ( 
.A(n_18263),
.B(n_6225),
.Y(n_18380)
);

NOR2x1_ASAP7_75t_L g18381 ( 
.A(n_18169),
.B(n_18120),
.Y(n_18381)
);

AND2x2_ASAP7_75t_L g18382 ( 
.A(n_18185),
.B(n_8609),
.Y(n_18382)
);

AND2x2_ASAP7_75t_L g18383 ( 
.A(n_18271),
.B(n_8609),
.Y(n_18383)
);

AND2x2_ASAP7_75t_L g18384 ( 
.A(n_18279),
.B(n_8623),
.Y(n_18384)
);

NOR3xp33_ASAP7_75t_SL g18385 ( 
.A(n_18242),
.B(n_18243),
.C(n_18128),
.Y(n_18385)
);

AND2x2_ASAP7_75t_L g18386 ( 
.A(n_18040),
.B(n_8623),
.Y(n_18386)
);

AND2x2_ASAP7_75t_L g18387 ( 
.A(n_18112),
.B(n_8623),
.Y(n_18387)
);

NAND2xp5_ASAP7_75t_L g18388 ( 
.A(n_18122),
.B(n_18265),
.Y(n_18388)
);

AOI21xp5_ASAP7_75t_L g18389 ( 
.A1(n_18250),
.A2(n_6958),
.B(n_7715),
.Y(n_18389)
);

INVx1_ASAP7_75t_L g18390 ( 
.A(n_18230),
.Y(n_18390)
);

INVxp67_ASAP7_75t_SL g18391 ( 
.A(n_18237),
.Y(n_18391)
);

AND2x2_ASAP7_75t_L g18392 ( 
.A(n_18245),
.B(n_8623),
.Y(n_18392)
);

XNOR2xp5_ASAP7_75t_L g18393 ( 
.A(n_18205),
.B(n_6225),
.Y(n_18393)
);

NAND2xp5_ASAP7_75t_L g18394 ( 
.A(n_18239),
.B(n_7945),
.Y(n_18394)
);

INVx1_ASAP7_75t_L g18395 ( 
.A(n_18206),
.Y(n_18395)
);

AND2x4_ASAP7_75t_L g18396 ( 
.A(n_18135),
.B(n_6231),
.Y(n_18396)
);

A2O1A1Ixp33_ASAP7_75t_SL g18397 ( 
.A1(n_18228),
.A2(n_7946),
.B(n_7975),
.C(n_7973),
.Y(n_18397)
);

INVx1_ASAP7_75t_L g18398 ( 
.A(n_18257),
.Y(n_18398)
);

INVx1_ASAP7_75t_L g18399 ( 
.A(n_18261),
.Y(n_18399)
);

NAND2xp5_ASAP7_75t_L g18400 ( 
.A(n_18248),
.B(n_7946),
.Y(n_18400)
);

NAND2xp5_ASAP7_75t_L g18401 ( 
.A(n_18145),
.B(n_18202),
.Y(n_18401)
);

CKINVDCx20_ASAP7_75t_L g18402 ( 
.A(n_18212),
.Y(n_18402)
);

INVx1_ASAP7_75t_L g18403 ( 
.A(n_18070),
.Y(n_18403)
);

INVx1_ASAP7_75t_L g18404 ( 
.A(n_18276),
.Y(n_18404)
);

AND2x2_ASAP7_75t_L g18405 ( 
.A(n_18102),
.B(n_8623),
.Y(n_18405)
);

INVx1_ASAP7_75t_L g18406 ( 
.A(n_18150),
.Y(n_18406)
);

INVx2_ASAP7_75t_L g18407 ( 
.A(n_18132),
.Y(n_18407)
);

AND2x2_ASAP7_75t_L g18408 ( 
.A(n_18095),
.B(n_8623),
.Y(n_18408)
);

XNOR2xp5_ASAP7_75t_L g18409 ( 
.A(n_18188),
.B(n_6231),
.Y(n_18409)
);

NOR2xp33_ASAP7_75t_L g18410 ( 
.A(n_18096),
.B(n_7421),
.Y(n_18410)
);

AND2x2_ASAP7_75t_L g18411 ( 
.A(n_18157),
.B(n_8623),
.Y(n_18411)
);

AND2x2_ASAP7_75t_L g18412 ( 
.A(n_18196),
.B(n_8623),
.Y(n_18412)
);

OR2x2_ASAP7_75t_L g18413 ( 
.A(n_18170),
.B(n_7967),
.Y(n_18413)
);

INVx1_ASAP7_75t_L g18414 ( 
.A(n_18174),
.Y(n_18414)
);

OR2x2_ASAP7_75t_L g18415 ( 
.A(n_18131),
.B(n_7967),
.Y(n_18415)
);

NOR3xp33_ASAP7_75t_SL g18416 ( 
.A(n_18198),
.B(n_6958),
.C(n_7587),
.Y(n_18416)
);

INVx1_ASAP7_75t_L g18417 ( 
.A(n_18155),
.Y(n_18417)
);

NOR3xp33_ASAP7_75t_SL g18418 ( 
.A(n_18199),
.B(n_7588),
.C(n_7445),
.Y(n_18418)
);

INVx1_ASAP7_75t_L g18419 ( 
.A(n_18166),
.Y(n_18419)
);

INVx2_ASAP7_75t_SL g18420 ( 
.A(n_18255),
.Y(n_18420)
);

INVx1_ASAP7_75t_L g18421 ( 
.A(n_18168),
.Y(n_18421)
);

NAND2xp5_ASAP7_75t_L g18422 ( 
.A(n_18141),
.B(n_7946),
.Y(n_18422)
);

INVx1_ASAP7_75t_L g18423 ( 
.A(n_18181),
.Y(n_18423)
);

AND2x2_ASAP7_75t_L g18424 ( 
.A(n_18164),
.B(n_8694),
.Y(n_18424)
);

NAND2xp5_ASAP7_75t_L g18425 ( 
.A(n_18142),
.B(n_7946),
.Y(n_18425)
);

INVx1_ASAP7_75t_L g18426 ( 
.A(n_18264),
.Y(n_18426)
);

BUFx2_ASAP7_75t_L g18427 ( 
.A(n_18133),
.Y(n_18427)
);

NOR4xp25_ASAP7_75t_SL g18428 ( 
.A(n_18260),
.B(n_18231),
.C(n_18229),
.D(n_18254),
.Y(n_18428)
);

INVx1_ASAP7_75t_L g18429 ( 
.A(n_18099),
.Y(n_18429)
);

NOR2x1_ASAP7_75t_L g18430 ( 
.A(n_18223),
.B(n_7061),
.Y(n_18430)
);

NOR3xp33_ASAP7_75t_SL g18431 ( 
.A(n_18138),
.B(n_7445),
.C(n_7444),
.Y(n_18431)
);

AND2x2_ASAP7_75t_L g18432 ( 
.A(n_18171),
.B(n_18186),
.Y(n_18432)
);

INVx1_ASAP7_75t_L g18433 ( 
.A(n_18213),
.Y(n_18433)
);

OR2x2_ASAP7_75t_L g18434 ( 
.A(n_18163),
.B(n_7967),
.Y(n_18434)
);

AOI221xp5_ASAP7_75t_L g18435 ( 
.A1(n_18165),
.A2(n_7450),
.B1(n_7455),
.B2(n_7422),
.C(n_7421),
.Y(n_18435)
);

AND2x2_ASAP7_75t_L g18436 ( 
.A(n_18259),
.B(n_8694),
.Y(n_18436)
);

INVx1_ASAP7_75t_L g18437 ( 
.A(n_18167),
.Y(n_18437)
);

NAND4xp25_ASAP7_75t_L g18438 ( 
.A(n_18043),
.B(n_6699),
.C(n_6713),
.D(n_6558),
.Y(n_18438)
);

NAND2xp5_ASAP7_75t_L g18439 ( 
.A(n_18235),
.B(n_7973),
.Y(n_18439)
);

INVx1_ASAP7_75t_SL g18440 ( 
.A(n_18063),
.Y(n_18440)
);

INVx1_ASAP7_75t_L g18441 ( 
.A(n_18273),
.Y(n_18441)
);

A2O1A1Ixp33_ASAP7_75t_L g18442 ( 
.A1(n_18253),
.A2(n_7920),
.B(n_8932),
.C(n_8928),
.Y(n_18442)
);

AND2x2_ASAP7_75t_L g18443 ( 
.A(n_18075),
.B(n_8694),
.Y(n_18443)
);

AOI21xp5_ASAP7_75t_L g18444 ( 
.A1(n_18241),
.A2(n_7766),
.B(n_7715),
.Y(n_18444)
);

INVx1_ASAP7_75t_L g18445 ( 
.A(n_18274),
.Y(n_18445)
);

BUFx6f_ASAP7_75t_L g18446 ( 
.A(n_18071),
.Y(n_18446)
);

INVx1_ASAP7_75t_L g18447 ( 
.A(n_18278),
.Y(n_18447)
);

INVx1_ASAP7_75t_L g18448 ( 
.A(n_18284),
.Y(n_18448)
);

INVx1_ASAP7_75t_L g18449 ( 
.A(n_18285),
.Y(n_18449)
);

NAND2xp5_ASAP7_75t_SL g18450 ( 
.A(n_18158),
.B(n_7422),
.Y(n_18450)
);

OAI22xp5_ASAP7_75t_L g18451 ( 
.A1(n_18154),
.A2(n_7966),
.B1(n_7886),
.B2(n_8137),
.Y(n_18451)
);

INVx1_ASAP7_75t_L g18452 ( 
.A(n_18105),
.Y(n_18452)
);

HB1xp67_ASAP7_75t_L g18453 ( 
.A(n_18084),
.Y(n_18453)
);

NOR4xp25_ASAP7_75t_L g18454 ( 
.A(n_18106),
.B(n_7975),
.C(n_7982),
.D(n_7973),
.Y(n_18454)
);

NOR2xp33_ASAP7_75t_L g18455 ( 
.A(n_18056),
.B(n_7422),
.Y(n_18455)
);

INVx1_ASAP7_75t_L g18456 ( 
.A(n_18107),
.Y(n_18456)
);

INVx1_ASAP7_75t_L g18457 ( 
.A(n_18111),
.Y(n_18457)
);

INVx2_ASAP7_75t_L g18458 ( 
.A(n_18090),
.Y(n_18458)
);

INVx1_ASAP7_75t_L g18459 ( 
.A(n_18238),
.Y(n_18459)
);

INVx1_ASAP7_75t_L g18460 ( 
.A(n_18068),
.Y(n_18460)
);

NAND2xp33_ASAP7_75t_R g18461 ( 
.A(n_18046),
.B(n_7863),
.Y(n_18461)
);

AOI221xp5_ASAP7_75t_L g18462 ( 
.A1(n_18123),
.A2(n_7455),
.B1(n_7464),
.B2(n_7450),
.C(n_7422),
.Y(n_18462)
);

INVx2_ASAP7_75t_L g18463 ( 
.A(n_18252),
.Y(n_18463)
);

INVx1_ASAP7_75t_L g18464 ( 
.A(n_18065),
.Y(n_18464)
);

INVx1_ASAP7_75t_L g18465 ( 
.A(n_18050),
.Y(n_18465)
);

INVx1_ASAP7_75t_L g18466 ( 
.A(n_18052),
.Y(n_18466)
);

AND2x2_ASAP7_75t_L g18467 ( 
.A(n_18217),
.B(n_18207),
.Y(n_18467)
);

INVx1_ASAP7_75t_L g18468 ( 
.A(n_18045),
.Y(n_18468)
);

AOI22xp5_ASAP7_75t_L g18469 ( 
.A1(n_18190),
.A2(n_7561),
.B1(n_7568),
.B2(n_7515),
.Y(n_18469)
);

INVx1_ASAP7_75t_L g18470 ( 
.A(n_18072),
.Y(n_18470)
);

NAND2xp5_ASAP7_75t_L g18471 ( 
.A(n_18246),
.B(n_7973),
.Y(n_18471)
);

INVx1_ASAP7_75t_L g18472 ( 
.A(n_18081),
.Y(n_18472)
);

INVx1_ASAP7_75t_L g18473 ( 
.A(n_18192),
.Y(n_18473)
);

OAI322xp33_ASAP7_75t_L g18474 ( 
.A1(n_18187),
.A2(n_8150),
.A3(n_8137),
.B1(n_8868),
.B2(n_7568),
.C1(n_7561),
.C2(n_7580),
.Y(n_18474)
);

AND2x2_ASAP7_75t_L g18475 ( 
.A(n_18203),
.B(n_8694),
.Y(n_18475)
);

HAxp5_ASAP7_75t_SL g18476 ( 
.A(n_18176),
.B(n_6729),
.CON(n_18476),
.SN(n_18476)
);

INVx2_ASAP7_75t_L g18477 ( 
.A(n_18251),
.Y(n_18477)
);

OAI21xp33_ASAP7_75t_L g18478 ( 
.A1(n_18267),
.A2(n_18061),
.B(n_18044),
.Y(n_18478)
);

INVx1_ASAP7_75t_L g18479 ( 
.A(n_18201),
.Y(n_18479)
);

AND2x2_ASAP7_75t_L g18480 ( 
.A(n_18256),
.B(n_8694),
.Y(n_18480)
);

NAND2xp5_ASAP7_75t_L g18481 ( 
.A(n_18227),
.B(n_7975),
.Y(n_18481)
);

NOR3xp33_ASAP7_75t_L g18482 ( 
.A(n_18137),
.B(n_6699),
.C(n_6558),
.Y(n_18482)
);

INVx1_ASAP7_75t_L g18483 ( 
.A(n_18204),
.Y(n_18483)
);

NAND2xp5_ASAP7_75t_L g18484 ( 
.A(n_18218),
.B(n_18225),
.Y(n_18484)
);

INVx1_ASAP7_75t_L g18485 ( 
.A(n_18208),
.Y(n_18485)
);

AND2x2_ASAP7_75t_L g18486 ( 
.A(n_18244),
.B(n_8694),
.Y(n_18486)
);

OAI21xp33_ASAP7_75t_L g18487 ( 
.A1(n_18258),
.A2(n_8868),
.B(n_8150),
.Y(n_18487)
);

OAI21xp5_ASAP7_75t_SL g18488 ( 
.A1(n_18194),
.A2(n_7450),
.B(n_7422),
.Y(n_18488)
);

INVx2_ASAP7_75t_L g18489 ( 
.A(n_18041),
.Y(n_18489)
);

NOR2x1_ASAP7_75t_L g18490 ( 
.A(n_18222),
.B(n_7061),
.Y(n_18490)
);

INVx4_ASAP7_75t_SL g18491 ( 
.A(n_18211),
.Y(n_18491)
);

INVx1_ASAP7_75t_L g18492 ( 
.A(n_18160),
.Y(n_18492)
);

NOR2x1p5_ASAP7_75t_L g18493 ( 
.A(n_18183),
.B(n_6231),
.Y(n_18493)
);

OAI22xp5_ASAP7_75t_L g18494 ( 
.A1(n_18287),
.A2(n_18219),
.B1(n_18266),
.B2(n_18149),
.Y(n_18494)
);

INVx1_ASAP7_75t_SL g18495 ( 
.A(n_18295),
.Y(n_18495)
);

NAND2xp5_ASAP7_75t_L g18496 ( 
.A(n_18293),
.B(n_18232),
.Y(n_18496)
);

AOI21xp5_ASAP7_75t_L g18497 ( 
.A1(n_18302),
.A2(n_18195),
.B(n_18094),
.Y(n_18497)
);

INVx2_ASAP7_75t_L g18498 ( 
.A(n_18307),
.Y(n_18498)
);

AOI211xp5_ASAP7_75t_L g18499 ( 
.A1(n_18305),
.A2(n_18281),
.B(n_18184),
.C(n_18211),
.Y(n_18499)
);

NOR2xp33_ASAP7_75t_L g18500 ( 
.A(n_18308),
.B(n_18108),
.Y(n_18500)
);

NOR2xp33_ASAP7_75t_L g18501 ( 
.A(n_18319),
.B(n_18108),
.Y(n_18501)
);

NOR3xp33_ASAP7_75t_L g18502 ( 
.A(n_18326),
.B(n_18121),
.C(n_18139),
.Y(n_18502)
);

AOI21xp5_ASAP7_75t_L g18503 ( 
.A1(n_18295),
.A2(n_18388),
.B(n_18359),
.Y(n_18503)
);

NOR2x1_ASAP7_75t_L g18504 ( 
.A(n_18329),
.B(n_18283),
.Y(n_18504)
);

XOR2xp5_ASAP7_75t_L g18505 ( 
.A(n_18380),
.B(n_18193),
.Y(n_18505)
);

NAND2xp5_ASAP7_75t_L g18506 ( 
.A(n_18312),
.B(n_18101),
.Y(n_18506)
);

AO22x2_ASAP7_75t_L g18507 ( 
.A1(n_18489),
.A2(n_18283),
.B1(n_18119),
.B2(n_18066),
.Y(n_18507)
);

NAND3xp33_ASAP7_75t_L g18508 ( 
.A(n_18345),
.B(n_18361),
.C(n_18385),
.Y(n_18508)
);

INVx2_ASAP7_75t_L g18509 ( 
.A(n_18374),
.Y(n_18509)
);

NAND2xp5_ASAP7_75t_L g18510 ( 
.A(n_18344),
.B(n_7975),
.Y(n_18510)
);

XNOR2x1_ASAP7_75t_L g18511 ( 
.A(n_18296),
.B(n_6344),
.Y(n_18511)
);

NOR2x1_ASAP7_75t_L g18512 ( 
.A(n_18381),
.B(n_6344),
.Y(n_18512)
);

OAI211xp5_ASAP7_75t_SL g18513 ( 
.A1(n_18366),
.A2(n_7776),
.B(n_7766),
.C(n_7444),
.Y(n_18513)
);

NAND2xp5_ASAP7_75t_SL g18514 ( 
.A(n_18430),
.B(n_7422),
.Y(n_18514)
);

OAI21xp5_ASAP7_75t_L g18515 ( 
.A1(n_18332),
.A2(n_7827),
.B(n_7818),
.Y(n_18515)
);

INVx1_ASAP7_75t_L g18516 ( 
.A(n_18491),
.Y(n_18516)
);

INVx2_ASAP7_75t_SL g18517 ( 
.A(n_18396),
.Y(n_18517)
);

NAND2xp5_ASAP7_75t_SL g18518 ( 
.A(n_18311),
.B(n_7422),
.Y(n_18518)
);

AOI21xp5_ASAP7_75t_L g18519 ( 
.A1(n_18376),
.A2(n_7776),
.B(n_7555),
.Y(n_18519)
);

NAND3xp33_ASAP7_75t_L g18520 ( 
.A(n_18318),
.B(n_7455),
.C(n_7450),
.Y(n_18520)
);

INVx1_ASAP7_75t_L g18521 ( 
.A(n_18491),
.Y(n_18521)
);

AO22x2_ASAP7_75t_L g18522 ( 
.A1(n_18320),
.A2(n_18420),
.B1(n_18355),
.B2(n_18370),
.Y(n_18522)
);

NAND2xp5_ASAP7_75t_SL g18523 ( 
.A(n_18297),
.B(n_7450),
.Y(n_18523)
);

AOI211xp5_ASAP7_75t_L g18524 ( 
.A1(n_18309),
.A2(n_7179),
.B(n_7274),
.C(n_7140),
.Y(n_18524)
);

AOI211x1_ASAP7_75t_L g18525 ( 
.A1(n_18288),
.A2(n_7559),
.B(n_7518),
.C(n_6982),
.Y(n_18525)
);

AOI22xp5_ASAP7_75t_L g18526 ( 
.A1(n_18391),
.A2(n_7561),
.B1(n_7568),
.B2(n_7515),
.Y(n_18526)
);

INVx1_ASAP7_75t_L g18527 ( 
.A(n_18352),
.Y(n_18527)
);

AOI211x1_ASAP7_75t_L g18528 ( 
.A1(n_18336),
.A2(n_7559),
.B(n_7518),
.C(n_6982),
.Y(n_18528)
);

AOI21xp5_ASAP7_75t_L g18529 ( 
.A1(n_18338),
.A2(n_7555),
.B(n_7548),
.Y(n_18529)
);

INVx1_ASAP7_75t_L g18530 ( 
.A(n_18409),
.Y(n_18530)
);

NOR2xp33_ASAP7_75t_L g18531 ( 
.A(n_18310),
.B(n_7450),
.Y(n_18531)
);

NAND2xp5_ASAP7_75t_L g18532 ( 
.A(n_18292),
.B(n_7982),
.Y(n_18532)
);

AOI211x1_ASAP7_75t_L g18533 ( 
.A1(n_18365),
.A2(n_6988),
.B(n_7067),
.C(n_7051),
.Y(n_18533)
);

AO22x2_ASAP7_75t_L g18534 ( 
.A1(n_18313),
.A2(n_7990),
.B1(n_8027),
.B2(n_7982),
.Y(n_18534)
);

NOR3xp33_ASAP7_75t_L g18535 ( 
.A(n_18348),
.B(n_7818),
.C(n_6699),
.Y(n_18535)
);

AOI21xp5_ASAP7_75t_L g18536 ( 
.A1(n_18315),
.A2(n_7548),
.B(n_6648),
.Y(n_18536)
);

NAND2xp5_ASAP7_75t_L g18537 ( 
.A(n_18396),
.B(n_7982),
.Y(n_18537)
);

NOR3xp33_ASAP7_75t_L g18538 ( 
.A(n_18368),
.B(n_6699),
.C(n_6558),
.Y(n_18538)
);

INVx1_ASAP7_75t_L g18539 ( 
.A(n_18346),
.Y(n_18539)
);

AOI211xp5_ASAP7_75t_L g18540 ( 
.A1(n_18327),
.A2(n_7274),
.B(n_7179),
.C(n_7920),
.Y(n_18540)
);

NAND2xp5_ASAP7_75t_L g18541 ( 
.A(n_18323),
.B(n_7990),
.Y(n_18541)
);

AOI21xp5_ASAP7_75t_SL g18542 ( 
.A1(n_18299),
.A2(n_6413),
.B(n_6344),
.Y(n_18542)
);

INVx1_ASAP7_75t_L g18543 ( 
.A(n_18490),
.Y(n_18543)
);

AND2x2_ASAP7_75t_L g18544 ( 
.A(n_18357),
.B(n_7967),
.Y(n_18544)
);

NAND2xp5_ASAP7_75t_L g18545 ( 
.A(n_18369),
.B(n_7990),
.Y(n_18545)
);

AOI22xp5_ASAP7_75t_L g18546 ( 
.A1(n_18378),
.A2(n_7580),
.B1(n_7515),
.B2(n_7455),
.Y(n_18546)
);

NAND2xp5_ASAP7_75t_L g18547 ( 
.A(n_18372),
.B(n_7990),
.Y(n_18547)
);

AOI22xp5_ASAP7_75t_L g18548 ( 
.A1(n_18322),
.A2(n_7580),
.B1(n_7515),
.B2(n_7455),
.Y(n_18548)
);

OAI211xp5_ASAP7_75t_SL g18549 ( 
.A1(n_18343),
.A2(n_6648),
.B(n_8150),
.C(n_8137),
.Y(n_18549)
);

OAI21xp5_ASAP7_75t_SL g18550 ( 
.A1(n_18363),
.A2(n_5734),
.B(n_7492),
.Y(n_18550)
);

AOI22xp5_ASAP7_75t_L g18551 ( 
.A1(n_18402),
.A2(n_7580),
.B1(n_7455),
.B2(n_7464),
.Y(n_18551)
);

AOI211xp5_ASAP7_75t_SL g18552 ( 
.A1(n_18398),
.A2(n_7051),
.B(n_7067),
.C(n_6988),
.Y(n_18552)
);

NAND4xp25_ASAP7_75t_L g18553 ( 
.A(n_18399),
.B(n_6713),
.C(n_6727),
.D(n_6699),
.Y(n_18553)
);

OAI211xp5_ASAP7_75t_SL g18554 ( 
.A1(n_18426),
.A2(n_8555),
.B(n_7275),
.C(n_7278),
.Y(n_18554)
);

AOI21xp5_ASAP7_75t_L g18555 ( 
.A1(n_18484),
.A2(n_7275),
.B(n_7253),
.Y(n_18555)
);

INVx2_ASAP7_75t_L g18556 ( 
.A(n_18291),
.Y(n_18556)
);

NAND2xp5_ASAP7_75t_L g18557 ( 
.A(n_18393),
.B(n_8027),
.Y(n_18557)
);

OA22x2_ASAP7_75t_L g18558 ( 
.A1(n_18488),
.A2(n_8032),
.B1(n_8036),
.B2(n_8027),
.Y(n_18558)
);

O2A1O1Ixp33_ASAP7_75t_SL g18559 ( 
.A1(n_18459),
.A2(n_7511),
.B(n_7579),
.C(n_7493),
.Y(n_18559)
);

INVx1_ASAP7_75t_L g18560 ( 
.A(n_18493),
.Y(n_18560)
);

OAI21xp33_ASAP7_75t_SL g18561 ( 
.A1(n_18290),
.A2(n_8577),
.B(n_8080),
.Y(n_18561)
);

AOI21xp33_ASAP7_75t_L g18562 ( 
.A1(n_18483),
.A2(n_6806),
.B(n_6729),
.Y(n_18562)
);

AOI211x1_ASAP7_75t_L g18563 ( 
.A1(n_18478),
.A2(n_7051),
.B(n_7067),
.C(n_7591),
.Y(n_18563)
);

AOI21xp5_ASAP7_75t_L g18564 ( 
.A1(n_18401),
.A2(n_7278),
.B(n_7253),
.Y(n_18564)
);

INVx1_ASAP7_75t_L g18565 ( 
.A(n_18467),
.Y(n_18565)
);

AOI211x1_ASAP7_75t_SL g18566 ( 
.A1(n_18477),
.A2(n_8032),
.B(n_8036),
.C(n_8027),
.Y(n_18566)
);

AOI22xp5_ASAP7_75t_L g18567 ( 
.A1(n_18392),
.A2(n_7455),
.B1(n_7464),
.B2(n_7450),
.Y(n_18567)
);

INVx1_ASAP7_75t_L g18568 ( 
.A(n_18328),
.Y(n_18568)
);

NAND2xp5_ASAP7_75t_L g18569 ( 
.A(n_18390),
.B(n_8032),
.Y(n_18569)
);

INVx1_ASAP7_75t_L g18570 ( 
.A(n_18373),
.Y(n_18570)
);

NAND4xp75_ASAP7_75t_L g18571 ( 
.A(n_18414),
.B(n_7991),
.C(n_8111),
.D(n_8069),
.Y(n_18571)
);

OAI211xp5_ASAP7_75t_SL g18572 ( 
.A1(n_18325),
.A2(n_18406),
.B(n_18419),
.C(n_18417),
.Y(n_18572)
);

AOI21xp5_ASAP7_75t_L g18573 ( 
.A1(n_18400),
.A2(n_7294),
.B(n_7278),
.Y(n_18573)
);

AO22x1_ASAP7_75t_L g18574 ( 
.A1(n_18301),
.A2(n_6729),
.B1(n_6869),
.B2(n_6806),
.Y(n_18574)
);

NOR3xp33_ASAP7_75t_L g18575 ( 
.A(n_18421),
.B(n_6713),
.C(n_6699),
.Y(n_18575)
);

AOI22xp5_ASAP7_75t_L g18576 ( 
.A1(n_18362),
.A2(n_7455),
.B1(n_7464),
.B2(n_7450),
.Y(n_18576)
);

AOI211x1_ASAP7_75t_L g18577 ( 
.A1(n_18450),
.A2(n_7591),
.B(n_7595),
.C(n_6860),
.Y(n_18577)
);

INVx2_ASAP7_75t_L g18578 ( 
.A(n_18342),
.Y(n_18578)
);

NAND2xp5_ASAP7_75t_L g18579 ( 
.A(n_18334),
.B(n_18367),
.Y(n_18579)
);

AND2x2_ASAP7_75t_SL g18580 ( 
.A(n_18423),
.B(n_5734),
.Y(n_18580)
);

OA22x2_ASAP7_75t_L g18581 ( 
.A1(n_18341),
.A2(n_8036),
.B1(n_8037),
.B2(n_8032),
.Y(n_18581)
);

NAND2xp5_ASAP7_75t_L g18582 ( 
.A(n_18432),
.B(n_8036),
.Y(n_18582)
);

AOI22xp5_ASAP7_75t_L g18583 ( 
.A1(n_18382),
.A2(n_18410),
.B1(n_18337),
.B2(n_18455),
.Y(n_18583)
);

OAI211xp5_ASAP7_75t_SL g18584 ( 
.A1(n_18335),
.A2(n_8555),
.B(n_7387),
.C(n_7394),
.Y(n_18584)
);

INVx1_ASAP7_75t_L g18585 ( 
.A(n_18317),
.Y(n_18585)
);

AOI22x1_ASAP7_75t_L g18586 ( 
.A1(n_18427),
.A2(n_5770),
.B1(n_5817),
.B2(n_5695),
.Y(n_18586)
);

OAI21xp5_ASAP7_75t_L g18587 ( 
.A1(n_18394),
.A2(n_7732),
.B(n_7791),
.Y(n_18587)
);

INVx1_ASAP7_75t_L g18588 ( 
.A(n_18371),
.Y(n_18588)
);

NOR2x1_ASAP7_75t_L g18589 ( 
.A(n_18404),
.B(n_6413),
.Y(n_18589)
);

AOI21xp5_ASAP7_75t_L g18590 ( 
.A1(n_18428),
.A2(n_7387),
.B(n_7294),
.Y(n_18590)
);

OA22x2_ASAP7_75t_L g18591 ( 
.A1(n_18463),
.A2(n_18395),
.B1(n_18429),
.B2(n_18294),
.Y(n_18591)
);

AOI21xp33_ASAP7_75t_SL g18592 ( 
.A1(n_18458),
.A2(n_7991),
.B(n_7906),
.Y(n_18592)
);

AOI211x1_ASAP7_75t_L g18593 ( 
.A1(n_18303),
.A2(n_7595),
.B(n_6860),
.C(n_7355),
.Y(n_18593)
);

AO22x1_ASAP7_75t_L g18594 ( 
.A1(n_18364),
.A2(n_6729),
.B1(n_6869),
.B2(n_6806),
.Y(n_18594)
);

INVx1_ASAP7_75t_L g18595 ( 
.A(n_18304),
.Y(n_18595)
);

INVx1_ASAP7_75t_L g18596 ( 
.A(n_18375),
.Y(n_18596)
);

AOI211x1_ASAP7_75t_L g18597 ( 
.A1(n_18356),
.A2(n_7355),
.B(n_7336),
.C(n_6820),
.Y(n_18597)
);

NOR3xp33_ASAP7_75t_L g18598 ( 
.A(n_18377),
.B(n_6727),
.C(n_6713),
.Y(n_18598)
);

AOI21xp5_ASAP7_75t_L g18599 ( 
.A1(n_18433),
.A2(n_7394),
.B(n_7387),
.Y(n_18599)
);

INVx2_ASAP7_75t_L g18600 ( 
.A(n_18286),
.Y(n_18600)
);

AOI21xp5_ASAP7_75t_L g18601 ( 
.A1(n_18440),
.A2(n_7395),
.B(n_7394),
.Y(n_18601)
);

NAND3xp33_ASAP7_75t_L g18602 ( 
.A(n_18407),
.B(n_7464),
.C(n_7455),
.Y(n_18602)
);

NOR2xp33_ASAP7_75t_SL g18603 ( 
.A(n_18403),
.B(n_6413),
.Y(n_18603)
);

AOI211xp5_ASAP7_75t_L g18604 ( 
.A1(n_18492),
.A2(n_7464),
.B(n_8577),
.C(n_7983),
.Y(n_18604)
);

INVx1_ASAP7_75t_L g18605 ( 
.A(n_18453),
.Y(n_18605)
);

OAI22xp5_ASAP7_75t_L g18606 ( 
.A1(n_18353),
.A2(n_8555),
.B1(n_7464),
.B2(n_7365),
.Y(n_18606)
);

AOI22xp33_ASAP7_75t_L g18607 ( 
.A1(n_18347),
.A2(n_7464),
.B1(n_7365),
.B2(n_7369),
.Y(n_18607)
);

INVx2_ASAP7_75t_L g18608 ( 
.A(n_18358),
.Y(n_18608)
);

NAND2xp5_ASAP7_75t_L g18609 ( 
.A(n_18331),
.B(n_8037),
.Y(n_18609)
);

NOR2x1_ASAP7_75t_L g18610 ( 
.A(n_18437),
.B(n_6416),
.Y(n_18610)
);

AOI21xp5_ASAP7_75t_L g18611 ( 
.A1(n_18485),
.A2(n_7447),
.B(n_7395),
.Y(n_18611)
);

NAND4xp75_ASAP7_75t_L g18612 ( 
.A(n_18452),
.B(n_18457),
.C(n_18456),
.D(n_18470),
.Y(n_18612)
);

INVx1_ASAP7_75t_L g18613 ( 
.A(n_18422),
.Y(n_18613)
);

INVx2_ASAP7_75t_SL g18614 ( 
.A(n_18425),
.Y(n_18614)
);

INVx1_ASAP7_75t_L g18615 ( 
.A(n_18446),
.Y(n_18615)
);

NAND2xp5_ASAP7_75t_L g18616 ( 
.A(n_18436),
.B(n_8037),
.Y(n_18616)
);

NOR3x1_ASAP7_75t_L g18617 ( 
.A(n_18472),
.B(n_18445),
.C(n_18441),
.Y(n_18617)
);

INVx1_ASAP7_75t_L g18618 ( 
.A(n_18446),
.Y(n_18618)
);

AOI211xp5_ASAP7_75t_L g18619 ( 
.A1(n_18447),
.A2(n_7464),
.B(n_7983),
.C(n_7961),
.Y(n_18619)
);

INVx1_ASAP7_75t_SL g18620 ( 
.A(n_18415),
.Y(n_18620)
);

NAND2xp5_ASAP7_75t_SL g18621 ( 
.A(n_18482),
.B(n_7127),
.Y(n_18621)
);

AOI21xp5_ASAP7_75t_L g18622 ( 
.A1(n_18448),
.A2(n_7447),
.B(n_7395),
.Y(n_18622)
);

NAND2xp5_ASAP7_75t_L g18623 ( 
.A(n_18431),
.B(n_8037),
.Y(n_18623)
);

OAI21xp33_ASAP7_75t_L g18624 ( 
.A1(n_18438),
.A2(n_7365),
.B(n_7283),
.Y(n_18624)
);

INVx1_ASAP7_75t_L g18625 ( 
.A(n_18446),
.Y(n_18625)
);

AOI22xp5_ASAP7_75t_L g18626 ( 
.A1(n_18480),
.A2(n_8111),
.B1(n_8069),
.B2(n_7583),
.Y(n_18626)
);

AOI22xp5_ASAP7_75t_L g18627 ( 
.A1(n_18461),
.A2(n_8111),
.B1(n_8069),
.B2(n_7583),
.Y(n_18627)
);

INVx1_ASAP7_75t_L g18628 ( 
.A(n_18460),
.Y(n_18628)
);

AO22x1_ASAP7_75t_L g18629 ( 
.A1(n_18449),
.A2(n_6806),
.B1(n_6869),
.B2(n_7015),
.Y(n_18629)
);

AOI22xp33_ASAP7_75t_L g18630 ( 
.A1(n_18487),
.A2(n_7365),
.B1(n_7369),
.B2(n_7283),
.Y(n_18630)
);

NAND3xp33_ASAP7_75t_L g18631 ( 
.A(n_18476),
.B(n_7991),
.C(n_5365),
.Y(n_18631)
);

NAND4xp25_ASAP7_75t_L g18632 ( 
.A(n_18468),
.B(n_6727),
.C(n_6875),
.D(n_6713),
.Y(n_18632)
);

AOI211x1_ASAP7_75t_L g18633 ( 
.A1(n_18289),
.A2(n_7336),
.B(n_6820),
.C(n_6818),
.Y(n_18633)
);

AND2x2_ASAP7_75t_L g18634 ( 
.A(n_18416),
.B(n_8006),
.Y(n_18634)
);

OAI21xp5_ASAP7_75t_SL g18635 ( 
.A1(n_18471),
.A2(n_7516),
.B(n_7492),
.Y(n_18635)
);

OAI21xp33_ASAP7_75t_L g18636 ( 
.A1(n_18413),
.A2(n_7369),
.B(n_7283),
.Y(n_18636)
);

INVx1_ASAP7_75t_L g18637 ( 
.A(n_18465),
.Y(n_18637)
);

INVx1_ASAP7_75t_L g18638 ( 
.A(n_18466),
.Y(n_18638)
);

OAI22xp5_ASAP7_75t_L g18639 ( 
.A1(n_18435),
.A2(n_7369),
.B1(n_7370),
.B2(n_7283),
.Y(n_18639)
);

NAND2xp5_ASAP7_75t_SL g18640 ( 
.A(n_18462),
.B(n_18454),
.Y(n_18640)
);

OAI21xp5_ASAP7_75t_L g18641 ( 
.A1(n_18349),
.A2(n_7732),
.B(n_7791),
.Y(n_18641)
);

AND2x2_ASAP7_75t_L g18642 ( 
.A(n_18418),
.B(n_8006),
.Y(n_18642)
);

OAI21xp5_ASAP7_75t_L g18643 ( 
.A1(n_18354),
.A2(n_7732),
.B(n_7791),
.Y(n_18643)
);

AOI21xp5_ASAP7_75t_L g18644 ( 
.A1(n_18473),
.A2(n_7471),
.B(n_7447),
.Y(n_18644)
);

INVx1_ASAP7_75t_L g18645 ( 
.A(n_18464),
.Y(n_18645)
);

NOR2x1_ASAP7_75t_L g18646 ( 
.A(n_18479),
.B(n_6416),
.Y(n_18646)
);

AND3x1_ASAP7_75t_L g18647 ( 
.A(n_18340),
.B(n_18351),
.C(n_18324),
.Y(n_18647)
);

NOR3x1_ASAP7_75t_L g18648 ( 
.A(n_18298),
.B(n_7983),
.C(n_7961),
.Y(n_18648)
);

AND2x2_ASAP7_75t_L g18649 ( 
.A(n_18330),
.B(n_8006),
.Y(n_18649)
);

NOR2xp33_ASAP7_75t_L g18650 ( 
.A(n_18481),
.B(n_6940),
.Y(n_18650)
);

NAND4xp75_ASAP7_75t_SL g18651 ( 
.A(n_18486),
.B(n_18411),
.C(n_18339),
.D(n_18408),
.Y(n_18651)
);

NAND2xp5_ASAP7_75t_L g18652 ( 
.A(n_18412),
.B(n_8038),
.Y(n_18652)
);

AOI22xp33_ASAP7_75t_L g18653 ( 
.A1(n_18387),
.A2(n_7378),
.B1(n_7386),
.B2(n_7370),
.Y(n_18653)
);

BUFx2_ASAP7_75t_L g18654 ( 
.A(n_18439),
.Y(n_18654)
);

INVx1_ASAP7_75t_L g18655 ( 
.A(n_18316),
.Y(n_18655)
);

OAI21xp33_ASAP7_75t_L g18656 ( 
.A1(n_18443),
.A2(n_7378),
.B(n_7370),
.Y(n_18656)
);

NOR2x1_ASAP7_75t_L g18657 ( 
.A(n_18360),
.B(n_6416),
.Y(n_18657)
);

NAND2xp5_ASAP7_75t_L g18658 ( 
.A(n_18424),
.B(n_18383),
.Y(n_18658)
);

INVx1_ASAP7_75t_L g18659 ( 
.A(n_18434),
.Y(n_18659)
);

NOR2xp33_ASAP7_75t_L g18660 ( 
.A(n_18384),
.B(n_6940),
.Y(n_18660)
);

NAND2xp5_ASAP7_75t_L g18661 ( 
.A(n_18386),
.B(n_8038),
.Y(n_18661)
);

OAI22xp5_ASAP7_75t_L g18662 ( 
.A1(n_18469),
.A2(n_7378),
.B1(n_7386),
.B2(n_7370),
.Y(n_18662)
);

NOR2xp33_ASAP7_75t_L g18663 ( 
.A(n_18405),
.B(n_6945),
.Y(n_18663)
);

NOR3xp33_ASAP7_75t_L g18664 ( 
.A(n_18389),
.B(n_6727),
.C(n_6713),
.Y(n_18664)
);

NAND2xp5_ASAP7_75t_SL g18665 ( 
.A(n_18475),
.B(n_7127),
.Y(n_18665)
);

NAND2xp5_ASAP7_75t_SL g18666 ( 
.A(n_18306),
.B(n_18333),
.Y(n_18666)
);

NAND2xp5_ASAP7_75t_L g18667 ( 
.A(n_18397),
.B(n_8038),
.Y(n_18667)
);

XNOR2x1_ASAP7_75t_SL g18668 ( 
.A(n_18350),
.B(n_5374),
.Y(n_18668)
);

NOR3xp33_ASAP7_75t_L g18669 ( 
.A(n_18474),
.B(n_6875),
.C(n_6727),
.Y(n_18669)
);

AOI22xp5_ASAP7_75t_L g18670 ( 
.A1(n_18451),
.A2(n_8111),
.B1(n_8069),
.B2(n_7583),
.Y(n_18670)
);

AO22x2_ASAP7_75t_L g18671 ( 
.A1(n_18444),
.A2(n_8041),
.B1(n_8056),
.B2(n_8038),
.Y(n_18671)
);

NOR3xp33_ASAP7_75t_L g18672 ( 
.A(n_18442),
.B(n_6875),
.C(n_6727),
.Y(n_18672)
);

OAI21xp5_ASAP7_75t_L g18673 ( 
.A1(n_18503),
.A2(n_18300),
.B(n_18321),
.Y(n_18673)
);

AOI22xp5_ASAP7_75t_L g18674 ( 
.A1(n_18527),
.A2(n_18314),
.B1(n_18379),
.B2(n_8111),
.Y(n_18674)
);

NAND2xp33_ASAP7_75t_SL g18675 ( 
.A(n_18498),
.B(n_7190),
.Y(n_18675)
);

INVx2_ASAP7_75t_SL g18676 ( 
.A(n_18512),
.Y(n_18676)
);

OAI22xp5_ASAP7_75t_L g18677 ( 
.A1(n_18508),
.A2(n_18495),
.B1(n_18631),
.B2(n_18565),
.Y(n_18677)
);

OR2x2_ASAP7_75t_L g18678 ( 
.A(n_18506),
.B(n_8006),
.Y(n_18678)
);

INVx1_ASAP7_75t_L g18679 ( 
.A(n_18516),
.Y(n_18679)
);

AOI21xp33_ASAP7_75t_L g18680 ( 
.A1(n_18521),
.A2(n_18504),
.B(n_18596),
.Y(n_18680)
);

INVx1_ASAP7_75t_L g18681 ( 
.A(n_18511),
.Y(n_18681)
);

CKINVDCx5p33_ASAP7_75t_R g18682 ( 
.A(n_18509),
.Y(n_18682)
);

OA21x2_ASAP7_75t_L g18683 ( 
.A1(n_18556),
.A2(n_7807),
.B(n_7801),
.Y(n_18683)
);

NAND5xp2_ASAP7_75t_L g18684 ( 
.A(n_18499),
.B(n_7419),
.C(n_7454),
.D(n_7401),
.E(n_7390),
.Y(n_18684)
);

OAI21xp33_ASAP7_75t_L g18685 ( 
.A1(n_18603),
.A2(n_7386),
.B(n_7378),
.Y(n_18685)
);

XNOR2xp5_ASAP7_75t_L g18686 ( 
.A(n_18505),
.B(n_6506),
.Y(n_18686)
);

OAI22x1_ASAP7_75t_L g18687 ( 
.A1(n_18517),
.A2(n_8307),
.B1(n_8111),
.B2(n_8304),
.Y(n_18687)
);

INVxp33_ASAP7_75t_L g18688 ( 
.A(n_18579),
.Y(n_18688)
);

INVx1_ASAP7_75t_L g18689 ( 
.A(n_18522),
.Y(n_18689)
);

AOI221x1_ASAP7_75t_L g18690 ( 
.A1(n_18572),
.A2(n_18522),
.B1(n_18500),
.B2(n_18502),
.C(n_18501),
.Y(n_18690)
);

OAI221xp5_ASAP7_75t_L g18691 ( 
.A1(n_18636),
.A2(n_8031),
.B1(n_8238),
.B2(n_8148),
.C(n_8002),
.Y(n_18691)
);

INVx1_ASAP7_75t_L g18692 ( 
.A(n_18589),
.Y(n_18692)
);

NAND2x1p5_ASAP7_75t_L g18693 ( 
.A(n_18543),
.B(n_6506),
.Y(n_18693)
);

AOI221x1_ASAP7_75t_L g18694 ( 
.A1(n_18497),
.A2(n_18494),
.B1(n_18615),
.B2(n_18625),
.C(n_18618),
.Y(n_18694)
);

OAI311xp33_ASAP7_75t_L g18695 ( 
.A1(n_18583),
.A2(n_6820),
.A3(n_6818),
.B1(n_7151),
.C1(n_7136),
.Y(n_18695)
);

AOI21xp5_ASAP7_75t_L g18696 ( 
.A1(n_18578),
.A2(n_7534),
.B(n_7471),
.Y(n_18696)
);

AOI322xp5_ASAP7_75t_L g18697 ( 
.A1(n_18531),
.A2(n_7585),
.A3(n_7511),
.B1(n_7592),
.B2(n_7579),
.C1(n_7493),
.C2(n_7257),
.Y(n_18697)
);

BUFx2_ASAP7_75t_L g18698 ( 
.A(n_18647),
.Y(n_18698)
);

OA21x2_ASAP7_75t_L g18699 ( 
.A1(n_18659),
.A2(n_7807),
.B(n_7801),
.Y(n_18699)
);

INVx1_ASAP7_75t_L g18700 ( 
.A(n_18668),
.Y(n_18700)
);

AOI22xp5_ASAP7_75t_L g18701 ( 
.A1(n_18605),
.A2(n_7582),
.B1(n_7191),
.B2(n_7242),
.Y(n_18701)
);

AOI222xp33_ASAP7_75t_L g18702 ( 
.A1(n_18523),
.A2(n_7530),
.B1(n_7516),
.B2(n_7538),
.C1(n_7525),
.C2(n_7492),
.Y(n_18702)
);

INVx1_ASAP7_75t_L g18703 ( 
.A(n_18610),
.Y(n_18703)
);

AOI22xp5_ASAP7_75t_L g18704 ( 
.A1(n_18530),
.A2(n_7191),
.B1(n_7242),
.B2(n_7202),
.Y(n_18704)
);

AOI21xp5_ASAP7_75t_L g18705 ( 
.A1(n_18666),
.A2(n_7534),
.B(n_7471),
.Y(n_18705)
);

INVx1_ASAP7_75t_SL g18706 ( 
.A(n_18651),
.Y(n_18706)
);

BUFx10_ASAP7_75t_L g18707 ( 
.A(n_18628),
.Y(n_18707)
);

AOI22xp5_ASAP7_75t_L g18708 ( 
.A1(n_18539),
.A2(n_7191),
.B1(n_7242),
.B2(n_7202),
.Y(n_18708)
);

OAI22xp33_ASAP7_75t_SL g18709 ( 
.A1(n_18514),
.A2(n_8056),
.B1(n_8059),
.B2(n_8041),
.Y(n_18709)
);

AOI221xp5_ASAP7_75t_L g18710 ( 
.A1(n_18559),
.A2(n_8059),
.B1(n_8062),
.B2(n_8056),
.C(n_8041),
.Y(n_18710)
);

O2A1O1Ixp33_ASAP7_75t_L g18711 ( 
.A1(n_18496),
.A2(n_18608),
.B(n_18638),
.C(n_18637),
.Y(n_18711)
);

INVx2_ASAP7_75t_L g18712 ( 
.A(n_18580),
.Y(n_18712)
);

INVxp67_ASAP7_75t_L g18713 ( 
.A(n_18658),
.Y(n_18713)
);

AOI221xp5_ASAP7_75t_L g18714 ( 
.A1(n_18562),
.A2(n_8059),
.B1(n_8062),
.B2(n_8056),
.C(n_8041),
.Y(n_18714)
);

NAND2xp5_ASAP7_75t_L g18715 ( 
.A(n_18646),
.B(n_8059),
.Y(n_18715)
);

AOI222xp33_ASAP7_75t_L g18716 ( 
.A1(n_18518),
.A2(n_7530),
.B1(n_7516),
.B2(n_7538),
.C1(n_7525),
.C2(n_7492),
.Y(n_18716)
);

AOI322xp5_ASAP7_75t_L g18717 ( 
.A1(n_18620),
.A2(n_7585),
.A3(n_7511),
.B1(n_7592),
.B2(n_7579),
.C1(n_7493),
.C2(n_7260),
.Y(n_18717)
);

INVxp67_ASAP7_75t_L g18718 ( 
.A(n_18654),
.Y(n_18718)
);

INVx2_ASAP7_75t_L g18719 ( 
.A(n_18544),
.Y(n_18719)
);

INVx1_ASAP7_75t_L g18720 ( 
.A(n_18510),
.Y(n_18720)
);

OAI22xp5_ASAP7_75t_L g18721 ( 
.A1(n_18520),
.A2(n_8073),
.B1(n_8074),
.B2(n_8062),
.Y(n_18721)
);

AOI221xp5_ASAP7_75t_L g18722 ( 
.A1(n_18560),
.A2(n_8074),
.B1(n_8077),
.B2(n_8073),
.C(n_8062),
.Y(n_18722)
);

AND2x2_ASAP7_75t_L g18723 ( 
.A(n_18600),
.B(n_8006),
.Y(n_18723)
);

AOI21xp5_ASAP7_75t_L g18724 ( 
.A1(n_18507),
.A2(n_7535),
.B(n_7534),
.Y(n_18724)
);

INVx1_ASAP7_75t_L g18725 ( 
.A(n_18541),
.Y(n_18725)
);

NOR4xp25_ASAP7_75t_L g18726 ( 
.A(n_18645),
.B(n_8074),
.C(n_8077),
.D(n_8073),
.Y(n_18726)
);

INVx2_ASAP7_75t_L g18727 ( 
.A(n_18581),
.Y(n_18727)
);

OAI211xp5_ASAP7_75t_SL g18728 ( 
.A1(n_18595),
.A2(n_7535),
.B(n_7136),
.C(n_7155),
.Y(n_18728)
);

CKINVDCx20_ASAP7_75t_R g18729 ( 
.A(n_18614),
.Y(n_18729)
);

INVx1_ASAP7_75t_L g18730 ( 
.A(n_18545),
.Y(n_18730)
);

INVx1_ASAP7_75t_L g18731 ( 
.A(n_18569),
.Y(n_18731)
);

OAI21xp5_ASAP7_75t_SL g18732 ( 
.A1(n_18570),
.A2(n_7516),
.B(n_7492),
.Y(n_18732)
);

OAI31xp33_ASAP7_75t_SL g18733 ( 
.A1(n_18657),
.A2(n_7712),
.A3(n_7903),
.B(n_7899),
.Y(n_18733)
);

NAND2xp5_ASAP7_75t_L g18734 ( 
.A(n_18588),
.B(n_8073),
.Y(n_18734)
);

NOR3xp33_ASAP7_75t_SL g18735 ( 
.A(n_18612),
.B(n_7535),
.C(n_6818),
.Y(n_18735)
);

NOR4xp25_ASAP7_75t_L g18736 ( 
.A(n_18568),
.B(n_8077),
.C(n_8087),
.D(n_8074),
.Y(n_18736)
);

AOI222xp33_ASAP7_75t_L g18737 ( 
.A1(n_18640),
.A2(n_7530),
.B1(n_7516),
.B2(n_7538),
.C1(n_7525),
.C2(n_7492),
.Y(n_18737)
);

NAND2xp5_ASAP7_75t_L g18738 ( 
.A(n_18613),
.B(n_18585),
.Y(n_18738)
);

AOI22xp33_ASAP7_75t_L g18739 ( 
.A1(n_18538),
.A2(n_7403),
.B1(n_7412),
.B2(n_7386),
.Y(n_18739)
);

INVx1_ASAP7_75t_L g18740 ( 
.A(n_18507),
.Y(n_18740)
);

O2A1O1Ixp33_ASAP7_75t_L g18741 ( 
.A1(n_18655),
.A2(n_6506),
.B(n_8031),
.C(n_8002),
.Y(n_18741)
);

HB1xp67_ASAP7_75t_L g18742 ( 
.A(n_18591),
.Y(n_18742)
);

INVx3_ASAP7_75t_L g18743 ( 
.A(n_18558),
.Y(n_18743)
);

NAND4xp25_ASAP7_75t_L g18744 ( 
.A(n_18617),
.B(n_6878),
.C(n_6895),
.D(n_6875),
.Y(n_18744)
);

INVx1_ASAP7_75t_L g18745 ( 
.A(n_18582),
.Y(n_18745)
);

NAND2xp5_ASAP7_75t_L g18746 ( 
.A(n_18660),
.B(n_8077),
.Y(n_18746)
);

NOR2x1_ASAP7_75t_L g18747 ( 
.A(n_18542),
.B(n_7061),
.Y(n_18747)
);

NAND2xp5_ASAP7_75t_L g18748 ( 
.A(n_18663),
.B(n_8087),
.Y(n_18748)
);

INVx1_ASAP7_75t_L g18749 ( 
.A(n_18557),
.Y(n_18749)
);

AOI211xp5_ASAP7_75t_SL g18750 ( 
.A1(n_18656),
.A2(n_6896),
.B(n_6937),
.C(n_6885),
.Y(n_18750)
);

BUFx3_ASAP7_75t_L g18751 ( 
.A(n_18650),
.Y(n_18751)
);

AOI21xp5_ASAP7_75t_L g18752 ( 
.A1(n_18621),
.A2(n_7807),
.B(n_7801),
.Y(n_18752)
);

OR2x2_ASAP7_75t_L g18753 ( 
.A(n_18623),
.B(n_8006),
.Y(n_18753)
);

INVx1_ASAP7_75t_L g18754 ( 
.A(n_18616),
.Y(n_18754)
);

AOI211xp5_ASAP7_75t_L g18755 ( 
.A1(n_18602),
.A2(n_8932),
.B(n_8951),
.C(n_8928),
.Y(n_18755)
);

INVxp67_ASAP7_75t_L g18756 ( 
.A(n_18665),
.Y(n_18756)
);

AOI221xp5_ASAP7_75t_L g18757 ( 
.A1(n_18669),
.A2(n_8090),
.B1(n_8095),
.B2(n_8089),
.C(n_8087),
.Y(n_18757)
);

OAI22xp33_ASAP7_75t_L g18758 ( 
.A1(n_18551),
.A2(n_7196),
.B1(n_7199),
.B2(n_7190),
.Y(n_18758)
);

AOI21xp5_ASAP7_75t_SL g18759 ( 
.A1(n_18590),
.A2(n_7991),
.B(n_7906),
.Y(n_18759)
);

AOI31xp33_ASAP7_75t_L g18760 ( 
.A1(n_18652),
.A2(n_7413),
.A3(n_7482),
.B(n_7398),
.Y(n_18760)
);

OA22x2_ASAP7_75t_L g18761 ( 
.A1(n_18550),
.A2(n_18635),
.B1(n_18661),
.B2(n_18537),
.Y(n_18761)
);

OAI21xp33_ASAP7_75t_L g18762 ( 
.A1(n_18624),
.A2(n_7412),
.B(n_7403),
.Y(n_18762)
);

AOI21xp5_ASAP7_75t_L g18763 ( 
.A1(n_18574),
.A2(n_7745),
.B(n_7741),
.Y(n_18763)
);

OAI21xp5_ASAP7_75t_SL g18764 ( 
.A1(n_18566),
.A2(n_7516),
.B(n_7492),
.Y(n_18764)
);

AOI22xp33_ASAP7_75t_L g18765 ( 
.A1(n_18598),
.A2(n_7412),
.B1(n_7430),
.B2(n_7403),
.Y(n_18765)
);

INVx1_ASAP7_75t_L g18766 ( 
.A(n_18667),
.Y(n_18766)
);

OAI31xp33_ASAP7_75t_L g18767 ( 
.A1(n_18642),
.A2(n_7028),
.A3(n_7082),
.B(n_7403),
.Y(n_18767)
);

OAI322xp33_ASAP7_75t_L g18768 ( 
.A1(n_18547),
.A2(n_8095),
.A3(n_8089),
.B1(n_8103),
.B2(n_8127),
.C1(n_8090),
.C2(n_8087),
.Y(n_18768)
);

INVx2_ASAP7_75t_L g18769 ( 
.A(n_18532),
.Y(n_18769)
);

XNOR2x1_ASAP7_75t_L g18770 ( 
.A(n_18594),
.B(n_8002),
.Y(n_18770)
);

NAND2xp5_ASAP7_75t_L g18771 ( 
.A(n_18533),
.B(n_8089),
.Y(n_18771)
);

INVx2_ASAP7_75t_L g18772 ( 
.A(n_18671),
.Y(n_18772)
);

AOI22xp33_ASAP7_75t_L g18773 ( 
.A1(n_18575),
.A2(n_7430),
.B1(n_7438),
.B2(n_7412),
.Y(n_18773)
);

HB1xp67_ASAP7_75t_L g18774 ( 
.A(n_18634),
.Y(n_18774)
);

OAI21xp33_ASAP7_75t_SL g18775 ( 
.A1(n_18553),
.A2(n_8080),
.B(n_8079),
.Y(n_18775)
);

AOI22xp5_ASAP7_75t_L g18776 ( 
.A1(n_18664),
.A2(n_18672),
.B1(n_18632),
.B2(n_18649),
.Y(n_18776)
);

INVx1_ASAP7_75t_SL g18777 ( 
.A(n_18609),
.Y(n_18777)
);

O2A1O1Ixp33_ASAP7_75t_L g18778 ( 
.A1(n_18662),
.A2(n_8031),
.B(n_8148),
.C(n_8002),
.Y(n_18778)
);

OAI21xp5_ASAP7_75t_L g18779 ( 
.A1(n_18519),
.A2(n_7645),
.B(n_7644),
.Y(n_18779)
);

INVx2_ASAP7_75t_SL g18780 ( 
.A(n_18671),
.Y(n_18780)
);

XNOR2x1_ASAP7_75t_L g18781 ( 
.A(n_18629),
.B(n_8002),
.Y(n_18781)
);

AOI22xp5_ASAP7_75t_SL g18782 ( 
.A1(n_18606),
.A2(n_7991),
.B1(n_8307),
.B2(n_7196),
.Y(n_18782)
);

AOI21xp5_ASAP7_75t_L g18783 ( 
.A1(n_18564),
.A2(n_7745),
.B(n_7741),
.Y(n_18783)
);

AOI21xp33_ASAP7_75t_L g18784 ( 
.A1(n_18586),
.A2(n_6869),
.B(n_6806),
.Y(n_18784)
);

OAI21xp5_ASAP7_75t_L g18785 ( 
.A1(n_18599),
.A2(n_7645),
.B(n_7644),
.Y(n_18785)
);

INVx2_ASAP7_75t_L g18786 ( 
.A(n_18633),
.Y(n_18786)
);

OAI21xp5_ASAP7_75t_L g18787 ( 
.A1(n_18555),
.A2(n_7645),
.B(n_7644),
.Y(n_18787)
);

AOI211xp5_ASAP7_75t_SL g18788 ( 
.A1(n_18548),
.A2(n_6896),
.B(n_6937),
.C(n_6885),
.Y(n_18788)
);

INVx1_ASAP7_75t_L g18789 ( 
.A(n_18577),
.Y(n_18789)
);

AOI31xp33_ASAP7_75t_L g18790 ( 
.A1(n_18552),
.A2(n_7398),
.A3(n_7482),
.B(n_7413),
.Y(n_18790)
);

NAND2xp5_ASAP7_75t_L g18791 ( 
.A(n_18593),
.B(n_8089),
.Y(n_18791)
);

AOI22xp5_ASAP7_75t_L g18792 ( 
.A1(n_18546),
.A2(n_7242),
.B1(n_7252),
.B2(n_7202),
.Y(n_18792)
);

AOI211x1_ASAP7_75t_L g18793 ( 
.A1(n_18611),
.A2(n_7126),
.B(n_7130),
.C(n_7117),
.Y(n_18793)
);

A2O1A1Ixp33_ASAP7_75t_L g18794 ( 
.A1(n_18561),
.A2(n_8932),
.B(n_8951),
.C(n_8928),
.Y(n_18794)
);

OAI22xp5_ASAP7_75t_L g18795 ( 
.A1(n_18607),
.A2(n_8095),
.B1(n_8103),
.B2(n_8090),
.Y(n_18795)
);

AOI221xp5_ASAP7_75t_L g18796 ( 
.A1(n_18563),
.A2(n_8103),
.B1(n_8127),
.B2(n_8095),
.C(n_8090),
.Y(n_18796)
);

AOI21xp33_ASAP7_75t_L g18797 ( 
.A1(n_18513),
.A2(n_6869),
.B(n_8103),
.Y(n_18797)
);

OAI22xp5_ASAP7_75t_L g18798 ( 
.A1(n_18526),
.A2(n_8154),
.B1(n_8171),
.B2(n_8127),
.Y(n_18798)
);

OAI32xp33_ASAP7_75t_L g18799 ( 
.A1(n_18639),
.A2(n_8171),
.A3(n_8212),
.B1(n_8154),
.B2(n_8127),
.Y(n_18799)
);

INVx1_ASAP7_75t_SL g18800 ( 
.A(n_18576),
.Y(n_18800)
);

INVx1_ASAP7_75t_L g18801 ( 
.A(n_18525),
.Y(n_18801)
);

AOI21xp5_ASAP7_75t_L g18802 ( 
.A1(n_18529),
.A2(n_7745),
.B(n_7741),
.Y(n_18802)
);

OAI21xp5_ASAP7_75t_SL g18803 ( 
.A1(n_18567),
.A2(n_7516),
.B(n_7492),
.Y(n_18803)
);

OAI21xp5_ASAP7_75t_SL g18804 ( 
.A1(n_18653),
.A2(n_7516),
.B(n_7492),
.Y(n_18804)
);

OAI22xp5_ASAP7_75t_L g18805 ( 
.A1(n_18630),
.A2(n_8171),
.B1(n_8212),
.B2(n_8154),
.Y(n_18805)
);

O2A1O1Ixp33_ASAP7_75t_L g18806 ( 
.A1(n_18554),
.A2(n_18592),
.B(n_18584),
.C(n_18536),
.Y(n_18806)
);

INVx1_ASAP7_75t_L g18807 ( 
.A(n_18528),
.Y(n_18807)
);

O2A1O1Ixp33_ASAP7_75t_L g18808 ( 
.A1(n_18601),
.A2(n_8031),
.B(n_8148),
.C(n_8002),
.Y(n_18808)
);

AOI22xp5_ASAP7_75t_L g18809 ( 
.A1(n_18524),
.A2(n_7252),
.B1(n_7257),
.B2(n_7202),
.Y(n_18809)
);

XNOR2x1_ASAP7_75t_L g18810 ( 
.A(n_18627),
.B(n_8031),
.Y(n_18810)
);

NAND2xp5_ASAP7_75t_L g18811 ( 
.A(n_18597),
.B(n_8154),
.Y(n_18811)
);

NAND4xp25_ASAP7_75t_L g18812 ( 
.A(n_18648),
.B(n_6878),
.C(n_6895),
.D(n_6875),
.Y(n_18812)
);

OAI321xp33_ASAP7_75t_L g18813 ( 
.A1(n_18626),
.A2(n_7200),
.A3(n_7196),
.B1(n_7209),
.B2(n_7199),
.C(n_7190),
.Y(n_18813)
);

AOI22xp5_ASAP7_75t_L g18814 ( 
.A1(n_18622),
.A2(n_7257),
.B1(n_7260),
.B2(n_7252),
.Y(n_18814)
);

NOR2x1_ASAP7_75t_L g18815 ( 
.A(n_18549),
.B(n_8253),
.Y(n_18815)
);

XNOR2x1_ASAP7_75t_L g18816 ( 
.A(n_18534),
.B(n_8031),
.Y(n_18816)
);

CKINVDCx20_ASAP7_75t_R g18817 ( 
.A(n_18644),
.Y(n_18817)
);

INVxp33_ASAP7_75t_L g18818 ( 
.A(n_18573),
.Y(n_18818)
);

INVx2_ASAP7_75t_SL g18819 ( 
.A(n_18534),
.Y(n_18819)
);

OAI21xp5_ASAP7_75t_SL g18820 ( 
.A1(n_18670),
.A2(n_7525),
.B(n_7516),
.Y(n_18820)
);

INVxp67_ASAP7_75t_L g18821 ( 
.A(n_18535),
.Y(n_18821)
);

INVx1_ASAP7_75t_L g18822 ( 
.A(n_18698),
.Y(n_18822)
);

OAI21xp5_ASAP7_75t_L g18823 ( 
.A1(n_18680),
.A2(n_18540),
.B(n_18587),
.Y(n_18823)
);

AOI21xp5_ASAP7_75t_L g18824 ( 
.A1(n_18711),
.A2(n_18641),
.B(n_18643),
.Y(n_18824)
);

NAND4xp25_ASAP7_75t_L g18825 ( 
.A(n_18690),
.B(n_18694),
.C(n_18706),
.D(n_18677),
.Y(n_18825)
);

NOR2x1p5_ASAP7_75t_L g18826 ( 
.A(n_18679),
.B(n_18571),
.Y(n_18826)
);

A2O1A1Ixp33_ASAP7_75t_L g18827 ( 
.A1(n_18689),
.A2(n_18740),
.B(n_18688),
.C(n_18676),
.Y(n_18827)
);

NAND2xp5_ASAP7_75t_L g18828 ( 
.A(n_18742),
.B(n_18619),
.Y(n_18828)
);

AOI22xp5_ASAP7_75t_L g18829 ( 
.A1(n_18729),
.A2(n_18682),
.B1(n_18718),
.B2(n_18713),
.Y(n_18829)
);

NAND2xp5_ASAP7_75t_L g18830 ( 
.A(n_18686),
.B(n_18747),
.Y(n_18830)
);

AOI22xp5_ASAP7_75t_L g18831 ( 
.A1(n_18723),
.A2(n_18604),
.B1(n_18515),
.B2(n_8307),
.Y(n_18831)
);

INVx1_ASAP7_75t_L g18832 ( 
.A(n_18707),
.Y(n_18832)
);

AOI322xp5_ASAP7_75t_L g18833 ( 
.A1(n_18681),
.A2(n_7592),
.A3(n_7585),
.B1(n_7252),
.B2(n_7298),
.C1(n_7260),
.C2(n_7323),
.Y(n_18833)
);

AOI221xp5_ASAP7_75t_L g18834 ( 
.A1(n_18673),
.A2(n_8214),
.B1(n_8248),
.B2(n_8212),
.C(n_8171),
.Y(n_18834)
);

AOI221xp5_ASAP7_75t_L g18835 ( 
.A1(n_18700),
.A2(n_8248),
.B1(n_8261),
.B2(n_8214),
.C(n_8212),
.Y(n_18835)
);

CKINVDCx5p33_ASAP7_75t_R g18836 ( 
.A(n_18707),
.Y(n_18836)
);

AOI221xp5_ASAP7_75t_L g18837 ( 
.A1(n_18675),
.A2(n_8261),
.B1(n_8278),
.B2(n_8248),
.C(n_8214),
.Y(n_18837)
);

INVx1_ASAP7_75t_SL g18838 ( 
.A(n_18692),
.Y(n_18838)
);

AOI221xp5_ASAP7_75t_L g18839 ( 
.A1(n_18756),
.A2(n_8261),
.B1(n_8278),
.B2(n_8248),
.C(n_8214),
.Y(n_18839)
);

AOI22xp33_ASAP7_75t_L g18840 ( 
.A1(n_18744),
.A2(n_7438),
.B1(n_7439),
.B2(n_7430),
.Y(n_18840)
);

INVx1_ASAP7_75t_SL g18841 ( 
.A(n_18817),
.Y(n_18841)
);

AOI321xp33_ASAP7_75t_L g18842 ( 
.A1(n_18738),
.A2(n_7430),
.A3(n_7439),
.B1(n_7476),
.B2(n_7470),
.C(n_7438),
.Y(n_18842)
);

NAND2xp5_ASAP7_75t_L g18843 ( 
.A(n_18774),
.B(n_8006),
.Y(n_18843)
);

AOI211xp5_ASAP7_75t_L g18844 ( 
.A1(n_18818),
.A2(n_8951),
.B(n_7994),
.C(n_7995),
.Y(n_18844)
);

NAND4xp25_ASAP7_75t_L g18845 ( 
.A(n_18776),
.B(n_6878),
.C(n_6895),
.D(n_6875),
.Y(n_18845)
);

OAI21xp5_ASAP7_75t_L g18846 ( 
.A1(n_18712),
.A2(n_7816),
.B(n_7712),
.Y(n_18846)
);

NOR3xp33_ASAP7_75t_L g18847 ( 
.A(n_18749),
.B(n_18703),
.C(n_18719),
.Y(n_18847)
);

AOI211xp5_ASAP7_75t_L g18848 ( 
.A1(n_18800),
.A2(n_7961),
.B(n_7995),
.C(n_7994),
.Y(n_18848)
);

AOI322xp5_ASAP7_75t_L g18849 ( 
.A1(n_18762),
.A2(n_7257),
.A3(n_7285),
.B1(n_7323),
.B2(n_7342),
.C1(n_7298),
.C2(n_7260),
.Y(n_18849)
);

OAI221xp5_ASAP7_75t_L g18850 ( 
.A1(n_18674),
.A2(n_8898),
.B1(n_8238),
.B2(n_8614),
.C(n_8148),
.Y(n_18850)
);

INVx1_ASAP7_75t_L g18851 ( 
.A(n_18766),
.Y(n_18851)
);

BUFx3_ASAP7_75t_L g18852 ( 
.A(n_18751),
.Y(n_18852)
);

NAND2xp5_ASAP7_75t_L g18853 ( 
.A(n_18767),
.B(n_8109),
.Y(n_18853)
);

INVx1_ASAP7_75t_SL g18854 ( 
.A(n_18777),
.Y(n_18854)
);

INVx1_ASAP7_75t_L g18855 ( 
.A(n_18780),
.Y(n_18855)
);

OAI211xp5_ASAP7_75t_L g18856 ( 
.A1(n_18821),
.A2(n_18727),
.B(n_18754),
.C(n_18745),
.Y(n_18856)
);

AOI221x1_ASAP7_75t_L g18857 ( 
.A1(n_18720),
.A2(n_8376),
.B1(n_8403),
.B2(n_8347),
.C(n_8308),
.Y(n_18857)
);

INVx1_ASAP7_75t_L g18858 ( 
.A(n_18772),
.Y(n_18858)
);

NOR3xp33_ASAP7_75t_SL g18859 ( 
.A(n_18725),
.B(n_7153),
.C(n_7425),
.Y(n_18859)
);

OAI221xp5_ASAP7_75t_SL g18860 ( 
.A1(n_18678),
.A2(n_18685),
.B1(n_18804),
.B2(n_18820),
.C(n_18803),
.Y(n_18860)
);

OAI22xp33_ASAP7_75t_SL g18861 ( 
.A1(n_18743),
.A2(n_8278),
.B1(n_8285),
.B2(n_8261),
.Y(n_18861)
);

AOI221xp5_ASAP7_75t_L g18862 ( 
.A1(n_18801),
.A2(n_8923),
.B1(n_8920),
.B2(n_8900),
.C(n_8287),
.Y(n_18862)
);

NAND4xp25_ASAP7_75t_L g18863 ( 
.A(n_18743),
.B(n_6895),
.C(n_6934),
.D(n_6878),
.Y(n_18863)
);

AOI221xp5_ASAP7_75t_L g18864 ( 
.A1(n_18807),
.A2(n_8923),
.B1(n_8920),
.B2(n_8900),
.C(n_8287),
.Y(n_18864)
);

AOI211xp5_ASAP7_75t_SL g18865 ( 
.A1(n_18730),
.A2(n_18731),
.B(n_18769),
.C(n_18790),
.Y(n_18865)
);

AOI21xp33_ASAP7_75t_L g18866 ( 
.A1(n_18761),
.A2(n_6869),
.B(n_8278),
.Y(n_18866)
);

AOI22xp5_ASAP7_75t_L g18867 ( 
.A1(n_18781),
.A2(n_8307),
.B1(n_7298),
.B2(n_7323),
.Y(n_18867)
);

OAI22xp33_ASAP7_75t_L g18868 ( 
.A1(n_18693),
.A2(n_7276),
.B1(n_7199),
.B2(n_7196),
.Y(n_18868)
);

AOI221xp5_ASAP7_75t_L g18869 ( 
.A1(n_18789),
.A2(n_8923),
.B1(n_8296),
.B2(n_8297),
.C(n_8287),
.Y(n_18869)
);

NOR4xp25_ASAP7_75t_L g18870 ( 
.A(n_18819),
.B(n_8287),
.C(n_8296),
.D(n_8285),
.Y(n_18870)
);

NAND3xp33_ASAP7_75t_SL g18871 ( 
.A(n_18786),
.B(n_5770),
.C(n_5695),
.Y(n_18871)
);

NOR2xp67_ASAP7_75t_L g18872 ( 
.A(n_18812),
.B(n_6878),
.Y(n_18872)
);

AOI222xp33_ASAP7_75t_L g18873 ( 
.A1(n_18715),
.A2(n_18775),
.B1(n_18734),
.B2(n_18757),
.C1(n_18732),
.C2(n_18748),
.Y(n_18873)
);

AOI211x1_ASAP7_75t_L g18874 ( 
.A1(n_18797),
.A2(n_7126),
.B(n_7130),
.C(n_7117),
.Y(n_18874)
);

OA22x2_ASAP7_75t_L g18875 ( 
.A1(n_18771),
.A2(n_8782),
.B1(n_8795),
.B2(n_8766),
.Y(n_18875)
);

AOI22xp5_ASAP7_75t_L g18876 ( 
.A1(n_18770),
.A2(n_8307),
.B1(n_7298),
.B2(n_7323),
.Y(n_18876)
);

AOI22xp5_ASAP7_75t_L g18877 ( 
.A1(n_18810),
.A2(n_7342),
.B1(n_7285),
.B2(n_7438),
.Y(n_18877)
);

AOI22xp5_ASAP7_75t_L g18878 ( 
.A1(n_18816),
.A2(n_7342),
.B1(n_7285),
.B2(n_7439),
.Y(n_18878)
);

INVx1_ASAP7_75t_L g18879 ( 
.A(n_18806),
.Y(n_18879)
);

OAI221xp5_ASAP7_75t_SL g18880 ( 
.A1(n_18753),
.A2(n_8238),
.B1(n_8614),
.B2(n_8148),
.C(n_8031),
.Y(n_18880)
);

OAI221xp5_ASAP7_75t_L g18881 ( 
.A1(n_18746),
.A2(n_8898),
.B1(n_8890),
.B2(n_8614),
.C(n_8792),
.Y(n_18881)
);

AOI221xp5_ASAP7_75t_L g18882 ( 
.A1(n_18760),
.A2(n_8900),
.B1(n_8920),
.B2(n_8865),
.C(n_8847),
.Y(n_18882)
);

O2A1O1Ixp33_ASAP7_75t_L g18883 ( 
.A1(n_18735),
.A2(n_8238),
.B(n_8614),
.C(n_8148),
.Y(n_18883)
);

NAND4xp75_ASAP7_75t_L g18884 ( 
.A(n_18724),
.B(n_7906),
.C(n_7863),
.D(n_8304),
.Y(n_18884)
);

AOI221xp5_ASAP7_75t_L g18885 ( 
.A1(n_18758),
.A2(n_8900),
.B1(n_8920),
.B2(n_8865),
.C(n_8847),
.Y(n_18885)
);

OAI21xp33_ASAP7_75t_L g18886 ( 
.A1(n_18684),
.A2(n_7470),
.B(n_7439),
.Y(n_18886)
);

NAND4xp25_ASAP7_75t_L g18887 ( 
.A(n_18778),
.B(n_6895),
.C(n_6934),
.D(n_6878),
.Y(n_18887)
);

AOI221x1_ASAP7_75t_L g18888 ( 
.A1(n_18709),
.A2(n_8865),
.B1(n_8620),
.B2(n_8672),
.C(n_8449),
.Y(n_18888)
);

INVx1_ASAP7_75t_L g18889 ( 
.A(n_18791),
.Y(n_18889)
);

AOI221xp5_ASAP7_75t_L g18890 ( 
.A1(n_18799),
.A2(n_8923),
.B1(n_8865),
.B2(n_8297),
.C(n_8308),
.Y(n_18890)
);

OAI21xp5_ASAP7_75t_SL g18891 ( 
.A1(n_18750),
.A2(n_7530),
.B(n_7525),
.Y(n_18891)
);

OAI22xp5_ASAP7_75t_L g18892 ( 
.A1(n_18708),
.A2(n_8296),
.B1(n_8297),
.B2(n_8285),
.Y(n_18892)
);

AOI22xp33_ASAP7_75t_L g18893 ( 
.A1(n_18784),
.A2(n_7476),
.B1(n_7503),
.B2(n_7470),
.Y(n_18893)
);

INVx1_ASAP7_75t_L g18894 ( 
.A(n_18811),
.Y(n_18894)
);

NOR3xp33_ASAP7_75t_L g18895 ( 
.A(n_18691),
.B(n_5770),
.C(n_5695),
.Y(n_18895)
);

AOI322xp5_ASAP7_75t_L g18896 ( 
.A1(n_18701),
.A2(n_7285),
.A3(n_7342),
.B1(n_7482),
.B2(n_7413),
.C1(n_7398),
.C2(n_7254),
.Y(n_18896)
);

NOR2xp33_ASAP7_75t_R g18897 ( 
.A(n_18773),
.B(n_6945),
.Y(n_18897)
);

A2O1A1Ixp33_ASAP7_75t_SL g18898 ( 
.A1(n_18788),
.A2(n_8736),
.B(n_8750),
.C(n_8730),
.Y(n_18898)
);

NOR4xp25_ASAP7_75t_L g18899 ( 
.A(n_18813),
.B(n_8296),
.C(n_8297),
.D(n_8285),
.Y(n_18899)
);

AOI22xp33_ASAP7_75t_L g18900 ( 
.A1(n_18699),
.A2(n_7476),
.B1(n_7503),
.B2(n_7470),
.Y(n_18900)
);

INVx1_ASAP7_75t_L g18901 ( 
.A(n_18683),
.Y(n_18901)
);

NOR3xp33_ASAP7_75t_L g18902 ( 
.A(n_18808),
.B(n_5770),
.C(n_5695),
.Y(n_18902)
);

O2A1O1Ixp33_ASAP7_75t_L g18903 ( 
.A1(n_18695),
.A2(n_8238),
.B(n_8614),
.C(n_8148),
.Y(n_18903)
);

NAND4xp25_ASAP7_75t_L g18904 ( 
.A(n_18741),
.B(n_6934),
.C(n_6963),
.D(n_6895),
.Y(n_18904)
);

AOI221xp5_ASAP7_75t_L g18905 ( 
.A1(n_18726),
.A2(n_8847),
.B1(n_8795),
.B2(n_8355),
.C(n_8376),
.Y(n_18905)
);

NAND4xp25_ASAP7_75t_SL g18906 ( 
.A(n_18809),
.B(n_8847),
.C(n_8795),
.D(n_8347),
.Y(n_18906)
);

INVx1_ASAP7_75t_L g18907 ( 
.A(n_18683),
.Y(n_18907)
);

O2A1O1Ixp33_ASAP7_75t_L g18908 ( 
.A1(n_18764),
.A2(n_8614),
.B(n_8792),
.C(n_8238),
.Y(n_18908)
);

INVx2_ASAP7_75t_SL g18909 ( 
.A(n_18792),
.Y(n_18909)
);

OAI221xp5_ASAP7_75t_L g18910 ( 
.A1(n_18759),
.A2(n_8898),
.B1(n_8890),
.B2(n_8792),
.C(n_8614),
.Y(n_18910)
);

AOI22xp5_ASAP7_75t_L g18911 ( 
.A1(n_18704),
.A2(n_7503),
.B1(n_7547),
.B2(n_7476),
.Y(n_18911)
);

NOR4xp25_ASAP7_75t_L g18912 ( 
.A(n_18728),
.B(n_8347),
.C(n_8355),
.D(n_8308),
.Y(n_18912)
);

AOI221xp5_ASAP7_75t_L g18913 ( 
.A1(n_18736),
.A2(n_8355),
.B1(n_8376),
.B2(n_8347),
.C(n_8308),
.Y(n_18913)
);

OAI211xp5_ASAP7_75t_L g18914 ( 
.A1(n_18814),
.A2(n_6963),
.B(n_6965),
.C(n_6934),
.Y(n_18914)
);

NAND4xp25_ASAP7_75t_L g18915 ( 
.A(n_18739),
.B(n_6963),
.C(n_6965),
.D(n_6934),
.Y(n_18915)
);

NAND2xp5_ASAP7_75t_L g18916 ( 
.A(n_18793),
.B(n_8109),
.Y(n_18916)
);

A2O1A1Ixp33_ASAP7_75t_L g18917 ( 
.A1(n_18705),
.A2(n_18782),
.B(n_18717),
.C(n_18697),
.Y(n_18917)
);

AOI221xp5_ASAP7_75t_L g18918 ( 
.A1(n_18765),
.A2(n_8384),
.B1(n_8388),
.B2(n_8376),
.C(n_8355),
.Y(n_18918)
);

XNOR2xp5_ASAP7_75t_L g18919 ( 
.A(n_18815),
.B(n_7028),
.Y(n_18919)
);

AOI211xp5_ASAP7_75t_L g18920 ( 
.A1(n_18696),
.A2(n_7994),
.B(n_7995),
.C(n_7833),
.Y(n_18920)
);

OAI221xp5_ASAP7_75t_L g18921 ( 
.A1(n_18733),
.A2(n_8890),
.B1(n_8898),
.B2(n_8792),
.C(n_8238),
.Y(n_18921)
);

AOI222xp33_ASAP7_75t_L g18922 ( 
.A1(n_18798),
.A2(n_7553),
.B1(n_7530),
.B2(n_7565),
.C1(n_7538),
.C2(n_7525),
.Y(n_18922)
);

AOI22xp33_ASAP7_75t_SL g18923 ( 
.A1(n_18699),
.A2(n_7196),
.B1(n_7199),
.B2(n_7190),
.Y(n_18923)
);

NAND2xp33_ASAP7_75t_SL g18924 ( 
.A(n_18687),
.B(n_7525),
.Y(n_18924)
);

NAND4xp25_ASAP7_75t_SL g18925 ( 
.A(n_18737),
.B(n_18714),
.C(n_18702),
.D(n_18716),
.Y(n_18925)
);

OAI222xp33_ASAP7_75t_L g18926 ( 
.A1(n_18752),
.A2(n_8402),
.B1(n_8388),
.B2(n_8403),
.C1(n_8397),
.C2(n_8384),
.Y(n_18926)
);

A2O1A1Ixp33_ASAP7_75t_L g18927 ( 
.A1(n_18710),
.A2(n_8079),
.B(n_8099),
.C(n_8093),
.Y(n_18927)
);

A2O1A1Ixp33_ASAP7_75t_L g18928 ( 
.A1(n_18763),
.A2(n_8079),
.B(n_8099),
.C(n_8093),
.Y(n_18928)
);

AOI21xp5_ASAP7_75t_L g18929 ( 
.A1(n_18794),
.A2(n_8890),
.B(n_8792),
.Y(n_18929)
);

O2A1O1Ixp33_ASAP7_75t_L g18930 ( 
.A1(n_18805),
.A2(n_8890),
.B(n_8898),
.C(n_8792),
.Y(n_18930)
);

NOR3x1_ASAP7_75t_L g18931 ( 
.A(n_18795),
.B(n_7903),
.C(n_7899),
.Y(n_18931)
);

NAND4xp25_ASAP7_75t_L g18932 ( 
.A(n_18722),
.B(n_6963),
.C(n_6965),
.D(n_6934),
.Y(n_18932)
);

AND2x4_ASAP7_75t_L g18933 ( 
.A(n_18779),
.B(n_6963),
.Y(n_18933)
);

A2O1A1Ixp33_ASAP7_75t_SL g18934 ( 
.A1(n_18787),
.A2(n_8766),
.B(n_8782),
.C(n_8750),
.Y(n_18934)
);

OAI22xp5_ASAP7_75t_L g18935 ( 
.A1(n_18721),
.A2(n_8388),
.B1(n_8397),
.B2(n_8384),
.Y(n_18935)
);

NOR2xp33_ASAP7_75t_L g18936 ( 
.A(n_18768),
.B(n_18783),
.Y(n_18936)
);

AOI221xp5_ASAP7_75t_L g18937 ( 
.A1(n_18796),
.A2(n_8782),
.B1(n_8795),
.B2(n_8766),
.C(n_8750),
.Y(n_18937)
);

NAND5xp2_ASAP7_75t_L g18938 ( 
.A(n_18802),
.B(n_7401),
.C(n_7475),
.D(n_7454),
.E(n_7390),
.Y(n_18938)
);

NAND4xp75_ASAP7_75t_L g18939 ( 
.A(n_18785),
.B(n_7906),
.C(n_7863),
.D(n_8304),
.Y(n_18939)
);

AOI221xp5_ASAP7_75t_L g18940 ( 
.A1(n_18755),
.A2(n_8782),
.B1(n_8766),
.B2(n_8750),
.C(n_8397),
.Y(n_18940)
);

AO221x1_ASAP7_75t_L g18941 ( 
.A1(n_18698),
.A2(n_7199),
.B1(n_7200),
.B2(n_7196),
.C(n_7190),
.Y(n_18941)
);

INVx1_ASAP7_75t_L g18942 ( 
.A(n_18698),
.Y(n_18942)
);

INVx1_ASAP7_75t_L g18943 ( 
.A(n_18698),
.Y(n_18943)
);

AOI21xp5_ASAP7_75t_L g18944 ( 
.A1(n_18680),
.A2(n_8890),
.B(n_8792),
.Y(n_18944)
);

NOR2xp33_ASAP7_75t_R g18945 ( 
.A(n_18729),
.B(n_6945),
.Y(n_18945)
);

A2O1A1Ixp33_ASAP7_75t_L g18946 ( 
.A1(n_18711),
.A2(n_8093),
.B(n_8100),
.C(n_8099),
.Y(n_18946)
);

AO22x2_ASAP7_75t_L g18947 ( 
.A1(n_18740),
.A2(n_8388),
.B1(n_8397),
.B2(n_8384),
.Y(n_18947)
);

NAND4xp25_ASAP7_75t_L g18948 ( 
.A(n_18690),
.B(n_6965),
.C(n_7050),
.D(n_6963),
.Y(n_18948)
);

INVx1_ASAP7_75t_L g18949 ( 
.A(n_18698),
.Y(n_18949)
);

OAI222xp33_ASAP7_75t_L g18950 ( 
.A1(n_18706),
.A2(n_8423),
.B1(n_8403),
.B2(n_8436),
.C1(n_8407),
.C2(n_8402),
.Y(n_18950)
);

HB1xp67_ASAP7_75t_L g18951 ( 
.A(n_18689),
.Y(n_18951)
);

AOI22xp33_ASAP7_75t_L g18952 ( 
.A1(n_18698),
.A2(n_7547),
.B1(n_7549),
.B2(n_7503),
.Y(n_18952)
);

AOI221xp5_ASAP7_75t_L g18953 ( 
.A1(n_18680),
.A2(n_8717),
.B1(n_8723),
.B2(n_8697),
.C(n_8696),
.Y(n_18953)
);

AOI22xp5_ASAP7_75t_L g18954 ( 
.A1(n_18729),
.A2(n_7549),
.B1(n_7569),
.B2(n_7547),
.Y(n_18954)
);

OAI221xp5_ASAP7_75t_SL g18955 ( 
.A1(n_18767),
.A2(n_8898),
.B1(n_8890),
.B2(n_7569),
.C(n_7549),
.Y(n_18955)
);

O2A1O1Ixp33_ASAP7_75t_L g18956 ( 
.A1(n_18680),
.A2(n_8898),
.B(n_8403),
.C(n_8407),
.Y(n_18956)
);

AOI221xp5_ASAP7_75t_SL g18957 ( 
.A1(n_18706),
.A2(n_7199),
.B1(n_7200),
.B2(n_7196),
.C(n_7190),
.Y(n_18957)
);

OAI211xp5_ASAP7_75t_SL g18958 ( 
.A1(n_18680),
.A2(n_7151),
.B(n_7155),
.C(n_7136),
.Y(n_18958)
);

AOI211xp5_ASAP7_75t_L g18959 ( 
.A1(n_18680),
.A2(n_7833),
.B(n_7530),
.C(n_7538),
.Y(n_18959)
);

AND2x2_ASAP7_75t_L g18960 ( 
.A(n_18698),
.B(n_8109),
.Y(n_18960)
);

OAI211xp5_ASAP7_75t_SL g18961 ( 
.A1(n_18680),
.A2(n_7151),
.B(n_7155),
.C(n_7136),
.Y(n_18961)
);

NOR2x1_ASAP7_75t_L g18962 ( 
.A(n_18825),
.B(n_6965),
.Y(n_18962)
);

NOR2x1_ASAP7_75t_L g18963 ( 
.A(n_18832),
.B(n_6965),
.Y(n_18963)
);

NAND4xp75_ASAP7_75t_L g18964 ( 
.A(n_18822),
.B(n_8304),
.C(n_7906),
.D(n_7863),
.Y(n_18964)
);

XOR2x1_ASAP7_75t_L g18965 ( 
.A(n_18826),
.B(n_7863),
.Y(n_18965)
);

NAND3xp33_ASAP7_75t_L g18966 ( 
.A(n_18827),
.B(n_5365),
.C(n_7212),
.Y(n_18966)
);

AOI21xp5_ASAP7_75t_L g18967 ( 
.A1(n_18942),
.A2(n_8723),
.B(n_8717),
.Y(n_18967)
);

NAND2xp5_ASAP7_75t_L g18968 ( 
.A(n_18943),
.B(n_8109),
.Y(n_18968)
);

OAI22xp5_ASAP7_75t_L g18969 ( 
.A1(n_18829),
.A2(n_8407),
.B1(n_8423),
.B2(n_8402),
.Y(n_18969)
);

OAI22xp5_ASAP7_75t_L g18970 ( 
.A1(n_18949),
.A2(n_8407),
.B1(n_8423),
.B2(n_8402),
.Y(n_18970)
);

INVx1_ASAP7_75t_L g18971 ( 
.A(n_18951),
.Y(n_18971)
);

INVx1_ASAP7_75t_L g18972 ( 
.A(n_18855),
.Y(n_18972)
);

NOR3xp33_ASAP7_75t_L g18973 ( 
.A(n_18856),
.B(n_5866),
.C(n_5817),
.Y(n_18973)
);

INVx1_ASAP7_75t_L g18974 ( 
.A(n_18836),
.Y(n_18974)
);

AND2x2_ASAP7_75t_L g18975 ( 
.A(n_18838),
.B(n_8109),
.Y(n_18975)
);

AOI22xp5_ASAP7_75t_L g18976 ( 
.A1(n_18847),
.A2(n_7549),
.B1(n_7569),
.B2(n_7547),
.Y(n_18976)
);

OA22x2_ASAP7_75t_L g18977 ( 
.A1(n_18879),
.A2(n_8436),
.B1(n_8440),
.B2(n_8423),
.Y(n_18977)
);

INVx1_ASAP7_75t_L g18978 ( 
.A(n_18858),
.Y(n_18978)
);

NOR2xp33_ASAP7_75t_SL g18979 ( 
.A(n_18841),
.B(n_6945),
.Y(n_18979)
);

NAND2xp5_ASAP7_75t_L g18980 ( 
.A(n_18854),
.B(n_8109),
.Y(n_18980)
);

NAND4xp75_ASAP7_75t_L g18981 ( 
.A(n_18828),
.B(n_8304),
.C(n_7906),
.D(n_7863),
.Y(n_18981)
);

OR2x2_ASAP7_75t_L g18982 ( 
.A(n_18948),
.B(n_18887),
.Y(n_18982)
);

NAND3x1_ASAP7_75t_L g18983 ( 
.A(n_18830),
.B(n_6896),
.C(n_6885),
.Y(n_18983)
);

NAND2x1p5_ASAP7_75t_L g18984 ( 
.A(n_18852),
.B(n_6290),
.Y(n_18984)
);

NAND2xp5_ASAP7_75t_L g18985 ( 
.A(n_18919),
.B(n_18865),
.Y(n_18985)
);

NAND3xp33_ASAP7_75t_SL g18986 ( 
.A(n_18823),
.B(n_5866),
.C(n_5817),
.Y(n_18986)
);

OA22x2_ASAP7_75t_SL g18987 ( 
.A1(n_18851),
.A2(n_8440),
.B1(n_8449),
.B2(n_8436),
.Y(n_18987)
);

AND2x2_ASAP7_75t_L g18988 ( 
.A(n_18960),
.B(n_8109),
.Y(n_18988)
);

INVx1_ASAP7_75t_L g18989 ( 
.A(n_18889),
.Y(n_18989)
);

XOR2xp5_ASAP7_75t_L g18990 ( 
.A(n_18909),
.B(n_6290),
.Y(n_18990)
);

NOR2x1_ASAP7_75t_SL g18991 ( 
.A(n_18901),
.B(n_7525),
.Y(n_18991)
);

NAND2xp5_ASAP7_75t_L g18992 ( 
.A(n_18894),
.B(n_8436),
.Y(n_18992)
);

NAND4xp75_ASAP7_75t_L g18993 ( 
.A(n_18824),
.B(n_8304),
.C(n_6595),
.D(n_6636),
.Y(n_18993)
);

NAND3xp33_ASAP7_75t_L g18994 ( 
.A(n_18873),
.B(n_5365),
.C(n_7212),
.Y(n_18994)
);

INVx1_ASAP7_75t_L g18995 ( 
.A(n_18907),
.Y(n_18995)
);

NAND2xp5_ASAP7_75t_L g18996 ( 
.A(n_18944),
.B(n_8440),
.Y(n_18996)
);

OAI22xp5_ASAP7_75t_L g18997 ( 
.A1(n_18850),
.A2(n_8440),
.B1(n_8489),
.B2(n_8449),
.Y(n_18997)
);

NOR2xp33_ASAP7_75t_L g18998 ( 
.A(n_18860),
.B(n_6945),
.Y(n_18998)
);

INVx1_ASAP7_75t_L g18999 ( 
.A(n_18936),
.Y(n_18999)
);

OAI22xp5_ASAP7_75t_L g19000 ( 
.A1(n_18877),
.A2(n_8449),
.B1(n_8504),
.B2(n_8489),
.Y(n_19000)
);

NAND2xp33_ASAP7_75t_L g19001 ( 
.A(n_18945),
.B(n_18897),
.Y(n_19001)
);

NAND2xp5_ASAP7_75t_L g19002 ( 
.A(n_18917),
.B(n_8489),
.Y(n_19002)
);

INVx1_ASAP7_75t_L g19003 ( 
.A(n_18925),
.Y(n_19003)
);

INVxp33_ASAP7_75t_SL g19004 ( 
.A(n_18878),
.Y(n_19004)
);

NOR3x1_ASAP7_75t_L g19005 ( 
.A(n_18843),
.B(n_7937),
.C(n_7927),
.Y(n_19005)
);

INVx1_ASAP7_75t_L g19006 ( 
.A(n_18831),
.Y(n_19006)
);

INVx1_ASAP7_75t_L g19007 ( 
.A(n_18895),
.Y(n_19007)
);

NOR3x2_ASAP7_75t_L g19008 ( 
.A(n_18884),
.B(n_6945),
.C(n_7212),
.Y(n_19008)
);

NOR2x1_ASAP7_75t_L g19009 ( 
.A(n_18872),
.B(n_7050),
.Y(n_19009)
);

INVxp67_ASAP7_75t_SL g19010 ( 
.A(n_18902),
.Y(n_19010)
);

AOI22xp5_ASAP7_75t_L g19011 ( 
.A1(n_18924),
.A2(n_18866),
.B1(n_18863),
.B2(n_18853),
.Y(n_19011)
);

NOR3xp33_ASAP7_75t_L g19012 ( 
.A(n_18955),
.B(n_5866),
.C(n_5817),
.Y(n_19012)
);

NAND3xp33_ASAP7_75t_L g19013 ( 
.A(n_18910),
.B(n_5365),
.C(n_7212),
.Y(n_19013)
);

NAND4xp25_ASAP7_75t_L g19014 ( 
.A(n_18883),
.B(n_7055),
.C(n_7064),
.D(n_7050),
.Y(n_19014)
);

NOR2xp33_ASAP7_75t_L g19015 ( 
.A(n_18904),
.B(n_7050),
.Y(n_19015)
);

NAND4xp25_ASAP7_75t_L g19016 ( 
.A(n_18908),
.B(n_7055),
.C(n_7064),
.D(n_7050),
.Y(n_19016)
);

NAND4xp75_ASAP7_75t_L g19017 ( 
.A(n_18874),
.B(n_6595),
.C(n_6636),
.D(n_6581),
.Y(n_19017)
);

NAND4xp25_ASAP7_75t_L g19018 ( 
.A(n_18880),
.B(n_7055),
.C(n_7064),
.D(n_7050),
.Y(n_19018)
);

NOR2xp33_ASAP7_75t_L g19019 ( 
.A(n_18933),
.B(n_7055),
.Y(n_19019)
);

NAND2xp5_ASAP7_75t_L g19020 ( 
.A(n_18933),
.B(n_8489),
.Y(n_19020)
);

INVx1_ASAP7_75t_L g19021 ( 
.A(n_18875),
.Y(n_19021)
);

NAND4xp25_ASAP7_75t_L g19022 ( 
.A(n_18956),
.B(n_7064),
.C(n_7083),
.D(n_7055),
.Y(n_19022)
);

NAND4xp75_ASAP7_75t_L g19023 ( 
.A(n_18957),
.B(n_6595),
.C(n_6636),
.D(n_6581),
.Y(n_19023)
);

AOI21xp5_ASAP7_75t_L g19024 ( 
.A1(n_18934),
.A2(n_8723),
.B(n_8717),
.Y(n_19024)
);

NAND3xp33_ASAP7_75t_SL g19025 ( 
.A(n_18899),
.B(n_5886),
.C(n_5866),
.Y(n_19025)
);

INVx1_ASAP7_75t_L g19026 ( 
.A(n_18861),
.Y(n_19026)
);

INVx1_ASAP7_75t_L g19027 ( 
.A(n_18871),
.Y(n_19027)
);

AOI22xp5_ASAP7_75t_L g19028 ( 
.A1(n_18906),
.A2(n_7569),
.B1(n_7199),
.B2(n_7200),
.Y(n_19028)
);

INVx1_ASAP7_75t_L g19029 ( 
.A(n_18891),
.Y(n_19029)
);

OR2x2_ASAP7_75t_L g19030 ( 
.A(n_18915),
.B(n_7781),
.Y(n_19030)
);

AOI22xp5_ASAP7_75t_L g19031 ( 
.A1(n_18845),
.A2(n_7199),
.B1(n_7200),
.B2(n_7190),
.Y(n_19031)
);

NOR2xp33_ASAP7_75t_L g19032 ( 
.A(n_18921),
.B(n_7055),
.Y(n_19032)
);

NAND4xp75_ASAP7_75t_L g19033 ( 
.A(n_18867),
.B(n_6595),
.C(n_6636),
.D(n_6581),
.Y(n_19033)
);

INVx1_ASAP7_75t_L g19034 ( 
.A(n_18941),
.Y(n_19034)
);

INVx1_ASAP7_75t_L g19035 ( 
.A(n_18916),
.Y(n_19035)
);

AND2x2_ASAP7_75t_L g19036 ( 
.A(n_18859),
.B(n_8694),
.Y(n_19036)
);

NOR3x1_ASAP7_75t_L g19037 ( 
.A(n_18914),
.B(n_7937),
.C(n_7927),
.Y(n_19037)
);

INVxp67_ASAP7_75t_L g19038 ( 
.A(n_18932),
.Y(n_19038)
);

NAND4xp75_ASAP7_75t_L g19039 ( 
.A(n_18876),
.B(n_6688),
.C(n_6691),
.D(n_6581),
.Y(n_19039)
);

NAND4xp75_ASAP7_75t_L g19040 ( 
.A(n_18888),
.B(n_6691),
.C(n_6694),
.D(n_6688),
.Y(n_19040)
);

NOR3x2_ASAP7_75t_L g19041 ( 
.A(n_18939),
.B(n_7233),
.C(n_7212),
.Y(n_19041)
);

INVx2_ASAP7_75t_L g19042 ( 
.A(n_18947),
.Y(n_19042)
);

NOR3x1_ASAP7_75t_L g19043 ( 
.A(n_18898),
.B(n_7937),
.C(n_7927),
.Y(n_19043)
);

AND2x2_ASAP7_75t_L g19044 ( 
.A(n_18893),
.B(n_8694),
.Y(n_19044)
);

NOR2x1_ASAP7_75t_L g19045 ( 
.A(n_18961),
.B(n_7064),
.Y(n_19045)
);

NOR3xp33_ASAP7_75t_L g19046 ( 
.A(n_18938),
.B(n_18958),
.C(n_18868),
.Y(n_19046)
);

NAND3xp33_ASAP7_75t_L g19047 ( 
.A(n_18923),
.B(n_5365),
.C(n_7212),
.Y(n_19047)
);

NOR3xp33_ASAP7_75t_SL g19048 ( 
.A(n_18886),
.B(n_7153),
.C(n_7425),
.Y(n_19048)
);

INVx1_ASAP7_75t_L g19049 ( 
.A(n_18870),
.Y(n_19049)
);

NAND4xp75_ASAP7_75t_L g19050 ( 
.A(n_18929),
.B(n_18931),
.C(n_18954),
.D(n_18911),
.Y(n_19050)
);

INVx3_ASAP7_75t_L g19051 ( 
.A(n_18947),
.Y(n_19051)
);

CKINVDCx16_ASAP7_75t_R g19052 ( 
.A(n_18912),
.Y(n_19052)
);

NAND4xp75_ASAP7_75t_L g19053 ( 
.A(n_18857),
.B(n_6691),
.C(n_6694),
.D(n_6688),
.Y(n_19053)
);

INVx1_ASAP7_75t_L g19054 ( 
.A(n_18930),
.Y(n_19054)
);

INVx2_ASAP7_75t_L g19055 ( 
.A(n_18935),
.Y(n_19055)
);

INVx1_ASAP7_75t_L g19056 ( 
.A(n_18842),
.Y(n_19056)
);

NAND3xp33_ASAP7_75t_L g19057 ( 
.A(n_18952),
.B(n_7233),
.C(n_7463),
.Y(n_19057)
);

INVx1_ASAP7_75t_L g19058 ( 
.A(n_18903),
.Y(n_19058)
);

NOR2xp33_ASAP7_75t_L g19059 ( 
.A(n_18881),
.B(n_7064),
.Y(n_19059)
);

NAND2xp5_ASAP7_75t_L g19060 ( 
.A(n_18896),
.B(n_8504),
.Y(n_19060)
);

NAND3xp33_ASAP7_75t_SL g19061 ( 
.A(n_18849),
.B(n_5886),
.C(n_5866),
.Y(n_19061)
);

NOR3xp33_ASAP7_75t_L g19062 ( 
.A(n_18950),
.B(n_5897),
.C(n_5886),
.Y(n_19062)
);

INVx1_ASAP7_75t_L g19063 ( 
.A(n_18892),
.Y(n_19063)
);

INVx1_ASAP7_75t_L g19064 ( 
.A(n_18927),
.Y(n_19064)
);

XNOR2xp5_ASAP7_75t_L g19065 ( 
.A(n_18840),
.B(n_18959),
.Y(n_19065)
);

NOR2xp33_ASAP7_75t_L g19066 ( 
.A(n_18926),
.B(n_7083),
.Y(n_19066)
);

NOR2x1_ASAP7_75t_L g19067 ( 
.A(n_18928),
.B(n_7083),
.Y(n_19067)
);

NAND4xp75_ASAP7_75t_L g19068 ( 
.A(n_18953),
.B(n_6691),
.C(n_6694),
.D(n_6688),
.Y(n_19068)
);

NOR2x1_ASAP7_75t_L g19069 ( 
.A(n_18946),
.B(n_18846),
.Y(n_19069)
);

INVx1_ASAP7_75t_L g19070 ( 
.A(n_18900),
.Y(n_19070)
);

NOR2x1_ASAP7_75t_L g19071 ( 
.A(n_18833),
.B(n_7083),
.Y(n_19071)
);

NAND4xp75_ASAP7_75t_L g19072 ( 
.A(n_18835),
.B(n_6706),
.C(n_6790),
.D(n_6694),
.Y(n_19072)
);

NOR3xp33_ASAP7_75t_L g19073 ( 
.A(n_18834),
.B(n_5897),
.C(n_5886),
.Y(n_19073)
);

NAND3xp33_ASAP7_75t_L g19074 ( 
.A(n_18862),
.B(n_18869),
.C(n_18864),
.Y(n_19074)
);

INVx2_ASAP7_75t_L g19075 ( 
.A(n_18940),
.Y(n_19075)
);

INVx1_ASAP7_75t_L g19076 ( 
.A(n_18922),
.Y(n_19076)
);

INVx1_ASAP7_75t_L g19077 ( 
.A(n_18920),
.Y(n_19077)
);

NAND2xp5_ASAP7_75t_L g19078 ( 
.A(n_18882),
.B(n_8504),
.Y(n_19078)
);

NAND3xp33_ASAP7_75t_SL g19079 ( 
.A(n_18848),
.B(n_5897),
.C(n_5886),
.Y(n_19079)
);

AOI221xp5_ASAP7_75t_L g19080 ( 
.A1(n_18998),
.A2(n_18885),
.B1(n_18890),
.B2(n_18837),
.C(n_18918),
.Y(n_19080)
);

AOI221xp5_ASAP7_75t_L g19081 ( 
.A1(n_18971),
.A2(n_18905),
.B1(n_18913),
.B2(n_18937),
.C(n_18839),
.Y(n_19081)
);

OAI22xp5_ASAP7_75t_L g19082 ( 
.A1(n_18966),
.A2(n_18972),
.B1(n_18978),
.B2(n_18994),
.Y(n_19082)
);

AOI211x1_ASAP7_75t_L g19083 ( 
.A1(n_19002),
.A2(n_18844),
.B(n_7131),
.C(n_7500),
.Y(n_19083)
);

NAND3xp33_ASAP7_75t_SL g19084 ( 
.A(n_19003),
.B(n_5942),
.C(n_5897),
.Y(n_19084)
);

AOI22xp5_ASAP7_75t_L g19085 ( 
.A1(n_18979),
.A2(n_18999),
.B1(n_18990),
.B2(n_18974),
.Y(n_19085)
);

AOI221xp5_ASAP7_75t_L g19086 ( 
.A1(n_19058),
.A2(n_8560),
.B1(n_8571),
.B2(n_8508),
.C(n_8504),
.Y(n_19086)
);

NAND4xp25_ASAP7_75t_SL g19087 ( 
.A(n_18962),
.B(n_8560),
.C(n_8571),
.D(n_8508),
.Y(n_19087)
);

NAND2xp5_ASAP7_75t_L g19088 ( 
.A(n_19034),
.B(n_8508),
.Y(n_19088)
);

AOI221xp5_ASAP7_75t_L g19089 ( 
.A1(n_19006),
.A2(n_8571),
.B1(n_8578),
.B2(n_8560),
.C(n_8508),
.Y(n_19089)
);

OAI221xp5_ASAP7_75t_SL g19090 ( 
.A1(n_19011),
.A2(n_8578),
.B1(n_8604),
.B2(n_8571),
.C(n_8560),
.Y(n_19090)
);

XNOR2x1_ASAP7_75t_L g19091 ( 
.A(n_18985),
.B(n_6290),
.Y(n_19091)
);

AND2x2_ASAP7_75t_L g19092 ( 
.A(n_18975),
.B(n_18984),
.Y(n_19092)
);

NAND3xp33_ASAP7_75t_SL g19093 ( 
.A(n_18989),
.B(n_5942),
.C(n_5897),
.Y(n_19093)
);

NAND4xp25_ASAP7_75t_SL g19094 ( 
.A(n_19046),
.B(n_8604),
.C(n_8615),
.D(n_8578),
.Y(n_19094)
);

NOR4xp25_ASAP7_75t_L g19095 ( 
.A(n_18995),
.B(n_8604),
.C(n_8615),
.D(n_8578),
.Y(n_19095)
);

NAND3xp33_ASAP7_75t_L g19096 ( 
.A(n_19001),
.B(n_7233),
.C(n_7463),
.Y(n_19096)
);

NAND4xp75_ASAP7_75t_L g19097 ( 
.A(n_19070),
.B(n_6706),
.C(n_6803),
.D(n_6790),
.Y(n_19097)
);

OAI211xp5_ASAP7_75t_SL g19098 ( 
.A1(n_19054),
.A2(n_8615),
.B(n_8620),
.C(n_8604),
.Y(n_19098)
);

NAND2xp5_ASAP7_75t_L g19099 ( 
.A(n_19052),
.B(n_8615),
.Y(n_19099)
);

OAI211xp5_ASAP7_75t_SL g19100 ( 
.A1(n_19038),
.A2(n_8630),
.B(n_8637),
.C(n_8620),
.Y(n_19100)
);

AOI221xp5_ASAP7_75t_L g19101 ( 
.A1(n_19064),
.A2(n_8637),
.B1(n_8654),
.B2(n_8630),
.C(n_8620),
.Y(n_19101)
);

AOI221xp5_ASAP7_75t_L g19102 ( 
.A1(n_19026),
.A2(n_8654),
.B1(n_8659),
.B2(n_8637),
.C(n_8630),
.Y(n_19102)
);

AOI211xp5_ASAP7_75t_L g19103 ( 
.A1(n_19056),
.A2(n_19027),
.B(n_19007),
.C(n_19077),
.Y(n_19103)
);

OR5x1_ASAP7_75t_L g19104 ( 
.A(n_19025),
.B(n_8708),
.C(n_8806),
.D(n_8942),
.E(n_8763),
.Y(n_19104)
);

AOI221xp5_ASAP7_75t_L g19105 ( 
.A1(n_19021),
.A2(n_8654),
.B1(n_8659),
.B2(n_8637),
.C(n_8630),
.Y(n_19105)
);

AOI221xp5_ASAP7_75t_L g19106 ( 
.A1(n_19035),
.A2(n_8665),
.B1(n_8672),
.B2(n_8659),
.C(n_8654),
.Y(n_19106)
);

NOR2xp67_ASAP7_75t_L g19107 ( 
.A(n_19051),
.B(n_5942),
.Y(n_19107)
);

NAND2xp5_ASAP7_75t_L g19108 ( 
.A(n_19032),
.B(n_8659),
.Y(n_19108)
);

OAI211xp5_ASAP7_75t_SL g19109 ( 
.A1(n_19076),
.A2(n_8672),
.B(n_8696),
.C(n_8665),
.Y(n_19109)
);

A2O1A1Ixp33_ASAP7_75t_L g19110 ( 
.A1(n_19049),
.A2(n_8725),
.B(n_8730),
.C(n_8723),
.Y(n_19110)
);

NAND3xp33_ASAP7_75t_SL g19111 ( 
.A(n_19029),
.B(n_5966),
.C(n_5942),
.Y(n_19111)
);

NAND4xp25_ASAP7_75t_L g19112 ( 
.A(n_19004),
.B(n_7128),
.C(n_7178),
.D(n_7083),
.Y(n_19112)
);

NOR3xp33_ASAP7_75t_L g19113 ( 
.A(n_19010),
.B(n_5966),
.C(n_5942),
.Y(n_19113)
);

NOR4xp25_ASAP7_75t_L g19114 ( 
.A(n_19063),
.B(n_8672),
.C(n_8696),
.D(n_8665),
.Y(n_19114)
);

NAND3xp33_ASAP7_75t_L g19115 ( 
.A(n_19075),
.B(n_7233),
.C(n_7463),
.Y(n_19115)
);

NOR3xp33_ASAP7_75t_L g19116 ( 
.A(n_19055),
.B(n_6028),
.C(n_5966),
.Y(n_19116)
);

AND5x1_ASAP7_75t_L g19117 ( 
.A(n_19059),
.B(n_7658),
.C(n_7781),
.D(n_7752),
.E(n_8708),
.Y(n_19117)
);

AOI211xp5_ASAP7_75t_L g19118 ( 
.A1(n_19065),
.A2(n_7530),
.B(n_7538),
.C(n_7525),
.Y(n_19118)
);

OAI211xp5_ASAP7_75t_SL g19119 ( 
.A1(n_18982),
.A2(n_8696),
.B(n_8697),
.C(n_8665),
.Y(n_19119)
);

O2A1O1Ixp5_ASAP7_75t_L g19120 ( 
.A1(n_19051),
.A2(n_8717),
.B(n_8725),
.C(n_8697),
.Y(n_19120)
);

NOR3xp33_ASAP7_75t_L g19121 ( 
.A(n_19050),
.B(n_6028),
.C(n_5966),
.Y(n_19121)
);

NOR4xp25_ASAP7_75t_L g19122 ( 
.A(n_19042),
.B(n_19074),
.C(n_18992),
.D(n_18968),
.Y(n_19122)
);

NAND3xp33_ASAP7_75t_L g19123 ( 
.A(n_18973),
.B(n_7233),
.C(n_7463),
.Y(n_19123)
);

NOR3x1_ASAP7_75t_L g19124 ( 
.A(n_18980),
.B(n_7833),
.C(n_7899),
.Y(n_19124)
);

NOR3xp33_ASAP7_75t_L g19125 ( 
.A(n_19069),
.B(n_6028),
.C(n_5966),
.Y(n_19125)
);

AOI322xp5_ASAP7_75t_L g19126 ( 
.A1(n_19015),
.A2(n_8697),
.A3(n_8736),
.B1(n_8725),
.B2(n_8730),
.C1(n_7095),
.C2(n_7116),
.Y(n_19126)
);

NAND3xp33_ASAP7_75t_SL g19127 ( 
.A(n_19012),
.B(n_6040),
.C(n_6028),
.Y(n_19127)
);

NOR3xp33_ASAP7_75t_L g19128 ( 
.A(n_19013),
.B(n_6040),
.C(n_6028),
.Y(n_19128)
);

OAI21xp5_ASAP7_75t_SL g19129 ( 
.A1(n_19009),
.A2(n_18963),
.B(n_19019),
.Y(n_19129)
);

NAND4xp25_ASAP7_75t_SL g19130 ( 
.A(n_18996),
.B(n_8730),
.C(n_8736),
.D(n_8725),
.Y(n_19130)
);

AOI221xp5_ASAP7_75t_L g19131 ( 
.A1(n_19061),
.A2(n_8736),
.B1(n_7209),
.B2(n_7228),
.C(n_7200),
.Y(n_19131)
);

OAI211xp5_ASAP7_75t_L g19132 ( 
.A1(n_19018),
.A2(n_7128),
.B(n_7178),
.C(n_7083),
.Y(n_19132)
);

NOR3xp33_ASAP7_75t_L g19133 ( 
.A(n_19014),
.B(n_6045),
.C(n_6040),
.Y(n_19133)
);

OAI221xp5_ASAP7_75t_L g19134 ( 
.A1(n_19066),
.A2(n_7186),
.B1(n_7227),
.B2(n_7178),
.C(n_7128),
.Y(n_19134)
);

OAI221xp5_ASAP7_75t_L g19135 ( 
.A1(n_19060),
.A2(n_7186),
.B1(n_7227),
.B2(n_7178),
.C(n_7128),
.Y(n_19135)
);

NAND3xp33_ASAP7_75t_SL g19136 ( 
.A(n_19073),
.B(n_6045),
.C(n_6040),
.Y(n_19136)
);

NAND4xp75_ASAP7_75t_L g19137 ( 
.A(n_19071),
.B(n_19067),
.C(n_19045),
.D(n_19044),
.Y(n_19137)
);

NAND4xp25_ASAP7_75t_L g19138 ( 
.A(n_19057),
.B(n_7178),
.C(n_7186),
.D(n_7128),
.Y(n_19138)
);

NAND2xp5_ASAP7_75t_L g19139 ( 
.A(n_18991),
.B(n_7530),
.Y(n_19139)
);

AOI211x1_ASAP7_75t_SL g19140 ( 
.A1(n_19079),
.A2(n_7200),
.B(n_7209),
.C(n_7190),
.Y(n_19140)
);

NAND5xp2_ASAP7_75t_L g19141 ( 
.A(n_18976),
.B(n_7401),
.C(n_7475),
.D(n_7454),
.E(n_7390),
.Y(n_19141)
);

NOR3xp33_ASAP7_75t_SL g19142 ( 
.A(n_19016),
.B(n_7131),
.C(n_7239),
.Y(n_19142)
);

NAND3xp33_ASAP7_75t_L g19143 ( 
.A(n_19047),
.B(n_7233),
.C(n_7463),
.Y(n_19143)
);

OAI211xp5_ASAP7_75t_L g19144 ( 
.A1(n_19022),
.A2(n_7178),
.B(n_7186),
.C(n_7128),
.Y(n_19144)
);

OAI211xp5_ASAP7_75t_SL g19145 ( 
.A1(n_19020),
.A2(n_7136),
.B(n_7155),
.C(n_7151),
.Y(n_19145)
);

NAND2xp5_ASAP7_75t_SL g19146 ( 
.A(n_19031),
.B(n_7530),
.Y(n_19146)
);

AOI22xp33_ASAP7_75t_L g19147 ( 
.A1(n_18986),
.A2(n_7553),
.B1(n_7565),
.B2(n_7538),
.Y(n_19147)
);

NAND4xp25_ASAP7_75t_L g19148 ( 
.A(n_19030),
.B(n_18967),
.C(n_19078),
.D(n_18997),
.Y(n_19148)
);

NOR3xp33_ASAP7_75t_SL g19149 ( 
.A(n_19033),
.B(n_7248),
.C(n_7239),
.Y(n_19149)
);

O2A1O1Ixp33_ASAP7_75t_L g19150 ( 
.A1(n_18969),
.A2(n_6666),
.B(n_6730),
.C(n_6626),
.Y(n_19150)
);

OAI221xp5_ASAP7_75t_L g19151 ( 
.A1(n_19062),
.A2(n_7235),
.B1(n_7265),
.B2(n_7227),
.C(n_7186),
.Y(n_19151)
);

AOI221xp5_ASAP7_75t_L g19152 ( 
.A1(n_19000),
.A2(n_7228),
.B1(n_7240),
.B2(n_7209),
.C(n_7200),
.Y(n_19152)
);

AOI211xp5_ASAP7_75t_L g19153 ( 
.A1(n_19036),
.A2(n_18970),
.B(n_18988),
.C(n_19008),
.Y(n_19153)
);

AOI22xp5_ASAP7_75t_L g19154 ( 
.A1(n_19039),
.A2(n_7209),
.B1(n_7228),
.B2(n_7200),
.Y(n_19154)
);

OAI221xp5_ASAP7_75t_SL g19155 ( 
.A1(n_19028),
.A2(n_7121),
.B1(n_7176),
.B2(n_7120),
.C(n_7099),
.Y(n_19155)
);

AND2x2_ASAP7_75t_L g19156 ( 
.A(n_19048),
.B(n_18965),
.Y(n_19156)
);

NAND2xp5_ASAP7_75t_L g19157 ( 
.A(n_19023),
.B(n_7538),
.Y(n_19157)
);

A2O1A1Ixp33_ASAP7_75t_L g19158 ( 
.A1(n_19024),
.A2(n_8681),
.B(n_8686),
.C(n_8675),
.Y(n_19158)
);

NAND3xp33_ASAP7_75t_L g19159 ( 
.A(n_19041),
.B(n_7596),
.C(n_7463),
.Y(n_19159)
);

NAND3xp33_ASAP7_75t_L g19160 ( 
.A(n_19040),
.B(n_7596),
.C(n_7553),
.Y(n_19160)
);

AOI322xp5_ASAP7_75t_L g19161 ( 
.A1(n_19017),
.A2(n_7013),
.A3(n_7093),
.B1(n_6899),
.B2(n_6873),
.C1(n_6790),
.C2(n_6803),
.Y(n_19161)
);

NOR3xp33_ASAP7_75t_L g19162 ( 
.A(n_19068),
.B(n_6045),
.C(n_6040),
.Y(n_19162)
);

NAND4xp25_ASAP7_75t_SL g19163 ( 
.A(n_19072),
.B(n_6953),
.C(n_6964),
.D(n_6928),
.Y(n_19163)
);

NAND4xp25_ASAP7_75t_L g19164 ( 
.A(n_19037),
.B(n_7227),
.C(n_7235),
.D(n_7186),
.Y(n_19164)
);

NAND2xp5_ASAP7_75t_L g19165 ( 
.A(n_19053),
.B(n_7538),
.Y(n_19165)
);

NOR5xp2_ASAP7_75t_L g19166 ( 
.A(n_18983),
.B(n_6856),
.C(n_6865),
.D(n_6853),
.E(n_6851),
.Y(n_19166)
);

NOR2xp33_ASAP7_75t_L g19167 ( 
.A(n_18977),
.B(n_7227),
.Y(n_19167)
);

NOR2xp67_ASAP7_75t_L g19168 ( 
.A(n_18987),
.B(n_6072),
.Y(n_19168)
);

OAI22xp5_ASAP7_75t_L g19169 ( 
.A1(n_18993),
.A2(n_7235),
.B1(n_7265),
.B2(n_7227),
.Y(n_19169)
);

INVxp33_ASAP7_75t_SL g19170 ( 
.A(n_19043),
.Y(n_19170)
);

BUFx2_ASAP7_75t_L g19171 ( 
.A(n_18981),
.Y(n_19171)
);

AOI211xp5_ASAP7_75t_L g19172 ( 
.A1(n_19005),
.A2(n_7565),
.B(n_7566),
.C(n_7553),
.Y(n_19172)
);

NAND2xp5_ASAP7_75t_L g19173 ( 
.A(n_18964),
.B(n_7553),
.Y(n_19173)
);

NOR2x1_ASAP7_75t_L g19174 ( 
.A(n_18971),
.B(n_7235),
.Y(n_19174)
);

AND2x4_ASAP7_75t_L g19175 ( 
.A(n_18971),
.B(n_7235),
.Y(n_19175)
);

AOI21xp5_ASAP7_75t_SL g19176 ( 
.A1(n_18971),
.A2(n_7565),
.B(n_7553),
.Y(n_19176)
);

AOI22xp5_ASAP7_75t_L g19177 ( 
.A1(n_18972),
.A2(n_7228),
.B1(n_7240),
.B2(n_7209),
.Y(n_19177)
);

NAND4xp25_ASAP7_75t_L g19178 ( 
.A(n_18972),
.B(n_7265),
.C(n_7266),
.D(n_7235),
.Y(n_19178)
);

AOI21xp5_ASAP7_75t_L g19179 ( 
.A1(n_18985),
.A2(n_7816),
.B(n_8253),
.Y(n_19179)
);

NAND3xp33_ASAP7_75t_SL g19180 ( 
.A(n_18971),
.B(n_6072),
.C(n_6045),
.Y(n_19180)
);

NOR3xp33_ASAP7_75t_SL g19181 ( 
.A(n_18971),
.B(n_7261),
.C(n_7248),
.Y(n_19181)
);

NOR2x1_ASAP7_75t_L g19182 ( 
.A(n_18971),
.B(n_7265),
.Y(n_19182)
);

OAI221xp5_ASAP7_75t_L g19183 ( 
.A1(n_18971),
.A2(n_7309),
.B1(n_7362),
.B2(n_7266),
.C(n_7265),
.Y(n_19183)
);

INVx1_ASAP7_75t_L g19184 ( 
.A(n_19175),
.Y(n_19184)
);

INVx1_ASAP7_75t_L g19185 ( 
.A(n_19175),
.Y(n_19185)
);

INVx1_ASAP7_75t_L g19186 ( 
.A(n_19091),
.Y(n_19186)
);

NOR2xp33_ASAP7_75t_L g19187 ( 
.A(n_19170),
.B(n_7265),
.Y(n_19187)
);

AOI22xp5_ASAP7_75t_L g19188 ( 
.A1(n_19082),
.A2(n_7228),
.B1(n_7240),
.B2(n_7209),
.Y(n_19188)
);

XNOR2xp5_ASAP7_75t_L g19189 ( 
.A(n_19103),
.B(n_5376),
.Y(n_19189)
);

XOR2x1_ASAP7_75t_L g19190 ( 
.A(n_19156),
.B(n_19092),
.Y(n_19190)
);

INVx1_ASAP7_75t_L g19191 ( 
.A(n_19099),
.Y(n_19191)
);

OAI21xp5_ASAP7_75t_L g19192 ( 
.A1(n_19085),
.A2(n_7816),
.B(n_7836),
.Y(n_19192)
);

NAND4xp75_ASAP7_75t_L g19193 ( 
.A(n_19088),
.B(n_6706),
.C(n_6803),
.D(n_6790),
.Y(n_19193)
);

NOR3xp33_ASAP7_75t_L g19194 ( 
.A(n_19148),
.B(n_6072),
.C(n_6045),
.Y(n_19194)
);

AOI22xp5_ASAP7_75t_L g19195 ( 
.A1(n_19121),
.A2(n_7228),
.B1(n_7240),
.B2(n_7209),
.Y(n_19195)
);

NAND4xp75_ASAP7_75t_L g19196 ( 
.A(n_19081),
.B(n_6706),
.C(n_6810),
.D(n_6803),
.Y(n_19196)
);

INVx1_ASAP7_75t_L g19197 ( 
.A(n_19171),
.Y(n_19197)
);

INVx1_ASAP7_75t_L g19198 ( 
.A(n_19137),
.Y(n_19198)
);

INVx1_ASAP7_75t_L g19199 ( 
.A(n_19129),
.Y(n_19199)
);

OAI21xp5_ASAP7_75t_L g19200 ( 
.A1(n_19122),
.A2(n_7836),
.B(n_7903),
.Y(n_19200)
);

NAND2xp5_ASAP7_75t_L g19201 ( 
.A(n_19107),
.B(n_7553),
.Y(n_19201)
);

AOI22xp33_ASAP7_75t_L g19202 ( 
.A1(n_19125),
.A2(n_7565),
.B1(n_7566),
.B2(n_7553),
.Y(n_19202)
);

NOR3xp33_ASAP7_75t_L g19203 ( 
.A(n_19153),
.B(n_19080),
.C(n_19127),
.Y(n_19203)
);

OAI22xp5_ASAP7_75t_L g19204 ( 
.A1(n_19096),
.A2(n_7565),
.B1(n_7566),
.B2(n_7553),
.Y(n_19204)
);

INVx1_ASAP7_75t_L g19205 ( 
.A(n_19168),
.Y(n_19205)
);

XNOR2xp5_ASAP7_75t_L g19206 ( 
.A(n_19115),
.B(n_5376),
.Y(n_19206)
);

INVx1_ASAP7_75t_L g19207 ( 
.A(n_19174),
.Y(n_19207)
);

INVx1_ASAP7_75t_L g19208 ( 
.A(n_19182),
.Y(n_19208)
);

INVx2_ASAP7_75t_SL g19209 ( 
.A(n_19173),
.Y(n_19209)
);

NAND4xp75_ASAP7_75t_L g19210 ( 
.A(n_19083),
.B(n_6810),
.C(n_6899),
.D(n_6873),
.Y(n_19210)
);

INVx3_ASAP7_75t_L g19211 ( 
.A(n_19139),
.Y(n_19211)
);

NOR3xp33_ASAP7_75t_L g19212 ( 
.A(n_19108),
.B(n_6119),
.C(n_6072),
.Y(n_19212)
);

NAND4xp75_ASAP7_75t_L g19213 ( 
.A(n_19165),
.B(n_6810),
.C(n_6899),
.D(n_6873),
.Y(n_19213)
);

INVx1_ASAP7_75t_L g19214 ( 
.A(n_19167),
.Y(n_19214)
);

INVx1_ASAP7_75t_L g19215 ( 
.A(n_19160),
.Y(n_19215)
);

NOR2x1_ASAP7_75t_L g19216 ( 
.A(n_19087),
.B(n_7266),
.Y(n_19216)
);

AOI22xp5_ASAP7_75t_L g19217 ( 
.A1(n_19128),
.A2(n_7228),
.B1(n_7240),
.B2(n_7209),
.Y(n_19217)
);

NAND4xp75_ASAP7_75t_L g19218 ( 
.A(n_19157),
.B(n_6810),
.C(n_6899),
.D(n_6873),
.Y(n_19218)
);

OAI221xp5_ASAP7_75t_L g19219 ( 
.A1(n_19172),
.A2(n_7362),
.B1(n_7427),
.B2(n_7309),
.C(n_7266),
.Y(n_19219)
);

XOR2x1_ASAP7_75t_L g19220 ( 
.A(n_19140),
.B(n_7596),
.Y(n_19220)
);

XNOR2x1_ASAP7_75t_L g19221 ( 
.A(n_19143),
.B(n_6290),
.Y(n_19221)
);

INVx1_ASAP7_75t_L g19222 ( 
.A(n_19084),
.Y(n_19222)
);

INVx1_ASAP7_75t_L g19223 ( 
.A(n_19164),
.Y(n_19223)
);

INVx1_ASAP7_75t_L g19224 ( 
.A(n_19123),
.Y(n_19224)
);

NAND2xp5_ASAP7_75t_L g19225 ( 
.A(n_19131),
.B(n_7565),
.Y(n_19225)
);

AND2x2_ASAP7_75t_L g19226 ( 
.A(n_19113),
.B(n_8708),
.Y(n_19226)
);

NOR2x1_ASAP7_75t_L g19227 ( 
.A(n_19176),
.B(n_7266),
.Y(n_19227)
);

AND2x4_ASAP7_75t_L g19228 ( 
.A(n_19159),
.B(n_7565),
.Y(n_19228)
);

AND2x2_ASAP7_75t_L g19229 ( 
.A(n_19142),
.B(n_8708),
.Y(n_19229)
);

XNOR2xp5_ASAP7_75t_L g19230 ( 
.A(n_19132),
.B(n_5376),
.Y(n_19230)
);

INVx1_ASAP7_75t_SL g19231 ( 
.A(n_19146),
.Y(n_19231)
);

INVx1_ASAP7_75t_L g19232 ( 
.A(n_19136),
.Y(n_19232)
);

INVx1_ASAP7_75t_L g19233 ( 
.A(n_19144),
.Y(n_19233)
);

INVx1_ASAP7_75t_L g19234 ( 
.A(n_19163),
.Y(n_19234)
);

NAND2xp5_ASAP7_75t_L g19235 ( 
.A(n_19116),
.B(n_7565),
.Y(n_19235)
);

INVx2_ASAP7_75t_L g19236 ( 
.A(n_19097),
.Y(n_19236)
);

INVx2_ASAP7_75t_L g19237 ( 
.A(n_19120),
.Y(n_19237)
);

AND2x4_ASAP7_75t_L g19238 ( 
.A(n_19133),
.B(n_7566),
.Y(n_19238)
);

OA22x2_ASAP7_75t_L g19239 ( 
.A1(n_19177),
.A2(n_8686),
.B1(n_8691),
.B2(n_8681),
.Y(n_19239)
);

NAND4xp75_ASAP7_75t_L g19240 ( 
.A(n_19124),
.B(n_6962),
.C(n_7013),
.D(n_7004),
.Y(n_19240)
);

NAND4xp75_ASAP7_75t_L g19241 ( 
.A(n_19149),
.B(n_6962),
.C(n_7013),
.D(n_7004),
.Y(n_19241)
);

AOI22xp5_ASAP7_75t_SL g19242 ( 
.A1(n_19141),
.A2(n_7240),
.B1(n_7246),
.B2(n_7228),
.Y(n_19242)
);

NOR2xp33_ASAP7_75t_L g19243 ( 
.A(n_19138),
.B(n_7266),
.Y(n_19243)
);

NOR2xp33_ASAP7_75t_L g19244 ( 
.A(n_19151),
.B(n_7309),
.Y(n_19244)
);

OAI22xp5_ASAP7_75t_L g19245 ( 
.A1(n_19134),
.A2(n_7586),
.B1(n_7566),
.B2(n_7362),
.Y(n_19245)
);

NOR2x1_ASAP7_75t_L g19246 ( 
.A(n_19093),
.B(n_7309),
.Y(n_19246)
);

NOR2xp33_ASAP7_75t_L g19247 ( 
.A(n_19180),
.B(n_7309),
.Y(n_19247)
);

XOR2xp5_ASAP7_75t_L g19248 ( 
.A(n_19094),
.B(n_6290),
.Y(n_19248)
);

INVx1_ASAP7_75t_L g19249 ( 
.A(n_19098),
.Y(n_19249)
);

INVx3_ASAP7_75t_L g19250 ( 
.A(n_19111),
.Y(n_19250)
);

OR2x2_ASAP7_75t_L g19251 ( 
.A(n_19155),
.B(n_7781),
.Y(n_19251)
);

NAND2xp5_ASAP7_75t_L g19252 ( 
.A(n_19181),
.B(n_19161),
.Y(n_19252)
);

NAND2xp5_ASAP7_75t_L g19253 ( 
.A(n_19126),
.B(n_7566),
.Y(n_19253)
);

OR3x1_ASAP7_75t_L g19254 ( 
.A(n_19109),
.B(n_4923),
.C(n_4918),
.Y(n_19254)
);

AND2x4_ASAP7_75t_L g19255 ( 
.A(n_19162),
.B(n_7566),
.Y(n_19255)
);

AO21x1_ASAP7_75t_L g19256 ( 
.A1(n_19118),
.A2(n_7362),
.B(n_7309),
.Y(n_19256)
);

XNOR2xp5_ASAP7_75t_L g19257 ( 
.A(n_19114),
.B(n_7028),
.Y(n_19257)
);

NAND4xp75_ASAP7_75t_L g19258 ( 
.A(n_19152),
.B(n_6962),
.C(n_7013),
.D(n_7004),
.Y(n_19258)
);

NAND2xp5_ASAP7_75t_L g19259 ( 
.A(n_19095),
.B(n_7566),
.Y(n_19259)
);

OAI21xp5_ASAP7_75t_L g19260 ( 
.A1(n_19090),
.A2(n_19135),
.B(n_19150),
.Y(n_19260)
);

INVx2_ASAP7_75t_L g19261 ( 
.A(n_19104),
.Y(n_19261)
);

XNOR2x1_ASAP7_75t_L g19262 ( 
.A(n_19169),
.B(n_6290),
.Y(n_19262)
);

INVx2_ASAP7_75t_SL g19263 ( 
.A(n_19154),
.Y(n_19263)
);

OR2x2_ASAP7_75t_L g19264 ( 
.A(n_19178),
.B(n_7781),
.Y(n_19264)
);

INVx1_ASAP7_75t_L g19265 ( 
.A(n_19110),
.Y(n_19265)
);

INVxp67_ASAP7_75t_L g19266 ( 
.A(n_19130),
.Y(n_19266)
);

NOR2xp67_ASAP7_75t_SL g19267 ( 
.A(n_19183),
.B(n_6290),
.Y(n_19267)
);

NAND2xp5_ASAP7_75t_L g19268 ( 
.A(n_19112),
.B(n_7566),
.Y(n_19268)
);

AND2x4_ASAP7_75t_L g19269 ( 
.A(n_19147),
.B(n_7586),
.Y(n_19269)
);

INVx2_ASAP7_75t_L g19270 ( 
.A(n_19166),
.Y(n_19270)
);

INVxp67_ASAP7_75t_L g19271 ( 
.A(n_19086),
.Y(n_19271)
);

INVx2_ASAP7_75t_L g19272 ( 
.A(n_19100),
.Y(n_19272)
);

INVx1_ASAP7_75t_L g19273 ( 
.A(n_19119),
.Y(n_19273)
);

AO211x2_ASAP7_75t_L g19274 ( 
.A1(n_19198),
.A2(n_19145),
.B(n_19179),
.C(n_19117),
.Y(n_19274)
);

INVx3_ASAP7_75t_L g19275 ( 
.A(n_19228),
.Y(n_19275)
);

AO211x2_ASAP7_75t_L g19276 ( 
.A1(n_19203),
.A2(n_19102),
.B(n_19105),
.C(n_19101),
.Y(n_19276)
);

CKINVDCx20_ASAP7_75t_R g19277 ( 
.A(n_19199),
.Y(n_19277)
);

INVx2_ASAP7_75t_L g19278 ( 
.A(n_19190),
.Y(n_19278)
);

INVx1_ASAP7_75t_L g19279 ( 
.A(n_19189),
.Y(n_19279)
);

NOR2x1_ASAP7_75t_L g19280 ( 
.A(n_19205),
.B(n_19158),
.Y(n_19280)
);

NAND2x1p5_ASAP7_75t_L g19281 ( 
.A(n_19197),
.B(n_19106),
.Y(n_19281)
);

AND2x4_ASAP7_75t_L g19282 ( 
.A(n_19191),
.B(n_19089),
.Y(n_19282)
);

NOR2x1_ASAP7_75t_L g19283 ( 
.A(n_19207),
.B(n_7362),
.Y(n_19283)
);

NAND2xp5_ASAP7_75t_L g19284 ( 
.A(n_19187),
.B(n_7586),
.Y(n_19284)
);

AND2x4_ASAP7_75t_SL g19285 ( 
.A(n_19224),
.B(n_4622),
.Y(n_19285)
);

NOR3xp33_ASAP7_75t_L g19286 ( 
.A(n_19214),
.B(n_6119),
.C(n_6072),
.Y(n_19286)
);

AOI21xp5_ASAP7_75t_L g19287 ( 
.A1(n_19209),
.A2(n_8253),
.B(n_7768),
.Y(n_19287)
);

AND3x2_ASAP7_75t_L g19288 ( 
.A(n_19208),
.B(n_7120),
.C(n_7099),
.Y(n_19288)
);

NOR2xp67_ASAP7_75t_L g19289 ( 
.A(n_19266),
.B(n_6119),
.Y(n_19289)
);

NOR3xp33_ASAP7_75t_L g19290 ( 
.A(n_19215),
.B(n_6133),
.C(n_6119),
.Y(n_19290)
);

NOR4xp25_ASAP7_75t_L g19291 ( 
.A(n_19231),
.B(n_7004),
.C(n_7037),
.D(n_6962),
.Y(n_19291)
);

NAND4xp25_ASAP7_75t_L g19292 ( 
.A(n_19234),
.B(n_6119),
.C(n_6140),
.D(n_6133),
.Y(n_19292)
);

NAND4xp25_ASAP7_75t_L g19293 ( 
.A(n_19186),
.B(n_6133),
.C(n_6143),
.D(n_6140),
.Y(n_19293)
);

INVx1_ASAP7_75t_L g19294 ( 
.A(n_19237),
.Y(n_19294)
);

OAI221xp5_ASAP7_75t_L g19295 ( 
.A1(n_19260),
.A2(n_7446),
.B1(n_7505),
.B2(n_7427),
.C(n_7362),
.Y(n_19295)
);

NOR5xp2_ASAP7_75t_L g19296 ( 
.A(n_19271),
.B(n_6971),
.C(n_7009),
.D(n_6948),
.E(n_6870),
.Y(n_19296)
);

NAND3xp33_ASAP7_75t_SL g19297 ( 
.A(n_19184),
.B(n_6140),
.C(n_6133),
.Y(n_19297)
);

NAND3xp33_ASAP7_75t_SL g19298 ( 
.A(n_19185),
.B(n_6140),
.C(n_6133),
.Y(n_19298)
);

OR5x1_ASAP7_75t_L g19299 ( 
.A(n_19263),
.B(n_8708),
.C(n_8806),
.D(n_8763),
.E(n_8631),
.Y(n_19299)
);

NAND4xp25_ASAP7_75t_L g19300 ( 
.A(n_19223),
.B(n_6140),
.C(n_6168),
.D(n_6143),
.Y(n_19300)
);

INVxp67_ASAP7_75t_SL g19301 ( 
.A(n_19211),
.Y(n_19301)
);

INVx1_ASAP7_75t_L g19302 ( 
.A(n_19270),
.Y(n_19302)
);

NOR2xp67_ASAP7_75t_L g19303 ( 
.A(n_19249),
.B(n_6143),
.Y(n_19303)
);

NOR3xp33_ASAP7_75t_L g19304 ( 
.A(n_19233),
.B(n_6168),
.C(n_6143),
.Y(n_19304)
);

OA22x2_ASAP7_75t_L g19305 ( 
.A1(n_19261),
.A2(n_19236),
.B1(n_19273),
.B2(n_19272),
.Y(n_19305)
);

INVx1_ASAP7_75t_L g19306 ( 
.A(n_19252),
.Y(n_19306)
);

NAND3x1_ASAP7_75t_L g19307 ( 
.A(n_19250),
.B(n_5221),
.C(n_5214),
.Y(n_19307)
);

AND2x2_ASAP7_75t_L g19308 ( 
.A(n_19220),
.B(n_7427),
.Y(n_19308)
);

NOR3xp33_ASAP7_75t_SL g19309 ( 
.A(n_19222),
.B(n_7267),
.C(n_7261),
.Y(n_19309)
);

INVx1_ASAP7_75t_L g19310 ( 
.A(n_19265),
.Y(n_19310)
);

AND5x1_ASAP7_75t_L g19311 ( 
.A(n_19244),
.B(n_7781),
.C(n_7658),
.D(n_7752),
.E(n_8708),
.Y(n_19311)
);

AND5x1_ASAP7_75t_L g19312 ( 
.A(n_19243),
.B(n_7781),
.C(n_7658),
.D(n_7752),
.E(n_8708),
.Y(n_19312)
);

INVx1_ASAP7_75t_L g19313 ( 
.A(n_19232),
.Y(n_19313)
);

NOR3xp33_ASAP7_75t_SL g19314 ( 
.A(n_19253),
.B(n_7269),
.C(n_7267),
.Y(n_19314)
);

NOR3xp33_ASAP7_75t_SL g19315 ( 
.A(n_19268),
.B(n_7304),
.C(n_7269),
.Y(n_19315)
);

OR3x2_ASAP7_75t_L g19316 ( 
.A(n_19251),
.B(n_6733),
.C(n_6599),
.Y(n_19316)
);

NAND4xp25_ASAP7_75t_SL g19317 ( 
.A(n_19201),
.B(n_6928),
.C(n_6964),
.D(n_6953),
.Y(n_19317)
);

NAND4xp75_ASAP7_75t_L g19318 ( 
.A(n_19216),
.B(n_7037),
.C(n_7095),
.D(n_7093),
.Y(n_19318)
);

XNOR2x1_ASAP7_75t_L g19319 ( 
.A(n_19221),
.B(n_6290),
.Y(n_19319)
);

NAND3xp33_ASAP7_75t_L g19320 ( 
.A(n_19267),
.B(n_7596),
.C(n_6320),
.Y(n_19320)
);

OR2x2_ASAP7_75t_L g19321 ( 
.A(n_19259),
.B(n_7781),
.Y(n_19321)
);

NAND2xp5_ASAP7_75t_L g19322 ( 
.A(n_19257),
.B(n_7586),
.Y(n_19322)
);

INVx1_ASAP7_75t_L g19323 ( 
.A(n_19227),
.Y(n_19323)
);

INVx6_ASAP7_75t_L g19324 ( 
.A(n_19255),
.Y(n_19324)
);

NOR4xp75_ASAP7_75t_L g19325 ( 
.A(n_19240),
.B(n_7402),
.C(n_7359),
.D(n_7304),
.Y(n_19325)
);

AOI22xp33_ASAP7_75t_SL g19326 ( 
.A1(n_19238),
.A2(n_7240),
.B1(n_7246),
.B2(n_7228),
.Y(n_19326)
);

AND2x4_ASAP7_75t_L g19327 ( 
.A(n_19246),
.B(n_7586),
.Y(n_19327)
);

NAND4xp25_ASAP7_75t_L g19328 ( 
.A(n_19194),
.B(n_19247),
.C(n_19225),
.D(n_19235),
.Y(n_19328)
);

NOR2x1_ASAP7_75t_L g19329 ( 
.A(n_19218),
.B(n_7427),
.Y(n_19329)
);

INVx1_ASAP7_75t_L g19330 ( 
.A(n_19230),
.Y(n_19330)
);

INVx1_ASAP7_75t_L g19331 ( 
.A(n_19262),
.Y(n_19331)
);

NAND4xp25_ASAP7_75t_SL g19332 ( 
.A(n_19256),
.B(n_6928),
.C(n_6964),
.D(n_6953),
.Y(n_19332)
);

NOR3x1_ASAP7_75t_L g19333 ( 
.A(n_19210),
.B(n_7836),
.C(n_7768),
.Y(n_19333)
);

AND2x4_ASAP7_75t_L g19334 ( 
.A(n_19212),
.B(n_7586),
.Y(n_19334)
);

NAND4xp25_ASAP7_75t_L g19335 ( 
.A(n_19217),
.B(n_6143),
.C(n_6196),
.D(n_6168),
.Y(n_19335)
);

NAND2x1p5_ASAP7_75t_L g19336 ( 
.A(n_19242),
.B(n_6311),
.Y(n_19336)
);

NOR5xp2_ASAP7_75t_L g19337 ( 
.A(n_19219),
.B(n_7027),
.C(n_7057),
.D(n_7005),
.E(n_6957),
.Y(n_19337)
);

INVx1_ASAP7_75t_L g19338 ( 
.A(n_19206),
.Y(n_19338)
);

NAND5xp2_ASAP7_75t_L g19339 ( 
.A(n_19195),
.B(n_7596),
.C(n_5804),
.D(n_7454),
.E(n_7401),
.Y(n_19339)
);

NAND4xp75_ASAP7_75t_L g19340 ( 
.A(n_19229),
.B(n_7093),
.C(n_7095),
.D(n_7037),
.Y(n_19340)
);

NAND4xp25_ASAP7_75t_L g19341 ( 
.A(n_19188),
.B(n_6168),
.C(n_6197),
.D(n_6196),
.Y(n_19341)
);

NOR3xp33_ASAP7_75t_L g19342 ( 
.A(n_19245),
.B(n_6196),
.C(n_6168),
.Y(n_19342)
);

NOR3xp33_ASAP7_75t_L g19343 ( 
.A(n_19241),
.B(n_6197),
.C(n_6196),
.Y(n_19343)
);

NAND2xp5_ASAP7_75t_L g19344 ( 
.A(n_19248),
.B(n_7586),
.Y(n_19344)
);

NAND5xp2_ASAP7_75t_L g19345 ( 
.A(n_19226),
.B(n_7596),
.C(n_7514),
.D(n_7536),
.E(n_7475),
.Y(n_19345)
);

NAND4xp75_ASAP7_75t_L g19346 ( 
.A(n_19200),
.B(n_7093),
.C(n_7095),
.D(n_7037),
.Y(n_19346)
);

NAND2xp5_ASAP7_75t_L g19347 ( 
.A(n_19254),
.B(n_7586),
.Y(n_19347)
);

NOR2x1_ASAP7_75t_L g19348 ( 
.A(n_19213),
.B(n_19258),
.Y(n_19348)
);

NAND5xp2_ASAP7_75t_L g19349 ( 
.A(n_19202),
.B(n_7514),
.C(n_7536),
.D(n_7475),
.E(n_7390),
.Y(n_19349)
);

NAND2xp5_ASAP7_75t_L g19350 ( 
.A(n_19269),
.B(n_7586),
.Y(n_19350)
);

AND2x2_ASAP7_75t_L g19351 ( 
.A(n_19264),
.B(n_7427),
.Y(n_19351)
);

NAND4xp25_ASAP7_75t_SL g19352 ( 
.A(n_19196),
.B(n_7045),
.C(n_7072),
.D(n_7054),
.Y(n_19352)
);

OR3x1_ASAP7_75t_L g19353 ( 
.A(n_19193),
.B(n_4923),
.C(n_4918),
.Y(n_19353)
);

INVx2_ASAP7_75t_L g19354 ( 
.A(n_19204),
.Y(n_19354)
);

NOR4xp75_ASAP7_75t_L g19355 ( 
.A(n_19192),
.B(n_19239),
.C(n_7402),
.D(n_7359),
.Y(n_19355)
);

AOI221x1_ASAP7_75t_L g19356 ( 
.A1(n_19203),
.A2(n_7256),
.B1(n_7264),
.B2(n_7246),
.C(n_7240),
.Y(n_19356)
);

AOI22xp33_ASAP7_75t_L g19357 ( 
.A1(n_19198),
.A2(n_6604),
.B1(n_6614),
.B2(n_6591),
.Y(n_19357)
);

NAND2xp5_ASAP7_75t_L g19358 ( 
.A(n_19187),
.B(n_7427),
.Y(n_19358)
);

NAND3xp33_ASAP7_75t_SL g19359 ( 
.A(n_19277),
.B(n_6197),
.C(n_6196),
.Y(n_19359)
);

OAI221xp5_ASAP7_75t_L g19360 ( 
.A1(n_19278),
.A2(n_7505),
.B1(n_7446),
.B2(n_6240),
.C(n_6241),
.Y(n_19360)
);

AOI32xp33_ASAP7_75t_L g19361 ( 
.A1(n_19302),
.A2(n_7505),
.A3(n_7446),
.B1(n_7028),
.B2(n_6236),
.Y(n_19361)
);

NAND2x1p5_ASAP7_75t_L g19362 ( 
.A(n_19313),
.B(n_6311),
.Y(n_19362)
);

OAI22x1_ASAP7_75t_L g19363 ( 
.A1(n_19301),
.A2(n_7505),
.B1(n_7446),
.B2(n_6236),
.Y(n_19363)
);

NOR4xp25_ASAP7_75t_L g19364 ( 
.A(n_19294),
.B(n_19306),
.C(n_19310),
.D(n_19323),
.Y(n_19364)
);

NOR2xp33_ASAP7_75t_L g19365 ( 
.A(n_19275),
.B(n_7446),
.Y(n_19365)
);

INVx1_ASAP7_75t_L g19366 ( 
.A(n_19305),
.Y(n_19366)
);

NAND2xp5_ASAP7_75t_L g19367 ( 
.A(n_19289),
.B(n_7446),
.Y(n_19367)
);

NAND3xp33_ASAP7_75t_SL g19368 ( 
.A(n_19281),
.B(n_6236),
.C(n_6197),
.Y(n_19368)
);

OAI22xp5_ASAP7_75t_L g19369 ( 
.A1(n_19322),
.A2(n_7505),
.B1(n_6604),
.B2(n_6614),
.Y(n_19369)
);

INVxp33_ASAP7_75t_SL g19370 ( 
.A(n_19280),
.Y(n_19370)
);

OAI21xp5_ASAP7_75t_L g19371 ( 
.A1(n_19279),
.A2(n_7660),
.B(n_7888),
.Y(n_19371)
);

AOI22xp5_ASAP7_75t_L g19372 ( 
.A1(n_19303),
.A2(n_6604),
.B1(n_6614),
.B2(n_6591),
.Y(n_19372)
);

AOI211xp5_ASAP7_75t_L g19373 ( 
.A1(n_19328),
.A2(n_6320),
.B(n_6338),
.C(n_6311),
.Y(n_19373)
);

OAI221xp5_ASAP7_75t_SL g19374 ( 
.A1(n_19330),
.A2(n_6730),
.B1(n_6821),
.B2(n_6666),
.C(n_6626),
.Y(n_19374)
);

NAND3xp33_ASAP7_75t_SL g19375 ( 
.A(n_19338),
.B(n_6236),
.C(n_6197),
.Y(n_19375)
);

INVxp33_ASAP7_75t_SL g19376 ( 
.A(n_19331),
.Y(n_19376)
);

NAND5xp2_ASAP7_75t_L g19377 ( 
.A(n_19308),
.B(n_7545),
.C(n_7571),
.D(n_7536),
.E(n_7514),
.Y(n_19377)
);

INVx1_ASAP7_75t_L g19378 ( 
.A(n_19316),
.Y(n_19378)
);

INVx1_ASAP7_75t_L g19379 ( 
.A(n_19324),
.Y(n_19379)
);

NAND5xp2_ASAP7_75t_L g19380 ( 
.A(n_19351),
.B(n_7545),
.C(n_7571),
.D(n_7536),
.E(n_7514),
.Y(n_19380)
);

AOI211x1_ASAP7_75t_SL g19381 ( 
.A1(n_19354),
.A2(n_6604),
.B(n_6614),
.C(n_6591),
.Y(n_19381)
);

NOR2x1p5_ASAP7_75t_L g19382 ( 
.A(n_19282),
.B(n_19340),
.Y(n_19382)
);

AOI22xp5_ASAP7_75t_L g19383 ( 
.A1(n_19324),
.A2(n_6604),
.B1(n_6614),
.B2(n_6591),
.Y(n_19383)
);

OAI22xp5_ASAP7_75t_L g19384 ( 
.A1(n_19344),
.A2(n_7505),
.B1(n_6604),
.B2(n_6614),
.Y(n_19384)
);

AO22x2_ASAP7_75t_L g19385 ( 
.A1(n_19282),
.A2(n_6240),
.B1(n_6241),
.B2(n_6236),
.Y(n_19385)
);

NAND3xp33_ASAP7_75t_L g19386 ( 
.A(n_19348),
.B(n_19320),
.C(n_19319),
.Y(n_19386)
);

AOI22xp5_ASAP7_75t_L g19387 ( 
.A1(n_19274),
.A2(n_6604),
.B1(n_6614),
.B2(n_6591),
.Y(n_19387)
);

NOR2x1p5_ASAP7_75t_L g19388 ( 
.A(n_19358),
.B(n_6240),
.Y(n_19388)
);

XOR2xp5_ASAP7_75t_L g19389 ( 
.A(n_19276),
.B(n_6311),
.Y(n_19389)
);

INVx2_ASAP7_75t_L g19390 ( 
.A(n_19327),
.Y(n_19390)
);

OAI211xp5_ASAP7_75t_SL g19391 ( 
.A1(n_19284),
.A2(n_7151),
.B(n_7155),
.C(n_7136),
.Y(n_19391)
);

INVx1_ASAP7_75t_L g19392 ( 
.A(n_19355),
.Y(n_19392)
);

INVx1_ASAP7_75t_L g19393 ( 
.A(n_19283),
.Y(n_19393)
);

AOI21xp5_ASAP7_75t_L g19394 ( 
.A1(n_19347),
.A2(n_8253),
.B(n_7768),
.Y(n_19394)
);

AND2x2_ASAP7_75t_L g19395 ( 
.A(n_19314),
.B(n_19285),
.Y(n_19395)
);

OAI221xp5_ASAP7_75t_L g19396 ( 
.A1(n_19350),
.A2(n_19342),
.B1(n_19336),
.B2(n_19329),
.C(n_19321),
.Y(n_19396)
);

INVx2_ASAP7_75t_L g19397 ( 
.A(n_19327),
.Y(n_19397)
);

OR2x2_ASAP7_75t_L g19398 ( 
.A(n_19345),
.B(n_7781),
.Y(n_19398)
);

OAI22xp5_ASAP7_75t_L g19399 ( 
.A1(n_19357),
.A2(n_6604),
.B1(n_6614),
.B2(n_6591),
.Y(n_19399)
);

NAND4xp25_ASAP7_75t_L g19400 ( 
.A(n_19339),
.B(n_6240),
.C(n_6244),
.D(n_6241),
.Y(n_19400)
);

NAND2xp5_ASAP7_75t_L g19401 ( 
.A(n_19334),
.B(n_19315),
.Y(n_19401)
);

INVx1_ASAP7_75t_L g19402 ( 
.A(n_19353),
.Y(n_19402)
);

OAI22xp5_ASAP7_75t_L g19403 ( 
.A1(n_19334),
.A2(n_6604),
.B1(n_6614),
.B2(n_6591),
.Y(n_19403)
);

AOI22xp5_ASAP7_75t_L g19404 ( 
.A1(n_19290),
.A2(n_6616),
.B1(n_6619),
.B2(n_6591),
.Y(n_19404)
);

INVx1_ASAP7_75t_L g19405 ( 
.A(n_19307),
.Y(n_19405)
);

AO22x2_ASAP7_75t_L g19406 ( 
.A1(n_19318),
.A2(n_6241),
.B1(n_6244),
.B2(n_6240),
.Y(n_19406)
);

AND2x4_ASAP7_75t_L g19407 ( 
.A(n_19325),
.B(n_19286),
.Y(n_19407)
);

OAI22xp5_ASAP7_75t_L g19408 ( 
.A1(n_19326),
.A2(n_6616),
.B1(n_6619),
.B2(n_6591),
.Y(n_19408)
);

NAND3xp33_ASAP7_75t_L g19409 ( 
.A(n_19304),
.B(n_6370),
.C(n_6320),
.Y(n_19409)
);

OAI221xp5_ASAP7_75t_L g19410 ( 
.A1(n_19335),
.A2(n_6254),
.B1(n_6278),
.B2(n_6244),
.C(n_6241),
.Y(n_19410)
);

INVx2_ASAP7_75t_L g19411 ( 
.A(n_19346),
.Y(n_19411)
);

NAND5xp2_ASAP7_75t_L g19412 ( 
.A(n_19295),
.B(n_7573),
.C(n_7576),
.D(n_7571),
.E(n_7545),
.Y(n_19412)
);

NAND4xp25_ASAP7_75t_L g19413 ( 
.A(n_19341),
.B(n_6244),
.C(n_6278),
.D(n_6254),
.Y(n_19413)
);

AND2x4_ASAP7_75t_L g19414 ( 
.A(n_19309),
.B(n_6244),
.Y(n_19414)
);

NAND5xp2_ASAP7_75t_L g19415 ( 
.A(n_19343),
.B(n_7573),
.C(n_7576),
.D(n_7571),
.E(n_7545),
.Y(n_19415)
);

OAI221xp5_ASAP7_75t_L g19416 ( 
.A1(n_19297),
.A2(n_19298),
.B1(n_19291),
.B2(n_19292),
.C(n_19300),
.Y(n_19416)
);

HB1xp67_ASAP7_75t_L g19417 ( 
.A(n_19332),
.Y(n_19417)
);

INVx1_ASAP7_75t_L g19418 ( 
.A(n_19352),
.Y(n_19418)
);

INVx1_ASAP7_75t_L g19419 ( 
.A(n_19317),
.Y(n_19419)
);

AND2x4_ASAP7_75t_L g19420 ( 
.A(n_19356),
.B(n_6254),
.Y(n_19420)
);

OAI211xp5_ASAP7_75t_SL g19421 ( 
.A1(n_19337),
.A2(n_7155),
.B(n_7156),
.C(n_7151),
.Y(n_19421)
);

AOI211xp5_ASAP7_75t_SL g19422 ( 
.A1(n_19288),
.A2(n_4880),
.B(n_4902),
.C(n_4869),
.Y(n_19422)
);

NAND4xp25_ASAP7_75t_SL g19423 ( 
.A(n_19349),
.B(n_19287),
.C(n_19296),
.D(n_19293),
.Y(n_19423)
);

NAND4xp25_ASAP7_75t_L g19424 ( 
.A(n_19333),
.B(n_6254),
.C(n_6313),
.D(n_6278),
.Y(n_19424)
);

AOI221xp5_ASAP7_75t_L g19425 ( 
.A1(n_19299),
.A2(n_6635),
.B1(n_6640),
.B2(n_6619),
.C(n_6616),
.Y(n_19425)
);

INVx2_ASAP7_75t_L g19426 ( 
.A(n_19311),
.Y(n_19426)
);

HB1xp67_ASAP7_75t_L g19427 ( 
.A(n_19312),
.Y(n_19427)
);

NOR3xp33_ASAP7_75t_SL g19428 ( 
.A(n_19302),
.B(n_7318),
.C(n_7307),
.Y(n_19428)
);

AOI22xp5_ASAP7_75t_L g19429 ( 
.A1(n_19277),
.A2(n_6619),
.B1(n_6635),
.B2(n_6616),
.Y(n_19429)
);

NOR4xp25_ASAP7_75t_L g19430 ( 
.A(n_19278),
.B(n_7116),
.C(n_6896),
.D(n_6937),
.Y(n_19430)
);

INVx1_ASAP7_75t_L g19431 ( 
.A(n_19278),
.Y(n_19431)
);

AO22x2_ASAP7_75t_L g19432 ( 
.A1(n_19278),
.A2(n_6278),
.B1(n_6313),
.B2(n_6254),
.Y(n_19432)
);

INVx2_ASAP7_75t_L g19433 ( 
.A(n_19278),
.Y(n_19433)
);

NAND3xp33_ASAP7_75t_SL g19434 ( 
.A(n_19277),
.B(n_6313),
.C(n_6278),
.Y(n_19434)
);

AOI221xp5_ASAP7_75t_L g19435 ( 
.A1(n_19364),
.A2(n_6616),
.B1(n_6640),
.B2(n_6635),
.C(n_6619),
.Y(n_19435)
);

OAI221xp5_ASAP7_75t_L g19436 ( 
.A1(n_19389),
.A2(n_6453),
.B1(n_6499),
.B2(n_6439),
.C(n_6313),
.Y(n_19436)
);

INVx1_ASAP7_75t_L g19437 ( 
.A(n_19362),
.Y(n_19437)
);

INVx2_ASAP7_75t_L g19438 ( 
.A(n_19433),
.Y(n_19438)
);

NAND4xp75_ASAP7_75t_L g19439 ( 
.A(n_19366),
.B(n_5837),
.C(n_5905),
.D(n_5846),
.Y(n_19439)
);

NAND2xp5_ASAP7_75t_L g19440 ( 
.A(n_19431),
.B(n_7752),
.Y(n_19440)
);

INVx1_ASAP7_75t_L g19441 ( 
.A(n_19379),
.Y(n_19441)
);

OAI22xp5_ASAP7_75t_L g19442 ( 
.A1(n_19370),
.A2(n_6619),
.B1(n_6635),
.B2(n_6616),
.Y(n_19442)
);

AOI21xp5_ASAP7_75t_L g19443 ( 
.A1(n_19376),
.A2(n_8253),
.B(n_7753),
.Y(n_19443)
);

NAND2xp5_ASAP7_75t_L g19444 ( 
.A(n_19365),
.B(n_7752),
.Y(n_19444)
);

OAI311xp33_ASAP7_75t_L g19445 ( 
.A1(n_19386),
.A2(n_7159),
.A3(n_7174),
.B1(n_7157),
.C1(n_7156),
.Y(n_19445)
);

XNOR2x1_ASAP7_75t_L g19446 ( 
.A(n_19382),
.B(n_6311),
.Y(n_19446)
);

AO22x2_ASAP7_75t_L g19447 ( 
.A1(n_19390),
.A2(n_6439),
.B1(n_6453),
.B2(n_6313),
.Y(n_19447)
);

HB1xp67_ASAP7_75t_L g19448 ( 
.A(n_19417),
.Y(n_19448)
);

NOR2xp33_ASAP7_75t_L g19449 ( 
.A(n_19418),
.B(n_6439),
.Y(n_19449)
);

AND2x4_ASAP7_75t_L g19450 ( 
.A(n_19388),
.B(n_7526),
.Y(n_19450)
);

AOI22xp5_ASAP7_75t_L g19451 ( 
.A1(n_19378),
.A2(n_6619),
.B1(n_6635),
.B2(n_6616),
.Y(n_19451)
);

AOI211xp5_ASAP7_75t_L g19452 ( 
.A1(n_19419),
.A2(n_6320),
.B(n_6338),
.C(n_6311),
.Y(n_19452)
);

AOI22xp5_ASAP7_75t_L g19453 ( 
.A1(n_19392),
.A2(n_6619),
.B1(n_6635),
.B2(n_6616),
.Y(n_19453)
);

OAI22xp5_ASAP7_75t_L g19454 ( 
.A1(n_19426),
.A2(n_6619),
.B1(n_6635),
.B2(n_6616),
.Y(n_19454)
);

INVx2_ASAP7_75t_L g19455 ( 
.A(n_19397),
.Y(n_19455)
);

A2O1A1Ixp33_ASAP7_75t_L g19456 ( 
.A1(n_19411),
.A2(n_19402),
.B(n_19393),
.C(n_19427),
.Y(n_19456)
);

INVx2_ASAP7_75t_L g19457 ( 
.A(n_19395),
.Y(n_19457)
);

AOI31xp33_ASAP7_75t_L g19458 ( 
.A1(n_19405),
.A2(n_5846),
.A3(n_5905),
.B(n_5837),
.Y(n_19458)
);

INVx3_ASAP7_75t_L g19459 ( 
.A(n_19407),
.Y(n_19459)
);

XNOR2x1_ASAP7_75t_L g19460 ( 
.A(n_19401),
.B(n_6311),
.Y(n_19460)
);

INVx2_ASAP7_75t_L g19461 ( 
.A(n_19420),
.Y(n_19461)
);

AOI22xp5_ASAP7_75t_L g19462 ( 
.A1(n_19423),
.A2(n_6640),
.B1(n_6644),
.B2(n_6635),
.Y(n_19462)
);

HB1xp67_ASAP7_75t_L g19463 ( 
.A(n_19396),
.Y(n_19463)
);

AOI22xp5_ASAP7_75t_L g19464 ( 
.A1(n_19416),
.A2(n_6640),
.B1(n_6644),
.B2(n_6635),
.Y(n_19464)
);

OAI321xp33_ASAP7_75t_L g19465 ( 
.A1(n_19424),
.A2(n_19367),
.A3(n_19413),
.B1(n_19400),
.B2(n_19368),
.C(n_19409),
.Y(n_19465)
);

INVx2_ASAP7_75t_L g19466 ( 
.A(n_19414),
.Y(n_19466)
);

AND2x2_ASAP7_75t_L g19467 ( 
.A(n_19428),
.B(n_8708),
.Y(n_19467)
);

NAND2xp5_ASAP7_75t_L g19468 ( 
.A(n_19422),
.B(n_7752),
.Y(n_19468)
);

OAI22x1_ASAP7_75t_L g19469 ( 
.A1(n_19387),
.A2(n_6453),
.B1(n_6499),
.B2(n_6439),
.Y(n_19469)
);

INVx2_ASAP7_75t_L g19470 ( 
.A(n_19406),
.Y(n_19470)
);

AOI22xp5_ASAP7_75t_L g19471 ( 
.A1(n_19375),
.A2(n_6644),
.B1(n_6645),
.B2(n_6640),
.Y(n_19471)
);

OAI211xp5_ASAP7_75t_L g19472 ( 
.A1(n_19421),
.A2(n_6453),
.B(n_6499),
.C(n_6439),
.Y(n_19472)
);

INVxp67_ASAP7_75t_L g19473 ( 
.A(n_19406),
.Y(n_19473)
);

OAI211xp5_ASAP7_75t_SL g19474 ( 
.A1(n_19381),
.A2(n_4880),
.B(n_4902),
.C(n_4869),
.Y(n_19474)
);

OAI211xp5_ASAP7_75t_SL g19475 ( 
.A1(n_19373),
.A2(n_4880),
.B(n_4902),
.C(n_4869),
.Y(n_19475)
);

NOR3xp33_ASAP7_75t_L g19476 ( 
.A(n_19359),
.B(n_6499),
.C(n_6453),
.Y(n_19476)
);

AOI21xp5_ASAP7_75t_L g19477 ( 
.A1(n_19434),
.A2(n_7753),
.B(n_7888),
.Y(n_19477)
);

NOR2xp33_ASAP7_75t_SL g19478 ( 
.A(n_19360),
.B(n_6499),
.Y(n_19478)
);

AND2x2_ASAP7_75t_L g19479 ( 
.A(n_19398),
.B(n_7397),
.Y(n_19479)
);

OAI221xp5_ASAP7_75t_L g19480 ( 
.A1(n_19430),
.A2(n_6504),
.B1(n_6338),
.B2(n_6341),
.C(n_6320),
.Y(n_19480)
);

INVx1_ASAP7_75t_L g19481 ( 
.A(n_19391),
.Y(n_19481)
);

INVx1_ASAP7_75t_L g19482 ( 
.A(n_19415),
.Y(n_19482)
);

AND2x2_ASAP7_75t_SL g19483 ( 
.A(n_19429),
.B(n_6504),
.Y(n_19483)
);

AOI22xp33_ASAP7_75t_L g19484 ( 
.A1(n_19363),
.A2(n_6644),
.B1(n_6645),
.B2(n_6640),
.Y(n_19484)
);

INVx1_ASAP7_75t_L g19485 ( 
.A(n_19412),
.Y(n_19485)
);

INVx2_ASAP7_75t_SL g19486 ( 
.A(n_19432),
.Y(n_19486)
);

AND2x4_ASAP7_75t_L g19487 ( 
.A(n_19383),
.B(n_19372),
.Y(n_19487)
);

NOR3xp33_ASAP7_75t_L g19488 ( 
.A(n_19377),
.B(n_6504),
.C(n_5501),
.Y(n_19488)
);

INVxp33_ASAP7_75t_L g19489 ( 
.A(n_19369),
.Y(n_19489)
);

NAND2xp5_ASAP7_75t_L g19490 ( 
.A(n_19361),
.B(n_7752),
.Y(n_19490)
);

INVx1_ASAP7_75t_L g19491 ( 
.A(n_19432),
.Y(n_19491)
);

O2A1O1Ixp33_ASAP7_75t_L g19492 ( 
.A1(n_19384),
.A2(n_6666),
.B(n_6730),
.C(n_6626),
.Y(n_19492)
);

AOI222xp33_ASAP7_75t_L g19493 ( 
.A1(n_19403),
.A2(n_7397),
.B1(n_7264),
.B2(n_7246),
.C1(n_7270),
.C2(n_7256),
.Y(n_19493)
);

INVx1_ASAP7_75t_L g19494 ( 
.A(n_19385),
.Y(n_19494)
);

INVx1_ASAP7_75t_L g19495 ( 
.A(n_19385),
.Y(n_19495)
);

XOR2x1_ASAP7_75t_L g19496 ( 
.A(n_19408),
.B(n_5837),
.Y(n_19496)
);

OAI22xp5_ASAP7_75t_L g19497 ( 
.A1(n_19404),
.A2(n_6644),
.B1(n_6645),
.B2(n_6640),
.Y(n_19497)
);

XNOR2xp5_ASAP7_75t_L g19498 ( 
.A(n_19448),
.B(n_19410),
.Y(n_19498)
);

INVx1_ASAP7_75t_L g19499 ( 
.A(n_19441),
.Y(n_19499)
);

XNOR2xp5_ASAP7_75t_L g19500 ( 
.A(n_19463),
.B(n_19399),
.Y(n_19500)
);

AO22x2_ASAP7_75t_L g19501 ( 
.A1(n_19438),
.A2(n_19371),
.B1(n_19394),
.B2(n_19380),
.Y(n_19501)
);

XNOR2xp5_ASAP7_75t_L g19502 ( 
.A(n_19459),
.B(n_19457),
.Y(n_19502)
);

INVx1_ASAP7_75t_L g19503 ( 
.A(n_19455),
.Y(n_19503)
);

INVx1_ASAP7_75t_L g19504 ( 
.A(n_19461),
.Y(n_19504)
);

INVx1_ASAP7_75t_L g19505 ( 
.A(n_19446),
.Y(n_19505)
);

INVx1_ASAP7_75t_L g19506 ( 
.A(n_19437),
.Y(n_19506)
);

INVx4_ASAP7_75t_L g19507 ( 
.A(n_19466),
.Y(n_19507)
);

OAI22xp5_ASAP7_75t_L g19508 ( 
.A1(n_19440),
.A2(n_19425),
.B1(n_19374),
.B2(n_6644),
.Y(n_19508)
);

INVxp67_ASAP7_75t_SL g19509 ( 
.A(n_19473),
.Y(n_19509)
);

INVx2_ASAP7_75t_L g19510 ( 
.A(n_19496),
.Y(n_19510)
);

XOR2x2_ASAP7_75t_L g19511 ( 
.A(n_19482),
.B(n_6504),
.Y(n_19511)
);

INVxp67_ASAP7_75t_L g19512 ( 
.A(n_19485),
.Y(n_19512)
);

INVx1_ASAP7_75t_L g19513 ( 
.A(n_19494),
.Y(n_19513)
);

INVx1_ASAP7_75t_L g19514 ( 
.A(n_19495),
.Y(n_19514)
);

XOR2xp5_ASAP7_75t_L g19515 ( 
.A(n_19460),
.B(n_6311),
.Y(n_19515)
);

AOI22x1_ASAP7_75t_L g19516 ( 
.A1(n_19470),
.A2(n_6504),
.B1(n_6320),
.B2(n_6341),
.Y(n_19516)
);

INVx1_ASAP7_75t_L g19517 ( 
.A(n_19491),
.Y(n_19517)
);

XNOR2xp5_ASAP7_75t_L g19518 ( 
.A(n_19481),
.B(n_4843),
.Y(n_19518)
);

XNOR2xp5_ASAP7_75t_L g19519 ( 
.A(n_19489),
.B(n_4843),
.Y(n_19519)
);

AOI22xp33_ASAP7_75t_L g19520 ( 
.A1(n_19449),
.A2(n_6644),
.B1(n_6645),
.B2(n_6640),
.Y(n_19520)
);

INVx1_ASAP7_75t_L g19521 ( 
.A(n_19456),
.Y(n_19521)
);

INVxp67_ASAP7_75t_SL g19522 ( 
.A(n_19486),
.Y(n_19522)
);

INVx1_ASAP7_75t_L g19523 ( 
.A(n_19487),
.Y(n_19523)
);

OA22x2_ASAP7_75t_L g19524 ( 
.A1(n_19479),
.A2(n_8686),
.B1(n_8691),
.B2(n_8681),
.Y(n_19524)
);

OAI22xp5_ASAP7_75t_L g19525 ( 
.A1(n_19490),
.A2(n_6644),
.B1(n_6645),
.B2(n_6640),
.Y(n_19525)
);

INVx1_ASAP7_75t_L g19526 ( 
.A(n_19465),
.Y(n_19526)
);

INVx1_ASAP7_75t_L g19527 ( 
.A(n_19483),
.Y(n_19527)
);

BUFx2_ASAP7_75t_L g19528 ( 
.A(n_19450),
.Y(n_19528)
);

HB1xp67_ASAP7_75t_L g19529 ( 
.A(n_19444),
.Y(n_19529)
);

INVx2_ASAP7_75t_L g19530 ( 
.A(n_19439),
.Y(n_19530)
);

OA22x2_ASAP7_75t_L g19531 ( 
.A1(n_19472),
.A2(n_19468),
.B1(n_19462),
.B2(n_19469),
.Y(n_19531)
);

NOR2x1_ASAP7_75t_L g19532 ( 
.A(n_19474),
.B(n_6338),
.Y(n_19532)
);

INVx1_ASAP7_75t_L g19533 ( 
.A(n_19488),
.Y(n_19533)
);

INVx1_ASAP7_75t_L g19534 ( 
.A(n_19476),
.Y(n_19534)
);

INVxp67_ASAP7_75t_SL g19535 ( 
.A(n_19478),
.Y(n_19535)
);

INVx1_ASAP7_75t_L g19536 ( 
.A(n_19467),
.Y(n_19536)
);

INVx1_ASAP7_75t_L g19537 ( 
.A(n_19458),
.Y(n_19537)
);

AOI22xp5_ASAP7_75t_L g19538 ( 
.A1(n_19435),
.A2(n_6645),
.B1(n_6652),
.B2(n_6644),
.Y(n_19538)
);

INVx1_ASAP7_75t_L g19539 ( 
.A(n_19475),
.Y(n_19539)
);

OAI22xp5_ASAP7_75t_L g19540 ( 
.A1(n_19464),
.A2(n_6652),
.B1(n_6663),
.B2(n_6645),
.Y(n_19540)
);

OAI22x1_ASAP7_75t_L g19541 ( 
.A1(n_19451),
.A2(n_7002),
.B1(n_6923),
.B2(n_6653),
.Y(n_19541)
);

XNOR2x2_ASAP7_75t_L g19542 ( 
.A(n_19442),
.B(n_19436),
.Y(n_19542)
);

NOR2x1_ASAP7_75t_L g19543 ( 
.A(n_19492),
.B(n_6338),
.Y(n_19543)
);

AOI22xp33_ASAP7_75t_L g19544 ( 
.A1(n_19454),
.A2(n_6652),
.B1(n_6663),
.B2(n_6645),
.Y(n_19544)
);

XNOR2x1_ASAP7_75t_L g19545 ( 
.A(n_19453),
.B(n_6320),
.Y(n_19545)
);

OAI22x1_ASAP7_75t_L g19546 ( 
.A1(n_19471),
.A2(n_7002),
.B1(n_6653),
.B2(n_6726),
.Y(n_19546)
);

OAI22x1_ASAP7_75t_L g19547 ( 
.A1(n_19502),
.A2(n_19445),
.B1(n_19452),
.B2(n_19493),
.Y(n_19547)
);

OR2x2_ASAP7_75t_L g19548 ( 
.A(n_19503),
.B(n_19497),
.Y(n_19548)
);

INVx1_ASAP7_75t_SL g19549 ( 
.A(n_19528),
.Y(n_19549)
);

INVx1_ASAP7_75t_L g19550 ( 
.A(n_19499),
.Y(n_19550)
);

OAI22xp33_ASAP7_75t_SL g19551 ( 
.A1(n_19521),
.A2(n_19480),
.B1(n_19477),
.B2(n_19443),
.Y(n_19551)
);

CKINVDCx20_ASAP7_75t_R g19552 ( 
.A(n_19512),
.Y(n_19552)
);

BUFx2_ASAP7_75t_L g19553 ( 
.A(n_19522),
.Y(n_19553)
);

INVx1_ASAP7_75t_L g19554 ( 
.A(n_19509),
.Y(n_19554)
);

AOI22xp5_ASAP7_75t_L g19555 ( 
.A1(n_19523),
.A2(n_19447),
.B1(n_19484),
.B2(n_6652),
.Y(n_19555)
);

INVx1_ASAP7_75t_SL g19556 ( 
.A(n_19513),
.Y(n_19556)
);

NAND2xp5_ASAP7_75t_L g19557 ( 
.A(n_19514),
.B(n_19447),
.Y(n_19557)
);

INVx2_ASAP7_75t_L g19558 ( 
.A(n_19511),
.Y(n_19558)
);

INVx1_ASAP7_75t_L g19559 ( 
.A(n_19517),
.Y(n_19559)
);

INVx2_ASAP7_75t_L g19560 ( 
.A(n_19507),
.Y(n_19560)
);

HB1xp67_ASAP7_75t_L g19561 ( 
.A(n_19506),
.Y(n_19561)
);

INVx1_ASAP7_75t_SL g19562 ( 
.A(n_19504),
.Y(n_19562)
);

BUFx2_ASAP7_75t_L g19563 ( 
.A(n_19501),
.Y(n_19563)
);

INVx1_ASAP7_75t_L g19564 ( 
.A(n_19501),
.Y(n_19564)
);

OAI22x1_ASAP7_75t_SL g19565 ( 
.A1(n_19526),
.A2(n_7002),
.B1(n_6653),
.B2(n_6726),
.Y(n_19565)
);

AOI22xp5_ASAP7_75t_L g19566 ( 
.A1(n_19498),
.A2(n_6652),
.B1(n_6663),
.B2(n_6645),
.Y(n_19566)
);

INVx1_ASAP7_75t_L g19567 ( 
.A(n_19500),
.Y(n_19567)
);

AO22x2_ASAP7_75t_L g19568 ( 
.A1(n_19536),
.A2(n_7397),
.B1(n_7116),
.B2(n_4986),
.Y(n_19568)
);

XOR2xp5_ASAP7_75t_L g19569 ( 
.A(n_19519),
.B(n_6320),
.Y(n_19569)
);

AO22x2_ASAP7_75t_L g19570 ( 
.A1(n_19510),
.A2(n_7397),
.B1(n_7116),
.B2(n_4986),
.Y(n_19570)
);

OAI22x1_ASAP7_75t_L g19571 ( 
.A1(n_19535),
.A2(n_4986),
.B1(n_5057),
.B2(n_4983),
.Y(n_19571)
);

OAI221xp5_ASAP7_75t_L g19572 ( 
.A1(n_19530),
.A2(n_6358),
.B1(n_6370),
.B2(n_6341),
.C(n_6338),
.Y(n_19572)
);

INVx1_ASAP7_75t_L g19573 ( 
.A(n_19531),
.Y(n_19573)
);

CKINVDCx20_ASAP7_75t_R g19574 ( 
.A(n_19529),
.Y(n_19574)
);

INVx2_ASAP7_75t_SL g19575 ( 
.A(n_19542),
.Y(n_19575)
);

NAND2xp5_ASAP7_75t_L g19576 ( 
.A(n_19537),
.B(n_19505),
.Y(n_19576)
);

HB1xp67_ASAP7_75t_L g19577 ( 
.A(n_19533),
.Y(n_19577)
);

AOI22xp5_ASAP7_75t_L g19578 ( 
.A1(n_19534),
.A2(n_6663),
.B1(n_6673),
.B2(n_6652),
.Y(n_19578)
);

OAI22x1_ASAP7_75t_L g19579 ( 
.A1(n_19527),
.A2(n_19518),
.B1(n_19539),
.B2(n_19515),
.Y(n_19579)
);

INVx1_ASAP7_75t_L g19580 ( 
.A(n_19508),
.Y(n_19580)
);

OAI222xp33_ASAP7_75t_L g19581 ( 
.A1(n_19549),
.A2(n_19543),
.B1(n_19525),
.B2(n_19532),
.C1(n_19516),
.C2(n_19538),
.Y(n_19581)
);

OAI221xp5_ASAP7_75t_L g19582 ( 
.A1(n_19575),
.A2(n_19545),
.B1(n_19520),
.B2(n_19544),
.C(n_19540),
.Y(n_19582)
);

OR2x2_ASAP7_75t_L g19583 ( 
.A(n_19553),
.B(n_19546),
.Y(n_19583)
);

AOI21xp5_ASAP7_75t_L g19584 ( 
.A1(n_19561),
.A2(n_19541),
.B(n_19524),
.Y(n_19584)
);

AOI22xp5_ASAP7_75t_L g19585 ( 
.A1(n_19554),
.A2(n_6341),
.B1(n_6358),
.B2(n_6338),
.Y(n_19585)
);

INVx1_ASAP7_75t_SL g19586 ( 
.A(n_19562),
.Y(n_19586)
);

NAND2x1p5_ASAP7_75t_SL g19587 ( 
.A(n_19560),
.B(n_5846),
.Y(n_19587)
);

XNOR2xp5_ASAP7_75t_L g19588 ( 
.A(n_19552),
.B(n_4843),
.Y(n_19588)
);

XNOR2x1_ASAP7_75t_L g19589 ( 
.A(n_19556),
.B(n_19573),
.Y(n_19589)
);

NOR3xp33_ASAP7_75t_L g19590 ( 
.A(n_19559),
.B(n_5501),
.C(n_5057),
.Y(n_19590)
);

NOR3xp33_ASAP7_75t_L g19591 ( 
.A(n_19550),
.B(n_5501),
.C(n_5057),
.Y(n_19591)
);

NOR3xp33_ASAP7_75t_SL g19592 ( 
.A(n_19564),
.B(n_4956),
.C(n_4943),
.Y(n_19592)
);

AOI22xp5_ASAP7_75t_SL g19593 ( 
.A1(n_19574),
.A2(n_19563),
.B1(n_19567),
.B2(n_19577),
.Y(n_19593)
);

NOR4xp25_ASAP7_75t_SL g19594 ( 
.A(n_19580),
.B(n_7120),
.C(n_7121),
.D(n_7099),
.Y(n_19594)
);

INVx1_ASAP7_75t_L g19595 ( 
.A(n_19576),
.Y(n_19595)
);

XNOR2xp5_ASAP7_75t_L g19596 ( 
.A(n_19579),
.B(n_4901),
.Y(n_19596)
);

AOI22xp5_ASAP7_75t_SL g19597 ( 
.A1(n_19551),
.A2(n_6341),
.B1(n_6358),
.B2(n_6338),
.Y(n_19597)
);

OAI222xp33_ASAP7_75t_L g19598 ( 
.A1(n_19548),
.A2(n_7002),
.B1(n_5159),
.B2(n_5057),
.C1(n_5170),
.C2(n_5136),
.Y(n_19598)
);

INVx1_ASAP7_75t_L g19599 ( 
.A(n_19557),
.Y(n_19599)
);

NAND3xp33_ASAP7_75t_SL g19600 ( 
.A(n_19558),
.B(n_5136),
.C(n_4983),
.Y(n_19600)
);

XNOR2xp5_ASAP7_75t_L g19601 ( 
.A(n_19547),
.B(n_4901),
.Y(n_19601)
);

NOR3xp33_ASAP7_75t_L g19602 ( 
.A(n_19555),
.B(n_19569),
.C(n_19566),
.Y(n_19602)
);

AOI22xp5_ASAP7_75t_L g19603 ( 
.A1(n_19571),
.A2(n_6358),
.B1(n_6370),
.B2(n_6341),
.Y(n_19603)
);

OAI221xp5_ASAP7_75t_L g19604 ( 
.A1(n_19586),
.A2(n_19578),
.B1(n_19572),
.B2(n_19568),
.C(n_19565),
.Y(n_19604)
);

INVx1_ASAP7_75t_SL g19605 ( 
.A(n_19589),
.Y(n_19605)
);

INVx1_ASAP7_75t_L g19606 ( 
.A(n_19593),
.Y(n_19606)
);

INVx3_ASAP7_75t_SL g19607 ( 
.A(n_19583),
.Y(n_19607)
);

OAI22xp5_ASAP7_75t_SL g19608 ( 
.A1(n_19595),
.A2(n_19568),
.B1(n_19570),
.B2(n_5540),
.Y(n_19608)
);

OAI22xp5_ASAP7_75t_L g19609 ( 
.A1(n_19601),
.A2(n_19570),
.B1(n_6358),
.B2(n_6370),
.Y(n_19609)
);

XNOR2x1_ASAP7_75t_L g19610 ( 
.A(n_19599),
.B(n_6341),
.Y(n_19610)
);

INVx2_ASAP7_75t_L g19611 ( 
.A(n_19596),
.Y(n_19611)
);

OAI22xp5_ASAP7_75t_L g19612 ( 
.A1(n_19582),
.A2(n_6358),
.B1(n_6370),
.B2(n_6341),
.Y(n_19612)
);

OAI22xp5_ASAP7_75t_SL g19613 ( 
.A1(n_19588),
.A2(n_5540),
.B1(n_5639),
.B2(n_5504),
.Y(n_19613)
);

XNOR2xp5_ASAP7_75t_L g19614 ( 
.A(n_19584),
.B(n_4901),
.Y(n_19614)
);

INVx1_ASAP7_75t_L g19615 ( 
.A(n_19602),
.Y(n_19615)
);

AO22x1_ASAP7_75t_L g19616 ( 
.A1(n_19590),
.A2(n_4820),
.B1(n_4848),
.B2(n_4529),
.Y(n_19616)
);

OAI22xp5_ASAP7_75t_L g19617 ( 
.A1(n_19591),
.A2(n_6370),
.B1(n_6393),
.B2(n_6358),
.Y(n_19617)
);

OR2x2_ASAP7_75t_L g19618 ( 
.A(n_19606),
.B(n_19587),
.Y(n_19618)
);

XNOR2xp5_ASAP7_75t_L g19619 ( 
.A(n_19605),
.B(n_19581),
.Y(n_19619)
);

XNOR2xp5_ASAP7_75t_L g19620 ( 
.A(n_19615),
.B(n_19600),
.Y(n_19620)
);

INVx2_ASAP7_75t_L g19621 ( 
.A(n_19610),
.Y(n_19621)
);

INVx1_ASAP7_75t_L g19622 ( 
.A(n_19607),
.Y(n_19622)
);

NOR2x1p5_ASAP7_75t_L g19623 ( 
.A(n_19611),
.B(n_19592),
.Y(n_19623)
);

AND2x2_ASAP7_75t_L g19624 ( 
.A(n_19614),
.B(n_19594),
.Y(n_19624)
);

XOR2xp5_ASAP7_75t_L g19625 ( 
.A(n_19608),
.B(n_19597),
.Y(n_19625)
);

OAI22xp5_ASAP7_75t_L g19626 ( 
.A1(n_19604),
.A2(n_19585),
.B1(n_19603),
.B2(n_19598),
.Y(n_19626)
);

OR3x1_ASAP7_75t_L g19627 ( 
.A(n_19609),
.B(n_19616),
.C(n_19613),
.Y(n_19627)
);

OAI22xp5_ASAP7_75t_L g19628 ( 
.A1(n_19612),
.A2(n_6370),
.B1(n_6393),
.B2(n_6358),
.Y(n_19628)
);

INVx1_ASAP7_75t_L g19629 ( 
.A(n_19617),
.Y(n_19629)
);

AOI22xp5_ASAP7_75t_SL g19630 ( 
.A1(n_19619),
.A2(n_6393),
.B1(n_6401),
.B2(n_6370),
.Y(n_19630)
);

INVx1_ASAP7_75t_L g19631 ( 
.A(n_19622),
.Y(n_19631)
);

OA21x2_ASAP7_75t_L g19632 ( 
.A1(n_19618),
.A2(n_7753),
.B(n_7780),
.Y(n_19632)
);

AOI21xp5_ASAP7_75t_L g19633 ( 
.A1(n_19620),
.A2(n_6401),
.B(n_6393),
.Y(n_19633)
);

NAND2xp5_ASAP7_75t_L g19634 ( 
.A(n_19621),
.B(n_19624),
.Y(n_19634)
);

AO21x2_ASAP7_75t_L g19635 ( 
.A1(n_19625),
.A2(n_7780),
.B(n_7888),
.Y(n_19635)
);

AOI22xp5_ASAP7_75t_L g19636 ( 
.A1(n_19623),
.A2(n_6401),
.B1(n_6432),
.B2(n_6393),
.Y(n_19636)
);

XNOR2xp5_ASAP7_75t_L g19637 ( 
.A(n_19631),
.B(n_19627),
.Y(n_19637)
);

OAI21xp5_ASAP7_75t_L g19638 ( 
.A1(n_19634),
.A2(n_19626),
.B(n_19629),
.Y(n_19638)
);

INVx2_ASAP7_75t_L g19639 ( 
.A(n_19632),
.Y(n_19639)
);

AOI22xp5_ASAP7_75t_L g19640 ( 
.A1(n_19633),
.A2(n_19628),
.B1(n_6401),
.B2(n_6432),
.Y(n_19640)
);

AOI21xp33_ASAP7_75t_L g19641 ( 
.A1(n_19636),
.A2(n_6401),
.B(n_6393),
.Y(n_19641)
);

NAND3xp33_ASAP7_75t_L g19642 ( 
.A(n_19638),
.B(n_19637),
.C(n_19639),
.Y(n_19642)
);

AOI21xp33_ASAP7_75t_L g19643 ( 
.A1(n_19640),
.A2(n_19630),
.B(n_19635),
.Y(n_19643)
);

NAND2xp5_ASAP7_75t_L g19644 ( 
.A(n_19641),
.B(n_6393),
.Y(n_19644)
);

NAND2xp5_ASAP7_75t_L g19645 ( 
.A(n_19637),
.B(n_6393),
.Y(n_19645)
);

AOI21xp5_ASAP7_75t_L g19646 ( 
.A1(n_19638),
.A2(n_6432),
.B(n_6401),
.Y(n_19646)
);

AOI21xp5_ASAP7_75t_L g19647 ( 
.A1(n_19638),
.A2(n_6432),
.B(n_6401),
.Y(n_19647)
);

AOI21xp5_ASAP7_75t_L g19648 ( 
.A1(n_19642),
.A2(n_6432),
.B(n_6401),
.Y(n_19648)
);

OAI21xp5_ASAP7_75t_L g19649 ( 
.A1(n_19645),
.A2(n_7780),
.B(n_7710),
.Y(n_19649)
);

XNOR2x1_ASAP7_75t_L g19650 ( 
.A(n_19643),
.B(n_6455),
.Y(n_19650)
);

NOR2x1_ASAP7_75t_L g19651 ( 
.A(n_19644),
.B(n_5136),
.Y(n_19651)
);

OAI22xp5_ASAP7_75t_L g19652 ( 
.A1(n_19646),
.A2(n_6455),
.B1(n_6476),
.B2(n_6432),
.Y(n_19652)
);

OAI21xp5_ASAP7_75t_L g19653 ( 
.A1(n_19647),
.A2(n_7710),
.B(n_7701),
.Y(n_19653)
);

INVx2_ASAP7_75t_SL g19654 ( 
.A(n_19650),
.Y(n_19654)
);

INVxp67_ASAP7_75t_L g19655 ( 
.A(n_19651),
.Y(n_19655)
);

INVx1_ASAP7_75t_L g19656 ( 
.A(n_19648),
.Y(n_19656)
);

INVx1_ASAP7_75t_L g19657 ( 
.A(n_19652),
.Y(n_19657)
);

INVx1_ASAP7_75t_L g19658 ( 
.A(n_19653),
.Y(n_19658)
);

INVx1_ASAP7_75t_L g19659 ( 
.A(n_19649),
.Y(n_19659)
);

INVx1_ASAP7_75t_L g19660 ( 
.A(n_19650),
.Y(n_19660)
);

OA21x2_ASAP7_75t_L g19661 ( 
.A1(n_19660),
.A2(n_8007),
.B(n_8000),
.Y(n_19661)
);

XNOR2x1_ASAP7_75t_L g19662 ( 
.A(n_19659),
.B(n_6432),
.Y(n_19662)
);

OAI221xp5_ASAP7_75t_L g19663 ( 
.A1(n_19662),
.A2(n_19655),
.B1(n_19654),
.B2(n_19657),
.C(n_19658),
.Y(n_19663)
);

AOI21xp33_ASAP7_75t_SL g19664 ( 
.A1(n_19663),
.A2(n_19656),
.B(n_19661),
.Y(n_19664)
);

AOI211xp5_ASAP7_75t_L g19665 ( 
.A1(n_19664),
.A2(n_6455),
.B(n_6476),
.C(n_6432),
.Y(n_19665)
);


endmodule