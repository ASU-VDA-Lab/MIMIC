module real_jpeg_24727_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_2),
.A2(n_43),
.B1(n_56),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_2),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_118),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_118),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_2),
.A2(n_63),
.B1(n_68),
.B2(n_118),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_3),
.A2(n_38),
.B1(n_63),
.B2(n_68),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

INVx8_ASAP7_75t_SL g49 ( 
.A(n_5),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_6),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_6),
.B(n_52),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_6),
.A2(n_29),
.B(n_32),
.C(n_245),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_183),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_6),
.B(n_63),
.C(n_66),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_183),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_6),
.A2(n_100),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_6),
.B(n_35),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_7),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_87),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_87),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_7),
.A2(n_63),
.B1(n_68),
.B2(n_87),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_32),
.B1(n_33),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_8),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_8),
.A2(n_44),
.B1(n_55),
.B2(n_173),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_8),
.A2(n_27),
.B1(n_28),
.B2(n_173),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_8),
.A2(n_63),
.B1(n_68),
.B2(n_173),
.Y(n_271)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_54),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_54),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_10),
.A2(n_54),
.B1(n_63),
.B2(n_68),
.Y(n_132)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_12),
.A2(n_55),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g79 ( 
.A(n_12),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_79),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_79),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_12),
.A2(n_63),
.B1(n_68),
.B2(n_79),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_13),
.A2(n_42),
.B1(n_55),
.B2(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_13),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_143),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_143),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_13),
.A2(n_63),
.B1(n_68),
.B2(n_143),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_45),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_14),
.A2(n_45),
.B1(n_63),
.B2(n_68),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_16),
.Y(n_103)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_16),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_16),
.A2(n_101),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_16),
.Y(n_205)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_16),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_16),
.A2(n_101),
.B1(n_270),
.B2(n_272),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_93),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_21),
.B(n_80),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_59),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_39),
.B1(n_57),
.B2(n_58),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_23),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_35),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_24),
.A2(n_35),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_24),
.A2(n_35),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_24),
.B(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_25),
.A2(n_26),
.B1(n_37),
.B2(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_25),
.A2(n_26),
.B1(n_91),
.B2(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_25),
.A2(n_26),
.B1(n_122),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_25),
.A2(n_210),
.B(n_211),
.Y(n_209)
);

OAI21xp33_ASAP7_75t_L g256 ( 
.A1(n_25),
.A2(n_211),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_26),
.A2(n_198),
.B(n_199),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_26),
.A2(n_139),
.B(n_199),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_28),
.B1(n_65),
.B2(n_66),
.Y(n_70)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_27),
.A2(n_30),
.B(n_183),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_28),
.B(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_52)
);

NAND3xp33_ASAP7_75t_SL g194 ( 
.A(n_32),
.B(n_49),
.C(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g193 ( 
.A1(n_33),
.A2(n_48),
.B(n_184),
.C(n_194),
.Y(n_193)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_35),
.B(n_200),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_51),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_43),
.B(n_183),
.Y(n_184)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_44),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_46),
.B(n_116),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_46),
.A2(n_145),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_46),
.A2(n_52),
.B1(n_142),
.B2(n_214),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_51),
.Y(n_46)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_76),
.B1(n_77),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_51),
.A2(n_86),
.B(n_115),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_51),
.B(n_117),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_51),
.A2(n_115),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_56),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_73),
.C(n_75),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_73),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_60),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_85),
.C(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_60),
.A2(n_84),
.B1(n_89),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B(n_71),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_69),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_61),
.A2(n_69),
.B1(n_109),
.B2(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_61),
.B(n_179),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_61),
.A2(n_69),
.B1(n_240),
.B2(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_62),
.A2(n_72),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_62),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_62),
.A2(n_124),
.B1(n_137),
.B2(n_177),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_62),
.B(n_183),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_62),
.A2(n_178),
.B(n_254),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_62)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_63),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_68),
.B(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_69),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_69),
.B(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_76),
.A2(n_141),
.B(n_144),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.C(n_88),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_81),
.A2(n_85),
.B1(n_155),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_85),
.A2(n_152),
.B1(n_153),
.B2(n_155),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_88),
.B(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_89),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI31xp33_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_156),
.A3(n_162),
.B(n_344),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_146),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_96),
.B(n_146),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_119),
.C(n_127),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_97),
.A2(n_119),
.B1(n_120),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_97),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_111),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g147 ( 
.A1(n_98),
.A2(n_99),
.B(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_99),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_99),
.A2(n_107),
.B1(n_108),
.B2(n_112),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_104),
.B(n_106),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_100),
.A2(n_106),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_100),
.A2(n_190),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_100),
.A2(n_132),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_100),
.A2(n_273),
.B(n_279),
.Y(n_293)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_101),
.B(n_248),
.Y(n_247)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_103),
.Y(n_105)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B(n_126),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_123),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_124),
.A2(n_239),
.B(n_241),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_124),
.A2(n_241),
.B(n_268),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_127),
.A2(n_128),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_138),
.C(n_140),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_129),
.A2(n_130),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_131),
.A2(n_134),
.B1(n_135),
.B2(n_316),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_131),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_133),
.B(n_183),
.Y(n_277)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_133),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_133),
.A2(n_247),
.B(n_271),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_138),
.B(n_140),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_149),
.C(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_157),
.A2(n_345),
.B(n_346),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_158),
.B(n_161),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_337),
.B(n_343),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_327),
.B(n_336),
.Y(n_163)
);

O2A1O1Ixp33_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_226),
.B(n_310),
.C(n_326),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_206),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_166),
.B(n_206),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_185),
.C(n_196),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_167),
.A2(n_168),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_180),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_175),
.B2(n_176),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_171),
.B(n_175),
.C(n_180),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B(n_184),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_185),
.A2(n_186),
.B1(n_196),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_192),
.B2(n_193),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_192),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_196),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_201),
.C(n_203),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_204),
.A2(n_205),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_215),
.B1(n_216),
.B2(n_225),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

BUFx24_ASAP7_75t_SL g348 ( 
.A(n_207),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.CI(n_212),
.CON(n_207),
.SN(n_207)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_208),
.B(n_209),
.C(n_212),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_224),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_217),
.B(n_224),
.C(n_225),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_218),
.B(n_223),
.Y(n_324)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_303),
.B(n_309),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_258),
.B(n_302),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_250),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_231),
.B(n_250),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_236),
.B2(n_249),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_232),
.B(n_238),
.C(n_242),
.Y(n_308)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_242),
.B2(n_243),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_244),
.B(n_246),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.C(n_255),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_251),
.B(n_298),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_252),
.A2(n_255),
.B1(n_256),
.B2(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_252),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_296),
.B(n_301),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_286),
.B(n_295),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_274),
.B(n_285),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_269),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_281),
.B(n_284),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_278),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_294),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_294),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_292),
.C(n_293),
.Y(n_300)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_300),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_308),
.Y(n_309)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_325),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_325),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_312),
.B(n_315),
.C(n_317),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_317),
.B2(n_318),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_322),
.C(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_329),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_331),
.B(n_332),
.C(n_335),
.Y(n_342)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_342),
.Y(n_343)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_339),
.Y(n_341)
);


endmodule