module real_aes_6416_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_1), .A2(n_137), .B(n_140), .C(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g164 ( .A1(n_2), .A2(n_165), .B(n_166), .Y(n_164) );
INVx1_ASAP7_75t_L g495 ( .A(n_3), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_4), .B(n_176), .Y(n_175) );
AOI21xp33_ASAP7_75t_L g472 ( .A1(n_5), .A2(n_165), .B(n_473), .Y(n_472) );
AND2x6_ASAP7_75t_L g137 ( .A(n_6), .B(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g240 ( .A(n_7), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_8), .B(n_40), .Y(n_102) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_8), .B(n_40), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_9), .A2(n_264), .B(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_10), .B(n_149), .Y(n_217) );
INVx1_ASAP7_75t_L g477 ( .A(n_11), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_12), .B(n_170), .Y(n_528) );
INVx1_ASAP7_75t_L g129 ( .A(n_13), .Y(n_129) );
INVx1_ASAP7_75t_L g540 ( .A(n_14), .Y(n_540) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_15), .A2(n_184), .B(n_225), .C(n_227), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_16), .B(n_176), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_17), .B(n_466), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_18), .B(n_165), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_19), .B(n_272), .Y(n_271) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_20), .A2(n_170), .B(n_201), .C(n_204), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_21), .B(n_176), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_22), .B(n_149), .Y(n_148) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_23), .A2(n_203), .B(n_227), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g185 ( .A(n_24), .B(n_149), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_25), .Y(n_131) );
INVx1_ASAP7_75t_L g182 ( .A(n_26), .Y(n_182) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_27), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_28), .Y(n_213) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_29), .A2(n_43), .B1(n_448), .B2(n_736), .C1(n_737), .C2(n_740), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_30), .B(n_149), .Y(n_496) );
INVx1_ASAP7_75t_L g269 ( .A(n_31), .Y(n_269) );
INVx1_ASAP7_75t_L g485 ( .A(n_32), .Y(n_485) );
INVx2_ASAP7_75t_L g135 ( .A(n_33), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_34), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g169 ( .A1(n_35), .A2(n_170), .B(n_171), .C(n_173), .Y(n_169) );
INVxp67_ASAP7_75t_L g270 ( .A(n_36), .Y(n_270) );
CKINVDCx14_ASAP7_75t_R g167 ( .A(n_37), .Y(n_167) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_38), .A2(n_140), .B(n_181), .C(n_188), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g506 ( .A1(n_39), .A2(n_137), .B(n_140), .C(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g484 ( .A(n_41), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g114 ( .A1(n_42), .A2(n_115), .B1(n_436), .B2(n_437), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_42), .Y(n_436) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_43), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_44), .A2(n_151), .B(n_238), .C(n_239), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_45), .B(n_149), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_46), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_47), .Y(n_266) );
INVx1_ASAP7_75t_L g199 ( .A(n_48), .Y(n_199) );
CKINVDCx16_ASAP7_75t_R g486 ( .A(n_49), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_50), .B(n_165), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g482 ( .A1(n_51), .A2(n_140), .B1(n_204), .B2(n_483), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_52), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g492 ( .A(n_53), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_54), .A2(n_100), .B1(n_108), .B2(n_744), .Y(n_99) );
CKINVDCx14_ASAP7_75t_R g236 ( .A(n_55), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g475 ( .A1(n_56), .A2(n_173), .B(n_238), .C(n_476), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_57), .Y(n_520) );
INVx1_ASAP7_75t_L g474 ( .A(n_58), .Y(n_474) );
INVx1_ASAP7_75t_L g138 ( .A(n_59), .Y(n_138) );
INVx1_ASAP7_75t_L g128 ( .A(n_60), .Y(n_128) );
INVx1_ASAP7_75t_SL g172 ( .A(n_61), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_62), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_63), .B(n_176), .Y(n_206) );
INVx1_ASAP7_75t_L g144 ( .A(n_64), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_SL g465 ( .A1(n_65), .A2(n_173), .B(n_466), .C(n_467), .Y(n_465) );
INVxp67_ASAP7_75t_L g468 ( .A(n_66), .Y(n_468) );
INVx1_ASAP7_75t_L g107 ( .A(n_67), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_68), .A2(n_165), .B(n_235), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g156 ( .A(n_69), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_70), .A2(n_165), .B(n_222), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_71), .Y(n_488) );
INVx1_ASAP7_75t_L g514 ( .A(n_72), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_73), .B(n_440), .Y(n_445) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_74), .A2(n_264), .B(n_265), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g179 ( .A(n_75), .Y(n_179) );
INVx1_ASAP7_75t_L g223 ( .A(n_76), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_77), .A2(n_137), .B(n_140), .C(n_516), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_78), .A2(n_165), .B(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g226 ( .A(n_79), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_80), .B(n_183), .Y(n_508) );
INVx2_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g216 ( .A(n_82), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_83), .B(n_466), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_84), .A2(n_137), .B(n_140), .C(n_494), .Y(n_493) );
NAND3xp33_ASAP7_75t_SL g103 ( .A(n_85), .B(n_104), .C(n_105), .Y(n_103) );
OR2x2_ASAP7_75t_L g441 ( .A(n_85), .B(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g452 ( .A(n_85), .Y(n_452) );
OR2x2_ASAP7_75t_L g735 ( .A(n_85), .B(n_443), .Y(n_735) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_86), .A2(n_140), .B(n_143), .C(n_153), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_87), .B(n_158), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_88), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g525 ( .A1(n_89), .A2(n_137), .B(n_140), .C(n_526), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_90), .Y(n_532) );
INVx1_ASAP7_75t_L g464 ( .A(n_91), .Y(n_464) );
CKINVDCx16_ASAP7_75t_R g537 ( .A(n_92), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_93), .B(n_183), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_94), .B(n_124), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_95), .B(n_124), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_96), .B(n_107), .Y(n_106) );
INVx2_ASAP7_75t_L g202 ( .A(n_97), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_98), .A2(n_165), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
BUFx2_ASAP7_75t_L g744 ( .A(n_101), .Y(n_744) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_103), .Y(n_101) );
AND2x2_ASAP7_75t_L g443 ( .A(n_104), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
AO21x2_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_113), .B(n_446), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
BUFx3_ASAP7_75t_L g743 ( .A(n_110), .Y(n_743) );
INVx2_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OAI21xp5_ASAP7_75t_SL g113 ( .A1(n_114), .A2(n_438), .B(n_445), .Y(n_113) );
INVx3_ASAP7_75t_L g437 ( .A(n_115), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_115), .A2(n_450), .B1(n_734), .B2(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_SL g115 ( .A(n_116), .B(n_391), .Y(n_115) );
NOR4xp25_ASAP7_75t_L g116 ( .A(n_117), .B(n_328), .C(n_362), .D(n_378), .Y(n_116) );
NAND4xp25_ASAP7_75t_SL g117 ( .A(n_118), .B(n_254), .C(n_292), .D(n_308), .Y(n_117) );
AOI222xp33_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_191), .B1(n_229), .B2(n_242), .C1(n_247), .C2(n_253), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI31xp33_ASAP7_75t_L g424 ( .A1(n_120), .A2(n_425), .A3(n_426), .B(n_428), .Y(n_424) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_159), .Y(n_120) );
AND2x2_ASAP7_75t_L g399 ( .A(n_121), .B(n_161), .Y(n_399) );
BUFx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_SL g246 ( .A(n_122), .Y(n_246) );
AND2x2_ASAP7_75t_L g253 ( .A(n_122), .B(n_177), .Y(n_253) );
AND2x2_ASAP7_75t_L g313 ( .A(n_122), .B(n_162), .Y(n_313) );
AO21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_130), .B(n_155), .Y(n_122) );
INVx3_ASAP7_75t_L g176 ( .A(n_123), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_123), .B(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_123), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_SL g510 ( .A(n_123), .B(n_511), .Y(n_510) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_124), .A2(n_462), .B(n_469), .Y(n_461) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g262 ( .A(n_125), .Y(n_262) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_126), .B(n_127), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B(n_139), .Y(n_130) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_132), .A2(n_158), .B(n_179), .C(n_180), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_132), .A2(n_213), .B(n_214), .Y(n_212) );
OAI22xp33_ASAP7_75t_L g481 ( .A1(n_132), .A2(n_154), .B1(n_482), .B2(n_486), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_132), .A2(n_492), .B(n_493), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g513 ( .A1(n_132), .A2(n_514), .B(n_515), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
AND2x4_ASAP7_75t_L g165 ( .A(n_133), .B(n_137), .Y(n_165) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g187 ( .A(n_134), .Y(n_187) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g205 ( .A(n_135), .Y(n_205) );
INVx1_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_136), .Y(n_147) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx3_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
INVx1_ASAP7_75t_L g466 ( .A(n_136), .Y(n_466) );
INVx4_ASAP7_75t_SL g154 ( .A(n_137), .Y(n_154) );
BUFx3_ASAP7_75t_L g188 ( .A(n_137), .Y(n_188) );
INVx5_ASAP7_75t_L g168 ( .A(n_140), .Y(n_168) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx3_ASAP7_75t_L g152 ( .A(n_141), .Y(n_152) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_148), .C(n_150), .Y(n_143) );
O2A1O1Ixp5_ASAP7_75t_L g215 ( .A1(n_145), .A2(n_150), .B(n_216), .C(n_217), .Y(n_215) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g483 ( .A1(n_146), .A2(n_147), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx4_ASAP7_75t_L g203 ( .A(n_147), .Y(n_203) );
INVx4_ASAP7_75t_L g170 ( .A(n_149), .Y(n_170) );
INVx2_ASAP7_75t_L g238 ( .A(n_149), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_150), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_150), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g227 ( .A(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp33_ASAP7_75t_L g166 ( .A1(n_154), .A2(n_167), .B(n_168), .C(n_169), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_SL g198 ( .A1(n_154), .A2(n_168), .B(n_199), .C(n_200), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_SL g222 ( .A1(n_154), .A2(n_168), .B(n_223), .C(n_224), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_154), .A2(n_168), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_SL g265 ( .A1(n_154), .A2(n_168), .B(n_266), .C(n_267), .Y(n_265) );
O2A1O1Ixp33_ASAP7_75t_L g463 ( .A1(n_154), .A2(n_168), .B(n_464), .C(n_465), .Y(n_463) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_154), .A2(n_168), .B(n_474), .C(n_475), .Y(n_473) );
O2A1O1Ixp33_ASAP7_75t_L g536 ( .A1(n_154), .A2(n_168), .B(n_537), .C(n_538), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx1_ASAP7_75t_L g272 ( .A(n_157), .Y(n_272) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_157), .A2(n_524), .B(n_531), .Y(n_523) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g211 ( .A(n_158), .Y(n_211) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_158), .A2(n_234), .B(n_241), .Y(n_233) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_158), .A2(n_535), .B(n_541), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_159), .B(n_343), .Y(n_342) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_160), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_160), .B(n_257), .Y(n_303) );
AND2x2_ASAP7_75t_L g396 ( .A(n_160), .B(n_336), .Y(n_396) );
OAI321xp33_ASAP7_75t_L g430 ( .A1(n_160), .A2(n_246), .A3(n_403), .B1(n_431), .B2(n_433), .C(n_434), .Y(n_430) );
NAND4xp25_ASAP7_75t_L g434 ( .A(n_160), .B(n_232), .C(n_343), .D(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_177), .Y(n_160) );
AND2x2_ASAP7_75t_L g298 ( .A(n_161), .B(n_244), .Y(n_298) );
AND2x2_ASAP7_75t_L g317 ( .A(n_161), .B(n_246), .Y(n_317) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g245 ( .A(n_162), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g273 ( .A(n_162), .B(n_177), .Y(n_273) );
AND2x2_ASAP7_75t_L g359 ( .A(n_162), .B(n_244), .Y(n_359) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_175), .Y(n_162) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_163), .A2(n_197), .B(n_206), .Y(n_196) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_163), .A2(n_221), .B(n_228), .Y(n_220) );
BUFx2_ASAP7_75t_L g264 ( .A(n_165), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_170), .B(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_174), .Y(n_529) );
OA21x2_ASAP7_75t_L g471 ( .A1(n_176), .A2(n_472), .B(n_478), .Y(n_471) );
INVx3_ASAP7_75t_SL g244 ( .A(n_177), .Y(n_244) );
AND2x2_ASAP7_75t_L g291 ( .A(n_177), .B(n_278), .Y(n_291) );
OR2x2_ASAP7_75t_L g324 ( .A(n_177), .B(n_246), .Y(n_324) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_177), .Y(n_331) );
AND2x2_ASAP7_75t_L g360 ( .A(n_177), .B(n_245), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_177), .B(n_333), .Y(n_375) );
AND2x2_ASAP7_75t_L g407 ( .A(n_177), .B(n_399), .Y(n_407) );
AND2x2_ASAP7_75t_L g416 ( .A(n_177), .B(n_258), .Y(n_416) );
OR2x6_ASAP7_75t_L g177 ( .A(n_178), .B(n_189), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_183), .B(n_185), .C(n_186), .Y(n_181) );
OAI22xp33_ASAP7_75t_L g268 ( .A1(n_183), .A2(n_203), .B1(n_269), .B2(n_270), .Y(n_268) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_183), .A2(n_495), .B(n_496), .C(n_497), .Y(n_494) );
INVx5_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_184), .B(n_240), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_184), .B(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_184), .B(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g267 ( .A(n_187), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_207), .Y(n_192) );
INVx1_ASAP7_75t_SL g384 ( .A(n_193), .Y(n_384) );
INVx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g249 ( .A(n_194), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g231 ( .A(n_195), .B(n_209), .Y(n_231) );
AND2x2_ASAP7_75t_L g320 ( .A(n_195), .B(n_233), .Y(n_320) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g290 ( .A(n_196), .B(n_220), .Y(n_290) );
OR2x2_ASAP7_75t_L g301 ( .A(n_196), .B(n_233), .Y(n_301) );
AND2x2_ASAP7_75t_L g327 ( .A(n_196), .B(n_233), .Y(n_327) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_196), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_203), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_203), .B(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g497 ( .A(n_204), .Y(n_497) );
INVx3_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_207), .B(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_207), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
OR2x2_ASAP7_75t_L g300 ( .A(n_208), .B(n_301), .Y(n_300) );
AOI322xp5_ASAP7_75t_L g386 ( .A1(n_208), .A2(n_290), .A3(n_296), .B1(n_327), .B2(n_377), .C1(n_387), .C2(n_389), .Y(n_386) );
OR2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_220), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_209), .B(n_232), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_209), .B(n_233), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_209), .B(n_250), .Y(n_307) );
AND2x2_ASAP7_75t_L g361 ( .A(n_209), .B(n_327), .Y(n_361) );
INVx1_ASAP7_75t_L g365 ( .A(n_209), .Y(n_365) );
AND2x2_ASAP7_75t_L g377 ( .A(n_209), .B(n_220), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_209), .B(n_249), .Y(n_409) );
INVx4_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g274 ( .A(n_210), .B(n_220), .Y(n_274) );
BUFx3_ASAP7_75t_L g288 ( .A(n_210), .Y(n_288) );
AND3x2_ASAP7_75t_L g370 ( .A(n_210), .B(n_350), .C(n_371), .Y(n_370) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_212), .B(n_218), .Y(n_210) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_211), .B(n_499), .Y(n_498) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_211), .B(n_520), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_211), .B(n_532), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g230 ( .A(n_220), .B(n_231), .C(n_232), .Y(n_230) );
INVx1_ASAP7_75t_SL g250 ( .A(n_220), .Y(n_250) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_220), .Y(n_355) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x2_ASAP7_75t_L g349 ( .A(n_231), .B(n_350), .Y(n_349) );
INVxp67_ASAP7_75t_L g356 ( .A(n_231), .Y(n_356) );
AND2x2_ASAP7_75t_L g394 ( .A(n_232), .B(n_372), .Y(n_394) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
BUFx3_ASAP7_75t_L g275 ( .A(n_233), .Y(n_275) );
AND2x2_ASAP7_75t_L g350 ( .A(n_233), .B(n_250), .Y(n_350) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
OR2x2_ASAP7_75t_L g294 ( .A(n_244), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g413 ( .A(n_244), .B(n_313), .Y(n_413) );
AND2x2_ASAP7_75t_L g427 ( .A(n_244), .B(n_246), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_245), .B(n_258), .Y(n_368) );
AND2x2_ASAP7_75t_L g415 ( .A(n_245), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g278 ( .A(n_246), .B(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g295 ( .A(n_246), .B(n_258), .Y(n_295) );
INVx1_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
AND2x2_ASAP7_75t_L g336 ( .A(n_246), .B(n_258), .Y(n_336) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OAI221xp5_ASAP7_75t_L g378 ( .A1(n_248), .A2(n_379), .B1(n_383), .B2(n_385), .C(n_386), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_249), .B(n_251), .Y(n_248) );
AND2x2_ASAP7_75t_L g282 ( .A(n_249), .B(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_252), .B(n_289), .Y(n_432) );
AOI322xp5_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_274), .A3(n_275), .B1(n_276), .B2(n_282), .C1(n_284), .C2(n_291), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_273), .Y(n_256) );
NAND2x1p5_ASAP7_75t_L g312 ( .A(n_257), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_257), .B(n_323), .Y(n_322) );
O2A1O1Ixp33_ASAP7_75t_L g346 ( .A1(n_257), .A2(n_273), .B(n_347), .C(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_257), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_257), .B(n_317), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_257), .B(n_399), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_257), .B(n_427), .Y(n_426) );
BUFx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_258), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_258), .B(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g388 ( .A(n_258), .B(n_275), .Y(n_388) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_263), .B(n_271), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_260), .A2(n_280), .B(n_281), .Y(n_279) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_260), .A2(n_513), .B(n_519), .Y(n_512) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AOI21xp5_ASAP7_75t_SL g504 ( .A1(n_261), .A2(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_262), .A2(n_481), .B(n_487), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_262), .B(n_488), .Y(n_487) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_262), .A2(n_491), .B(n_498), .Y(n_490) );
INVx1_ASAP7_75t_L g280 ( .A(n_263), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_271), .Y(n_281) );
INVx1_ASAP7_75t_L g363 ( .A(n_273), .Y(n_363) );
OAI31xp33_ASAP7_75t_L g373 ( .A1(n_273), .A2(n_298), .A3(n_374), .B(n_376), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_273), .B(n_279), .Y(n_425) );
INVx1_ASAP7_75t_SL g286 ( .A(n_274), .Y(n_286) );
AND2x2_ASAP7_75t_L g319 ( .A(n_274), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g400 ( .A(n_274), .B(n_401), .Y(n_400) );
OR2x2_ASAP7_75t_L g285 ( .A(n_275), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g310 ( .A(n_275), .Y(n_310) );
AND2x2_ASAP7_75t_L g337 ( .A(n_275), .B(n_290), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_275), .B(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g429 ( .A(n_275), .B(n_377), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_277), .B(n_347), .Y(n_420) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g316 ( .A(n_279), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g334 ( .A(n_279), .Y(n_334) );
NAND2xp33_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
OAI211xp5_ASAP7_75t_SL g328 ( .A1(n_286), .A2(n_329), .B(n_335), .C(n_351), .Y(n_328) );
OR2x2_ASAP7_75t_L g403 ( .A(n_286), .B(n_384), .Y(n_403) );
OR2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_288), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_288), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g309 ( .A(n_290), .B(n_310), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_296), .B(n_299), .C(n_302), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_SL g343 ( .A(n_295), .Y(n_343) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_298), .B(n_336), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_298), .Y(n_347) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g306 ( .A(n_301), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g339 ( .A(n_301), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g401 ( .A(n_301), .Y(n_401) );
AOI21xp33_ASAP7_75t_SL g302 ( .A1(n_303), .A2(n_304), .B(n_306), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_304), .A2(n_315), .B(n_318), .Y(n_314) );
AOI211xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B(n_314), .C(n_321), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_309), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_312), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_SL g325 ( .A(n_313), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_315), .A2(n_381), .B(n_382), .Y(n_380) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_320), .B(n_333), .Y(n_332) );
INVx1_ASAP7_75t_SL g345 ( .A(n_320), .Y(n_345) );
AOI21xp33_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_325), .B(n_326), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g376 ( .A(n_327), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_333), .B(n_359), .Y(n_385) );
AND2x2_ASAP7_75t_L g398 ( .A(n_333), .B(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g412 ( .A(n_333), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g422 ( .A(n_333), .B(n_360), .Y(n_422) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_337), .B(n_338), .C(n_346), .Y(n_335) );
INVx1_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
OAI22xp33_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_341), .B1(n_342), .B2(n_344), .Y(n_338) );
OR2x2_ASAP7_75t_L g344 ( .A(n_340), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_340), .B(n_401), .Y(n_423) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g417 ( .A(n_350), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_357), .B1(n_360), .B2(n_361), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g435 ( .A(n_355), .Y(n_435) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g381 ( .A(n_359), .Y(n_381) );
OAI211xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_364), .B(n_366), .C(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVxp67_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_381), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR5xp2_ASAP7_75t_L g391 ( .A(n_392), .B(n_410), .C(n_418), .D(n_424), .E(n_430), .Y(n_391) );
OAI211xp5_ASAP7_75t_SL g392 ( .A1(n_393), .A2(n_395), .B(n_397), .C(n_404), .Y(n_392) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B(n_402), .Y(n_397) );
OAI21xp33_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_407), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_407), .B(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .B(n_417), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g433 ( .A(n_413), .Y(n_433) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_421), .B(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_437), .A2(n_450), .B1(n_453), .B2(n_734), .Y(n_449) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2x2_ASAP7_75t_L g739 ( .A(n_442), .B(n_452), .Y(n_739) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g451 ( .A(n_443), .B(n_452), .Y(n_451) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_445), .A2(n_447), .B(n_743), .Y(n_446) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g742 ( .A(n_453), .Y(n_742) );
INVx3_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND4x1_ASAP7_75t_L g454 ( .A(n_455), .B(n_652), .C(n_699), .D(n_719), .Y(n_454) );
NOR3xp33_ASAP7_75t_SL g455 ( .A(n_456), .B(n_582), .C(n_607), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_457), .A2(n_500), .B(n_542), .C(n_572), .Y(n_456) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_479), .Y(n_458) );
INVx3_ASAP7_75t_SL g624 ( .A(n_459), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_459), .B(n_555), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_459), .B(n_489), .Y(n_705) );
AND2x2_ASAP7_75t_L g728 ( .A(n_459), .B(n_594), .Y(n_728) );
AND2x4_ASAP7_75t_L g459 ( .A(n_460), .B(n_470), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g546 ( .A(n_461), .B(n_471), .Y(n_546) );
INVx3_ASAP7_75t_L g559 ( .A(n_461), .Y(n_559) );
AND2x2_ASAP7_75t_L g564 ( .A(n_461), .B(n_470), .Y(n_564) );
OR2x2_ASAP7_75t_L g615 ( .A(n_461), .B(n_556), .Y(n_615) );
BUFx2_ASAP7_75t_L g635 ( .A(n_461), .Y(n_635) );
AND2x2_ASAP7_75t_L g645 ( .A(n_461), .B(n_556), .Y(n_645) );
AND2x2_ASAP7_75t_L g651 ( .A(n_461), .B(n_480), .Y(n_651) );
INVx1_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_471), .B(n_556), .Y(n_570) );
INVx2_ASAP7_75t_L g580 ( .A(n_471), .Y(n_580) );
AND2x2_ASAP7_75t_L g593 ( .A(n_471), .B(n_559), .Y(n_593) );
OR2x2_ASAP7_75t_L g604 ( .A(n_471), .B(n_556), .Y(n_604) );
AND2x2_ASAP7_75t_SL g650 ( .A(n_471), .B(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g662 ( .A(n_471), .Y(n_662) );
AND2x2_ASAP7_75t_L g708 ( .A(n_471), .B(n_480), .Y(n_708) );
INVx3_ASAP7_75t_SL g581 ( .A(n_479), .Y(n_581) );
OR2x2_ASAP7_75t_L g634 ( .A(n_479), .B(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g479 ( .A(n_480), .B(n_489), .Y(n_479) );
INVx3_ASAP7_75t_L g556 ( .A(n_480), .Y(n_556) );
AND2x2_ASAP7_75t_L g623 ( .A(n_480), .B(n_490), .Y(n_623) );
HB1xp67_ASAP7_75t_L g691 ( .A(n_480), .Y(n_691) );
AOI33xp33_ASAP7_75t_L g695 ( .A1(n_480), .A2(n_624), .A3(n_631), .B1(n_640), .B2(n_696), .B3(n_697), .Y(n_695) );
INVx1_ASAP7_75t_L g544 ( .A(n_489), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_489), .B(n_559), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g618 ( .A(n_489), .B(n_619), .C(n_621), .Y(n_618) );
AND2x2_ASAP7_75t_L g644 ( .A(n_489), .B(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_489), .B(n_651), .Y(n_654) );
AND2x2_ASAP7_75t_L g707 ( .A(n_489), .B(n_708), .Y(n_707) );
INVx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx3_ASAP7_75t_L g563 ( .A(n_490), .Y(n_563) );
OR2x2_ASAP7_75t_L g657 ( .A(n_490), .B(n_556), .Y(n_657) );
OR2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_521), .Y(n_500) );
AOI32xp33_ASAP7_75t_L g608 ( .A1(n_501), .A2(n_609), .A3(n_611), .B1(n_613), .B2(n_616), .Y(n_608) );
NOR2xp67_ASAP7_75t_L g681 ( .A(n_501), .B(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g711 ( .A(n_501), .Y(n_711) );
INVx4_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g643 ( .A(n_502), .B(n_627), .Y(n_643) );
AND2x2_ASAP7_75t_L g663 ( .A(n_502), .B(n_589), .Y(n_663) );
AND2x2_ASAP7_75t_L g731 ( .A(n_502), .B(n_649), .Y(n_731) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_512), .Y(n_502) );
INVx3_ASAP7_75t_L g552 ( .A(n_503), .Y(n_552) );
AND2x2_ASAP7_75t_L g566 ( .A(n_503), .B(n_550), .Y(n_566) );
OR2x2_ASAP7_75t_L g571 ( .A(n_503), .B(n_549), .Y(n_571) );
INVx1_ASAP7_75t_L g578 ( .A(n_503), .Y(n_578) );
AND2x2_ASAP7_75t_L g586 ( .A(n_503), .B(n_560), .Y(n_586) );
AND2x2_ASAP7_75t_L g588 ( .A(n_503), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_503), .B(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g641 ( .A(n_503), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_503), .B(n_726), .Y(n_725) );
OR2x6_ASAP7_75t_L g503 ( .A(n_504), .B(n_510), .Y(n_503) );
INVx2_ASAP7_75t_L g550 ( .A(n_512), .Y(n_550) );
AND2x2_ASAP7_75t_L g596 ( .A(n_512), .B(n_522), .Y(n_596) );
AND2x2_ASAP7_75t_L g606 ( .A(n_512), .B(n_534), .Y(n_606) );
INVx2_ASAP7_75t_L g726 ( .A(n_521), .Y(n_726) );
OR2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_533), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_522), .B(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g567 ( .A(n_522), .Y(n_567) );
AND2x2_ASAP7_75t_L g611 ( .A(n_522), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g627 ( .A(n_522), .B(n_590), .Y(n_627) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g575 ( .A(n_523), .Y(n_575) );
AND2x2_ASAP7_75t_L g589 ( .A(n_523), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g640 ( .A(n_523), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_523), .B(n_550), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_530), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
AND2x2_ASAP7_75t_L g551 ( .A(n_533), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g612 ( .A(n_533), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_533), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g649 ( .A(n_533), .Y(n_649) );
INVx1_ASAP7_75t_L g682 ( .A(n_533), .Y(n_682) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g560 ( .A(n_534), .B(n_550), .Y(n_560) );
INVx1_ASAP7_75t_L g590 ( .A(n_534), .Y(n_590) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_547), .B1(n_553), .B2(n_560), .C(n_561), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_544), .B(n_564), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_544), .B(n_627), .Y(n_704) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_546), .B(n_594), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_546), .B(n_555), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_546), .B(n_569), .Y(n_698) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_551), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g620 ( .A(n_550), .Y(n_620) );
AND2x2_ASAP7_75t_L g595 ( .A(n_551), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g673 ( .A(n_551), .Y(n_673) );
AND2x2_ASAP7_75t_L g605 ( .A(n_552), .B(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_552), .B(n_575), .Y(n_621) );
AND2x2_ASAP7_75t_L g685 ( .A(n_552), .B(n_611), .Y(n_685) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g594 ( .A(n_556), .B(n_563), .Y(n_594) );
AND2x2_ASAP7_75t_L g690 ( .A(n_557), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_559), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_560), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_560), .B(n_567), .Y(n_655) );
AND2x2_ASAP7_75t_L g675 ( .A(n_560), .B(n_575), .Y(n_675) );
AND2x2_ASAP7_75t_L g696 ( .A(n_560), .B(n_640), .Y(n_696) );
OAI32xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_565), .A3(n_567), .B1(n_568), .B2(n_571), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_SL g569 ( .A(n_563), .Y(n_569) );
NAND2x1_ASAP7_75t_L g610 ( .A(n_563), .B(n_593), .Y(n_610) );
OR2x2_ASAP7_75t_L g614 ( .A(n_563), .B(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_563), .B(n_662), .Y(n_715) );
INVx1_ASAP7_75t_L g583 ( .A(n_564), .Y(n_583) );
OAI221xp5_ASAP7_75t_SL g701 ( .A1(n_565), .A2(n_656), .B1(n_702), .B2(n_705), .C(n_706), .Y(n_701) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g573 ( .A(n_566), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g616 ( .A(n_566), .B(n_589), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_566), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g694 ( .A(n_566), .B(n_627), .Y(n_694) );
INVxp67_ASAP7_75t_L g630 ( .A(n_567), .Y(n_630) );
OR2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
AND2x2_ASAP7_75t_L g700 ( .A(n_569), .B(n_687), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_569), .B(n_650), .Y(n_723) );
INVx1_ASAP7_75t_L g598 ( .A(n_571), .Y(n_598) );
NAND2xp5_ASAP7_75t_SL g679 ( .A(n_571), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g716 ( .A(n_571), .B(n_717), .Y(n_716) );
OAI21xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_576), .B(n_579), .Y(n_572) );
AND2x2_ASAP7_75t_L g585 ( .A(n_574), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x2_ASAP7_75t_L g669 ( .A(n_578), .B(n_589), .Y(n_669) );
AND2x2_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
AND2x2_ASAP7_75t_L g687 ( .A(n_580), .B(n_645), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_580), .B(n_644), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_581), .B(n_593), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_584), .B(n_587), .C(n_597), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_583), .A2(n_618), .B1(n_622), .B2(n_625), .C(n_628), .Y(n_617) );
AOI31xp33_ASAP7_75t_L g712 ( .A1(n_583), .A2(n_713), .A3(n_714), .B(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_591), .B1(n_593), .B2(n_595), .Y(n_587) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g713 ( .A(n_593), .Y(n_713) );
INVx1_ASAP7_75t_L g676 ( .A(n_594), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g719 ( .A1(n_596), .A2(n_720), .B(n_722), .C(n_724), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B1(n_601), .B2(n_605), .Y(n_597) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_602), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI221xp5_ASAP7_75t_SL g692 ( .A1(n_604), .A2(n_638), .B1(n_657), .B2(n_693), .C(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g688 ( .A(n_605), .Y(n_688) );
INVx1_ASAP7_75t_L g642 ( .A(n_606), .Y(n_642) );
NAND3xp33_ASAP7_75t_SL g607 ( .A(n_608), .B(n_617), .C(n_632), .Y(n_607) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_609), .A2(n_659), .B(n_663), .Y(n_658) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_611), .B(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g718 ( .A(n_612), .Y(n_718) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g656 ( .A(n_619), .B(n_639), .Y(n_656) );
INVx1_ASAP7_75t_L g631 ( .A(n_620), .Y(n_631) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g629 ( .A(n_623), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_623), .B(n_661), .Y(n_660) );
NOR4xp25_ASAP7_75t_L g628 ( .A(n_624), .B(n_629), .C(n_630), .D(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_637), .B1(n_643), .B2(n_644), .C1(n_646), .C2(n_650), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx1_ASAP7_75t_L g730 ( .A(n_634), .Y(n_730) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_646), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_651), .A2(n_707), .B(n_709), .Y(n_706) );
NOR4xp25_ASAP7_75t_L g652 ( .A(n_653), .B(n_664), .C(n_677), .D(n_692), .Y(n_652) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_655), .B1(n_656), .B2(n_657), .C(n_658), .Y(n_653) );
INVx1_ASAP7_75t_L g733 ( .A(n_654), .Y(n_733) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_661), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
OAI222xp33_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_668), .B1(n_670), .B2(n_671), .C1(n_674), .C2(n_676), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_669), .A2(n_700), .B(n_701), .C(n_712), .Y(n_699) );
OR2x2_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
INVx1_ASAP7_75t_SL g674 ( .A(n_675), .Y(n_674) );
OAI222xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_683), .B1(n_684), .B2(n_686), .C1(n_688), .C2(n_689), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_694), .A2(n_697), .B1(n_730), .B2(n_731), .Y(n_729) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OAI211xp5_ASAP7_75t_SL g724 ( .A1(n_725), .A2(n_727), .B(n_729), .C(n_732), .Y(n_724) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx2_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
endmodule