module real_jpeg_23889_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_0),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_0),
.B(n_41),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_0),
.B(n_50),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_0),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_0),
.B(n_85),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_0),
.B(n_99),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_0),
.B(n_226),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_1),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_1),
.B(n_41),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_50),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_1),
.B(n_47),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_1),
.B(n_85),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_1),
.B(n_99),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_1),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_1),
.B(n_204),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_3),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_3),
.B(n_41),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_3),
.B(n_50),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_3),
.B(n_47),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_3),
.B(n_85),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_3),
.B(n_99),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_3),
.B(n_131),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_3),
.B(n_204),
.Y(n_374)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_5),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_41),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_5),
.B(n_50),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_5),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_5),
.B(n_99),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_5),
.B(n_131),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_5),
.B(n_204),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_7),
.B(n_119),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_7),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_7),
.B(n_50),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_47),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_7),
.B(n_85),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_7),
.B(n_99),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_7),
.B(n_131),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_7),
.B(n_204),
.Y(n_361)
);

INVx8_ASAP7_75t_SL g132 ( 
.A(n_8),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_10),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_10),
.B(n_17),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_10),
.B(n_50),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_10),
.B(n_47),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_10),
.B(n_85),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_10),
.B(n_99),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_10),
.B(n_131),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_10),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_11),
.B(n_41),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_11),
.B(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_11),
.B(n_47),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_11),
.B(n_85),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_11),
.B(n_99),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_11),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_11),
.B(n_226),
.Y(n_272)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_12),
.Y(n_163)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_13),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_13),
.B(n_50),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_13),
.B(n_85),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_13),
.B(n_99),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_13),
.B(n_162),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_15),
.B(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_15),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_15),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_15),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_15),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_16),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_85),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_16),
.B(n_99),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_16),
.B(n_131),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_16),
.B(n_204),
.Y(n_203)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_17),
.Y(n_111)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_380),
.B(n_381),
.C(n_385),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_370),
.C(n_379),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_355),
.C(n_356),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_333),
.C(n_334),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_303),
.C(n_304),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_278),
.C(n_279),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_246),
.C(n_247),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_208),
.C(n_209),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_169),
.C(n_170),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_136),
.C(n_137),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_113),
.C(n_114),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_90),
.C(n_91),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_67),
.C(n_68),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_52),
.C(n_57),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_44),
.B2(n_45),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_46),
.C(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_36),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_36),
.Y(n_43)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_43),
.Y(n_71)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_41),
.Y(n_200)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_47),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.C(n_62),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_60),
.B(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_66),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_66),
.B(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_73),
.C(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_73)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_79),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_89),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_84),
.Y(n_88)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_85),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_88),
.C(n_89),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_102),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_94),
.C(n_102),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_105),
.C(n_106),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_112),
.Y(n_106)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_107),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_108),
.B(n_112),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_128),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_129),
.C(n_135),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_124),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_123),
.C(n_124),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_120),
.B(n_122),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g391 ( 
.A(n_124),
.Y(n_391)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_126),
.CI(n_127),
.CON(n_124),
.SN(n_124)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_126),
.C(n_127),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_135),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_129),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_133),
.CI(n_134),
.CON(n_129),
.SN(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_131),
.Y(n_221)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_152),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_140),
.B(n_141),
.C(n_152),
.Y(n_169)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_148),
.C(n_151),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g389 ( 
.A(n_143),
.Y(n_389)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.CI(n_146),
.CON(n_143),
.SN(n_143)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_144),
.B(n_145),
.C(n_146),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_159),
.C(n_167),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_159),
.B1(n_167),
.B2(n_168),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B(n_158),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_158),
.B(n_195),
.C(n_196),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_164),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_165),
.C(n_166),
.Y(n_190)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_172),
.B1(n_191),
.B2(n_207),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_192),
.C(n_193),
.Y(n_208)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_175),
.C(n_184),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_184),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_176),
.B(n_180),
.C(n_183),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_178),
.B(n_231),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_182),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_190),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_189),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_186),
.B(n_189),
.C(n_190),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_188),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_201),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_200),
.B(n_231),
.Y(n_256)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_244),
.B2(n_245),
.Y(n_209)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_211),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_235),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_235),
.C(n_244),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_222),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_213),
.B(n_223),
.C(n_224),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_214),
.B(n_217),
.C(n_219),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_215),
.B(n_221),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_221),
.B(n_231),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_227),
.B1(n_228),
.B2(n_234),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_225),
.Y(n_234)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_229),
.A2(n_230),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_233),
.C(n_234),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_229),
.B(n_253),
.C(n_256),
.Y(n_301)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_238),
.C(n_239),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_250),
.C(n_277),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_264),
.B2(n_277),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_258),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_259),
.C(n_260),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_256),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_256),
.A2(n_257),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_SL g318 ( 
.A(n_256),
.B(n_283),
.C(n_286),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_260),
.Y(n_387)
);

FAx1_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.CI(n_263),
.CON(n_260),
.SN(n_260)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_267),
.C(n_268),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_271),
.B2(n_276),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_269),
.B(n_272),
.C(n_274),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_272),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_273),
.A2(n_274),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_300),
.C(n_301),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_302),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_293),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_293),
.C(n_302),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_288),
.C(n_289),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_285),
.A2(n_286),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_SL g344 ( 
.A(n_286),
.B(n_311),
.C(n_313),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_289),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.CI(n_292),
.CON(n_289),
.SN(n_289)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_291),
.C(n_292),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_296),
.C(n_297),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_299),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_307),
.C(n_320),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_319),
.B2(n_320),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_315),
.B2(n_316),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_317),
.C(n_318),
.Y(n_336)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_313),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_313),
.A2(n_314),
.B1(n_348),
.B2(n_349),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_313),
.B(n_349),
.C(n_350),
.Y(n_362)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_323),
.C(n_326),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_323),
.A2(n_324),
.B1(n_325),
.B2(n_326),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_327),
.B(n_329),
.C(n_332),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_330),
.B1(n_331),
.B2(n_332),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_330),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_331),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_352),
.B1(n_353),
.B2(n_354),
.Y(n_334)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_337),
.C(n_354),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_343),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_344),
.C(n_345),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_359),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_339),
.B(n_357),
.C(n_359),
.Y(n_379)
);

FAx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.CI(n_342),
.CON(n_339),
.SN(n_339)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_346),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_347),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_348),
.A2(n_349),
.B1(n_366),
.B2(n_367),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_349),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_349),
.B(n_366),
.C(n_369),
.Y(n_372)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_352),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_362),
.C(n_363),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_368),
.B2(n_369),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_365),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_366),
.A2(n_367),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_SL g386 ( 
.A(n_367),
.B(n_374),
.C(n_377),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_368),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_378),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_372),
.B(n_373),
.C(n_378),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_376),
.A2(n_377),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_377),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_383),
.B(n_386),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_384),
.Y(n_385)
);


endmodule