module fake_jpeg_7470_n_257 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_257);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_257;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_6),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_0),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_39),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_51),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_19),
.B1(n_18),
.B2(n_33),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_50),
.A2(n_52),
.B1(n_30),
.B2(n_22),
.Y(n_88)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_19),
.B1(n_18),
.B2(n_31),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_19),
.B1(n_18),
.B2(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_53),
.A2(n_27),
.B1(n_31),
.B2(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_59),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_39),
.B(n_27),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_37),
.A2(n_18),
.B1(n_34),
.B2(n_26),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_60),
.A2(n_27),
.B1(n_20),
.B2(n_30),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_21),
.B(n_20),
.C(n_26),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_29),
.Y(n_69)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_59),
.B(n_22),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_55),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_24),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_74),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_43),
.B1(n_24),
.B2(n_33),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_73),
.A2(n_88),
.B1(n_32),
.B2(n_17),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_65),
.B(n_24),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_78),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_81),
.B1(n_63),
.B2(n_46),
.Y(n_99)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g83 ( 
.A(n_57),
.B(n_22),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_17),
.A3(n_28),
.B1(n_3),
.B2(n_4),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_43),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_85),
.B(n_90),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_91),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_SL g89 ( 
.A1(n_61),
.A2(n_17),
.B(n_32),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_22),
.B(n_32),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_61),
.B(n_51),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_28),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_101),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_109),
.B(n_111),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_55),
.C(n_62),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_107),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_87),
.A2(n_63),
.B1(n_64),
.B2(n_54),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_97),
.A2(n_104),
.B1(n_70),
.B2(n_72),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_102),
.B1(n_78),
.B2(n_75),
.Y(n_125)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_67),
.B1(n_46),
.B2(n_64),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_28),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_86),
.Y(n_135)
);

AO22x2_ASAP7_75t_L g104 ( 
.A1(n_83),
.A2(n_54),
.B1(n_36),
.B2(n_58),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_58),
.C(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_0),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_115),
.B(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_28),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_73),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_117),
.B(n_77),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_120),
.A2(n_112),
.B(n_107),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_123),
.Y(n_168)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_104),
.A2(n_86),
.B1(n_89),
.B2(n_71),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_127),
.A2(n_128),
.B1(n_103),
.B2(n_80),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_104),
.A2(n_117),
.B1(n_105),
.B2(n_108),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_133),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_131),
.A2(n_135),
.B(n_143),
.Y(n_148)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_136),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_92),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_104),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_108),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_116),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_118),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_28),
.Y(n_161)
);

NAND2x1p5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_86),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_134),
.A2(n_111),
.B1(n_101),
.B2(n_109),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_158),
.B(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_156),
.Y(n_173)
);

A2O1A1O1Ixp25_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_106),
.B(n_7),
.C(n_8),
.D(n_9),
.Y(n_189)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_150),
.B(n_155),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_135),
.C(n_140),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_154),
.Y(n_183)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_160),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_96),
.C(n_76),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_143),
.B(n_112),
.C(n_72),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_143),
.B(n_103),
.C(n_80),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_162),
.Y(n_177)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_142),
.Y(n_160)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_81),
.Y(n_162)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_106),
.B(n_118),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_165),
.B(n_167),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_138),
.A2(n_1),
.B(n_2),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_155),
.A2(n_130),
.B1(n_131),
.B2(n_129),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_180),
.B1(n_188),
.B2(n_6),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_163),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_166),
.B1(n_158),
.B2(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_126),
.B1(n_123),
.B2(n_122),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_120),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_184),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_122),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_182),
.B(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_4),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_185),
.A2(n_187),
.B(n_178),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_157),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_106),
.B1(n_7),
.B2(n_8),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_189),
.B(n_159),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_154),
.C(n_151),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_203),
.C(n_207),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_176),
.A2(n_148),
.B1(n_150),
.B2(n_164),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_183),
.B(n_148),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_198),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_156),
.C(n_149),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_185),
.B(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_201),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_161),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_6),
.C(n_7),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_189),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_9),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_9),
.C(n_10),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_11),
.C(n_12),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_184),
.Y(n_221)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_179),
.B(n_186),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_210),
.A2(n_214),
.B(n_217),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_192),
.A2(n_172),
.B(n_175),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_196),
.A2(n_169),
.B(n_171),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_199),
.B(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_187),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_220),
.B(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_221),
.B(n_203),
.C(n_174),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_191),
.A2(n_190),
.B(n_171),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_222),
.A2(n_170),
.B(n_205),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_194),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_211),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_218),
.B(n_216),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_190),
.B1(n_208),
.B2(n_207),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_226),
.A2(n_212),
.B1(n_222),
.B2(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_231),
.C(n_221),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_11),
.Y(n_231)
);

O2A1O1Ixp33_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_232),
.B(n_13),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_233),
.A2(n_239),
.B1(n_232),
.B2(n_236),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_234),
.B(n_235),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_237),
.A2(n_240),
.B(n_229),
.Y(n_246)
);

A2O1A1Ixp33_ASAP7_75t_SL g238 ( 
.A1(n_223),
.A2(n_215),
.B(n_14),
.C(n_15),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_215),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_223),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_243),
.Y(n_247)
);

O2A1O1Ixp5_ASAP7_75t_L g243 ( 
.A1(n_238),
.A2(n_231),
.B(n_225),
.C(n_228),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_245),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_226),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_241),
.C(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_239),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_16),
.C(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_16),
.C(n_247),
.Y(n_252)
);

FAx1_ASAP7_75t_SL g254 ( 
.A(n_253),
.B(n_252),
.CI(n_242),
.CON(n_254),
.SN(n_254)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_254),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_256),
.B(n_255),
.Y(n_257)
);


endmodule