module real_jpeg_8836_n_15 (n_5, n_4, n_8, n_0, n_12, n_70, n_1, n_11, n_14, n_2, n_13, n_71, n_6, n_72, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_70;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_71;
input n_6;
input n_72;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_17;
wire n_57;
wire n_43;
wire n_37;
wire n_21;
wire n_54;
wire n_65;
wire n_35;
wire n_38;
wire n_33;
wire n_50;
wire n_29;
wire n_55;
wire n_58;
wire n_31;
wire n_67;
wire n_49;
wire n_52;
wire n_63;
wire n_68;
wire n_24;
wire n_66;
wire n_34;
wire n_28;
wire n_60;
wire n_44;
wire n_46;
wire n_62;
wire n_59;
wire n_64;
wire n_23;
wire n_47;
wire n_45;
wire n_61;
wire n_25;
wire n_51;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_40;
wire n_39;
wire n_36;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_48;
wire n_30;
wire n_56;
wire n_16;

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_0),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_0),
.A2(n_35),
.B1(n_37),
.B2(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_1),
.B(n_70),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_3),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_2),
.B(n_3),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_4),
.A2(n_17),
.B1(n_45),
.B2(n_46),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_4),
.A2(n_45),
.B1(n_61),
.B2(n_67),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_8),
.B(n_71),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_8),
.B(n_72),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_9),
.B(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

AOI321xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_47),
.A3(n_57),
.B1(n_58),
.B2(n_60),
.C(n_68),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_17),
.Y(n_46)
);

OAI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_30),
.B1(n_34),
.B2(n_38),
.C(n_40),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_19),
.A2(n_28),
.B(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B(n_22),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_20),
.A2(n_29),
.B(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_29),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NAND3xp33_ASAP7_75t_SL g34 ( 
.A(n_22),
.B(n_35),
.C(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_26),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_29),
.B(n_65),
.Y(n_64)
);

OAI221xp5_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_34),
.B1(n_40),
.B2(n_62),
.C(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_57),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_57),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_53),
.B(n_56),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B(n_52),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_63),
.B(n_66),
.Y(n_65)
);


endmodule