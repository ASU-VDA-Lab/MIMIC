module fake_netlist_6_1786_n_574 (n_52, n_16, n_1, n_91, n_46, n_18, n_21, n_88, n_3, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_77, n_92, n_42, n_96, n_8, n_90, n_24, n_54, n_0, n_87, n_32, n_66, n_85, n_78, n_84, n_13, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_45, n_34, n_70, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_61, n_81, n_59, n_76, n_36, n_26, n_55, n_94, n_97, n_58, n_64, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_86, n_95, n_9, n_10, n_71, n_74, n_6, n_14, n_72, n_89, n_60, n_35, n_12, n_69, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_574);

input n_52;
input n_16;
input n_1;
input n_91;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_77;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_54;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_78;
input n_84;
input n_13;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_45;
input n_34;
input n_70;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_61;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_55;
input n_94;
input n_97;
input n_58;
input n_64;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_86;
input n_95;
input n_9;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_72;
input n_89;
input n_60;
input n_35;
input n_12;
input n_69;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_574;

wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_507;
wire n_209;
wire n_367;
wire n_465;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_144;
wire n_365;
wire n_125;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_106;
wire n_358;
wire n_160;
wire n_449;
wire n_131;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_396;
wire n_495;
wire n_350;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_108;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_114;
wire n_198;
wire n_104;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_111;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_119;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_428;
wire n_432;
wire n_101;
wire n_167;
wire n_174;
wire n_127;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_129;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_109;
wire n_529;
wire n_445;
wire n_425;
wire n_122;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_112;
wire n_172;
wire n_472;
wire n_270;
wire n_239;
wire n_126;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_118;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_460;
wire n_107;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_103;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_98;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_356;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_105;
wire n_227;
wire n_132;
wire n_570;
wire n_406;
wire n_483;
wire n_102;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_130;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_100;
wire n_121;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_244;
wire n_399;
wire n_243;
wire n_124;
wire n_548;
wire n_282;
wire n_436;
wire n_116;
wire n_211;
wire n_523;
wire n_175;
wire n_117;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_123;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_115;
wire n_550;
wire n_487;
wire n_128;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_113;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_99;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_120;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_110;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_295;
wire n_385;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_64),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_2),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NOR2xp67_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_43),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_13),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_47),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_21),
.Y(n_112)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_66),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_42),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_36),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_61),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_12),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_11),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_52),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_80),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_34),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_38),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_24),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_51),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_5),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_77),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_9),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g137 ( 
.A(n_48),
.B(n_4),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_32),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_7),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_2),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_97),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_17),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_15),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_49),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_27),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_63),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_15),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_12),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_17),
.Y(n_152)
);

INVxp67_ASAP7_75t_SL g153 ( 
.A(n_57),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_56),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_53),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_73),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_85),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_44),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_16),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_65),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_28),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

BUFx4f_ASAP7_75t_SL g164 ( 
.A(n_50),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_86),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_23),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_6),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_93),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_26),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_96),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_19),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_1),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_41),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_3),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_30),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_31),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_54),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_20),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_76),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_0),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_78),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g183 ( 
.A(n_5),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_59),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_33),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_19),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_11),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_60),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_82),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_115),
.A2(n_173),
.B1(n_147),
.B2(n_182),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_178),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_178),
.Y(n_194)
);

OA21x2_ASAP7_75t_L g195 ( 
.A1(n_142),
.A2(n_1),
.B(n_3),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_178),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_159),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g200 ( 
.A1(n_142),
.A2(n_151),
.B(n_123),
.Y(n_200)
);

OAI21x1_ASAP7_75t_L g201 ( 
.A1(n_111),
.A2(n_4),
.B(n_8),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

NAND2xp33_ASAP7_75t_L g203 ( 
.A(n_172),
.B(n_8),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_172),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_106),
.B(n_9),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g206 ( 
.A(n_149),
.B(n_35),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_10),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_135),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_172),
.Y(n_210)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_29),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_10),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_172),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_122),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_115),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_215)
);

AND3x2_ASAP7_75t_L g216 ( 
.A(n_151),
.B(n_14),
.C(n_18),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_130),
.B(n_67),
.Y(n_218)
);

AOI22x1_ASAP7_75t_SL g219 ( 
.A1(n_135),
.A2(n_18),
.B1(n_25),
.B2(n_37),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_99),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_62),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g222 ( 
.A1(n_107),
.A2(n_87),
.B(n_90),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_136),
.A2(n_94),
.B(n_160),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_133),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_154),
.B(n_174),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_186),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_130),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_154),
.Y(n_232)
);

NAND2xp33_ASAP7_75t_L g233 ( 
.A(n_139),
.B(n_140),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_111),
.B(n_128),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_128),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_137),
.A2(n_152),
.B1(n_167),
.B2(n_187),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_138),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_138),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_148),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_138),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_129),
.Y(n_241)
);

AND2x4_ASAP7_75t_L g242 ( 
.A(n_129),
.B(n_120),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_113),
.B(n_183),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_100),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_102),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_144),
.B(n_188),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_104),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_143),
.Y(n_248)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_113),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_101),
.A2(n_171),
.B1(n_161),
.B2(n_157),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_105),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_112),
.B(n_118),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_101),
.A2(n_157),
.B1(n_161),
.B2(n_171),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_108),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_116),
.A2(n_189),
.B1(n_126),
.B2(n_109),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_110),
.B(n_155),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_121),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_125),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_127),
.B(n_169),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_131),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_132),
.B(n_184),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_141),
.Y(n_262)
);

AND2x4_ASAP7_75t_L g263 ( 
.A(n_145),
.B(n_179),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_98),
.Y(n_264)
);

NOR3xp33_ASAP7_75t_L g265 ( 
.A(n_207),
.B(n_163),
.C(n_150),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_146),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

NOR2x1p5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_185),
.Y(n_269)
);

NAND3xp33_ASAP7_75t_L g270 ( 
.A(n_205),
.B(n_162),
.C(n_119),
.Y(n_270)
);

NOR2x1p5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_153),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_250),
.B(n_180),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_213),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_200),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_L g278 ( 
.A1(n_191),
.A2(n_164),
.B1(n_103),
.B2(n_134),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_206),
.B(n_177),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_192),
.Y(n_280)
);

INVx4_ASAP7_75t_SL g281 ( 
.A(n_218),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_192),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_225),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_246),
.B(n_124),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_212),
.A2(n_261),
.B1(n_256),
.B2(n_235),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_225),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_200),
.Y(n_289)
);

OR2x2_ASAP7_75t_SL g290 ( 
.A(n_195),
.B(n_164),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g291 ( 
.A(n_206),
.B(n_156),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_258),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_158),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_243),
.B(n_166),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_258),
.Y(n_295)
);

CKINVDCx11_ASAP7_75t_R g296 ( 
.A(n_208),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_168),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_262),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_237),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_248),
.B(n_170),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_206),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_253),
.B(n_176),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_218),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_212),
.A2(n_261),
.B1(n_256),
.B2(n_235),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_255),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_238),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_192),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_235),
.A2(n_242),
.B1(n_243),
.B2(n_263),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_196),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_238),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_R g316 ( 
.A(n_239),
.B(n_224),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_221),
.B(n_233),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_215),
.A2(n_239),
.B1(n_234),
.B2(n_232),
.Y(n_318)
);

AND2x6_ASAP7_75t_L g319 ( 
.A(n_211),
.B(n_240),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_241),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_293),
.A2(n_233),
.B1(n_211),
.B2(n_203),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_273),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_317),
.B(n_211),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_263),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_277),
.B(n_263),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_259),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_266),
.B(n_259),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_298),
.B(n_232),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_313),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_287),
.B(n_242),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_307),
.A2(n_219),
.B1(n_208),
.B2(n_203),
.Y(n_331)
);

AND3x1_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_265),
.C(n_284),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_306),
.B(n_202),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_311),
.B(n_198),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_244),
.Y(n_335)
);

NOR2xp67_ASAP7_75t_L g336 ( 
.A(n_270),
.B(n_247),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_257),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_241),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_320),
.B(n_241),
.Y(n_339)
);

OR2x6_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_201),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_267),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_274),
.B(n_278),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_268),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_320),
.B(n_241),
.Y(n_344)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_272),
.Y(n_346)
);

AND2x6_ASAP7_75t_SL g347 ( 
.A(n_296),
.B(n_220),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_314),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_274),
.B(n_254),
.Y(n_349)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_279),
.C(n_264),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_275),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g353 ( 
.A(n_264),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_251),
.C(n_229),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_224),
.B1(n_201),
.B2(n_260),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_272),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_276),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_292),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_193),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g362 ( 
.A(n_288),
.B(n_228),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_295),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_194),
.Y(n_364)
);

NAND2x1p5_ASAP7_75t_L g365 ( 
.A(n_305),
.B(n_222),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_307),
.A2(n_228),
.B1(n_223),
.B2(n_222),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_280),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_319),
.B(n_271),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_299),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_288),
.B(n_260),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_362),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_328),
.B(n_303),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_303),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_290),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_350),
.B(n_296),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_345),
.B(n_218),
.Y(n_377)
);

OAI22x1_ASAP7_75t_L g378 ( 
.A1(n_321),
.A2(n_224),
.B1(n_223),
.B2(n_216),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g379 ( 
.A1(n_324),
.A2(n_218),
.B1(n_319),
.B2(n_260),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_341),
.Y(n_380)
);

O2A1O1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_333),
.A2(n_194),
.B(n_197),
.C(n_199),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_330),
.A2(n_300),
.B1(n_260),
.B2(n_245),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_325),
.B1(n_326),
.B2(n_335),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_343),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_337),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_361),
.A2(n_282),
.B(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_331),
.Y(n_389)
);

BUFx8_ASAP7_75t_L g390 ( 
.A(n_347),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_371),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_245),
.Y(n_392)
);

NOR2x1_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_336),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_281),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_361),
.A2(n_283),
.B(n_312),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_340),
.A2(n_245),
.B1(n_281),
.B2(n_283),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_334),
.B(n_283),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_340),
.B(n_369),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_364),
.A2(n_309),
.B(n_315),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_348),
.B(n_309),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_366),
.A2(n_315),
.B1(n_308),
.B2(n_304),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_L g403 ( 
.A1(n_356),
.A2(n_304),
.B(n_297),
.C(n_217),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_364),
.A2(n_297),
.B(n_209),
.C(n_217),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_352),
.B(n_196),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_367),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_339),
.A2(n_196),
.B(n_209),
.C(n_217),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_L g408 ( 
.A1(n_322),
.A2(n_196),
.B1(n_209),
.B2(n_217),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_365),
.A2(n_209),
.B(n_217),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_339),
.A2(n_209),
.B(n_227),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_346),
.B(n_227),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_351),
.A2(n_240),
.B1(n_227),
.B2(n_230),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_344),
.A2(n_227),
.B(n_230),
.Y(n_413)
);

OAI21xp33_ASAP7_75t_L g414 ( 
.A1(n_357),
.A2(n_227),
.B(n_230),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_358),
.B(n_230),
.Y(n_415)
);

OR2x6_ASAP7_75t_SL g416 ( 
.A(n_329),
.B(n_230),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_329),
.A2(n_240),
.B(n_355),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_341),
.Y(n_419)
);

A2O1A1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_321),
.A2(n_317),
.B(n_323),
.C(n_327),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_274),
.Y(n_421)
);

OR2x6_ASAP7_75t_L g422 ( 
.A(n_330),
.B(n_250),
.Y(n_422)
);

AND2x4_ASAP7_75t_L g423 ( 
.A(n_353),
.B(n_341),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_323),
.B(n_324),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_323),
.A2(n_321),
.B1(n_317),
.B2(n_302),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_323),
.B(n_324),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_321),
.A2(n_317),
.B1(n_323),
.B2(n_324),
.Y(n_427)
);

INVx3_ASAP7_75t_SL g428 ( 
.A(n_362),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_323),
.B(n_324),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_422),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_427),
.B(n_420),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_L g432 ( 
.A1(n_375),
.A2(n_426),
.B(n_424),
.C(n_429),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_372),
.Y(n_433)
);

BUFx4f_ASAP7_75t_L g434 ( 
.A(n_428),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_389),
.A2(n_373),
.B1(n_422),
.B2(n_374),
.Y(n_435)
);

AOI22xp33_ASAP7_75t_L g436 ( 
.A1(n_422),
.A2(n_394),
.B1(n_392),
.B2(n_397),
.Y(n_436)
);

AO31x2_ASAP7_75t_L g437 ( 
.A1(n_384),
.A2(n_409),
.A3(n_398),
.B(n_407),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_380),
.Y(n_438)
);

INVx3_ASAP7_75t_SL g439 ( 
.A(n_423),
.Y(n_439)
);

AND2x4_ASAP7_75t_L g440 ( 
.A(n_423),
.B(n_419),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_386),
.A2(n_402),
.B1(n_393),
.B2(n_400),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_383),
.B(n_411),
.Y(n_442)
);

CKINVDCx6p67_ASAP7_75t_R g443 ( 
.A(n_416),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

AO31x2_ASAP7_75t_L g446 ( 
.A1(n_399),
.A2(n_405),
.A3(n_388),
.B(n_395),
.Y(n_446)
);

NAND3xp33_ASAP7_75t_SL g447 ( 
.A(n_376),
.B(n_382),
.C(n_396),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_379),
.A2(n_414),
.B1(n_377),
.B2(n_401),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_404),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_417),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_410),
.A2(n_413),
.B(n_408),
.Y(n_453)
);

BUFx4_ASAP7_75t_SL g454 ( 
.A(n_390),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_412),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_390),
.A2(n_289),
.B(n_338),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_427),
.A2(n_375),
.B(n_420),
.C(n_317),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g458 ( 
.A(n_422),
.Y(n_458)
);

AO32x2_ASAP7_75t_L g459 ( 
.A1(n_425),
.A2(n_366),
.A3(n_385),
.B1(n_384),
.B2(n_255),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_424),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_427),
.B(n_420),
.Y(n_461)
);

NOR2xp67_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_350),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_427),
.B(n_420),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g464 ( 
.A(n_428),
.Y(n_464)
);

BUFx10_ASAP7_75t_L g465 ( 
.A(n_376),
.Y(n_465)
);

AO31x2_ASAP7_75t_L g466 ( 
.A1(n_403),
.A2(n_420),
.A3(n_425),
.B(n_378),
.Y(n_466)
);

AO31x2_ASAP7_75t_L g467 ( 
.A1(n_403),
.A2(n_420),
.A3(n_425),
.B(n_378),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_375),
.B(n_387),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_391),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_391),
.Y(n_470)
);

NOR2x1_ASAP7_75t_L g471 ( 
.A(n_424),
.B(n_426),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_391),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_427),
.B(n_420),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_418),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_375),
.B(n_387),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_471),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_433),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_457),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_464),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_439),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_449),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_438),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_431),
.A2(n_473),
.B(n_463),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_431),
.A2(n_463),
.B(n_461),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_440),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_440),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_435),
.B(n_445),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_432),
.B(n_436),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_441),
.A2(n_435),
.B(n_468),
.C(n_476),
.Y(n_491)
);

BUFx8_ASAP7_75t_L g492 ( 
.A(n_430),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_469),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_444),
.Y(n_494)
);

OR2x2_ASAP7_75t_L g495 ( 
.A(n_442),
.B(n_464),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_474),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_456),
.B(n_472),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_453),
.A2(n_448),
.B(n_447),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_451),
.A2(n_441),
.B(n_448),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_470),
.A2(n_450),
.B1(n_455),
.B2(n_458),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_466),
.Y(n_501)
);

OA21x2_ASAP7_75t_L g502 ( 
.A1(n_466),
.A2(n_467),
.B(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_483),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_492),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_R g505 ( 
.A(n_494),
.B(n_434),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_501),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_477),
.Y(n_507)
);

OA21x2_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_467),
.B(n_446),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_484),
.Y(n_509)
);

AOI22xp33_ASAP7_75t_SL g510 ( 
.A1(n_490),
.A2(n_465),
.B1(n_434),
.B2(n_459),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_494),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g512 ( 
.A(n_479),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_480),
.B(n_437),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_437),
.Y(n_514)
);

INVx3_ASAP7_75t_SL g515 ( 
.A(n_482),
.Y(n_515)
);

AOI22xp33_ASAP7_75t_L g516 ( 
.A1(n_489),
.A2(n_465),
.B1(n_475),
.B2(n_443),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_437),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_506),
.Y(n_518)
);

NOR2x1_ASAP7_75t_L g519 ( 
.A(n_507),
.B(n_478),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_515),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_514),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_511),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_511),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_512),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_510),
.B(n_485),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_513),
.B(n_490),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_510),
.B(n_486),
.Y(n_527)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_491),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_514),
.A2(n_500),
.B1(n_479),
.B2(n_495),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_512),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_503),
.B(n_499),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_521),
.B(n_517),
.Y(n_533)
);

NAND2x1_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_497),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_522),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_521),
.B(n_517),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_518),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g538 ( 
.A(n_520),
.B(n_515),
.Y(n_538)
);

INVxp67_ASAP7_75t_SL g539 ( 
.A(n_530),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_532),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_508),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_518),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_537),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_540),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_538),
.A2(n_528),
.B1(n_525),
.B2(n_527),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_528),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_536),
.B(n_531),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_541),
.B(n_525),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_535),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_544),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_549),
.B(n_539),
.Y(n_551)
);

NAND2x1_ASAP7_75t_L g552 ( 
.A(n_544),
.B(n_542),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_543),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_536),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_541),
.Y(n_555)
);

INVxp67_ASAP7_75t_L g556 ( 
.A(n_548),
.Y(n_556)
);

AOI222xp33_ASAP7_75t_L g557 ( 
.A1(n_556),
.A2(n_545),
.B1(n_527),
.B2(n_529),
.C1(n_524),
.C2(n_546),
.Y(n_557)
);

AOI31xp33_ASAP7_75t_L g558 ( 
.A1(n_556),
.A2(n_550),
.A3(n_551),
.B(n_548),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g559 ( 
.A1(n_554),
.A2(n_516),
.B(n_524),
.Y(n_559)
);

NAND3xp33_ASAP7_75t_SL g560 ( 
.A(n_552),
.B(n_534),
.C(n_495),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_560),
.A2(n_504),
.B1(n_547),
.B2(n_555),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_561),
.B(n_559),
.C(n_557),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_562),
.A2(n_558),
.B(n_553),
.Y(n_563)
);

NOR2x1_ASAP7_75t_L g564 ( 
.A(n_563),
.B(n_504),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_564),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_564),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_565),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_481),
.Y(n_568)
);

OAI22x1_ASAP7_75t_SL g569 ( 
.A1(n_567),
.A2(n_454),
.B1(n_566),
.B2(n_515),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_569),
.A2(n_568),
.B(n_505),
.Y(n_570)
);

AOI221xp5_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_523),
.B1(n_504),
.B2(n_488),
.C(n_487),
.Y(n_571)
);

AO21x2_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_496),
.B(n_493),
.Y(n_572)
);

OR2x6_ASAP7_75t_L g573 ( 
.A(n_572),
.B(n_488),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_492),
.B1(n_487),
.B2(n_475),
.Y(n_574)
);


endmodule