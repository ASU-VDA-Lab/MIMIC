module fake_jpeg_30474_n_85 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_3),
.B(n_16),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_0),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_8),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_44),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_1),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_29),
.B(n_1),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_30),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_51),
.C(n_52),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_41),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_22),
.B(n_31),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_24),
.A2(n_36),
.B1(n_38),
.B2(n_26),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_23),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_22),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_63),
.B(n_57),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_54),
.B1(n_56),
.B2(n_51),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_67),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_72),
.B1(n_65),
.B2(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_74),
.C(n_73),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_79),
.A2(n_70),
.B(n_77),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_78),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_49),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_83),
.B(n_61),
.C(n_64),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_64),
.B(n_59),
.Y(n_85)
);


endmodule