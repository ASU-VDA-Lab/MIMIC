module fake_jpeg_17935_n_152 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_152);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_28),
.B(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_30),
.B(n_31),
.Y(n_51)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_17),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_25),
.B1(n_23),
.B2(n_17),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_37),
.A2(n_25),
.B1(n_32),
.B2(n_30),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_38),
.B(n_42),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx12_ASAP7_75t_R g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_41),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_20),
.C(n_21),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_58),
.B1(n_60),
.B2(n_47),
.Y(n_80)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_63),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_32),
.B1(n_33),
.B2(n_15),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_34),
.B1(n_33),
.B2(n_28),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_28),
.B(n_3),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_51),
.A3(n_41),
.B1(n_44),
.B2(n_37),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_65),
.A3(n_18),
.B1(n_57),
.B2(n_27),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_70),
.B(n_73),
.Y(n_93)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_64),
.B(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_43),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_81),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_59),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_77),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_59),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_56),
.B(n_61),
.Y(n_82)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_88),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_68),
.B(n_79),
.Y(n_98)
);

INVxp33_ASAP7_75t_SL g86 ( 
.A(n_75),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_80),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_18),
.C(n_39),
.Y(n_108)
);

OA21x2_ASAP7_75t_L g88 ( 
.A1(n_74),
.A2(n_43),
.B(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_46),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_76),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_90),
.B(n_95),
.Y(n_102)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_99),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_98),
.A2(n_14),
.B(n_15),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_93),
.B(n_77),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_63),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_108),
.C(n_91),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_88),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_104),
.B(n_105),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_72),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_94),
.A2(n_71),
.B(n_3),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_71),
.B(n_19),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_19),
.B(n_26),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_85),
.B(n_12),
.C(n_10),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_8),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_100),
.A2(n_82),
.B1(n_88),
.B2(n_95),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_109),
.B(n_104),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_82),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_113),
.C(n_108),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_116),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_90),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_104),
.A2(n_91),
.B1(n_92),
.B2(n_45),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_126),
.C(n_127),
.Y(n_130)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_122),
.A2(n_21),
.B(n_24),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_103),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_124),
.A2(n_112),
.B(n_125),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_106),
.C(n_96),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_26),
.CI(n_24),
.CON(n_127),
.SN(n_127)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_123),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_124),
.A2(n_128),
.B(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_127),
.B(n_92),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_133),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_112),
.B(n_4),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_34),
.B1(n_48),
.B2(n_2),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_120),
.C(n_126),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_144),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_140),
.A2(n_135),
.B1(n_9),
.B2(n_4),
.Y(n_144)
);

NOR2xp67_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_136),
.Y(n_145)
);

AOI21x1_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_146),
.B(n_142),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_141),
.A2(n_137),
.B(n_138),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_147),
.A2(n_9),
.B(n_2),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_148),
.B(n_149),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_2),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_4),
.Y(n_152)
);


endmodule