module fake_netlist_6_2097_n_1751 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1751);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1751;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_19),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_30),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_20),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_24),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_50),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_28),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_163),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_32),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_105),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_41),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_32),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_42),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_150),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_101),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_4),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_44),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_54),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_42),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_73),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_100),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_39),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_61),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_2),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_119),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_126),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_143),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_130),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_72),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_122),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_142),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_16),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_75),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_128),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_132),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_169),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_148),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_31),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_21),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_174),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_131),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_76),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_90),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_153),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_134),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_39),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_104),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_28),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_117),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_109),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g233 ( 
.A(n_87),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_107),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_135),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_77),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_57),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_94),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_62),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_66),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_154),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_138),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_83),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_26),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_16),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_164),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_103),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_65),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_111),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_8),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_161),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_110),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_48),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_129),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_137),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_70),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_159),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_157),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_147),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_74),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_50),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_141),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_22),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_78),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_19),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_80),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_56),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_88),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_171),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_112),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_45),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_13),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_53),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_158),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_55),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_69),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_24),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_160),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_82),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_84),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_6),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_36),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_96),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_152),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_98),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_38),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_12),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_166),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_97),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_12),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_41),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_95),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_58),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_64),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_11),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_120),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_29),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_18),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_168),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_4),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_91),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_145),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_165),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_63),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_29),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_33),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_57),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_23),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_27),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_37),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_113),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_58),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_5),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_151),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_89),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_48),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_124),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_15),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_149),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_79),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_30),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_43),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_33),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_46),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_81),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_47),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_54),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_108),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_36),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_55),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_102),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_93),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_23),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_99),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_37),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_52),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_52),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_139),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_5),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_116),
.Y(n_342)
);

CKINVDCx11_ASAP7_75t_R g343 ( 
.A(n_43),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_38),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_7),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_3),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_121),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_0),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_118),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_14),
.Y(n_350)
);

NOR2xp67_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_0),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_213),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_236),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_253),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_343),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_273),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_273),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_182),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_183),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_251),
.B(n_2),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_273),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_346),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_187),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_231),
.B(n_3),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_279),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_295),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_231),
.B(n_210),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_252),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_346),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_192),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_199),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_230),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_346),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_346),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_295),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_204),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_298),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_298),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_230),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_205),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_240),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_185),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_185),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_299),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_206),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_177),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_177),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_208),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_209),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_184),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_211),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_214),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_285),
.B(n_6),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_240),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_184),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_215),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_186),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_216),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_233),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_191),
.B(n_7),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_217),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_186),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_188),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_220),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_188),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_240),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_243),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_221),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_222),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_194),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_194),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_201),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_224),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_227),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_201),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_203),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_203),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_232),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_246),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_234),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_235),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_246),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_238),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_239),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_248),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_191),
.B(n_8),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_262),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_262),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_207),
.B(n_9),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_249),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_255),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_356),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_356),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_357),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g441 ( 
.A(n_351),
.B(n_275),
.Y(n_441)
);

CKINVDCx8_ASAP7_75t_R g442 ( 
.A(n_405),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_400),
.B(n_243),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_355),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_387),
.B(n_256),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_357),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_358),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_358),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_362),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_362),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_363),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_363),
.Y(n_454)
);

AND2x6_ASAP7_75t_L g455 ( 
.A(n_387),
.B(n_275),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_376),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_364),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_364),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_361),
.B(n_233),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_365),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_372),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_372),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_373),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_370),
.B(n_233),
.Y(n_466)
);

NAND2xp33_ASAP7_75t_R g467 ( 
.A(n_367),
.B(n_176),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_377),
.Y(n_469)
);

NAND2xp33_ASAP7_75t_L g470 ( 
.A(n_387),
.B(n_198),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_378),
.B(n_243),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_392),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_382),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_382),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_412),
.B(n_270),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_416),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_413),
.B(n_258),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_388),
.B(n_270),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_389),
.B(n_267),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_406),
.B(n_269),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_383),
.Y(n_484)
);

NOR2x1_ASAP7_75t_L g485 ( 
.A(n_381),
.B(n_275),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_383),
.B(n_270),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_393),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_369),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_393),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_396),
.B(n_259),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_352),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_401),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_401),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_380),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_403),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_403),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_408),
.B(n_202),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_409),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_411),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_417),
.Y(n_509)
);

CKINVDCx11_ASAP7_75t_R g510 ( 
.A(n_353),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_399),
.B(n_244),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_371),
.B(n_260),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g513 ( 
.A(n_432),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_418),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_359),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_444),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_446),
.B(n_360),
.Y(n_517)
);

OR2x2_ASAP7_75t_L g518 ( 
.A(n_456),
.B(n_366),
.Y(n_518)
);

BUFx4f_ASAP7_75t_L g519 ( 
.A(n_455),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_438),
.Y(n_520)
);

INVx3_ASAP7_75t_L g521 ( 
.A(n_449),
.Y(n_521)
);

AOI22xp33_ASAP7_75t_L g522 ( 
.A1(n_513),
.A2(n_435),
.B1(n_294),
.B2(n_309),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_449),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_443),
.B(n_418),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_374),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_444),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_444),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_452),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_485),
.B(n_274),
.Y(n_529)
);

BUFx4f_ASAP7_75t_L g530 ( 
.A(n_455),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_511),
.B(n_375),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_501),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_456),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_512),
.B(n_391),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_455),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_513),
.B(n_395),
.C(n_394),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_455),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_512),
.B(n_397),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_452),
.Y(n_541)
);

BUFx6f_ASAP7_75t_SL g542 ( 
.A(n_481),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_467),
.A2(n_319),
.B1(n_296),
.B2(n_301),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_452),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_466),
.B(n_398),
.Y(n_545)
);

AND2x2_ASAP7_75t_SL g546 ( 
.A(n_483),
.B(n_202),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_480),
.B(n_404),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_439),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_495),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_463),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_440),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_449),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_480),
.B(n_483),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_485),
.B(n_202),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_463),
.Y(n_555)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_473),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_460),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_R g558 ( 
.A(n_489),
.B(n_407),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_443),
.B(n_477),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_443),
.B(n_410),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_460),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_501),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_466),
.A2(n_345),
.B1(n_274),
.B2(n_282),
.Y(n_563)
);

BUFx10_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_463),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_440),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_464),
.Y(n_567)
);

AND2x6_ASAP7_75t_L g568 ( 
.A(n_441),
.B(n_290),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_449),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_464),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_467),
.A2(n_385),
.B1(n_402),
.B2(n_420),
.Y(n_571)
);

INVxp67_ASAP7_75t_SL g572 ( 
.A(n_449),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_447),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_464),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_447),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_459),
.B(n_414),
.Y(n_576)
);

AND3x1_ASAP7_75t_L g577 ( 
.A(n_478),
.B(n_294),
.C(n_282),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_501),
.Y(n_578)
);

INVxp33_ASAP7_75t_SL g579 ( 
.A(n_478),
.Y(n_579)
);

INVx8_ASAP7_75t_L g580 ( 
.A(n_455),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_477),
.A2(n_459),
.B1(n_481),
.B2(n_494),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_477),
.B(n_421),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_448),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_468),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_482),
.B(n_415),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_468),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_510),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_482),
.A2(n_178),
.B1(n_283),
.B2(n_288),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_448),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_449),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_468),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_450),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_450),
.Y(n_593)
);

AND3x2_ASAP7_75t_L g594 ( 
.A(n_489),
.B(n_290),
.C(n_284),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_449),
.Y(n_595)
);

AND2x4_ASAP7_75t_SL g596 ( 
.A(n_495),
.B(n_354),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_451),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_449),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_455),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_490),
.B(n_419),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_490),
.B(n_424),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_473),
.B(n_429),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_473),
.B(n_430),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_442),
.B(n_431),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_510),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_453),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_453),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_451),
.Y(n_608)
);

INVxp67_ASAP7_75t_SL g609 ( 
.A(n_470),
.Y(n_609)
);

BUFx6f_ASAP7_75t_SL g610 ( 
.A(n_481),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_462),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_457),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_L g613 ( 
.A1(n_481),
.A2(n_494),
.B1(n_441),
.B2(n_473),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_453),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_501),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_490),
.B(n_436),
.Y(n_616)
);

INVx5_ASAP7_75t_L g617 ( 
.A(n_455),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_462),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_442),
.B(n_437),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_502),
.B(n_426),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_457),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_462),
.Y(n_623)
);

INVx4_ASAP7_75t_L g624 ( 
.A(n_455),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_486),
.B(n_207),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_442),
.B(n_427),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_453),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_486),
.B(n_223),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_458),
.B(n_461),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_470),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_489),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_465),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_458),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_462),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_503),
.B(n_290),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_455),
.Y(n_636)
);

INVx1_ASAP7_75t_SL g637 ( 
.A(n_499),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_501),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_461),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_494),
.A2(n_309),
.B1(n_325),
.B2(n_311),
.Y(n_640)
);

AO22x2_ASAP7_75t_L g641 ( 
.A1(n_503),
.A2(n_311),
.B1(n_325),
.B2(n_345),
.Y(n_641)
);

INVx6_ASAP7_75t_L g642 ( 
.A(n_494),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_445),
.B(n_233),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_469),
.B(n_271),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_499),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_465),
.Y(n_646)
);

OR2x6_ASAP7_75t_L g647 ( 
.A(n_503),
.B(n_223),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_469),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_501),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_502),
.B(n_505),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_465),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_474),
.B(n_421),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_462),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_462),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_471),
.B(n_277),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_445),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_465),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_455),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_SL g659 ( 
.A(n_474),
.B(n_193),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_472),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_494),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_502),
.B(n_198),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_479),
.B(n_225),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_501),
.B(n_281),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g665 ( 
.A(n_479),
.Y(n_665)
);

BUFx5_ASAP7_75t_L g666 ( 
.A(n_636),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_546),
.A2(n_289),
.B1(n_226),
.B2(n_229),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_545),
.A2(n_368),
.B1(n_303),
.B2(n_286),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_546),
.A2(n_641),
.B1(n_559),
.B2(n_553),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_556),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_652),
.Y(n_671)
);

A2O1A1Ixp33_ASAP7_75t_L g672 ( 
.A1(n_525),
.A2(n_259),
.B(n_284),
.C(n_329),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_560),
.A2(n_502),
.B(n_509),
.C(n_505),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_652),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_531),
.B(n_502),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_576),
.B(n_293),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_563),
.B(n_180),
.C(n_179),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_620),
.B(n_505),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_621),
.B(n_300),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_556),
.Y(n_680)
);

OAI221xp5_ASAP7_75t_L g681 ( 
.A1(n_522),
.A2(n_514),
.B1(n_488),
.B2(n_508),
.C(n_507),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_516),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_581),
.A2(n_329),
.B1(n_347),
.B2(n_241),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_620),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_524),
.B(n_488),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_641),
.A2(n_250),
.B1(n_305),
.B2(n_312),
.Y(n_686)
);

AO221x1_ASAP7_75t_L g687 ( 
.A1(n_588),
.A2(n_198),
.B1(n_225),
.B2(n_226),
.C(n_229),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_536),
.B(n_505),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_613),
.A2(n_347),
.B1(n_261),
.B2(n_263),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_520),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_609),
.B(n_505),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_L g692 ( 
.A(n_571),
.B(n_492),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_547),
.B(n_509),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_630),
.B(n_509),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_600),
.B(n_302),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_515),
.B(n_509),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_517),
.B(n_509),
.Y(n_697)
);

A2O1A1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_650),
.A2(n_349),
.B(n_247),
.C(n_250),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_601),
.B(n_315),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_616),
.B(n_316),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_656),
.B(n_197),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_554),
.A2(n_336),
.B1(n_340),
.B2(n_334),
.Y(n_702)
);

NAND3xp33_ASAP7_75t_L g703 ( 
.A(n_659),
.B(n_189),
.C(n_181),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_526),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_556),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_527),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_524),
.B(n_318),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_533),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_564),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_554),
.A2(n_326),
.B1(n_321),
.B2(n_342),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_582),
.B(n_585),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_665),
.B(n_492),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_533),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_582),
.B(n_501),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_534),
.B(n_190),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_561),
.B(n_498),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_625),
.A2(n_628),
.B(n_530),
.C(n_519),
.Y(n_717)
);

AOI22xp5_ASAP7_75t_L g718 ( 
.A1(n_554),
.A2(n_333),
.B1(n_241),
.B2(n_247),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_561),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_L g720 ( 
.A(n_554),
.B(n_198),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_656),
.B(n_498),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_661),
.B(n_506),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_661),
.B(n_506),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_641),
.A2(n_333),
.B1(n_257),
.B2(n_261),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_631),
.B(n_257),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_579),
.B(n_506),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_520),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_579),
.B(n_506),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_529),
.A2(n_200),
.B1(n_245),
.B2(n_272),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_549),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_518),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_527),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_537),
.B(n_506),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_539),
.B(n_195),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_543),
.B(n_196),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_556),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_606),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_540),
.B(n_506),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_540),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_554),
.A2(n_280),
.B1(n_312),
.B2(n_320),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_606),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_625),
.A2(n_263),
.B(n_265),
.C(n_280),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_548),
.B(n_551),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_518),
.B(n_506),
.Y(n_744)
);

INVxp67_ASAP7_75t_L g745 ( 
.A(n_577),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_594),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_SL g747 ( 
.A(n_643),
.B(n_278),
.Y(n_747)
);

BUFx8_ASAP7_75t_L g748 ( 
.A(n_554),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_637),
.B(n_504),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_554),
.A2(n_297),
.B1(n_349),
.B2(n_320),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_548),
.B(n_506),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_551),
.B(n_471),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_566),
.B(n_487),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_566),
.B(n_487),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_573),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_607),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_573),
.B(n_487),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_529),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_519),
.A2(n_530),
.B(n_572),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_575),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_557),
.B(n_504),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_529),
.A2(n_327),
.B1(n_350),
.B2(n_338),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_575),
.B(n_487),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_583),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_625),
.B(n_507),
.Y(n_765)
);

BUFx3_ASAP7_75t_L g766 ( 
.A(n_596),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_628),
.B(n_508),
.Y(n_767)
);

NOR2x1p5_ASAP7_75t_L g768 ( 
.A(n_587),
.B(n_212),
.Y(n_768)
);

OR2x6_ASAP7_75t_L g769 ( 
.A(n_645),
.B(n_265),
.Y(n_769)
);

BUFx8_ASAP7_75t_L g770 ( 
.A(n_542),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_614),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_549),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_589),
.B(n_454),
.Y(n_773)
);

NOR3xp33_ASAP7_75t_L g774 ( 
.A(n_659),
.B(n_289),
.C(n_297),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_592),
.B(n_593),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_602),
.B(n_218),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_603),
.B(n_198),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_L g778 ( 
.A1(n_529),
.A2(n_305),
.B1(n_304),
.B2(n_500),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_641),
.A2(n_304),
.B1(n_500),
.B2(n_497),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_592),
.B(n_454),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_593),
.Y(n_781)
);

NOR3xp33_ASAP7_75t_L g782 ( 
.A(n_604),
.B(n_422),
.C(n_423),
.Y(n_782)
);

OAI21xp5_ASAP7_75t_L g783 ( 
.A1(n_519),
.A2(n_454),
.B(n_472),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_644),
.B(n_219),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_530),
.B(n_497),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_597),
.B(n_454),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_580),
.Y(n_787)
);

OAI22xp33_ASAP7_75t_L g788 ( 
.A1(n_647),
.A2(n_237),
.B1(n_228),
.B2(n_242),
.Y(n_788)
);

AND2x2_ASAP7_75t_L g789 ( 
.A(n_628),
.B(n_422),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_635),
.A2(n_500),
.B1(n_497),
.B2(n_423),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_564),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_608),
.B(n_454),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_608),
.B(n_500),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_612),
.B(n_493),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_612),
.B(n_493),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_617),
.B(n_254),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_493),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_617),
.B(n_264),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_655),
.B(n_266),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_633),
.B(n_639),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_580),
.A2(n_538),
.B(n_535),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_617),
.B(n_268),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_633),
.B(n_493),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_639),
.B(n_493),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_617),
.B(n_276),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_648),
.B(n_493),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_647),
.B(n_287),
.Y(n_807)
);

HB1xp67_ASAP7_75t_L g808 ( 
.A(n_647),
.Y(n_808)
);

INVxp67_ASAP7_75t_L g809 ( 
.A(n_558),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_648),
.B(n_493),
.Y(n_810)
);

OAI221xp5_ASAP7_75t_L g811 ( 
.A1(n_640),
.A2(n_425),
.B1(n_428),
.B2(n_433),
.C(n_434),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_642),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_663),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_642),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_635),
.B(n_493),
.Y(n_815)
);

BUFx6f_ASAP7_75t_SL g816 ( 
.A(n_663),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_535),
.B(n_496),
.Y(n_817)
);

NOR3xp33_ASAP7_75t_L g818 ( 
.A(n_619),
.B(n_434),
.C(n_433),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_596),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_663),
.B(n_642),
.Y(n_820)
);

INVxp67_ASAP7_75t_L g821 ( 
.A(n_663),
.Y(n_821)
);

AND2x4_ASAP7_75t_L g822 ( 
.A(n_636),
.B(n_658),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_635),
.B(n_496),
.Y(n_823)
);

OAI22xp5_ASAP7_75t_L g824 ( 
.A1(n_642),
.A2(n_332),
.B1(n_292),
.B2(n_306),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_629),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_822),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_684),
.Y(n_827)
);

NOR3xp33_ASAP7_75t_L g828 ( 
.A(n_729),
.B(n_626),
.C(n_605),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_801),
.A2(n_580),
.B(n_535),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_669),
.A2(n_658),
.B1(n_538),
.B2(n_599),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_825),
.B(n_635),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_759),
.A2(n_580),
.B(n_538),
.Y(n_832)
);

OAI21xp5_ASAP7_75t_L g833 ( 
.A1(n_673),
.A2(n_693),
.B(n_717),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_809),
.B(n_599),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_675),
.B(n_635),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_690),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_SL g837 ( 
.A(n_701),
.B(n_587),
.Y(n_837)
);

INVx2_ASAP7_75t_SL g838 ( 
.A(n_749),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_787),
.A2(n_599),
.B(n_624),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_809),
.B(n_542),
.Y(n_840)
);

A2O1A1Ixp33_ASAP7_75t_L g841 ( 
.A1(n_693),
.A2(n_598),
.B(n_521),
.C(n_523),
.Y(n_841)
);

NAND3xp33_ASAP7_75t_L g842 ( 
.A(n_715),
.B(n_335),
.C(n_348),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_667),
.A2(n_624),
.B1(n_610),
.B2(n_552),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_721),
.B(n_564),
.Y(n_844)
);

AOI21x1_ASAP7_75t_L g845 ( 
.A1(n_785),
.A2(n_664),
.B(n_555),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_787),
.A2(n_615),
.B(n_578),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_713),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_691),
.A2(n_694),
.B(n_783),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_727),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_817),
.A2(n_615),
.B(n_578),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_711),
.B(n_635),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_667),
.A2(n_610),
.B1(n_595),
.B2(n_598),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_817),
.A2(n_615),
.B(n_578),
.Y(n_853)
);

INVx3_ASAP7_75t_L g854 ( 
.A(n_822),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_685),
.B(n_635),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_790),
.A2(n_578),
.B(n_615),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_765),
.B(n_568),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_790),
.A2(n_578),
.B(n_615),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_739),
.Y(n_859)
);

INVxp67_ASAP7_75t_L g860 ( 
.A(n_761),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_708),
.Y(n_861)
);

OAI21xp33_ASAP7_75t_L g862 ( 
.A1(n_735),
.A2(n_323),
.B(n_339),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_682),
.Y(n_863)
);

BUFx2_ASAP7_75t_L g864 ( 
.A(n_713),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_767),
.B(n_425),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_670),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_755),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_745),
.B(n_291),
.Y(n_868)
);

OAI21xp33_ASAP7_75t_L g869 ( 
.A1(n_735),
.A2(n_322),
.B(n_331),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_745),
.B(n_307),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_731),
.B(n_308),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_760),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_784),
.B(n_568),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_784),
.B(n_568),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_715),
.A2(n_523),
.B(n_552),
.C(n_521),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_696),
.A2(n_627),
.B(n_660),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_686),
.A2(n_568),
.B1(n_662),
.B2(n_574),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_686),
.A2(n_568),
.B1(n_662),
.B2(n_574),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_719),
.B(n_310),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_SL g880 ( 
.A1(n_672),
.A2(n_598),
.B(n_595),
.C(n_590),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_799),
.B(n_568),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_719),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_764),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_799),
.B(n_568),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_722),
.A2(n_638),
.B(n_562),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_709),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_697),
.A2(n_632),
.B(n_660),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_716),
.B(n_428),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_776),
.B(n_313),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_729),
.B(n_314),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_688),
.A2(n_618),
.B1(n_623),
.B2(n_654),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_781),
.B(n_523),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_723),
.A2(n_562),
.B(n_532),
.Y(n_893)
);

O2A1O1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_689),
.A2(n_567),
.B(n_528),
.C(n_541),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_680),
.A2(n_678),
.B(n_815),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_709),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_709),
.B(n_532),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_683),
.A2(n_567),
.B(n_528),
.C(n_541),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_680),
.A2(n_532),
.B(n_562),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_791),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_776),
.B(n_743),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_734),
.B(n_317),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_766),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_823),
.A2(n_562),
.B(n_638),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_734),
.A2(n_569),
.B(n_590),
.C(n_595),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_688),
.A2(n_611),
.B1(n_623),
.B2(n_654),
.Y(n_906)
);

AND2x6_ASAP7_75t_L g907 ( 
.A(n_791),
.B(n_562),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_775),
.B(n_569),
.Y(n_908)
);

INVxp67_ASAP7_75t_L g909 ( 
.A(n_789),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_800),
.B(n_590),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_670),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_714),
.A2(n_638),
.B(n_649),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_705),
.A2(n_638),
.B(n_649),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_730),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_L g915 ( 
.A1(n_698),
.A2(n_565),
.B(n_544),
.C(n_550),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_753),
.A2(n_632),
.B(n_657),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_820),
.A2(n_623),
.B(n_611),
.C(n_654),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_725),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_704),
.Y(n_919)
);

BUFx4f_ASAP7_75t_L g920 ( 
.A(n_758),
.Y(n_920)
);

AOI22xp33_ASAP7_75t_L g921 ( 
.A1(n_724),
.A2(n_662),
.B1(n_555),
.B2(n_550),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_705),
.A2(n_649),
.B(n_638),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_820),
.A2(n_634),
.B1(n_611),
.B2(n_653),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_808),
.Y(n_924)
);

BUFx3_ASAP7_75t_L g925 ( 
.A(n_819),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_736),
.A2(n_649),
.B(n_634),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_791),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_736),
.A2(n_634),
.B(n_618),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_671),
.B(n_618),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_674),
.B(n_653),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_744),
.A2(n_653),
.B(n_570),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_767),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_706),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_712),
.B(n_570),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_812),
.A2(n_584),
.B(n_591),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_814),
.A2(n_584),
.B(n_591),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_772),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_732),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_720),
.A2(n_586),
.B(n_657),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_712),
.B(n_666),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_754),
.A2(n_651),
.B(n_646),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_692),
.A2(n_662),
.B1(n_651),
.B2(n_646),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_757),
.A2(n_662),
.B(n_472),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_762),
.B(n_324),
.Y(n_944)
);

AO21x1_ASAP7_75t_L g945 ( 
.A1(n_774),
.A2(n_472),
.B(n_491),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_752),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_763),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_666),
.B(n_484),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_762),
.B(n_788),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_758),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_666),
.B(n_484),
.Y(n_951)
);

NAND2x1_ASAP7_75t_L g952 ( 
.A(n_737),
.B(n_662),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_666),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_741),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_808),
.Y(n_955)
);

NAND2x1p5_ASAP7_75t_L g956 ( 
.A(n_726),
.B(n_496),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_668),
.B(n_344),
.Y(n_957)
);

INVxp67_ASAP7_75t_L g958 ( 
.A(n_707),
.Y(n_958)
);

NOR2xp67_ASAP7_75t_L g959 ( 
.A(n_703),
.B(n_71),
.Y(n_959)
);

BUFx2_ASAP7_75t_L g960 ( 
.A(n_725),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_777),
.A2(n_462),
.B(n_491),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_788),
.B(n_476),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_793),
.A2(n_475),
.B(n_491),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_782),
.A2(n_341),
.B(n_330),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_821),
.B(n_337),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_807),
.B(n_328),
.Y(n_966)
);

OAI21xp33_ASAP7_75t_L g967 ( 
.A1(n_782),
.A2(n_818),
.B(n_774),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_724),
.A2(n_484),
.B1(n_476),
.B2(n_475),
.Y(n_968)
);

OAI22xp33_ASAP7_75t_L g969 ( 
.A1(n_758),
.A2(n_476),
.B1(n_475),
.B2(n_496),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_687),
.A2(n_779),
.B1(n_750),
.B2(n_740),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_666),
.B(n_475),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_733),
.A2(n_496),
.B(n_173),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_666),
.B(n_496),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_725),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_813),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_813),
.B(n_496),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_738),
.A2(n_496),
.B(n_172),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_695),
.B(n_9),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_756),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_821),
.B(n_10),
.Y(n_980)
);

O2A1O1Ixp5_ASAP7_75t_L g981 ( 
.A1(n_751),
.A2(n_792),
.B(n_786),
.C(n_773),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_780),
.A2(n_170),
.B(n_167),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_771),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_769),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_699),
.B(n_10),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_794),
.Y(n_986)
);

OAI22xp5_ASAP7_75t_L g987 ( 
.A1(n_779),
.A2(n_162),
.B1(n_156),
.B2(n_146),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_778),
.A2(n_11),
.B(n_14),
.C(n_15),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_700),
.B(n_17),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_795),
.A2(n_144),
.B(n_133),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_807),
.B(n_769),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_747),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_992)
);

OAI21xp33_ASAP7_75t_L g993 ( 
.A1(n_818),
.A2(n_22),
.B(n_25),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_797),
.A2(n_127),
.B(n_123),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_803),
.A2(n_115),
.B(n_114),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_728),
.B(n_676),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_804),
.A2(n_106),
.B(n_92),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_806),
.A2(n_86),
.B(n_85),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_679),
.A2(n_68),
.B1(n_67),
.B2(n_27),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_L g1000 ( 
.A(n_702),
.B(n_25),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_810),
.A2(n_26),
.B(n_31),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_796),
.A2(n_34),
.B(n_35),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_681),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_769),
.B(n_34),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_888),
.B(n_768),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_902),
.B(n_816),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_889),
.B(n_816),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_914),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_901),
.B(n_824),
.Y(n_1009)
);

NAND2xp33_ASAP7_75t_SL g1010 ( 
.A(n_950),
.B(n_746),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_946),
.B(n_742),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_L g1012 ( 
.A(n_886),
.B(n_826),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_889),
.B(n_860),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_836),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_826),
.B(n_770),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_953),
.A2(n_805),
.B(n_802),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_847),
.B(n_864),
.Y(n_1017)
);

INVx6_ASAP7_75t_L g1018 ( 
.A(n_903),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_949),
.A2(n_718),
.B1(n_710),
.B2(n_811),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_953),
.A2(n_832),
.B(n_829),
.Y(n_1020)
);

OAI22xp5_ASAP7_75t_SL g1021 ( 
.A1(n_949),
.A2(n_677),
.B1(n_770),
.B2(n_748),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_848),
.A2(n_830),
.B(n_895),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_SL g1023 ( 
.A1(n_962),
.A2(n_798),
.B(n_748),
.C(n_45),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_896),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_849),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_882),
.B(n_35),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_838),
.B(n_40),
.Y(n_1027)
);

AO32x1_ASAP7_75t_L g1028 ( 
.A1(n_999),
.A2(n_46),
.A3(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_854),
.B(n_49),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_896),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_839),
.A2(n_60),
.B(n_53),
.Y(n_1031)
);

OAI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_921),
.A2(n_51),
.B1(n_56),
.B2(n_59),
.Y(n_1032)
);

NOR2xp67_ASAP7_75t_SL g1033 ( 
.A(n_896),
.B(n_900),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_896),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_860),
.B(n_59),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_861),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_909),
.B(n_60),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_909),
.B(n_944),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_937),
.B(n_924),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_924),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_955),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_992),
.A2(n_1000),
.B(n_985),
.C(n_989),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_947),
.B(n_986),
.Y(n_1043)
);

O2A1O1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_978),
.A2(n_967),
.B(n_993),
.C(n_944),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_950),
.B(n_932),
.Y(n_1045)
);

CKINVDCx16_ASAP7_75t_R g1046 ( 
.A(n_837),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1003),
.B(n_940),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_854),
.B(n_859),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_867),
.B(n_872),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_835),
.A2(n_951),
.B(n_948),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_862),
.A2(n_869),
.B(n_988),
.C(n_890),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_883),
.B(n_966),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_L g1053 ( 
.A(n_842),
.B(n_958),
.Y(n_1053)
);

AND2x4_ASAP7_75t_L g1054 ( 
.A(n_950),
.B(n_865),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_958),
.A2(n_874),
.B(n_873),
.C(n_884),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_900),
.Y(n_1056)
);

OAI21xp33_ASAP7_75t_SL g1057 ( 
.A1(n_921),
.A2(n_878),
.B(n_877),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_954),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_934),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_SL g1060 ( 
.A1(n_1004),
.A2(n_960),
.B1(n_974),
.B2(n_918),
.Y(n_1060)
);

CKINVDCx11_ASAP7_75t_R g1061 ( 
.A(n_950),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_955),
.Y(n_1062)
);

NAND3xp33_ASAP7_75t_L g1063 ( 
.A(n_868),
.B(n_870),
.C(n_965),
.Y(n_1063)
);

OA22x2_ASAP7_75t_L g1064 ( 
.A1(n_975),
.A2(n_984),
.B1(n_957),
.B2(n_991),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_868),
.B(n_870),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_865),
.B(n_827),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_855),
.A2(n_971),
.B(n_881),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_996),
.A2(n_840),
.B1(n_828),
.B2(n_857),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_900),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_900),
.B(n_927),
.Y(n_1070)
);

AOI22x1_ASAP7_75t_L g1071 ( 
.A1(n_833),
.A2(n_956),
.B1(n_885),
.B2(n_893),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_954),
.Y(n_1072)
);

INVx3_ASAP7_75t_SL g1073 ( 
.A(n_925),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_879),
.B(n_871),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_879),
.B(n_908),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_929),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_927),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_927),
.B(n_920),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_831),
.A2(n_843),
.B(n_910),
.Y(n_1079)
);

BUFx4f_ASAP7_75t_L g1080 ( 
.A(n_927),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_930),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_886),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_938),
.Y(n_1083)
);

INVx6_ASAP7_75t_L g1084 ( 
.A(n_976),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_877),
.A2(n_878),
.B1(n_970),
.B2(n_976),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_920),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_L g1087 ( 
.A(n_965),
.B(n_980),
.C(n_871),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_L g1088 ( 
.A(n_984),
.B(n_964),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_970),
.A2(n_976),
.B1(n_987),
.B2(n_968),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1004),
.B(n_834),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_938),
.B(n_863),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_851),
.B(n_866),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_968),
.A2(n_969),
.B1(n_998),
.B2(n_990),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_969),
.A2(n_858),
.B1(n_856),
.B2(n_852),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_979),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_844),
.A2(n_911),
.B1(n_866),
.B2(n_959),
.Y(n_1096)
);

INVx6_ASAP7_75t_L g1097 ( 
.A(n_979),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_919),
.B(n_933),
.Y(n_1098)
);

NOR2xp67_ASAP7_75t_L g1099 ( 
.A(n_911),
.B(n_983),
.Y(n_1099)
);

AO32x2_ASAP7_75t_L g1100 ( 
.A1(n_923),
.A2(n_945),
.A3(n_880),
.B1(n_841),
.B2(n_905),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_979),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_892),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_904),
.A2(n_973),
.B(n_846),
.Y(n_1103)
);

CKINVDCx6p67_ASAP7_75t_R g1104 ( 
.A(n_907),
.Y(n_1104)
);

OAI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_917),
.A2(n_956),
.B1(n_891),
.B2(n_906),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_907),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_897),
.B(n_907),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_907),
.Y(n_1108)
);

OAI22x1_ASAP7_75t_L g1109 ( 
.A1(n_942),
.A2(n_845),
.B1(n_997),
.B2(n_1002),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_899),
.A2(n_850),
.B(n_853),
.Y(n_1110)
);

BUFx3_ASAP7_75t_L g1111 ( 
.A(n_907),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1001),
.A2(n_943),
.B1(n_931),
.B2(n_916),
.Y(n_1112)
);

CKINVDCx6p67_ASAP7_75t_R g1113 ( 
.A(n_982),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_952),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_994),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_913),
.A2(n_922),
.B(n_876),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_887),
.B(n_875),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_963),
.A2(n_936),
.B1(n_935),
.B2(n_928),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_981),
.A2(n_894),
.B(n_915),
.C(n_898),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_981),
.B(n_977),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_939),
.A2(n_912),
.B1(n_941),
.B2(n_926),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_961),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_995),
.A2(n_889),
.B(n_902),
.C(n_949),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_SL g1124 ( 
.A(n_972),
.B(n_901),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_836),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_953),
.A2(n_801),
.B(n_759),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_901),
.B(n_946),
.Y(n_1127)
);

O2A1O1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_902),
.A2(n_889),
.B(n_949),
.C(n_992),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_954),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_949),
.A2(n_667),
.B1(n_669),
.B2(n_686),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_847),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_901),
.B(n_946),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_902),
.B(n_809),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_901),
.B(n_946),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_861),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_954),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_902),
.A2(n_889),
.B(n_949),
.C(n_992),
.Y(n_1137)
);

NOR3xp33_ASAP7_75t_SL g1138 ( 
.A(n_949),
.B(n_762),
.C(n_729),
.Y(n_1138)
);

NOR2xp67_ASAP7_75t_L g1139 ( 
.A(n_842),
.B(n_838),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_953),
.A2(n_801),
.B(n_759),
.Y(n_1140)
);

BUFx6f_ASAP7_75t_L g1141 ( 
.A(n_896),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_902),
.B(n_809),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_953),
.A2(n_801),
.B(n_759),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_901),
.B(n_809),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_836),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_902),
.B(n_809),
.Y(n_1146)
);

AND2x4_ASAP7_75t_L g1147 ( 
.A(n_950),
.B(n_909),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_847),
.Y(n_1148)
);

OAI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_949),
.A2(n_667),
.B1(n_669),
.B2(n_686),
.Y(n_1149)
);

INVxp67_ASAP7_75t_L g1150 ( 
.A(n_847),
.Y(n_1150)
);

CKINVDCx8_ASAP7_75t_R g1151 ( 
.A(n_914),
.Y(n_1151)
);

AOI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_902),
.A2(n_889),
.B1(n_949),
.B2(n_545),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_953),
.A2(n_801),
.B(n_759),
.Y(n_1153)
);

O2A1O1Ixp5_ASAP7_75t_SL g1154 ( 
.A1(n_1124),
.A2(n_1093),
.B(n_1121),
.C(n_1144),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1014),
.Y(n_1155)
);

AOI221x1_ASAP7_75t_L g1156 ( 
.A1(n_1123),
.A2(n_1149),
.B1(n_1130),
.B2(n_1093),
.C(n_1063),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1143),
.A2(n_1153),
.B(n_1103),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1134),
.B(n_1127),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1127),
.B(n_1132),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1110),
.A2(n_1116),
.B(n_1071),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1054),
.B(n_1147),
.Y(n_1161)
);

AOI211x1_ASAP7_75t_L g1162 ( 
.A1(n_1130),
.A2(n_1149),
.B(n_1132),
.C(n_1032),
.Y(n_1162)
);

OAI22x1_ASAP7_75t_L g1163 ( 
.A1(n_1152),
.A2(n_1074),
.B1(n_1063),
.B2(n_1087),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1065),
.B(n_1138),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_1128),
.A2(n_1137),
.B(n_1042),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1025),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_SL g1167 ( 
.A1(n_1009),
.A2(n_1013),
.B(n_1075),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1054),
.B(n_1147),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1121),
.A2(n_1022),
.B(n_1050),
.Y(n_1169)
);

CKINVDCx11_ASAP7_75t_R g1170 ( 
.A(n_1151),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1087),
.A2(n_1044),
.B(n_1133),
.C(n_1142),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1079),
.A2(n_1067),
.B(n_1055),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1051),
.A2(n_1146),
.B(n_1038),
.C(n_1090),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1094),
.A2(n_1016),
.B(n_1112),
.Y(n_1174)
);

AOI211x1_ASAP7_75t_L g1175 ( 
.A1(n_1032),
.A2(n_1043),
.B(n_1085),
.C(n_1089),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1109),
.A2(n_1094),
.A3(n_1105),
.B(n_1089),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1117),
.A2(n_1105),
.B(n_1120),
.Y(n_1177)
);

INVx5_ASAP7_75t_L g1178 ( 
.A(n_1106),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1125),
.Y(n_1179)
);

INVx1_ASAP7_75t_SL g1180 ( 
.A(n_1131),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1148),
.B(n_1052),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1119),
.A2(n_1118),
.B(n_1092),
.Y(n_1182)
);

INVx4_ASAP7_75t_L g1183 ( 
.A(n_1080),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1043),
.A2(n_1057),
.B(n_1047),
.Y(n_1184)
);

AO21x1_ASAP7_75t_L g1185 ( 
.A1(n_1068),
.A2(n_1031),
.B(n_1019),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1122),
.A2(n_1047),
.B(n_1107),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_1088),
.A2(n_1053),
.B(n_1007),
.C(n_1006),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1115),
.A2(n_1011),
.B(n_1102),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1019),
.A2(n_1011),
.B(n_1059),
.C(n_1139),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1076),
.B(n_1081),
.Y(n_1190)
);

O2A1O1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1029),
.A2(n_1035),
.B(n_1027),
.C(n_1026),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1049),
.B(n_1145),
.Y(n_1192)
);

AOI221x1_ASAP7_75t_L g1193 ( 
.A1(n_1021),
.A2(n_1060),
.B1(n_1028),
.B2(n_1010),
.C(n_1037),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_SL g1194 ( 
.A1(n_1070),
.A2(n_1048),
.B(n_1114),
.C(n_1098),
.Y(n_1194)
);

AO32x2_ASAP7_75t_L g1195 ( 
.A1(n_1028),
.A2(n_1023),
.A3(n_1064),
.B1(n_1100),
.B2(n_1082),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1048),
.A2(n_1096),
.B(n_1091),
.Y(n_1196)
);

NOR4xp25_ASAP7_75t_L g1197 ( 
.A(n_1015),
.B(n_1028),
.C(n_1066),
.D(n_1005),
.Y(n_1197)
);

INVxp67_ASAP7_75t_SL g1198 ( 
.A(n_1033),
.Y(n_1198)
);

AO21x2_ASAP7_75t_L g1199 ( 
.A1(n_1099),
.A2(n_1100),
.B(n_1072),
.Y(n_1199)
);

CKINVDCx16_ASAP7_75t_R g1200 ( 
.A(n_1078),
.Y(n_1200)
);

BUFx10_ASAP7_75t_L g1201 ( 
.A(n_1018),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1058),
.A2(n_1083),
.B(n_1129),
.C(n_1136),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_L g1203 ( 
.A1(n_1101),
.A2(n_1012),
.B(n_1069),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1045),
.B(n_1150),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1101),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1045),
.B(n_1062),
.Y(n_1206)
);

BUFx3_ASAP7_75t_L g1207 ( 
.A(n_1073),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1106),
.A2(n_1113),
.B(n_1082),
.Y(n_1208)
);

NOR2x1_ASAP7_75t_SL g1209 ( 
.A(n_1111),
.B(n_1141),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1095),
.A2(n_1069),
.B(n_1030),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1100),
.A2(n_1041),
.B(n_1040),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1084),
.B(n_1135),
.Y(n_1212)
);

O2A1O1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1036),
.A2(n_1030),
.B(n_1084),
.C(n_1008),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1024),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1086),
.B(n_1095),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1104),
.A2(n_1097),
.B(n_1095),
.C(n_1056),
.Y(n_1216)
);

INVxp67_ASAP7_75t_SL g1217 ( 
.A(n_1024),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1061),
.A2(n_1097),
.B1(n_1034),
.B2(n_1056),
.Y(n_1218)
);

BUFx8_ASAP7_75t_L g1219 ( 
.A(n_1024),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1034),
.A2(n_1056),
.B(n_1077),
.C(n_1141),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1034),
.A2(n_1077),
.B(n_1141),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1077),
.Y(n_1222)
);

OR2x6_ASAP7_75t_L g1223 ( 
.A(n_1084),
.B(n_758),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1152),
.A2(n_1123),
.B(n_1128),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1134),
.B(n_1127),
.Y(n_1225)
);

AND2x2_ASAP7_75t_L g1226 ( 
.A(n_1065),
.B(n_888),
.Y(n_1226)
);

CKINVDCx11_ASAP7_75t_R g1227 ( 
.A(n_1151),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_1061),
.Y(n_1228)
);

INVx3_ASAP7_75t_L g1229 ( 
.A(n_1106),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1126),
.A2(n_953),
.B(n_1140),
.Y(n_1230)
);

CKINVDCx6p67_ASAP7_75t_R g1231 ( 
.A(n_1073),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1020),
.A2(n_1153),
.B(n_1140),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1093),
.A2(n_1109),
.A3(n_1094),
.B(n_1123),
.Y(n_1233)
);

AOI221x1_ASAP7_75t_L g1234 ( 
.A1(n_1123),
.A2(n_1149),
.B1(n_1130),
.B2(n_1093),
.C(n_1063),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1014),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_1008),
.Y(n_1236)
);

BUFx2_ASAP7_75t_SL g1237 ( 
.A(n_1151),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1093),
.A2(n_1109),
.A3(n_1094),
.B(n_1123),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_SL g1239 ( 
.A1(n_1152),
.A2(n_949),
.B(n_1074),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1131),
.Y(n_1240)
);

INVx2_ASAP7_75t_SL g1241 ( 
.A(n_1018),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1065),
.B(n_888),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1106),
.Y(n_1243)
);

BUFx10_ASAP7_75t_L g1244 ( 
.A(n_1017),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1134),
.B(n_1127),
.Y(n_1245)
);

INVx2_ASAP7_75t_SL g1246 ( 
.A(n_1018),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1061),
.Y(n_1247)
);

NAND2x1_ASAP7_75t_L g1248 ( 
.A(n_1033),
.B(n_907),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1152),
.A2(n_1123),
.B(n_1128),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1152),
.A2(n_1130),
.B1(n_1149),
.B2(n_1085),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1126),
.A2(n_953),
.B(n_1140),
.Y(n_1251)
);

INVx1_ASAP7_75t_SL g1252 ( 
.A(n_1039),
.Y(n_1252)
);

A2O1A1Ixp33_ASAP7_75t_L g1253 ( 
.A1(n_1152),
.A2(n_1128),
.B(n_1137),
.C(n_1074),
.Y(n_1253)
);

OAI22x1_ASAP7_75t_L g1254 ( 
.A1(n_1152),
.A2(n_949),
.B1(n_1074),
.B2(n_1063),
.Y(n_1254)
);

BUFx10_ASAP7_75t_L g1255 ( 
.A(n_1017),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1080),
.Y(n_1256)
);

BUFx10_ASAP7_75t_L g1257 ( 
.A(n_1017),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1126),
.A2(n_953),
.B(n_1140),
.Y(n_1258)
);

INVxp67_ASAP7_75t_L g1259 ( 
.A(n_1017),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1134),
.B(n_1127),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1093),
.A2(n_1109),
.A3(n_1094),
.B(n_1123),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_SL g1262 ( 
.A1(n_1123),
.A2(n_1152),
.B(n_1137),
.C(n_1128),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1061),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1134),
.B(n_1127),
.Y(n_1264)
);

O2A1O1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1074),
.A2(n_1128),
.B(n_1137),
.C(n_902),
.Y(n_1265)
);

NAND3xp33_ASAP7_75t_SL g1266 ( 
.A(n_1152),
.B(n_1074),
.C(n_1128),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_SL g1267 ( 
.A1(n_1123),
.A2(n_1152),
.B(n_1137),
.C(n_1128),
.Y(n_1267)
);

INVxp67_ASAP7_75t_SL g1268 ( 
.A(n_1033),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1152),
.B(n_1074),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1014),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1020),
.A2(n_1153),
.B(n_1140),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_SL g1272 ( 
.A1(n_1123),
.A2(n_1152),
.B(n_1137),
.C(n_1128),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1020),
.A2(n_1153),
.B(n_1140),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1126),
.A2(n_953),
.B(n_1140),
.Y(n_1274)
);

NOR2xp33_ASAP7_75t_L g1275 ( 
.A(n_1152),
.B(n_1074),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1074),
.A2(n_1128),
.B(n_1137),
.C(n_902),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1126),
.A2(n_953),
.B(n_1140),
.Y(n_1277)
);

AOI221xp5_ASAP7_75t_L g1278 ( 
.A1(n_1074),
.A2(n_949),
.B1(n_944),
.B2(n_370),
.C(n_513),
.Y(n_1278)
);

OAI21xp33_ASAP7_75t_L g1279 ( 
.A1(n_1074),
.A2(n_1152),
.B(n_949),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_1017),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1022),
.A2(n_1055),
.B(n_833),
.Y(n_1281)
);

AO31x2_ASAP7_75t_L g1282 ( 
.A1(n_1093),
.A2(n_1109),
.A3(n_1094),
.B(n_1123),
.Y(n_1282)
);

AOI221x1_ASAP7_75t_L g1283 ( 
.A1(n_1123),
.A2(n_1149),
.B1(n_1130),
.B2(n_1093),
.C(n_1063),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1134),
.B(n_1127),
.Y(n_1284)
);

O2A1O1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1074),
.A2(n_1128),
.B(n_1137),
.C(n_902),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1152),
.A2(n_1123),
.B(n_1128),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1152),
.B(n_1074),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1152),
.A2(n_1130),
.B1(n_1149),
.B2(n_1085),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1134),
.B(n_1127),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1061),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1018),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1123),
.A2(n_953),
.B(n_1093),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1093),
.A2(n_1109),
.A3(n_1094),
.B(n_1123),
.Y(n_1293)
);

INVx2_ASAP7_75t_SL g1294 ( 
.A(n_1201),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1201),
.Y(n_1295)
);

AOI22x1_ASAP7_75t_SL g1296 ( 
.A1(n_1236),
.A2(n_1183),
.B1(n_1256),
.B2(n_1198),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_SL g1297 ( 
.A1(n_1275),
.A2(n_1287),
.B(n_1278),
.Y(n_1297)
);

CKINVDCx11_ASAP7_75t_R g1298 ( 
.A(n_1170),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1207),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1250),
.A2(n_1288),
.B1(n_1224),
.B2(n_1286),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1155),
.Y(n_1301)
);

OAI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1239),
.A2(n_1269),
.B1(n_1250),
.B2(n_1288),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1279),
.A2(n_1266),
.B1(n_1254),
.B2(n_1163),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1239),
.A2(n_1234),
.B1(n_1283),
.B2(n_1156),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1224),
.A2(n_1286),
.B1(n_1249),
.B2(n_1164),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1279),
.A2(n_1249),
.B1(n_1165),
.B2(n_1185),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1166),
.Y(n_1307)
);

OAI21xp33_ASAP7_75t_L g1308 ( 
.A1(n_1253),
.A2(n_1173),
.B(n_1265),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1179),
.Y(n_1309)
);

CKINVDCx10_ASAP7_75t_R g1310 ( 
.A(n_1200),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1227),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_SL g1312 ( 
.A1(n_1228),
.A2(n_1263),
.B1(n_1247),
.B2(n_1290),
.Y(n_1312)
);

BUFx8_ASAP7_75t_L g1313 ( 
.A(n_1228),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1226),
.A2(n_1242),
.B1(n_1225),
.B2(n_1284),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_SL g1315 ( 
.A1(n_1175),
.A2(n_1237),
.B1(n_1159),
.B2(n_1264),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1158),
.A2(n_1260),
.B1(n_1245),
.B2(n_1289),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1270),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_SL g1318 ( 
.A(n_1228),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1192),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1252),
.A2(n_1259),
.B1(n_1181),
.B2(n_1174),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1190),
.Y(n_1321)
);

AO22x2_ASAP7_75t_L g1322 ( 
.A1(n_1175),
.A2(n_1193),
.B1(n_1162),
.B2(n_1172),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1184),
.A2(n_1180),
.B1(n_1161),
.B2(n_1168),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1231),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1247),
.Y(n_1325)
);

BUFx12f_ASAP7_75t_L g1326 ( 
.A(n_1263),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1162),
.A2(n_1263),
.B1(n_1290),
.B2(n_1262),
.Y(n_1327)
);

CKINVDCx6p67_ASAP7_75t_R g1328 ( 
.A(n_1290),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1276),
.A2(n_1285),
.B1(n_1187),
.B2(n_1191),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1267),
.A2(n_1272),
.B1(n_1281),
.B2(n_1292),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1218),
.A2(n_1206),
.B1(n_1223),
.B2(n_1204),
.Y(n_1331)
);

CKINVDCx11_ASAP7_75t_R g1332 ( 
.A(n_1244),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1244),
.A2(n_1255),
.B1(n_1280),
.B2(n_1257),
.Y(n_1333)
);

OAI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1171),
.A2(n_1189),
.B1(n_1223),
.B2(n_1218),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1211),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1219),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1280),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1188),
.A2(n_1281),
.B1(n_1196),
.B2(n_1223),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1212),
.B(n_1215),
.Y(n_1339)
);

CKINVDCx11_ASAP7_75t_R g1340 ( 
.A(n_1183),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1211),
.A2(n_1209),
.B1(n_1268),
.B2(n_1256),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1182),
.A2(n_1199),
.B1(n_1186),
.B2(n_1169),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1178),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1199),
.A2(n_1214),
.B1(n_1222),
.B2(n_1243),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1208),
.A2(n_1160),
.B1(n_1167),
.B2(n_1229),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1202),
.Y(n_1346)
);

BUFx4f_ASAP7_75t_SL g1347 ( 
.A(n_1241),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_SL g1348 ( 
.A1(n_1176),
.A2(n_1197),
.B1(n_1293),
.B2(n_1238),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1243),
.A2(n_1205),
.B1(n_1217),
.B2(n_1230),
.Y(n_1349)
);

BUFx4f_ASAP7_75t_SL g1350 ( 
.A(n_1246),
.Y(n_1350)
);

OAI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1177),
.A2(n_1248),
.B1(n_1291),
.B2(n_1210),
.Y(n_1351)
);

INVx3_ASAP7_75t_SL g1352 ( 
.A(n_1213),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1176),
.A2(n_1197),
.B1(n_1293),
.B2(n_1282),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1176),
.A2(n_1238),
.B1(n_1282),
.B2(n_1261),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1221),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1203),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1216),
.Y(n_1357)
);

OAI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1233),
.A2(n_1293),
.B1(n_1282),
.B2(n_1261),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1220),
.Y(n_1359)
);

INVx1_ASAP7_75t_SL g1360 ( 
.A(n_1251),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1195),
.Y(n_1361)
);

CKINVDCx11_ASAP7_75t_R g1362 ( 
.A(n_1154),
.Y(n_1362)
);

BUFx12f_ASAP7_75t_L g1363 ( 
.A(n_1194),
.Y(n_1363)
);

OAI22x1_ASAP7_75t_L g1364 ( 
.A1(n_1195),
.A2(n_1238),
.B1(n_1157),
.B2(n_1232),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1195),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1258),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1274),
.A2(n_1277),
.B1(n_1271),
.B2(n_1273),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1368)
);

BUFx8_ASAP7_75t_L g1369 ( 
.A(n_1228),
.Y(n_1369)
);

AOI22xp33_ASAP7_75t_SL g1370 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1130),
.B2(n_1149),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1235),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1240),
.Y(n_1373)
);

BUFx8_ASAP7_75t_L g1374 ( 
.A(n_1228),
.Y(n_1374)
);

OAI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1275),
.A2(n_1152),
.B1(n_1130),
.B2(n_1149),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1130),
.B2(n_1149),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1269),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1201),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1235),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_SL g1384 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_949),
.B2(n_1046),
.Y(n_1384)
);

NAND2x1p5_ASAP7_75t_L g1385 ( 
.A(n_1178),
.B(n_1033),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1236),
.Y(n_1386)
);

BUFx2_ASAP7_75t_SL g1387 ( 
.A(n_1201),
.Y(n_1387)
);

NOR2x1_ASAP7_75t_L g1388 ( 
.A(n_1158),
.B(n_1225),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1201),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1275),
.B(n_1287),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1235),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1152),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1170),
.Y(n_1395)
);

BUFx4f_ASAP7_75t_SL g1396 ( 
.A(n_1231),
.Y(n_1396)
);

CKINVDCx11_ASAP7_75t_R g1397 ( 
.A(n_1170),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1279),
.B2(n_1269),
.Y(n_1398)
);

BUFx6f_ASAP7_75t_L g1399 ( 
.A(n_1178),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1130),
.B2(n_1149),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_R g1401 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_949),
.B2(n_944),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1130),
.B2(n_1149),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1275),
.A2(n_1287),
.B1(n_1130),
.B2(n_1149),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1170),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1298),
.Y(n_1405)
);

INVx3_ASAP7_75t_L g1406 ( 
.A(n_1356),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1335),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1305),
.B(n_1300),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1305),
.B(n_1300),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1322),
.B(n_1370),
.Y(n_1410)
);

INVx3_ASAP7_75t_L g1411 ( 
.A(n_1360),
.Y(n_1411)
);

NOR2x1_ASAP7_75t_R g1412 ( 
.A(n_1395),
.B(n_1397),
.Y(n_1412)
);

OA21x2_ASAP7_75t_L g1413 ( 
.A1(n_1342),
.A2(n_1306),
.B(n_1365),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1366),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1364),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1322),
.B(n_1370),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1361),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1361),
.Y(n_1418)
);

A2O1A1Ixp33_ASAP7_75t_SL g1419 ( 
.A1(n_1303),
.A2(n_1329),
.B(n_1381),
.C(n_1383),
.Y(n_1419)
);

BUFx4f_ASAP7_75t_SL g1420 ( 
.A(n_1325),
.Y(n_1420)
);

INVx2_ASAP7_75t_L g1421 ( 
.A(n_1322),
.Y(n_1421)
);

AOI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1334),
.A2(n_1346),
.B(n_1359),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1301),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1307),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1342),
.A2(n_1345),
.B(n_1338),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1376),
.B(n_1400),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1358),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1401),
.A2(n_1376),
.B1(n_1403),
.B2(n_1400),
.Y(n_1428)
);

BUFx2_ASAP7_75t_SL g1429 ( 
.A(n_1318),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1358),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1297),
.A2(n_1308),
.B(n_1391),
.Y(n_1431)
);

INVxp67_ASAP7_75t_SL g1432 ( 
.A(n_1316),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1354),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1354),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1402),
.A2(n_1403),
.B1(n_1380),
.B2(n_1371),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1345),
.B(n_1317),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1309),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1368),
.A2(n_1379),
.B(n_1394),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1402),
.B(n_1348),
.Y(n_1439)
);

INVxp67_ASAP7_75t_L g1440 ( 
.A(n_1388),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1373),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1348),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1353),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1355),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1344),
.A2(n_1323),
.B(n_1349),
.Y(n_1445)
);

INVx3_ASAP7_75t_L g1446 ( 
.A(n_1363),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_L g1447 ( 
.A(n_1362),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1353),
.B(n_1377),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1392),
.B(n_1384),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1377),
.B(n_1398),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1389),
.A2(n_1375),
.B1(n_1398),
.B2(n_1302),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1375),
.A2(n_1302),
.B1(n_1327),
.B2(n_1304),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1304),
.B(n_1320),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1315),
.B(n_1327),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1382),
.Y(n_1455)
);

AOI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1393),
.A2(n_1321),
.B(n_1319),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1367),
.A2(n_1316),
.B(n_1351),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1314),
.B(n_1315),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1330),
.B(n_1372),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1330),
.B(n_1331),
.Y(n_1460)
);

BUFx4f_ASAP7_75t_L g1461 ( 
.A(n_1385),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1351),
.Y(n_1462)
);

INVx11_ASAP7_75t_L g1463 ( 
.A(n_1313),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1352),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1336),
.A2(n_1333),
.B1(n_1337),
.B2(n_1339),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1310),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1367),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1341),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1341),
.A2(n_1357),
.B(n_1343),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_SL g1470 ( 
.A1(n_1312),
.A2(n_1296),
.B1(n_1318),
.B2(n_1336),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1399),
.Y(n_1471)
);

INVx3_ASAP7_75t_L g1472 ( 
.A(n_1336),
.Y(n_1472)
);

HB1xp67_ASAP7_75t_L g1473 ( 
.A(n_1294),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1340),
.A2(n_1332),
.B(n_1328),
.Y(n_1474)
);

AO21x2_ASAP7_75t_L g1475 ( 
.A1(n_1387),
.A2(n_1390),
.B(n_1295),
.Y(n_1475)
);

BUFx12f_ASAP7_75t_L g1476 ( 
.A(n_1313),
.Y(n_1476)
);

OAI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1378),
.A2(n_1396),
.B1(n_1299),
.B2(n_1390),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1396),
.A2(n_1374),
.B(n_1369),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1347),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1469),
.B(n_1326),
.Y(n_1480)
);

INVx5_ASAP7_75t_SL g1481 ( 
.A(n_1463),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1431),
.A2(n_1324),
.B(n_1311),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1437),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1431),
.A2(n_1404),
.B1(n_1386),
.B2(n_1350),
.C(n_1347),
.Y(n_1484)
);

AO22x2_ASAP7_75t_L g1485 ( 
.A1(n_1427),
.A2(n_1350),
.B1(n_1386),
.B2(n_1430),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1438),
.A2(n_1451),
.B(n_1419),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_1466),
.Y(n_1487)
);

NOR2x1_ASAP7_75t_SL g1488 ( 
.A(n_1475),
.B(n_1457),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1428),
.A2(n_1452),
.B1(n_1435),
.B2(n_1408),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1437),
.Y(n_1490)
);

NAND2x1p5_ASAP7_75t_L g1491 ( 
.A(n_1411),
.B(n_1469),
.Y(n_1491)
);

OAI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1438),
.A2(n_1449),
.B(n_1450),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1408),
.A2(n_1409),
.B1(n_1426),
.B2(n_1453),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1450),
.A2(n_1432),
.B(n_1460),
.Y(n_1494)
);

CKINVDCx16_ASAP7_75t_R g1495 ( 
.A(n_1405),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1432),
.B(n_1410),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1467),
.A2(n_1425),
.B(n_1457),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1410),
.B(n_1416),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1409),
.A2(n_1426),
.B1(n_1454),
.B2(n_1439),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1475),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1464),
.A2(n_1460),
.B(n_1414),
.C(n_1453),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1454),
.A2(n_1458),
.B1(n_1439),
.B2(n_1447),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1464),
.B(n_1465),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1445),
.A2(n_1448),
.B(n_1461),
.C(n_1468),
.Y(n_1504)
);

AND2x4_ASAP7_75t_L g1505 ( 
.A(n_1417),
.B(n_1418),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1422),
.A2(n_1445),
.B(n_1440),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1465),
.A2(n_1470),
.B1(n_1477),
.B2(n_1447),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1444),
.B(n_1441),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1444),
.A2(n_1462),
.B(n_1411),
.Y(n_1509)
);

O2A1O1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1477),
.A2(n_1441),
.B(n_1411),
.C(n_1473),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1461),
.A2(n_1447),
.B(n_1474),
.C(n_1446),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1423),
.B(n_1424),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1456),
.A2(n_1461),
.B(n_1436),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1447),
.A2(n_1474),
.B(n_1446),
.C(n_1478),
.Y(n_1514)
);

AOI221xp5_ASAP7_75t_L g1515 ( 
.A1(n_1442),
.A2(n_1443),
.B1(n_1427),
.B2(n_1430),
.C(n_1433),
.Y(n_1515)
);

AO32x2_ASAP7_75t_L g1516 ( 
.A1(n_1421),
.A2(n_1471),
.A3(n_1443),
.B1(n_1442),
.B2(n_1433),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1483),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1490),
.Y(n_1518)
);

NOR2xp33_ASAP7_75t_R g1519 ( 
.A(n_1487),
.B(n_1476),
.Y(n_1519)
);

AOI22xp33_ASAP7_75t_L g1520 ( 
.A1(n_1486),
.A2(n_1447),
.B1(n_1434),
.B2(n_1421),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1498),
.B(n_1415),
.Y(n_1521)
);

NOR2xp67_ASAP7_75t_L g1522 ( 
.A(n_1500),
.B(n_1407),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1495),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1482),
.B(n_1472),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1512),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1512),
.Y(n_1526)
);

OAI221xp5_ASAP7_75t_SL g1527 ( 
.A1(n_1501),
.A2(n_1434),
.B1(n_1459),
.B2(n_1479),
.C(n_1446),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1497),
.B(n_1413),
.Y(n_1528)
);

INVxp67_ASAP7_75t_SL g1529 ( 
.A(n_1509),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1497),
.B(n_1413),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1480),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_SL g1532 ( 
.A(n_1508),
.B(n_1459),
.Y(n_1532)
);

NAND2x1_ASAP7_75t_L g1533 ( 
.A(n_1480),
.B(n_1406),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1516),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1491),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1516),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1516),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1482),
.B(n_1472),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1528),
.B(n_1530),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1517),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1542)
);

OAI33xp33_ASAP7_75t_L g1543 ( 
.A1(n_1534),
.A2(n_1489),
.A3(n_1493),
.B1(n_1502),
.B2(n_1496),
.B3(n_1455),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1528),
.B(n_1505),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1533),
.A2(n_1506),
.B(n_1513),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_SL g1546 ( 
.A1(n_1529),
.A2(n_1492),
.B1(n_1486),
.B2(n_1489),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1536),
.B(n_1496),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1521),
.B(n_1492),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1535),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1537),
.B(n_1506),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1520),
.A2(n_1494),
.B1(n_1499),
.B2(n_1502),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1530),
.B(n_1491),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1524),
.A2(n_1494),
.B1(n_1499),
.B2(n_1493),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1518),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1518),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1537),
.B(n_1515),
.Y(n_1556)
);

AND2x2_ASAP7_75t_SL g1557 ( 
.A(n_1531),
.B(n_1447),
.Y(n_1557)
);

OR2x6_ASAP7_75t_L g1558 ( 
.A(n_1535),
.B(n_1513),
.Y(n_1558)
);

OA21x2_ASAP7_75t_L g1559 ( 
.A1(n_1522),
.A2(n_1504),
.B(n_1509),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1539),
.B(n_1529),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1550),
.B(n_1532),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1542),
.B(n_1549),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1539),
.B(n_1531),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1550),
.B(n_1532),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1541),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1548),
.B(n_1521),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1548),
.B(n_1525),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1541),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1541),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1549),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1554),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1542),
.B(n_1549),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1556),
.B(n_1525),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1556),
.B(n_1547),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1540),
.B(n_1535),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1556),
.B(n_1526),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1540),
.B(n_1535),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1542),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1555),
.Y(n_1579)
);

INVxp67_ASAP7_75t_SL g1580 ( 
.A(n_1573),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1578),
.B(n_1552),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1565),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1578),
.A2(n_1546),
.B1(n_1551),
.B2(n_1543),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1569),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1578),
.B(n_1552),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1569),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1567),
.B(n_1546),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1561),
.B(n_1550),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1570),
.B(n_1511),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1562),
.B(n_1542),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1563),
.B(n_1552),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1561),
.A2(n_1553),
.B(n_1551),
.C(n_1503),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1562),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1567),
.B(n_1553),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1579),
.Y(n_1595)
);

NOR2x1p5_ASAP7_75t_L g1596 ( 
.A(n_1561),
.B(n_1476),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1562),
.B(n_1542),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1579),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1552),
.Y(n_1599)
);

INVx3_ASAP7_75t_SL g1600 ( 
.A(n_1570),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1563),
.B(n_1540),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1568),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1568),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1566),
.B(n_1547),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1564),
.A2(n_1557),
.B(n_1542),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1562),
.B(n_1540),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1571),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1571),
.Y(n_1611)
);

OAI21xp5_ASAP7_75t_SL g1612 ( 
.A1(n_1564),
.A2(n_1507),
.B(n_1484),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1562),
.B(n_1542),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1564),
.B(n_1550),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1572),
.B(n_1542),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1576),
.B(n_1544),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1602),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1602),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1582),
.Y(n_1619)
);

AOI32xp33_ASAP7_75t_L g1620 ( 
.A1(n_1583),
.A2(n_1484),
.A3(n_1560),
.B1(n_1485),
.B2(n_1574),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1604),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1604),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1587),
.B(n_1594),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1600),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1589),
.B(n_1572),
.Y(n_1625)
);

OR2x6_ASAP7_75t_L g1626 ( 
.A(n_1596),
.B(n_1429),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1607),
.Y(n_1627)
);

XOR2xp5_ASAP7_75t_L g1628 ( 
.A(n_1590),
.B(n_1523),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1607),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1589),
.B(n_1572),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1589),
.B(n_1593),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1589),
.B(n_1572),
.Y(n_1632)
);

AND2x4_ASAP7_75t_L g1633 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1610),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1610),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1590),
.B(n_1570),
.Y(n_1636)
);

INVxp67_ASAP7_75t_SL g1637 ( 
.A(n_1593),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1600),
.Y(n_1638)
);

NAND2x1_ASAP7_75t_L g1639 ( 
.A(n_1590),
.B(n_1575),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1591),
.B(n_1575),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1611),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1612),
.B(n_1592),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1591),
.B(n_1575),
.Y(n_1643)
);

NAND2x1p5_ASAP7_75t_L g1644 ( 
.A(n_1590),
.B(n_1559),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1582),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1606),
.B(n_1560),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1599),
.B(n_1577),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1600),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1584),
.Y(n_1649)
);

AOI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1580),
.A2(n_1559),
.B(n_1538),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1560),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1599),
.B(n_1577),
.Y(n_1652)
);

OAI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1642),
.A2(n_1608),
.B(n_1545),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_SL g1654 ( 
.A1(n_1623),
.A2(n_1559),
.B1(n_1557),
.B2(n_1597),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1620),
.A2(n_1412),
.B(n_1543),
.Y(n_1655)
);

AOI222xp33_ASAP7_75t_L g1656 ( 
.A1(n_1620),
.A2(n_1605),
.B1(n_1557),
.B2(n_1585),
.C1(n_1581),
.C2(n_1586),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_SL g1657 ( 
.A1(n_1628),
.A2(n_1586),
.B(n_1584),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1631),
.B(n_1581),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1646),
.B(n_1616),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1638),
.B(n_1585),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1617),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1628),
.A2(n_1527),
.B1(n_1559),
.B2(n_1558),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1617),
.Y(n_1663)
);

NOR2xp67_ASAP7_75t_SL g1664 ( 
.A(n_1624),
.B(n_1476),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1631),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1638),
.B(n_1601),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1650),
.A2(n_1624),
.B(n_1637),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1633),
.A2(n_1527),
.B1(n_1559),
.B2(n_1558),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1648),
.B(n_1601),
.Y(n_1669)
);

NOR3xp33_ASAP7_75t_L g1670 ( 
.A(n_1648),
.B(n_1412),
.C(n_1514),
.Y(n_1670)
);

OAI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1633),
.A2(n_1559),
.B1(n_1558),
.B2(n_1557),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1640),
.Y(n_1672)
);

NAND2xp33_ASAP7_75t_SL g1673 ( 
.A(n_1639),
.B(n_1519),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1633),
.B(n_1420),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1651),
.B(n_1588),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1618),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1640),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1625),
.B(n_1609),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1661),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1663),
.Y(n_1680)
);

AOI21xp33_ASAP7_75t_L g1681 ( 
.A1(n_1656),
.A2(n_1626),
.B(n_1639),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1658),
.B(n_1633),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1676),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1665),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1665),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1658),
.B(n_1626),
.Y(n_1686)
);

NOR3xp33_ASAP7_75t_SL g1687 ( 
.A(n_1673),
.B(n_1621),
.C(n_1618),
.Y(n_1687)
);

OAI211xp5_ASAP7_75t_L g1688 ( 
.A1(n_1655),
.A2(n_1649),
.B(n_1630),
.C(n_1625),
.Y(n_1688)
);

OAI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1667),
.A2(n_1626),
.B1(n_1644),
.B2(n_1588),
.C(n_1614),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1652),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1678),
.B(n_1672),
.Y(n_1691)
);

A2O1A1Ixp33_ASAP7_75t_L g1692 ( 
.A1(n_1670),
.A2(n_1474),
.B(n_1510),
.C(n_1614),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1654),
.A2(n_1626),
.B1(n_1644),
.B2(n_1557),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1662),
.A2(n_1626),
.B1(n_1597),
.B2(n_1630),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1674),
.B(n_1463),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1672),
.Y(n_1696)
);

OAI211xp5_ASAP7_75t_L g1697 ( 
.A1(n_1673),
.A2(n_1632),
.B(n_1622),
.C(n_1627),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1678),
.Y(n_1698)
);

XNOR2xp5_ASAP7_75t_L g1699 ( 
.A(n_1682),
.B(n_1666),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1682),
.A2(n_1664),
.B1(n_1674),
.B2(n_1677),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1691),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1691),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1688),
.A2(n_1668),
.B(n_1653),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1698),
.A2(n_1677),
.B1(n_1669),
.B2(n_1632),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1684),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1695),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1684),
.Y(n_1707)
);

OAI211xp5_ASAP7_75t_SL g1708 ( 
.A1(n_1687),
.A2(n_1657),
.B(n_1675),
.C(n_1659),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1698),
.B(n_1643),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1685),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1702),
.Y(n_1711)
);

INVx1_ASAP7_75t_SL g1712 ( 
.A(n_1709),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1701),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1699),
.B(n_1696),
.Y(n_1714)
);

O2A1O1Ixp33_ASAP7_75t_L g1715 ( 
.A1(n_1708),
.A2(n_1692),
.B(n_1681),
.C(n_1689),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1704),
.B(n_1690),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1710),
.B(n_1700),
.Y(n_1717)
);

NOR4xp25_ASAP7_75t_L g1718 ( 
.A(n_1708),
.B(n_1683),
.C(n_1679),
.D(n_1680),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1705),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1718),
.A2(n_1703),
.B1(n_1692),
.B2(n_1693),
.C(n_1697),
.Y(n_1720)
);

NAND3xp33_ASAP7_75t_L g1721 ( 
.A(n_1715),
.B(n_1707),
.C(n_1706),
.Y(n_1721)
);

AOI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1712),
.A2(n_1686),
.B(n_1683),
.C(n_1671),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1717),
.A2(n_1694),
.B(n_1686),
.C(n_1644),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1714),
.A2(n_1636),
.B1(n_1597),
.B2(n_1647),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1720),
.B(n_1713),
.Y(n_1725)
);

OAI211xp5_ASAP7_75t_L g1726 ( 
.A1(n_1721),
.A2(n_1713),
.B(n_1716),
.C(n_1711),
.Y(n_1726)
);

OAI211xp5_ASAP7_75t_L g1727 ( 
.A1(n_1723),
.A2(n_1719),
.B(n_1478),
.C(n_1641),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1724),
.Y(n_1728)
);

NAND5xp2_ASAP7_75t_L g1729 ( 
.A(n_1722),
.B(n_1615),
.C(n_1613),
.D(n_1652),
.E(n_1643),
.Y(n_1729)
);

OAI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1720),
.A2(n_1634),
.B1(n_1629),
.B2(n_1622),
.C(n_1621),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1728),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1726),
.Y(n_1732)
);

NOR2xp67_ASAP7_75t_L g1733 ( 
.A(n_1727),
.B(n_1627),
.Y(n_1733)
);

NAND4xp75_ASAP7_75t_L g1734 ( 
.A(n_1725),
.B(n_1629),
.C(n_1641),
.D(n_1635),
.Y(n_1734)
);

INVxp67_ASAP7_75t_SL g1735 ( 
.A(n_1730),
.Y(n_1735)
);

A2O1A1Ixp33_ASAP7_75t_L g1736 ( 
.A1(n_1732),
.A2(n_1735),
.B(n_1733),
.C(n_1731),
.Y(n_1736)
);

OR3x2_ASAP7_75t_L g1737 ( 
.A(n_1734),
.B(n_1729),
.C(n_1429),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1733),
.B(n_1636),
.Y(n_1738)
);

OAI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1634),
.B1(n_1635),
.B2(n_1619),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1737),
.B1(n_1736),
.B2(n_1636),
.Y(n_1740)
);

AND2x4_ASAP7_75t_L g1741 ( 
.A(n_1740),
.B(n_1636),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1740),
.Y(n_1742)
);

OAI22x1_ASAP7_75t_L g1743 ( 
.A1(n_1742),
.A2(n_1741),
.B1(n_1479),
.B2(n_1645),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1645),
.B1(n_1619),
.B2(n_1598),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1743),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1744),
.A2(n_1645),
.B(n_1619),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1745),
.B(n_1481),
.Y(n_1747)
);

AOI21xp33_ASAP7_75t_L g1748 ( 
.A1(n_1747),
.A2(n_1746),
.B(n_1478),
.Y(n_1748)
);

XNOR2xp5_ASAP7_75t_L g1749 ( 
.A(n_1748),
.B(n_1479),
.Y(n_1749)
);

OAI221xp5_ASAP7_75t_R g1750 ( 
.A1(n_1749),
.A2(n_1481),
.B1(n_1595),
.B2(n_1598),
.C(n_1597),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1750),
.A2(n_1473),
.B(n_1481),
.C(n_1595),
.Y(n_1751)
);


endmodule