module fake_jpeg_20045_n_176 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_176);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_176;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_10),
.B(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_18),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_46),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_40),
.B(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_32),
.B(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_29),
.B(n_28),
.C(n_14),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_48),
.B(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_32),
.B(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_26),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_31),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_54),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_21),
.B1(n_37),
.B2(n_36),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_57),
.B(n_58),
.Y(n_89)
);

NOR2x1_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_34),
.Y(n_59)
);

OR2x4_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_30),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_61),
.B(n_70),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_67),
.Y(n_79)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_27),
.B1(n_15),
.B2(n_23),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_69),
.Y(n_86)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_44),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_39),
.B(n_33),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_40),
.B1(n_33),
.B2(n_36),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_75),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_36),
.B1(n_47),
.B2(n_37),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_78),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_70),
.A2(n_42),
.B1(n_51),
.B2(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_80),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_14),
.B1(n_21),
.B2(n_16),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_65),
.A2(n_14),
.B1(n_40),
.B2(n_21),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_64),
.A2(n_35),
.B1(n_22),
.B2(n_27),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_88),
.B(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_49),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_55),
.B(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_87),
.B(n_60),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_35),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_101),
.Y(n_117)
);

AND2x6_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_60),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_91),
.B(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_72),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_106),
.B1(n_73),
.B2(n_85),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_97),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_69),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_58),
.C(n_62),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_77),
.C(n_88),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_71),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_79),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_110),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_88),
.B1(n_86),
.B2(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_114),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_106),
.C(n_99),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_86),
.B(n_89),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_86),
.B1(n_68),
.B2(n_67),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_119),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_15),
.A3(n_20),
.B1(n_24),
.B2(n_28),
.C1(n_12),
.C2(n_7),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_120),
.C(n_103),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_62),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_74),
.B1(n_62),
.B2(n_53),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g120 ( 
.A1(n_98),
.A2(n_0),
.B(n_1),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_100),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_113),
.C(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_130),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_118),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_132),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_98),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_117),
.Y(n_135)
);

OA21x2_ASAP7_75t_SL g149 ( 
.A1(n_136),
.A2(n_125),
.B(n_120),
.Y(n_149)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_90),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_139),
.Y(n_148)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_128),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_125),
.C(n_127),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_114),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_28),
.C(n_24),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_107),
.B(n_115),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_127),
.B(n_119),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_152),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_143),
.A2(n_146),
.B1(n_133),
.B2(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_154),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_140),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_SL g157 ( 
.A1(n_147),
.A2(n_145),
.B(n_138),
.C(n_142),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_151),
.A2(n_144),
.B(n_141),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_161),
.Y(n_165)
);

NAND4xp25_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_8),
.C(n_13),
.D(n_53),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_2),
.B(n_3),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_8),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_152),
.C(n_154),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

INVx11_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_157),
.A2(n_151),
.B(n_3),
.C(n_4),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_2),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_165),
.B(n_155),
.C(n_20),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_167),
.A2(n_168),
.B1(n_166),
.B2(n_163),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_169),
.A2(n_2),
.B(n_4),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_167),
.B(n_170),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_173),
.A3(n_170),
.B1(n_168),
.B2(n_6),
.C1(n_5),
.C2(n_24),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_175),
.B(n_20),
.Y(n_176)
);


endmodule