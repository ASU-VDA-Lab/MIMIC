module fake_netlist_6_4034_n_722 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_722);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_722;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_344;
wire n_581;
wire n_428;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_681;
wire n_151;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_17),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_25),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_51),
.Y(n_151)
);

NOR2xp67_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_21),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_6),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_134),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_23),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_11),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_37),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_121),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_20),
.Y(n_163)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_49),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_40),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_70),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_8),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_17),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_12),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_5),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_6),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_0),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_39),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_34),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_89),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_38),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_53),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_62),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_67),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_30),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_18),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_119),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_84),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_0),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_74),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_28),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_114),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_42),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_15),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_111),
.B(n_9),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_105),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_83),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_147),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_193),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_146),
.B(n_1),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_1),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_193),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_145),
.B(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_171),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_168),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_185),
.Y(n_211)
);

AND2x6_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_22),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

CKINVDCx11_ASAP7_75t_R g214 ( 
.A(n_185),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_160),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_193),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_145),
.B(n_2),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_150),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_179),
.B(n_3),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_163),
.B(n_3),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_149),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_157),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_170),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_158),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_165),
.Y(n_234)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_187),
.B(n_4),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_7),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_191),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_222),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_195),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_187),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_216),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_219),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_220),
.Y(n_250)
);

OR2x6_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_152),
.Y(n_251)
);

AND2x4_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_197),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_161),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_164),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_224),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_223),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_235),
.B(n_211),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_223),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_221),
.B(n_180),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_205),
.Y(n_267)
);

CKINVDCx8_ASAP7_75t_R g268 ( 
.A(n_210),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_198),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_222),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_205),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_225),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_206),
.Y(n_273)
);

INVx8_ASAP7_75t_L g274 ( 
.A(n_200),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_154),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_222),
.B(n_198),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_203),
.B(n_210),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_225),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_218),
.B(n_151),
.Y(n_279)
);

AND2x6_ASAP7_75t_L g280 ( 
.A(n_222),
.B(n_24),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_159),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_L g282 ( 
.A(n_207),
.B(n_173),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_218),
.B(n_162),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_206),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_230),
.B(n_161),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_214),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_217),
.B(n_166),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_209),
.B(n_174),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_247),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_238),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_200),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_251),
.A2(n_232),
.B1(n_192),
.B2(n_186),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_251),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_200),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_230),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_246),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_200),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_255),
.B(n_228),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_267),
.B(n_200),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_248),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_231),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_231),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_271),
.B(n_233),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_271),
.B(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_255),
.B(n_175),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_277),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_248),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_246),
.B(n_233),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_254),
.B(n_186),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_266),
.B(n_237),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_266),
.B(n_237),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_240),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_252),
.B(n_178),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_249),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_276),
.B(n_240),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_242),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_269),
.B(n_242),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_243),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_270),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_288),
.B(n_236),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_252),
.B(n_182),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g331 ( 
.A1(n_251),
.A2(n_212),
.B1(n_236),
.B2(n_215),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_252),
.B(n_183),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_252),
.B(n_189),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_250),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_251),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_251),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_270),
.Y(n_337)
);

OR2x6_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_204),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_253),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_279),
.B(n_236),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_272),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_283),
.B(n_239),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_244),
.B(n_213),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_268),
.B(n_213),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_278),
.B(n_215),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_226),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_291),
.A2(n_282),
.B1(n_192),
.B2(n_190),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_346),
.Y(n_349)
);

AOI21x1_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_309),
.B(n_308),
.Y(n_350)
);

OAI21x1_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_259),
.B(n_257),
.Y(n_351)
);

NOR3xp33_ASAP7_75t_L g352 ( 
.A(n_291),
.B(n_286),
.C(n_188),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_302),
.B(n_262),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_314),
.A2(n_262),
.B(n_264),
.C(n_284),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_292),
.A2(n_274),
.B(n_259),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_L g357 ( 
.A1(n_312),
.A2(n_268),
.B1(n_194),
.B2(n_286),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_298),
.A2(n_274),
.B(n_260),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_303),
.A2(n_274),
.B(n_260),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_305),
.A2(n_274),
.B(n_264),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_325),
.A2(n_289),
.B(n_284),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_345),
.B(n_304),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_294),
.B(n_241),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

NOR3xp33_ASAP7_75t_L g365 ( 
.A(n_316),
.B(n_208),
.C(n_273),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_226),
.Y(n_366)
);

AO22x1_ASAP7_75t_L g367 ( 
.A1(n_293),
.A2(n_212),
.B1(n_280),
.B2(n_208),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_315),
.A2(n_289),
.B(n_273),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_329),
.A2(n_261),
.B(n_258),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_314),
.A2(n_261),
.B(n_258),
.C(n_234),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_R g371 ( 
.A(n_335),
.B(n_241),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_320),
.B(n_226),
.Y(n_372)
);

AOI22x1_ASAP7_75t_L g373 ( 
.A1(n_295),
.A2(n_234),
.B1(n_229),
.B2(n_226),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_323),
.B(n_229),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_297),
.B(n_280),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_329),
.A2(n_234),
.B(n_229),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_336),
.A2(n_234),
.B1(n_229),
.B2(n_280),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_307),
.A2(n_234),
.B(n_229),
.C(n_212),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_307),
.A2(n_212),
.B(n_280),
.C(n_10),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_326),
.A2(n_280),
.B1(n_212),
.B2(n_72),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_317),
.A2(n_280),
.B(n_212),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_311),
.B(n_8),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_342),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_331),
.A2(n_280),
.B1(n_10),
.B2(n_11),
.Y(n_384)
);

OAI22xp33_ASAP7_75t_L g385 ( 
.A1(n_319),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_311),
.B(n_301),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_340),
.A2(n_75),
.B(n_141),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_341),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_338),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_327),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_296),
.A2(n_73),
.B(n_140),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_300),
.A2(n_71),
.B(n_139),
.Y(n_393)
);

NOR3xp33_ASAP7_75t_L g394 ( 
.A(n_301),
.B(n_13),
.C(n_14),
.Y(n_394)
);

O2A1O1Ixp33_ASAP7_75t_SL g395 ( 
.A1(n_321),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_338),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_L g397 ( 
.A1(n_343),
.A2(n_16),
.B(n_18),
.C(n_19),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_321),
.B(n_19),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_306),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_330),
.A2(n_332),
.B(n_333),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_306),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_332),
.A2(n_26),
.B(n_27),
.Y(n_403)
);

NOR2x1_ASAP7_75t_L g404 ( 
.A(n_338),
.B(n_29),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_328),
.A2(n_337),
.B(n_347),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_344),
.B(n_31),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

OR2x6_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_297),
.Y(n_408)
);

OA22x2_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_297),
.B1(n_331),
.B2(n_339),
.Y(n_409)
);

NOR2xp67_ASAP7_75t_SL g410 ( 
.A(n_349),
.B(n_407),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_353),
.A2(n_327),
.B(n_334),
.Y(n_411)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_362),
.Y(n_412)
);

OAI21x1_ASAP7_75t_L g413 ( 
.A1(n_351),
.A2(n_318),
.B(n_313),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_402),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_313),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_363),
.B(n_318),
.Y(n_416)
);

AO31x2_ASAP7_75t_L g417 ( 
.A1(n_370),
.A2(n_299),
.A3(n_290),
.B(n_322),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_401),
.B(n_290),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_348),
.B(n_299),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_32),
.B(n_33),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_350),
.A2(n_35),
.B(n_36),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_349),
.B(n_41),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_43),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_366),
.B(n_44),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_381),
.A2(n_45),
.B(n_46),
.Y(n_425)
);

AO31x2_ASAP7_75t_L g426 ( 
.A1(n_398),
.A2(n_47),
.A3(n_48),
.B(n_50),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_372),
.A2(n_52),
.B(n_54),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_382),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_428)
);

OAI21x1_ASAP7_75t_SL g429 ( 
.A1(n_403),
.A2(n_59),
.B(n_60),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_374),
.B(n_61),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_364),
.B(n_63),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_406),
.B(n_64),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_381),
.A2(n_65),
.B(n_66),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_384),
.A2(n_69),
.B1(n_76),
.B2(n_79),
.Y(n_434)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_360),
.A2(n_80),
.B(n_81),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_371),
.Y(n_436)
);

BUFx12f_ASAP7_75t_L g437 ( 
.A(n_391),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_365),
.B(n_82),
.Y(n_439)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_355),
.A2(n_85),
.B(n_86),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_383),
.B(n_87),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_387),
.A2(n_88),
.B(n_90),
.C(n_91),
.Y(n_442)
);

OAI21x1_ASAP7_75t_L g443 ( 
.A1(n_358),
.A2(n_142),
.B(n_94),
.Y(n_443)
);

OR2x6_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_92),
.Y(n_444)
);

OAI21x1_ASAP7_75t_L g445 ( 
.A1(n_359),
.A2(n_95),
.B(n_96),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_352),
.B(n_97),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_368),
.A2(n_138),
.B(n_99),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_369),
.A2(n_98),
.B(n_100),
.C(n_104),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_389),
.A2(n_107),
.B(n_108),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_L g450 ( 
.A(n_407),
.B(n_110),
.Y(n_450)
);

OAI21x1_ASAP7_75t_L g451 ( 
.A1(n_389),
.A2(n_135),
.B(n_112),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_399),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_361),
.B(n_115),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_400),
.A2(n_117),
.B(n_120),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_376),
.A2(n_122),
.B(n_123),
.Y(n_455)
);

OAI22xp33_ASAP7_75t_L g456 ( 
.A1(n_412),
.A2(n_375),
.B1(n_380),
.B2(n_385),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_423),
.A2(n_394),
.B1(n_375),
.B2(n_395),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_425),
.A2(n_354),
.B(n_378),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_416),
.B(n_397),
.Y(n_460)
);

OAI222xp33_ASAP7_75t_L g461 ( 
.A1(n_434),
.A2(n_377),
.B1(n_393),
.B2(n_392),
.C1(n_367),
.C2(n_356),
.Y(n_461)
);

AOI22xp33_ASAP7_75t_L g462 ( 
.A1(n_409),
.A2(n_388),
.B1(n_373),
.B2(n_379),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_439),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_463)
);

O2A1O1Ixp33_ASAP7_75t_SL g464 ( 
.A1(n_442),
.A2(n_128),
.B(n_130),
.C(n_131),
.Y(n_464)
);

OR2x2_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_132),
.Y(n_465)
);

AO21x1_ASAP7_75t_L g466 ( 
.A1(n_432),
.A2(n_133),
.B(n_433),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_418),
.A2(n_415),
.B(n_411),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_454),
.A2(n_435),
.B(n_440),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_424),
.A2(n_430),
.B(n_453),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_421),
.A2(n_422),
.B(n_441),
.Y(n_470)
);

OA21x2_ASAP7_75t_L g471 ( 
.A1(n_420),
.A2(n_443),
.B(n_445),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_414),
.Y(n_472)
);

OAI21x1_ASAP7_75t_L g473 ( 
.A1(n_447),
.A2(n_451),
.B(n_449),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_452),
.B(n_419),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_437),
.Y(n_475)
);

AND2x2_ASAP7_75t_L g476 ( 
.A(n_408),
.B(n_439),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

BUFx4f_ASAP7_75t_SL g478 ( 
.A(n_446),
.Y(n_478)
);

OAI22xp33_ASAP7_75t_L g479 ( 
.A1(n_444),
.A2(n_428),
.B1(n_431),
.B2(n_438),
.Y(n_479)
);

AO31x2_ASAP7_75t_L g480 ( 
.A1(n_448),
.A2(n_427),
.A3(n_455),
.B(n_417),
.Y(n_480)
);

AND2x4_ASAP7_75t_SL g481 ( 
.A(n_438),
.B(n_444),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_438),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_426),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_450),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_426),
.A2(n_418),
.B(n_415),
.Y(n_485)
);

AO31x2_ASAP7_75t_L g486 ( 
.A1(n_442),
.A2(n_398),
.A3(n_370),
.B(n_378),
.Y(n_486)
);

INVx3_ASAP7_75t_SL g487 ( 
.A(n_436),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_412),
.B(n_408),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_425),
.A2(n_433),
.B(n_302),
.Y(n_489)
);

AO31x2_ASAP7_75t_L g490 ( 
.A1(n_442),
.A2(n_398),
.A3(n_370),
.B(n_378),
.Y(n_490)
);

OAI21x1_ASAP7_75t_SL g491 ( 
.A1(n_429),
.A2(n_403),
.B(n_425),
.Y(n_491)
);

OAI21x1_ASAP7_75t_L g492 ( 
.A1(n_413),
.A2(n_351),
.B(n_411),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_415),
.B(n_302),
.Y(n_493)
);

O2A1O1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_423),
.A2(n_291),
.B(n_312),
.C(n_398),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_418),
.A2(n_415),
.B(n_353),
.Y(n_495)
);

AO21x2_ASAP7_75t_L g496 ( 
.A1(n_421),
.A2(n_430),
.B(n_424),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_437),
.Y(n_497)
);

NAND2x1p5_ASAP7_75t_L g498 ( 
.A(n_410),
.B(n_438),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_472),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_474),
.Y(n_501)
);

AOI222xp33_ASAP7_75t_L g502 ( 
.A1(n_489),
.A2(n_460),
.B1(n_478),
.B2(n_476),
.C1(n_463),
.C2(n_493),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_492),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_493),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_498),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_498),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_488),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_480),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_475),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_467),
.Y(n_511)
);

AOI22xp33_ASAP7_75t_L g512 ( 
.A1(n_489),
.A2(n_466),
.B1(n_457),
.B2(n_491),
.Y(n_512)
);

BUFx2_ASAP7_75t_L g513 ( 
.A(n_482),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_488),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_457),
.B(n_481),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_465),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_467),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_462),
.B(n_486),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_456),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_480),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_486),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_479),
.A2(n_470),
.B1(n_495),
.B2(n_485),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_486),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_495),
.B(n_485),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_490),
.Y(n_526)
);

BUFx2_ASAP7_75t_L g527 ( 
.A(n_497),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_490),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_490),
.B(n_459),
.Y(n_529)
);

OAI21x1_ASAP7_75t_L g530 ( 
.A1(n_459),
.A2(n_470),
.B(n_469),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_464),
.Y(n_531)
);

AOI221xp5_ASAP7_75t_L g532 ( 
.A1(n_461),
.A2(n_487),
.B1(n_469),
.B2(n_496),
.C(n_471),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_496),
.A2(n_468),
.B(n_473),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_460),
.B(n_493),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_458),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_458),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_505),
.Y(n_537)
);

INVxp33_ASAP7_75t_SL g538 ( 
.A(n_527),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_505),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_534),
.B(n_504),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_534),
.B(n_504),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_520),
.B(n_499),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_502),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_513),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_499),
.B(n_519),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_519),
.B(n_515),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_515),
.B(n_529),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_524),
.Y(n_549)
);

OR2x2_ASAP7_75t_L g550 ( 
.A(n_511),
.B(n_517),
.Y(n_550)
);

NAND2x1p5_ASAP7_75t_L g551 ( 
.A(n_511),
.B(n_517),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_513),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_529),
.B(n_500),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_500),
.B(n_535),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_522),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_535),
.B(n_536),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_527),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_526),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_526),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_512),
.A2(n_516),
.B1(n_523),
.B2(n_514),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_518),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_528),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_528),
.B(n_525),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_509),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_506),
.B(n_507),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_506),
.B(n_507),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_509),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_510),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_508),
.B(n_531),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_521),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_521),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_530),
.B(n_532),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_530),
.B(n_503),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_533),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_541),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_571),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_541),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_549),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_549),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_558),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_544),
.B(n_542),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_548),
.B(n_547),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_548),
.B(n_547),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_544),
.B(n_542),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_558),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_545),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_553),
.B(n_546),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_553),
.B(n_546),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_559),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_571),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_540),
.B(n_543),
.Y(n_592)
);

INVxp67_ASAP7_75t_SL g593 ( 
.A(n_563),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_545),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_540),
.B(n_554),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_543),
.B(n_560),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_557),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_559),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_556),
.B(n_554),
.Y(n_599)
);

HB1xp67_ASAP7_75t_L g600 ( 
.A(n_557),
.Y(n_600)
);

OR2x2_ASAP7_75t_L g601 ( 
.A(n_562),
.B(n_555),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_557),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_564),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_562),
.B(n_555),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_561),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_564),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_556),
.B(n_572),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_572),
.B(n_550),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_607),
.B(n_551),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_607),
.B(n_551),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_608),
.B(n_551),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_608),
.B(n_573),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_581),
.B(n_550),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_575),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_577),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_585),
.B(n_593),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_588),
.B(n_567),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_595),
.B(n_561),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_601),
.B(n_573),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_595),
.B(n_561),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_582),
.B(n_538),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_577),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_605),
.B(n_568),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_578),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_588),
.B(n_567),
.Y(n_626)
);

OR2x2_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_574),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_578),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_587),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_592),
.B(n_568),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_589),
.B(n_571),
.Y(n_631)
);

OR2x2_ASAP7_75t_L g632 ( 
.A(n_604),
.B(n_574),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_579),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_589),
.B(n_570),
.Y(n_634)
);

BUFx2_ASAP7_75t_SL g635 ( 
.A(n_605),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_597),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_583),
.B(n_570),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_579),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_580),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_639),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_612),
.B(n_604),
.Y(n_641)
);

NOR2x1_ASAP7_75t_L g642 ( 
.A(n_617),
.B(n_568),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_636),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_614),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_639),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_619),
.Y(n_646)
);

NAND2x1_ASAP7_75t_L g647 ( 
.A(n_614),
.B(n_591),
.Y(n_647)
);

OR2x2_ASAP7_75t_L g648 ( 
.A(n_612),
.B(n_620),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_613),
.B(n_594),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_609),
.B(n_584),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_629),
.B(n_584),
.Y(n_651)
);

NOR2x1_ASAP7_75t_L g652 ( 
.A(n_635),
.B(n_569),
.Y(n_652)
);

NAND3xp33_ASAP7_75t_L g653 ( 
.A(n_624),
.B(n_596),
.C(n_602),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_609),
.B(n_583),
.Y(n_654)
);

AOI222xp33_ASAP7_75t_L g655 ( 
.A1(n_630),
.A2(n_599),
.B1(n_566),
.B2(n_565),
.C1(n_598),
.C2(n_590),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_627),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_633),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_633),
.Y(n_658)
);

NAND2x1_ASAP7_75t_SL g659 ( 
.A(n_611),
.B(n_600),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_615),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_616),
.Y(n_661)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_648),
.B(n_620),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_644),
.Y(n_663)
);

INVxp67_ASAP7_75t_L g664 ( 
.A(n_642),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_640),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_656),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_645),
.Y(n_667)
);

AOI222xp33_ASAP7_75t_L g668 ( 
.A1(n_653),
.A2(n_622),
.B1(n_621),
.B2(n_618),
.C1(n_626),
.C2(n_611),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_660),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_652),
.B(n_610),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_661),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_656),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_644),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_668),
.B(n_646),
.Y(n_674)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_670),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_664),
.B(n_643),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_662),
.B(n_654),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_664),
.B(n_654),
.Y(n_678)
);

AOI221xp5_ASAP7_75t_L g679 ( 
.A1(n_672),
.A2(n_651),
.B1(n_649),
.B2(n_650),
.C(n_610),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_675),
.B(n_655),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_678),
.Y(n_681)
);

OAI21xp5_ASAP7_75t_L g682 ( 
.A1(n_674),
.A2(n_671),
.B(n_669),
.Y(n_682)
);

OAI21xp5_ASAP7_75t_SL g683 ( 
.A1(n_676),
.A2(n_666),
.B(n_631),
.Y(n_683)
);

AOI221xp5_ASAP7_75t_L g684 ( 
.A1(n_679),
.A2(n_667),
.B1(n_665),
.B2(n_666),
.C(n_673),
.Y(n_684)
);

OAI32xp33_ASAP7_75t_L g685 ( 
.A1(n_677),
.A2(n_641),
.A3(n_663),
.B1(n_627),
.B2(n_632),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_681),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_680),
.Y(n_687)
);

OAI21xp33_ASAP7_75t_L g688 ( 
.A1(n_682),
.A2(n_684),
.B(n_683),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_685),
.B(n_650),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_682),
.B(n_641),
.Y(n_690)
);

OAI211xp5_ASAP7_75t_L g691 ( 
.A1(n_688),
.A2(n_659),
.B(n_647),
.C(n_623),
.Y(n_691)
);

AND3x1_ASAP7_75t_L g692 ( 
.A(n_687),
.B(n_631),
.C(n_618),
.Y(n_692)
);

CKINVDCx20_ASAP7_75t_R g693 ( 
.A(n_691),
.Y(n_693)
);

NOR2x1_ASAP7_75t_L g694 ( 
.A(n_692),
.B(n_686),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_692),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_694),
.B(n_690),
.Y(n_696)
);

AND3x4_ASAP7_75t_L g697 ( 
.A(n_693),
.B(n_695),
.C(n_689),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_693),
.B(n_658),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_693),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_695),
.B(n_637),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_695),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_697),
.A2(n_696),
.B1(n_699),
.B2(n_701),
.Y(n_702)
);

AOI211xp5_ASAP7_75t_L g703 ( 
.A1(n_696),
.A2(n_698),
.B(n_700),
.C(n_566),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_699),
.Y(n_704)
);

NAND4xp25_ASAP7_75t_L g705 ( 
.A(n_699),
.B(n_565),
.C(n_632),
.D(n_638),
.Y(n_705)
);

NAND3xp33_ASAP7_75t_L g706 ( 
.A(n_701),
.B(n_628),
.C(n_625),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_SL g707 ( 
.A(n_696),
.B(n_658),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_704),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_702),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_707),
.A2(n_635),
.B1(n_576),
.B2(n_591),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_709),
.A2(n_703),
.B1(n_705),
.B2(n_657),
.Y(n_712)
);

AOI32xp33_ASAP7_75t_L g713 ( 
.A1(n_708),
.A2(n_626),
.A3(n_637),
.B1(n_657),
.B2(n_634),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_711),
.B(n_634),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_714),
.A2(n_710),
.B(n_539),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_712),
.A2(n_537),
.B(n_539),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_L g717 ( 
.A1(n_713),
.A2(n_537),
.B(n_598),
.Y(n_717)
);

AO21x2_ASAP7_75t_L g718 ( 
.A1(n_716),
.A2(n_580),
.B(n_590),
.Y(n_718)
);

AOI22xp5_ASAP7_75t_L g719 ( 
.A1(n_715),
.A2(n_586),
.B1(n_576),
.B2(n_591),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_719),
.A2(n_717),
.B(n_586),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_720),
.B(n_718),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_721),
.A2(n_576),
.B1(n_603),
.B2(n_606),
.Y(n_722)
);


endmodule