module fake_jpeg_18403_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx5_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx6_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OR2x2_ASAP7_75t_SL g27 ( 
.A(n_17),
.B(n_19),
.Y(n_27)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_20),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_26),
.B(n_17),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_32),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_17),
.C(n_23),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_27),
.B1(n_18),
.B2(n_28),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

NOR2xp67_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_25),
.Y(n_39)
);

MAJx2_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_34),
.C(n_35),
.Y(n_38)
);

A2O1A1O1Ixp25_ASAP7_75t_L g40 ( 
.A1(n_38),
.A2(n_39),
.B(n_35),
.C(n_34),
.D(n_17),
.Y(n_40)
);

AOI322xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.A3(n_8),
.B1(n_12),
.B2(n_15),
.C1(n_28),
.C2(n_21),
.Y(n_42)
);

AOI322xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_18),
.A3(n_23),
.B1(n_14),
.B2(n_15),
.C1(n_10),
.C2(n_22),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_16),
.B(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_43),
.Y(n_44)
);


endmodule