module fake_jpeg_26343_n_172 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_0),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

BUFx2_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_18),
.B1(n_26),
.B2(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_41),
.B1(n_48),
.B2(n_33),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_41)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_24),
.Y(n_45)
);

OR2x4_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_28),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_32),
.A2(n_25),
.B1(n_23),
.B2(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_37),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_52),
.A2(n_64),
.B(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_46),
.A2(n_32),
.B1(n_29),
.B2(n_37),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_56),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_49),
.B(n_15),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_55),
.B(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_33),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_34),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_34),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_19),
.B1(n_28),
.B2(n_15),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_29),
.B1(n_37),
.B2(n_14),
.Y(n_64)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_68),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_33),
.B(n_34),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_70),
.B(n_47),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_77),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_38),
.C(n_40),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_73),
.B(n_59),
.C(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_44),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_0),
.Y(n_87)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_88),
.A2(n_67),
.B1(n_40),
.B2(n_71),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_20),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_91),
.A2(n_66),
.B(n_58),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_103),
.B1(n_97),
.B2(n_95),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_106),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_102),
.B(n_103),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_99),
.Y(n_115)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_91),
.C(n_92),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_27),
.Y(n_101)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

AND2x6_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_12),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_20),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_62),
.A3(n_59),
.B1(n_65),
.B2(n_68),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_105),
.B(n_75),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_27),
.B(n_16),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_1),
.Y(n_108)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_2),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_109),
.B(n_110),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_2),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_120),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_116),
.B(n_118),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_90),
.B(n_84),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_100),
.B(n_73),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_122),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_72),
.B(n_81),
.C(n_87),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_99),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_76),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_123),
.A2(n_91),
.B1(n_102),
.B2(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_81),
.C(n_74),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_108),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_128),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_93),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_124),
.B(n_103),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_130),
.A2(n_118),
.B(n_125),
.C(n_111),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_93),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_136),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_112),
.B1(n_114),
.B2(n_121),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_76),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_120),
.B1(n_129),
.B2(n_78),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_145),
.B(n_146),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_116),
.B(n_130),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_149),
.A2(n_144),
.B1(n_140),
.B2(n_142),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g150 ( 
.A(n_141),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_89),
.C(n_74),
.Y(n_158)
);

NOR3xp33_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_134),
.C(n_136),
.Y(n_151)
);

AOI31xp67_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_154),
.A3(n_131),
.B(n_147),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_82),
.B(n_78),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_118),
.B(n_133),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_153),
.A2(n_147),
.B(n_131),
.Y(n_156)
);

AOI31xp67_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_118),
.A3(n_128),
.B(n_111),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_155),
.B(n_158),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_160),
.C(n_3),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_89),
.C(n_85),
.Y(n_160)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_13),
.A3(n_12),
.B1(n_83),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_162)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_162),
.A2(n_3),
.B(n_6),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_161),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_167),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_163),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_166),
.B(n_9),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_168),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_9),
.Y(n_172)
);


endmodule