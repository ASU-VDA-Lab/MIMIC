module fake_netlist_5_2563_n_1696 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1696);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1696;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_368;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_33),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_15),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_44),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_53),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_58),
.Y(n_165)
);

INVx2_ASAP7_75t_SL g166 ( 
.A(n_45),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_51),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_81),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_37),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_111),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_89),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_25),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_103),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_73),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_70),
.Y(n_178)
);

BUFx8_ASAP7_75t_SL g179 ( 
.A(n_40),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_27),
.Y(n_180)
);

INVxp67_ASAP7_75t_SL g181 ( 
.A(n_85),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_97),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_12),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_158),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_50),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_87),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_139),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_55),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_55),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_155),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_9),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_3),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_156),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_24),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_18),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_122),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_52),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_13),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_82),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_45),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_147),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_78),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_90),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_84),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_19),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_50),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_52),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_53),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_40),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_76),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_31),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_115),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_18),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_66),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_15),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_12),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_77),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_47),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_37),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_68),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_2),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_127),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_23),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_28),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_99),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_56),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_9),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_48),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_116),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_159),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_74),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_137),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_69),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_121),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_10),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_10),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_119),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_32),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_136),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_107),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_148),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_49),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_22),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_109),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_6),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_28),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_130),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_17),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_32),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_16),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_31),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_6),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_48),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_106),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_8),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_95),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_113),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_123),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_91),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_36),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_128),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_33),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_47),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_36),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_98),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_140),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_13),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_64),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_86),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_23),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_135),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_65),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_1),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_1),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_112),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_96),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_27),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g290 ( 
.A(n_146),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_54),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_63),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_92),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_54),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_42),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_42),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_154),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_94),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_59),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_80),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_35),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_3),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_24),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_61),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_16),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_14),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_120),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_117),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_79),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_104),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_72),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_41),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_101),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_129),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_14),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_44),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_151),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_75),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_22),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_179),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_163),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_163),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_164),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_164),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_168),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_168),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_184),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_170),
.Y(n_329)
);

BUFx2_ASAP7_75t_SL g330 ( 
.A(n_204),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_167),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_170),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_206),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_221),
.B(n_0),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_175),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_289),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_169),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_175),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_162),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_206),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_171),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_172),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_190),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_276),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_190),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_176),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_177),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_178),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_194),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_182),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_194),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_197),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_185),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_197),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_205),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_205),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_230),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_187),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_276),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_233),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_267),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_188),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_213),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_213),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_214),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_193),
.Y(n_366)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_294),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_196),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_268),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_214),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_201),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_227),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_172),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_265),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_227),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_172),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_199),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_209),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_210),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_311),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_180),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_165),
.B(n_0),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_219),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_229),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_229),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_236),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_311),
.B(n_2),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_220),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_222),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_290),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_236),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_225),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_237),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_186),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_234),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_323),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_373),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_373),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_340),
.B(n_311),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_344),
.B(n_238),
.Y(n_404)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_326),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_359),
.B(n_202),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_326),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_242),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_334),
.B(n_189),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_339),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_367),
.B(n_224),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_336),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_243),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_327),
.Y(n_418)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_330),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_165),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_367),
.B(n_186),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_333),
.B(n_244),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_333),
.B(n_202),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_378),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_342),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_377),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_377),
.B(n_173),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_333),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_343),
.B(n_250),
.Y(n_432)
);

OA21x2_ASAP7_75t_L g433 ( 
.A1(n_321),
.A2(n_255),
.B(n_237),
.Y(n_433)
);

AND2x4_ASAP7_75t_L g434 ( 
.A(n_343),
.B(n_173),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_351),
.B(n_174),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_321),
.Y(n_436)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_351),
.B(n_174),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_355),
.B(n_183),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_355),
.B(n_251),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_329),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_322),
.B(n_183),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_322),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_332),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_378),
.A2(n_231),
.B1(n_261),
.B2(n_278),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_328),
.B(n_228),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_324),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_332),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_335),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_335),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_338),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_338),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_345),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_345),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_349),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_324),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_383),
.B(n_254),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_352),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_352),
.B(n_172),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_354),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_354),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_356),
.Y(n_463)
);

CKINVDCx6p67_ASAP7_75t_R g464 ( 
.A(n_374),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_356),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_363),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_363),
.B(n_200),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_403),
.B(n_395),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_424),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_424),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_425),
.B(n_331),
.Y(n_471)
);

BUFx8_ASAP7_75t_SL g472 ( 
.A(n_431),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_425),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_433),
.Y(n_474)
);

BUFx3_ASAP7_75t_L g475 ( 
.A(n_431),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_413),
.B(n_337),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_455),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_433),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_455),
.Y(n_480)
);

BUFx3_ASAP7_75t_L g481 ( 
.A(n_431),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_413),
.B(n_341),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_396),
.B(n_346),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_455),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_433),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_424),
.Y(n_487)
);

AOI22xp33_ASAP7_75t_L g488 ( 
.A1(n_434),
.A2(n_166),
.B1(n_319),
.B2(n_255),
.Y(n_488)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_414),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_408),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_419),
.B(n_347),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_455),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_433),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_434),
.A2(n_166),
.B1(n_319),
.B2(n_263),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_433),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_455),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_455),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_447),
.B(n_391),
.Y(n_499)
);

INVx4_ASAP7_75t_L g500 ( 
.A(n_455),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_420),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

AND3x2_ASAP7_75t_L g503 ( 
.A(n_414),
.B(n_266),
.C(n_293),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_403),
.B(n_364),
.Y(n_504)
);

BUFx2_ASAP7_75t_L g505 ( 
.A(n_416),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_412),
.B(n_348),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_408),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_464),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

AND2x6_ASAP7_75t_L g510 ( 
.A(n_403),
.B(n_172),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_434),
.B(n_330),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_408),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_412),
.B(n_350),
.Y(n_513)
);

INVx2_ASAP7_75t_SL g514 ( 
.A(n_423),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_434),
.B(n_435),
.Y(n_515)
);

NAND2xp33_ASAP7_75t_SL g516 ( 
.A(n_447),
.B(n_306),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_456),
.Y(n_517)
);

BUFx2_ASAP7_75t_L g518 ( 
.A(n_416),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_419),
.B(n_353),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_464),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_434),
.B(n_364),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_456),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_446),
.B(n_358),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_406),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_396),
.B(n_362),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g526 ( 
.A(n_446),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_417),
.B(n_366),
.Y(n_527)
);

OR2x2_ASAP7_75t_L g528 ( 
.A(n_457),
.B(n_382),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_457),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_464),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_432),
.B(n_368),
.Y(n_531)
);

AO22x2_ASAP7_75t_L g532 ( 
.A1(n_435),
.A2(n_263),
.B1(n_286),
.B2(n_315),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_420),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_435),
.B(n_365),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_458),
.B(n_371),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_420),
.Y(n_536)
);

INVx4_ASAP7_75t_SL g537 ( 
.A(n_460),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_420),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_432),
.B(n_376),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_458),
.B(n_379),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_440),
.B(n_380),
.Y(n_541)
);

BUFx8_ASAP7_75t_SL g542 ( 
.A(n_440),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_437),
.B(n_365),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_417),
.B(n_384),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_456),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_404),
.B(n_389),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_456),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_428),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_456),
.Y(n_549)
);

AND2x6_ASAP7_75t_L g550 ( 
.A(n_437),
.B(n_235),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_445),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_404),
.B(n_390),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_L g553 ( 
.A(n_423),
.B(n_393),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_428),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_415),
.B(n_382),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_437),
.B(n_211),
.C(n_200),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_406),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_456),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_456),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_438),
.B(n_271),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_428),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_438),
.B(n_451),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_438),
.B(n_370),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_415),
.B(n_320),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_442),
.B(n_370),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_421),
.B(n_357),
.Y(n_566)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_406),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g568 ( 
.A(n_445),
.Y(n_568)
);

BUFx8_ASAP7_75t_SL g569 ( 
.A(n_467),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_428),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_467),
.B(n_235),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_442),
.B(n_372),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_451),
.B(n_428),
.Y(n_573)
);

BUFx10_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_452),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_406),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_452),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_452),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_451),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

AND2x6_ASAP7_75t_L g581 ( 
.A(n_467),
.B(n_235),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_451),
.B(n_207),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_421),
.B(n_360),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_467),
.B(n_270),
.Y(n_584)
);

AO21x2_ASAP7_75t_L g585 ( 
.A1(n_442),
.A2(n_258),
.B(n_256),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_406),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_406),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g588 ( 
.A1(n_397),
.A2(n_369),
.B1(n_361),
.B2(n_195),
.Y(n_588)
);

OAI22xp33_ASAP7_75t_L g589 ( 
.A1(n_397),
.A2(n_305),
.B1(n_253),
.B2(n_316),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_398),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_400),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_460),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_400),
.A2(n_260),
.B1(n_259),
.B2(n_257),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_402),
.B(n_240),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_402),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_407),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_466),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_410),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_407),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_460),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_409),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_409),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_418),
.B(n_372),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_410),
.Y(n_605)
);

INVxp33_ASAP7_75t_L g606 ( 
.A(n_418),
.Y(n_606)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_429),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_466),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_429),
.B(n_375),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_405),
.B(n_241),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_439),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_405),
.B(n_299),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_405),
.B(n_272),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_439),
.B(n_161),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_410),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_466),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_603),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_603),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_514),
.B(n_466),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_515),
.B(n_490),
.Y(n_620)
);

BUFx5_ASAP7_75t_L g621 ( 
.A(n_474),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_535),
.A2(n_181),
.B1(n_307),
.B2(n_277),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_473),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_609),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_575),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_540),
.B(n_466),
.Y(n_626)
);

OAI22xp33_ASAP7_75t_L g627 ( 
.A1(n_560),
.A2(n_279),
.B1(n_269),
.B2(n_283),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_526),
.B(n_191),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_484),
.B(n_525),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_515),
.A2(n_286),
.B(n_295),
.C(n_302),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_609),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_490),
.B(n_235),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_546),
.B(n_466),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_596),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_577),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_577),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_599),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_578),
.Y(n_639)
);

BUFx4f_ASAP7_75t_L g640 ( 
.A(n_511),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_599),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_552),
.B(n_192),
.Y(n_642)
);

NOR2xp67_ASAP7_75t_SL g643 ( 
.A(n_592),
.B(n_600),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_507),
.B(n_235),
.Y(n_644)
);

INVx8_ASAP7_75t_L g645 ( 
.A(n_511),
.Y(n_645)
);

INVxp33_ASAP7_75t_SL g646 ( 
.A(n_473),
.Y(n_646)
);

AND3x1_ASAP7_75t_L g647 ( 
.A(n_560),
.B(n_302),
.C(n_295),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_534),
.B(n_441),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_507),
.B(n_436),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_512),
.B(n_318),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_578),
.Y(n_651)
);

AO221x1_ASAP7_75t_L g652 ( 
.A1(n_532),
.A2(n_318),
.B1(n_312),
.B2(n_315),
.C(n_258),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_512),
.B(n_436),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_591),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_474),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_521),
.B(n_602),
.Y(n_656)
);

O2A1O1Ixp33_ASAP7_75t_L g657 ( 
.A1(n_562),
.A2(n_453),
.B(n_441),
.C(n_444),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_574),
.B(n_318),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_521),
.B(n_436),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_468),
.A2(n_297),
.B1(n_280),
.B2(n_282),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_602),
.B(n_436),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_469),
.B(n_436),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_607),
.B(n_444),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_469),
.A2(n_211),
.B1(n_217),
.B2(n_239),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_574),
.B(n_318),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_470),
.B(n_448),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_470),
.B(n_448),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_506),
.B(n_198),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_479),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_468),
.A2(n_308),
.B1(n_287),
.B2(n_288),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_487),
.B(n_448),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_487),
.B(n_448),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_504),
.B(n_459),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_504),
.B(n_459),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_607),
.B(n_459),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_534),
.B(n_459),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_479),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_574),
.B(n_318),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_543),
.B(n_461),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_574),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_543),
.B(n_461),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_563),
.B(n_461),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_573),
.B(n_292),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_563),
.B(n_461),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_553),
.A2(n_309),
.B1(n_298),
.B2(n_300),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_565),
.B(n_449),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_513),
.B(n_462),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_475),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_527),
.B(n_462),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_505),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_544),
.B(n_462),
.Y(n_691)
);

AOI22xp5_ASAP7_75t_L g692 ( 
.A1(n_531),
.A2(n_304),
.B1(n_310),
.B2(n_314),
.Y(n_692)
);

BUFx6f_ASAP7_75t_SL g693 ( 
.A(n_529),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_483),
.B(n_217),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_582),
.B(n_462),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_565),
.B(n_463),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_570),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_483),
.B(n_239),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_585),
.A2(n_313),
.B1(n_247),
.B2(n_317),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_475),
.Y(n_700)
);

O2A1O1Ixp33_ASAP7_75t_L g701 ( 
.A1(n_486),
.A2(n_495),
.B(n_493),
.C(n_590),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_572),
.B(n_463),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_486),
.B(n_247),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_595),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_493),
.B(n_249),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_572),
.B(n_463),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_530),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_595),
.B(n_601),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_495),
.B(n_249),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_601),
.B(n_463),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_501),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_611),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_611),
.B(n_465),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_570),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_501),
.B(n_465),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_502),
.B(n_256),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_530),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_505),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_533),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_533),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_536),
.B(n_538),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_481),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_536),
.B(n_465),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_538),
.B(n_269),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_548),
.B(n_465),
.Y(n_725)
);

AO221x1_ASAP7_75t_L g726 ( 
.A1(n_532),
.A2(n_312),
.B1(n_279),
.B2(n_283),
.C(n_285),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_471),
.B(n_203),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_548),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_554),
.B(n_405),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_523),
.B(n_212),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_554),
.B(n_405),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_476),
.B(n_215),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_561),
.B(n_579),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_518),
.B(n_449),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_579),
.B(n_313),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_481),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_529),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_580),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_482),
.B(n_216),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_580),
.B(n_317),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_606),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_594),
.B(n_450),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_528),
.B(n_450),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_529),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_529),
.B(n_453),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_550),
.B(n_454),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_511),
.A2(n_454),
.B1(n_296),
.B2(n_301),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_550),
.B(n_399),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_610),
.B(n_410),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_585),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_550),
.B(n_399),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_539),
.B(n_218),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_585),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_550),
.B(n_399),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_541),
.B(n_223),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_550),
.B(n_399),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_511),
.A2(n_262),
.B1(n_252),
.B2(n_248),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_556),
.A2(n_460),
.B1(n_443),
.B2(n_186),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_489),
.B(n_186),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_489),
.B(n_195),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_532),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_550),
.B(n_411),
.Y(n_762)
);

OAI221xp5_ASAP7_75t_L g763 ( 
.A1(n_488),
.A2(n_394),
.B1(n_392),
.B2(n_387),
.C(n_386),
.Y(n_763)
);

NOR3xp33_ASAP7_75t_L g764 ( 
.A(n_499),
.B(n_226),
.C(n_303),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_550),
.B(n_411),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_612),
.B(n_411),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_477),
.B(n_410),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_478),
.Y(n_768)
);

NOR2x1p5_ASAP7_75t_L g769 ( 
.A(n_555),
.B(n_528),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_532),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_510),
.B(n_411),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_478),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_491),
.B(n_232),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_510),
.B(n_443),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_510),
.B(n_443),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_510),
.B(n_443),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_480),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_510),
.B(n_430),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_711),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_629),
.B(n_614),
.Y(n_780)
);

A2O1A1Ixp33_ASAP7_75t_L g781 ( 
.A1(n_642),
.A2(n_583),
.B(n_566),
.C(n_556),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_633),
.A2(n_557),
.B(n_613),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_675),
.B(n_511),
.Y(n_783)
);

BUFx8_ASAP7_75t_L g784 ( 
.A(n_693),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_626),
.A2(n_500),
.B(n_547),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_621),
.B(n_510),
.Y(n_786)
);

CKINVDCx10_ASAP7_75t_R g787 ( 
.A(n_693),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_656),
.B(n_519),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_687),
.A2(n_500),
.B(n_547),
.Y(n_789)
);

A2O1A1Ixp33_ASAP7_75t_L g790 ( 
.A1(n_668),
.A2(n_564),
.B(n_568),
.C(n_551),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_663),
.B(n_494),
.Y(n_791)
);

O2A1O1Ixp5_ASAP7_75t_L g792 ( 
.A1(n_694),
.A2(n_584),
.B(n_480),
.C(n_608),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_742),
.B(n_496),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_689),
.A2(n_547),
.B(n_500),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_691),
.A2(n_695),
.B(n_749),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_700),
.B(n_588),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_623),
.B(n_551),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_736),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_688),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_645),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_749),
.A2(n_547),
.B(n_500),
.Y(n_801)
);

A2O1A1Ixp33_ASAP7_75t_L g802 ( 
.A1(n_732),
.A2(n_555),
.B(n_516),
.C(n_608),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_707),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_766),
.A2(n_567),
.B(n_615),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_646),
.B(n_542),
.Y(n_805)
);

NAND2x1p5_ASAP7_75t_L g806 ( 
.A(n_680),
.B(n_592),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_648),
.B(n_496),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_640),
.A2(n_753),
.B1(n_750),
.B2(n_655),
.Y(n_808)
);

AOI21x1_ASAP7_75t_L g809 ( 
.A1(n_767),
.A2(n_616),
.B(n_492),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_648),
.B(n_496),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_619),
.A2(n_731),
.B(n_729),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_673),
.A2(n_567),
.B(n_615),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_719),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_700),
.B(n_589),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_674),
.A2(n_567),
.B(n_605),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_SL g816 ( 
.A1(n_646),
.A2(n_508),
.B1(n_520),
.B2(n_245),
.Y(n_816)
);

HB1xp67_ASAP7_75t_L g817 ( 
.A(n_722),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_SL g818 ( 
.A1(n_694),
.A2(n_703),
.B(n_705),
.C(n_698),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_676),
.A2(n_567),
.B(n_605),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_679),
.A2(n_524),
.B(n_605),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_690),
.B(n_472),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_686),
.B(n_509),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_681),
.A2(n_509),
.B(n_524),
.Y(n_823)
);

AO21x1_ASAP7_75t_L g824 ( 
.A1(n_698),
.A2(n_616),
.B(n_604),
.Y(n_824)
);

INVxp67_ASAP7_75t_L g825 ( 
.A(n_734),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_741),
.B(n_593),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_682),
.A2(n_509),
.B(n_524),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_718),
.B(n_569),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_728),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_736),
.B(n_503),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_686),
.B(n_621),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_L g832 ( 
.A(n_628),
.B(n_246),
.C(n_264),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_621),
.B(n_576),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_621),
.B(n_576),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_730),
.B(n_576),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_761),
.Y(n_836)
);

NOR3xp33_ASAP7_75t_L g837 ( 
.A(n_739),
.B(n_273),
.C(n_274),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_684),
.A2(n_586),
.B(n_587),
.Y(n_838)
);

BUFx4f_ASAP7_75t_L g839 ( 
.A(n_770),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_659),
.A2(n_586),
.B(n_587),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_621),
.B(n_586),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_195),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_625),
.Y(n_843)
);

AO21x1_ASAP7_75t_L g844 ( 
.A1(n_703),
.A2(n_604),
.B(n_597),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_620),
.A2(n_571),
.B1(n_581),
.B2(n_597),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_752),
.A2(n_485),
.B(n_492),
.C(n_497),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_743),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_737),
.B(n_592),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_645),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_621),
.B(n_620),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_696),
.A2(n_587),
.B(n_598),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_625),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_755),
.A2(n_517),
.B(n_498),
.C(n_497),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_702),
.A2(n_598),
.B(n_545),
.Y(n_854)
);

OR2x2_ASAP7_75t_L g855 ( 
.A(n_769),
.B(n_759),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_621),
.B(n_598),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_737),
.B(n_592),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_634),
.B(n_275),
.Y(n_858)
);

INVx5_ASAP7_75t_L g859 ( 
.A(n_680),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_654),
.B(n_522),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_635),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_704),
.B(n_545),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_706),
.A2(n_559),
.B(n_549),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_712),
.B(n_708),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_655),
.B(n_669),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_669),
.B(n_677),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_635),
.Y(n_867)
);

BUFx8_ASAP7_75t_SL g868 ( 
.A(n_707),
.Y(n_868)
);

OAI321xp33_ASAP7_75t_L g869 ( 
.A1(n_627),
.A2(n_727),
.A3(n_664),
.B1(n_773),
.B2(n_757),
.C(n_747),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_662),
.A2(n_721),
.B(n_653),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_R g871 ( 
.A(n_717),
.B(n_281),
.Y(n_871)
);

OAI321xp33_ASAP7_75t_L g872 ( 
.A1(n_699),
.A2(n_387),
.A3(n_394),
.B1(n_392),
.B2(n_375),
.C(n_385),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_677),
.B(n_558),
.Y(n_873)
);

AOI21x1_ASAP7_75t_L g874 ( 
.A1(n_767),
.A2(n_549),
.B(n_559),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_637),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_617),
.B(n_581),
.Y(n_876)
);

OAI21xp5_ASAP7_75t_L g877 ( 
.A1(n_701),
.A2(n_581),
.B(n_571),
.Y(n_877)
);

INVxp67_ASAP7_75t_L g878 ( 
.A(n_647),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_649),
.A2(n_600),
.B(n_592),
.Y(n_879)
);

O2A1O1Ixp33_ASAP7_75t_SL g880 ( 
.A1(n_705),
.A2(n_422),
.B(n_385),
.C(n_386),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_760),
.B(n_284),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_618),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_636),
.B(n_537),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_744),
.B(n_600),
.Y(n_884)
);

HB1xp67_ASAP7_75t_L g885 ( 
.A(n_624),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_709),
.A2(n_581),
.B(n_571),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_631),
.B(n_720),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_744),
.B(n_291),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_714),
.A2(n_683),
.B1(n_697),
.B2(n_638),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_666),
.A2(n_672),
.B(n_667),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_709),
.A2(n_581),
.B(n_571),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_671),
.A2(n_600),
.B(n_592),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_733),
.A2(n_571),
.B(n_600),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_680),
.B(n_640),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_639),
.B(n_571),
.Y(n_895)
);

BUFx2_ASAP7_75t_SL g896 ( 
.A(n_693),
.Y(n_896)
);

AOI21xp33_ASAP7_75t_L g897 ( 
.A1(n_622),
.A2(n_4),
.B(n_5),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_733),
.A2(n_571),
.B(n_427),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_683),
.A2(n_460),
.B1(n_422),
.B2(n_537),
.Y(n_899)
);

CKINVDCx8_ASAP7_75t_R g900 ( 
.A(n_717),
.Y(n_900)
);

CKINVDCx8_ASAP7_75t_R g901 ( 
.A(n_645),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_639),
.B(n_427),
.Y(n_902)
);

NAND3xp33_ASAP7_75t_L g903 ( 
.A(n_660),
.B(n_430),
.C(n_426),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_658),
.A2(n_401),
.B(n_410),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_665),
.A2(n_401),
.B(n_410),
.Y(n_905)
);

NOR2xp67_ASAP7_75t_L g906 ( 
.A(n_692),
.B(n_670),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_651),
.B(n_427),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_651),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_641),
.B(n_685),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_738),
.B(n_427),
.Y(n_910)
);

AOI21xp33_ASAP7_75t_L g911 ( 
.A1(n_657),
.A2(n_4),
.B(n_5),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_665),
.A2(n_401),
.B(n_410),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_661),
.B(n_426),
.Y(n_913)
);

CKINVDCx10_ASAP7_75t_R g914 ( 
.A(n_764),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_678),
.A2(n_401),
.B(n_430),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_716),
.B(n_7),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_715),
.A2(n_401),
.B(n_430),
.Y(n_917)
);

OAI21xp33_ASAP7_75t_L g918 ( 
.A1(n_630),
.A2(n_195),
.B(n_430),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_723),
.A2(n_401),
.B(n_430),
.Y(n_919)
);

AOI22xp33_ASAP7_75t_L g920 ( 
.A1(n_726),
.A2(n_652),
.B1(n_724),
.B2(n_716),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_725),
.A2(n_401),
.B(n_430),
.Y(n_921)
);

NOR2x1_ASAP7_75t_R g922 ( 
.A(n_724),
.B(n_8),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_645),
.A2(n_537),
.B1(n_71),
.B2(n_83),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_778),
.A2(n_460),
.B(n_62),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_746),
.B(n_67),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_632),
.B(n_460),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_768),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_632),
.B(n_11),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_644),
.B(n_11),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_768),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_777),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_644),
.B(n_460),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_777),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_650),
.B(n_460),
.Y(n_934)
);

OR2x2_ASAP7_75t_L g935 ( 
.A(n_740),
.B(n_630),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_771),
.A2(n_460),
.B(n_93),
.Y(n_936)
);

NOR2x1p5_ASAP7_75t_L g937 ( 
.A(n_772),
.B(n_17),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_710),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_650),
.B(n_20),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_713),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_748),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_735),
.A2(n_20),
.B(n_21),
.C(n_26),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_751),
.A2(n_102),
.B(n_157),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_735),
.B(n_21),
.Y(n_944)
);

INVx5_ASAP7_75t_L g945 ( 
.A(n_643),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_774),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_775),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_758),
.B(n_26),
.Y(n_948)
);

NOR3xp33_ASAP7_75t_L g949 ( 
.A(n_763),
.B(n_29),
.C(n_30),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_868),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_798),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_883),
.Y(n_952)
);

O2A1O1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_781),
.A2(n_776),
.B(n_765),
.C(n_762),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_818),
.A2(n_756),
.B(n_754),
.Y(n_954)
);

AO22x2_ASAP7_75t_L g955 ( 
.A1(n_949),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_955)
);

INVx3_ASAP7_75t_L g956 ( 
.A(n_883),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_780),
.A2(n_34),
.B(n_35),
.C(n_38),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_786),
.A2(n_114),
.B(n_153),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_831),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_837),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_837),
.A2(n_118),
.B1(n_150),
.B2(n_149),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_790),
.B(n_43),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_800),
.Y(n_963)
);

AOI21x1_ASAP7_75t_L g964 ( 
.A1(n_783),
.A2(n_108),
.B(n_145),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_825),
.B(n_46),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_842),
.B(n_49),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_897),
.A2(n_51),
.B(n_57),
.C(n_60),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_825),
.B(n_105),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_869),
.A2(n_131),
.B(n_132),
.C(n_142),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_782),
.A2(n_144),
.B(n_160),
.Y(n_970)
);

OAI21xp33_ASAP7_75t_L g971 ( 
.A1(n_881),
.A2(n_858),
.B(n_797),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_800),
.B(n_849),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_938),
.B(n_940),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_864),
.B(n_807),
.Y(n_974)
);

OAI22xp5_ASAP7_75t_L g975 ( 
.A1(n_791),
.A2(n_839),
.B1(n_878),
.B2(n_866),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_799),
.Y(n_976)
);

A2O1A1Ixp33_ASAP7_75t_SL g977 ( 
.A1(n_835),
.A2(n_832),
.B(n_888),
.C(n_909),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_788),
.B(n_878),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_796),
.A2(n_814),
.B(n_802),
.C(n_832),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_800),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_870),
.A2(n_811),
.B(n_890),
.Y(n_981)
);

AOI22x1_ASAP7_75t_L g982 ( 
.A1(n_795),
.A2(n_935),
.B1(n_863),
.B2(n_854),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_816),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_803),
.B(n_855),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_908),
.Y(n_985)
);

O2A1O1Ixp5_ASAP7_75t_L g986 ( 
.A1(n_792),
.A2(n_844),
.B(n_824),
.C(n_877),
.Y(n_986)
);

NAND3xp33_ASAP7_75t_SL g987 ( 
.A(n_871),
.B(n_805),
.C(n_949),
.Y(n_987)
);

BUFx12f_ASAP7_75t_L g988 ( 
.A(n_784),
.Y(n_988)
);

OAI21xp33_ASAP7_75t_SL g989 ( 
.A1(n_850),
.A2(n_887),
.B(n_865),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_847),
.B(n_799),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_839),
.A2(n_906),
.B1(n_882),
.B2(n_836),
.Y(n_991)
);

BUFx12f_ASAP7_75t_L g992 ( 
.A(n_784),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_810),
.B(n_822),
.Y(n_993)
);

INVx2_ASAP7_75t_SL g994 ( 
.A(n_817),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_916),
.A2(n_929),
.B(n_928),
.C(n_939),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_SL g996 ( 
.A(n_882),
.B(n_826),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_947),
.B(n_793),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_847),
.B(n_817),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_885),
.B(n_858),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_829),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_885),
.B(n_836),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_813),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_916),
.A2(n_929),
.B(n_944),
.C(n_792),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_911),
.A2(n_942),
.B(n_944),
.C(n_808),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_946),
.B(n_843),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_927),
.Y(n_1006)
);

O2A1O1Ixp5_ASAP7_75t_SL g1007 ( 
.A1(n_925),
.A2(n_875),
.B(n_867),
.C(n_852),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_821),
.B(n_828),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_900),
.B(n_830),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_830),
.B(n_941),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_861),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_922),
.Y(n_1012)
);

AOI221xp5_ASAP7_75t_L g1013 ( 
.A1(n_942),
.A2(n_948),
.B1(n_872),
.B2(n_880),
.C(n_918),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_833),
.A2(n_856),
.B(n_841),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_834),
.A2(n_785),
.B(n_945),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_941),
.B(n_849),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_930),
.B(n_931),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_896),
.Y(n_1018)
);

OA22x2_ASAP7_75t_L g1019 ( 
.A1(n_889),
.A2(n_923),
.B1(n_876),
.B2(n_845),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_920),
.A2(n_901),
.B1(n_894),
.B2(n_859),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_894),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_859),
.B(n_945),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_933),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_945),
.A2(n_789),
.B(n_794),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_945),
.A2(n_801),
.B(n_815),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_920),
.A2(n_859),
.B1(n_873),
.B2(n_862),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_937),
.Y(n_1027)
);

INVx3_ASAP7_75t_SL g1028 ( 
.A(n_787),
.Y(n_1028)
);

OAI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_846),
.A2(n_853),
.B(n_851),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_SL g1030 ( 
.A(n_943),
.B(n_914),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_860),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_902),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_806),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_848),
.B(n_884),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_857),
.B(n_895),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_898),
.B(n_934),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_SL g1037 ( 
.A(n_924),
.B(n_936),
.C(n_903),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_907),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_806),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_899),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_812),
.A2(n_819),
.B(n_804),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_926),
.B(n_932),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_910),
.B(n_840),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_820),
.B(n_838),
.Y(n_1044)
);

INVx6_ASAP7_75t_L g1045 ( 
.A(n_809),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_913),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_823),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_827),
.A2(n_886),
.B(n_891),
.C(n_893),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_879),
.A2(n_892),
.B(n_921),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_917),
.A2(n_919),
.B1(n_905),
.B2(n_912),
.Y(n_1050)
);

NAND3xp33_ASAP7_75t_L g1051 ( 
.A(n_904),
.B(n_629),
.C(n_642),
.Y(n_1051)
);

OAI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_915),
.A2(n_629),
.B1(n_780),
.B2(n_560),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_786),
.A2(n_629),
.B(n_782),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_781),
.A2(n_629),
.B(n_780),
.C(n_790),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_780),
.B(n_629),
.Y(n_1055)
);

INVxp67_ASAP7_75t_L g1056 ( 
.A(n_799),
.Y(n_1056)
);

NAND2x1p5_ASAP7_75t_L g1057 ( 
.A(n_800),
.B(n_849),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_SL g1058 ( 
.A(n_837),
.B(n_629),
.C(n_425),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_SL g1059 ( 
.A1(n_781),
.A2(n_790),
.B(n_780),
.C(n_925),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_SL g1060 ( 
.A(n_837),
.B(n_629),
.C(n_425),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_779),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_842),
.B(n_473),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_799),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_795),
.A2(n_629),
.B(n_870),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_790),
.B(n_629),
.Y(n_1065)
);

A2O1A1Ixp33_ASAP7_75t_L g1066 ( 
.A1(n_781),
.A2(n_629),
.B(n_780),
.C(n_642),
.Y(n_1066)
);

INVxp67_ASAP7_75t_L g1067 ( 
.A(n_799),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_809),
.A2(n_874),
.B(n_863),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_818),
.A2(n_629),
.B(n_870),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_800),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_790),
.B(n_629),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_780),
.B(n_629),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_800),
.Y(n_1073)
);

O2A1O1Ixp5_ASAP7_75t_L g1074 ( 
.A1(n_781),
.A2(n_629),
.B(n_642),
.C(n_780),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_780),
.B(n_629),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_779),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_781),
.A2(n_629),
.B(n_780),
.C(n_790),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_781),
.A2(n_629),
.B(n_780),
.C(n_790),
.Y(n_1078)
);

AO31x2_ASAP7_75t_L g1079 ( 
.A1(n_1026),
.A2(n_1003),
.A3(n_1066),
.B(n_1069),
.Y(n_1079)
);

OAI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1074),
.A2(n_995),
.B(n_1072),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_981),
.A2(n_1053),
.B(n_1064),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1075),
.A2(n_1077),
.B(n_1054),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1064),
.A2(n_1069),
.B(n_1024),
.Y(n_1083)
);

AO31x2_ASAP7_75t_L g1084 ( 
.A1(n_1026),
.A2(n_1050),
.A3(n_1043),
.B(n_1041),
.Y(n_1084)
);

INVx3_ASAP7_75t_L g1085 ( 
.A(n_1021),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_1001),
.Y(n_1086)
);

AO31x2_ASAP7_75t_L g1087 ( 
.A1(n_1050),
.A2(n_1041),
.A3(n_1044),
.B(n_1020),
.Y(n_1087)
);

OAI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_1078),
.A2(n_1055),
.B(n_1004),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_950),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_1025),
.A2(n_1015),
.B(n_989),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_1055),
.B(n_1058),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_971),
.B(n_1062),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_1028),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_976),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1065),
.A2(n_1071),
.B(n_979),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_978),
.B(n_973),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_1010),
.B(n_951),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_1044),
.A2(n_1020),
.A3(n_1049),
.B(n_1014),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_962),
.A2(n_975),
.A3(n_954),
.B(n_1035),
.Y(n_1099)
);

AO31x2_ASAP7_75t_L g1100 ( 
.A1(n_991),
.A2(n_970),
.A3(n_997),
.B(n_993),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_973),
.B(n_999),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_974),
.B(n_1046),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1060),
.A2(n_977),
.B(n_996),
.C(n_987),
.Y(n_1103)
);

AO32x2_ASAP7_75t_L g1104 ( 
.A1(n_959),
.A2(n_955),
.A3(n_986),
.B1(n_1059),
.B2(n_1007),
.Y(n_1104)
);

INVxp67_ASAP7_75t_L g1105 ( 
.A(n_1063),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_997),
.A2(n_993),
.A3(n_1034),
.B(n_959),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1023),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_994),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_1056),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_974),
.A2(n_1042),
.A3(n_958),
.B(n_1032),
.Y(n_1110)
);

OAI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1051),
.A2(n_1052),
.B(n_953),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_969),
.A2(n_967),
.B(n_1013),
.C(n_1048),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_988),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1029),
.A2(n_982),
.B(n_1047),
.Y(n_1114)
);

O2A1O1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_957),
.A2(n_965),
.B(n_1012),
.C(n_1030),
.Y(n_1115)
);

AO21x2_ASAP7_75t_L g1116 ( 
.A1(n_1068),
.A2(n_1037),
.B(n_964),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_984),
.B(n_990),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_960),
.A2(n_966),
.B1(n_955),
.B2(n_1040),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_1013),
.A2(n_961),
.B(n_1031),
.C(n_1005),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1022),
.A2(n_1019),
.B(n_1016),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1005),
.A2(n_1039),
.B(n_1038),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_998),
.B(n_1067),
.Y(n_1122)
);

AND2x2_ASAP7_75t_SL g1123 ( 
.A(n_983),
.B(n_1008),
.Y(n_1123)
);

AOI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_955),
.A2(n_1027),
.B1(n_968),
.B2(n_1061),
.Y(n_1124)
);

AOI21xp33_ASAP7_75t_L g1125 ( 
.A1(n_1036),
.A2(n_1002),
.B(n_1011),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_952),
.B(n_956),
.Y(n_1126)
);

NAND3x1_ASAP7_75t_L g1127 ( 
.A(n_1009),
.B(n_992),
.C(n_980),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_952),
.B(n_956),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1018),
.B(n_985),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1039),
.A2(n_1033),
.B(n_1017),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1000),
.B(n_1076),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1039),
.A2(n_1033),
.B(n_1017),
.Y(n_1132)
);

NOR2x1_ASAP7_75t_SL g1133 ( 
.A(n_1039),
.B(n_963),
.Y(n_1133)
);

BUFx8_ASAP7_75t_L g1134 ( 
.A(n_963),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_972),
.A2(n_1057),
.B(n_1006),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_972),
.A2(n_1057),
.B(n_1045),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_1070),
.A2(n_629),
.B1(n_1075),
.B2(n_1072),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_1073),
.B(n_1010),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_1054),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1140)
);

INVx5_ASAP7_75t_L g1141 ( 
.A(n_963),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1072),
.A2(n_629),
.B1(n_780),
.B2(n_560),
.Y(n_1142)
);

CKINVDCx11_ASAP7_75t_R g1143 ( 
.A(n_1028),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1147)
);

A2O1A1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_1054),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1066),
.A2(n_629),
.B(n_1074),
.Y(n_1150)
);

NOR2xp67_ASAP7_75t_SL g1151 ( 
.A(n_988),
.B(n_900),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_976),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1001),
.Y(n_1154)
);

BUFx10_ASAP7_75t_L g1155 ( 
.A(n_950),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_781),
.Y(n_1156)
);

AO32x2_ASAP7_75t_L g1157 ( 
.A1(n_1026),
.A2(n_1020),
.A3(n_959),
.B1(n_975),
.B2(n_991),
.Y(n_1157)
);

AOI221x1_ASAP7_75t_L g1158 ( 
.A1(n_1066),
.A2(n_629),
.B1(n_995),
.B2(n_781),
.C(n_955),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1159)
);

OR2x2_ASAP7_75t_L g1160 ( 
.A(n_1055),
.B(n_797),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1161)
);

A2O1A1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_1054),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1058),
.A2(n_629),
.B1(n_1060),
.B2(n_642),
.Y(n_1164)
);

AO32x2_ASAP7_75t_L g1165 ( 
.A1(n_1026),
.A2(n_1020),
.A3(n_959),
.B1(n_975),
.B2(n_991),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_976),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1001),
.Y(n_1167)
);

INVx3_ASAP7_75t_SL g1168 ( 
.A(n_950),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1066),
.A2(n_629),
.B(n_1074),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1062),
.B(n_473),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1172)
);

AOI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1024),
.A2(n_1069),
.B(n_1015),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_963),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_781),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1001),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1068),
.A2(n_1025),
.B(n_1024),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_976),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1181)
);

A2O1A1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_1054),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_1054),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_L g1185 ( 
.A(n_1072),
.B(n_629),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1066),
.A2(n_629),
.B(n_1074),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1066),
.A2(n_629),
.B(n_1074),
.Y(n_1188)
);

BUFx12f_ASAP7_75t_L g1189 ( 
.A(n_988),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1066),
.A2(n_629),
.B(n_1074),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_971),
.B(n_629),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_950),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1072),
.A2(n_629),
.B1(n_1075),
.B2(n_780),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_SL g1195 ( 
.A1(n_979),
.A2(n_969),
.B(n_973),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1062),
.B(n_473),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1066),
.A2(n_629),
.B(n_1074),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1001),
.Y(n_1199)
);

INVxp67_ASAP7_75t_SL g1200 ( 
.A(n_1056),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_971),
.B(n_629),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1026),
.A2(n_1003),
.A3(n_1066),
.B(n_1069),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_981),
.A2(n_629),
.B(n_1053),
.Y(n_1204)
);

INVx1_ASAP7_75t_SL g1205 ( 
.A(n_976),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_L g1206 ( 
.A1(n_1072),
.A2(n_1075),
.B1(n_629),
.B2(n_1060),
.C(n_1058),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1072),
.B(n_1075),
.Y(n_1207)
);

OAI22x1_ASAP7_75t_L g1208 ( 
.A1(n_962),
.A2(n_629),
.B1(n_1075),
.B2(n_1072),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_781),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1021),
.Y(n_1210)
);

A2O1A1Ixp33_ASAP7_75t_L g1211 ( 
.A1(n_1072),
.A2(n_629),
.B(n_1075),
.C(n_1054),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1072),
.B(n_629),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_L g1213 ( 
.A(n_1070),
.B(n_952),
.Y(n_1213)
);

AOI22xp5_ASAP7_75t_L g1214 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1193),
.B2(n_1206),
.Y(n_1214)
);

INVx1_ASAP7_75t_SL g1215 ( 
.A(n_1205),
.Y(n_1215)
);

BUFx12f_ASAP7_75t_L g1216 ( 
.A(n_1143),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_1093),
.Y(n_1217)
);

OAI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1101),
.A2(n_1202),
.B1(n_1207),
.B2(n_1181),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1192),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1118),
.A2(n_1191),
.B1(n_1201),
.B2(n_1096),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1107),
.Y(n_1221)
);

OAI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1118),
.A2(n_1175),
.B1(n_1147),
.B2(n_1163),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1208),
.A2(n_1164),
.B1(n_1142),
.B2(n_1091),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1089),
.Y(n_1224)
);

OAI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1137),
.A2(n_1158),
.B1(n_1160),
.B2(n_1102),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1139),
.A2(n_1211),
.B1(n_1184),
.B2(n_1162),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1166),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1148),
.B(n_1182),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1189),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1141),
.Y(n_1230)
);

NAND2x1p5_ASAP7_75t_L g1231 ( 
.A(n_1141),
.B(n_1136),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1097),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1082),
.A2(n_1080),
.B1(n_1088),
.B2(n_1123),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1092),
.A2(n_1195),
.B1(n_1186),
.B2(n_1150),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1179),
.Y(n_1235)
);

INVx6_ASAP7_75t_L g1236 ( 
.A(n_1134),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1137),
.A2(n_1117),
.B1(n_1171),
.B2(n_1196),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1086),
.Y(n_1238)
);

BUFx2_ASAP7_75t_R g1239 ( 
.A(n_1168),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1169),
.A2(n_1198),
.B1(n_1190),
.B2(n_1188),
.Y(n_1240)
);

BUFx2_ASAP7_75t_SL g1241 ( 
.A(n_1097),
.Y(n_1241)
);

CKINVDCx11_ASAP7_75t_R g1242 ( 
.A(n_1155),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1095),
.A2(n_1124),
.B1(n_1111),
.B2(n_1114),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1155),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1174),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1124),
.A2(n_1125),
.B1(n_1109),
.B2(n_1122),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1113),
.Y(n_1247)
);

INVx2_ASAP7_75t_SL g1248 ( 
.A(n_1108),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1154),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1205),
.A2(n_1105),
.B1(n_1094),
.B2(n_1200),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1167),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1156),
.B(n_1176),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_1134),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1177),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1153),
.Y(n_1255)
);

AOI22xp33_ASAP7_75t_L g1256 ( 
.A1(n_1120),
.A2(n_1199),
.B1(n_1129),
.B2(n_1138),
.Y(n_1256)
);

BUFx8_ASAP7_75t_L g1257 ( 
.A(n_1138),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1128),
.A2(n_1151),
.B1(n_1172),
.B2(n_1183),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1144),
.A2(n_1204),
.B1(n_1197),
.B2(n_1194),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1157),
.Y(n_1260)
);

OAI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1126),
.A2(n_1115),
.B1(n_1209),
.B2(n_1121),
.Y(n_1261)
);

AND2x6_ASAP7_75t_L g1262 ( 
.A(n_1085),
.B(n_1210),
.Y(n_1262)
);

OAI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1083),
.A2(n_1187),
.B1(n_1180),
.B2(n_1081),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1103),
.A2(n_1112),
.B(n_1119),
.Y(n_1264)
);

BUFx10_ASAP7_75t_L g1265 ( 
.A(n_1127),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1157),
.A2(n_1165),
.B1(n_1133),
.B2(n_1104),
.Y(n_1266)
);

CKINVDCx6p67_ASAP7_75t_R g1267 ( 
.A(n_1213),
.Y(n_1267)
);

CKINVDCx11_ASAP7_75t_R g1268 ( 
.A(n_1213),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1090),
.A2(n_1165),
.B1(n_1157),
.B2(n_1130),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1099),
.B(n_1165),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1135),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1116),
.A2(n_1132),
.B1(n_1178),
.B2(n_1170),
.Y(n_1272)
);

HB1xp67_ASAP7_75t_L g1273 ( 
.A(n_1087),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1099),
.B(n_1106),
.Y(n_1274)
);

BUFx4_ASAP7_75t_SL g1275 ( 
.A(n_1100),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1087),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1104),
.A2(n_1079),
.B1(n_1203),
.B2(n_1084),
.Y(n_1277)
);

NAND2x1p5_ASAP7_75t_L g1278 ( 
.A(n_1140),
.B(n_1145),
.Y(n_1278)
);

CKINVDCx14_ASAP7_75t_R g1279 ( 
.A(n_1100),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1087),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1104),
.A2(n_1203),
.B1(n_1079),
.B2(n_1173),
.Y(n_1281)
);

INVx5_ASAP7_75t_L g1282 ( 
.A(n_1110),
.Y(n_1282)
);

OAI22x1_ASAP7_75t_L g1283 ( 
.A1(n_1203),
.A2(n_1110),
.B1(n_1084),
.B2(n_1098),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1146),
.A2(n_1161),
.B1(n_1149),
.B2(n_1152),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1084),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1098),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_SL g1287 ( 
.A1(n_1098),
.A2(n_629),
.B1(n_1212),
.B2(n_1185),
.Y(n_1287)
);

OAI22xp33_ASAP7_75t_L g1288 ( 
.A1(n_1110),
.A2(n_1185),
.B1(n_1212),
.B2(n_629),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1159),
.A2(n_629),
.B1(n_1185),
.B2(n_1212),
.Y(n_1289)
);

BUFx2_ASAP7_75t_SL g1290 ( 
.A(n_1093),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_1143),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1141),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1131),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_SL g1294 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_425),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1153),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1139),
.B(n_1148),
.Y(n_1296)
);

BUFx2_ASAP7_75t_SL g1297 ( 
.A(n_1093),
.Y(n_1297)
);

CKINVDCx8_ASAP7_75t_R g1298 ( 
.A(n_1089),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1131),
.Y(n_1299)
);

OAI22xp5_ASAP7_75t_L g1300 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1072),
.B2(n_1075),
.Y(n_1300)
);

INVxp67_ASAP7_75t_SL g1301 ( 
.A(n_1114),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1166),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1305)
);

BUFx3_ASAP7_75t_L g1306 ( 
.A(n_1166),
.Y(n_1306)
);

CKINVDCx6p67_ASAP7_75t_R g1307 ( 
.A(n_1143),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1072),
.B2(n_1075),
.Y(n_1309)
);

INVx6_ASAP7_75t_L g1310 ( 
.A(n_1134),
.Y(n_1310)
);

BUFx10_ASAP7_75t_L g1311 ( 
.A(n_1089),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_629),
.B2(n_1193),
.Y(n_1313)
);

OAI22xp5_ASAP7_75t_L g1314 ( 
.A1(n_1185),
.A2(n_1212),
.B1(n_1072),
.B2(n_1075),
.Y(n_1314)
);

BUFx2_ASAP7_75t_L g1315 ( 
.A(n_1166),
.Y(n_1315)
);

INVx4_ASAP7_75t_L g1316 ( 
.A(n_1141),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1141),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1143),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1205),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1143),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1185),
.A2(n_629),
.B1(n_1212),
.B2(n_1060),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1278),
.A2(n_1284),
.B(n_1272),
.Y(n_1325)
);

INVxp33_ASAP7_75t_L g1326 ( 
.A(n_1227),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1271),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1276),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1280),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1257),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1278),
.A2(n_1259),
.B(n_1286),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1263),
.A2(n_1301),
.B(n_1240),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1270),
.B(n_1287),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1295),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1274),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1225),
.B(n_1218),
.Y(n_1336)
);

OA21x2_ASAP7_75t_L g1337 ( 
.A1(n_1243),
.A2(n_1285),
.B(n_1301),
.Y(n_1337)
);

OAI211xp5_ASAP7_75t_SL g1338 ( 
.A1(n_1294),
.A2(n_1324),
.B(n_1312),
.C(n_1302),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1273),
.Y(n_1339)
);

BUFx6f_ASAP7_75t_L g1340 ( 
.A(n_1231),
.Y(n_1340)
);

INVx2_ASAP7_75t_L g1341 ( 
.A(n_1283),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1214),
.A2(n_1264),
.B(n_1226),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1273),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1287),
.B(n_1266),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1257),
.Y(n_1345)
);

OAI21xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1233),
.A2(n_1260),
.B(n_1228),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1225),
.B(n_1218),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1275),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1230),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1275),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1269),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1295),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1279),
.B(n_1277),
.Y(n_1353)
);

AO21x2_ASAP7_75t_L g1354 ( 
.A1(n_1263),
.A2(n_1288),
.B(n_1281),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_1260),
.Y(n_1355)
);

BUFx4f_ASAP7_75t_L g1356 ( 
.A(n_1262),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1269),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1304),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1215),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1282),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1221),
.Y(n_1361)
);

AOI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1252),
.A2(n_1226),
.B(n_1228),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1222),
.B(n_1313),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1288),
.A2(n_1281),
.B(n_1296),
.Y(n_1364)
);

OAI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1313),
.A2(n_1303),
.B(n_1308),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1262),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1315),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1222),
.B(n_1289),
.Y(n_1368)
);

HB1xp67_ASAP7_75t_L g1369 ( 
.A(n_1321),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1262),
.Y(n_1370)
);

BUFx2_ASAP7_75t_L g1371 ( 
.A(n_1255),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1234),
.B(n_1223),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1293),
.B(n_1299),
.Y(n_1373)
);

BUFx3_ASAP7_75t_L g1374 ( 
.A(n_1262),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1230),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1238),
.Y(n_1376)
);

AO21x1_ASAP7_75t_L g1377 ( 
.A1(n_1220),
.A2(n_1261),
.B(n_1300),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1249),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1251),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1254),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1258),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_SL g1382 ( 
.A(n_1239),
.Y(n_1382)
);

INVx2_ASAP7_75t_SL g1383 ( 
.A(n_1230),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1241),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1246),
.B(n_1237),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1256),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1294),
.A2(n_1322),
.B1(n_1305),
.B2(n_1320),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1250),
.Y(n_1388)
);

INVx1_ASAP7_75t_SL g1389 ( 
.A(n_1235),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1306),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1317),
.A2(n_1309),
.B(n_1300),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1309),
.A2(n_1314),
.B1(n_1310),
.B2(n_1253),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1314),
.A2(n_1267),
.B(n_1265),
.Y(n_1393)
);

NAND2x1p5_ASAP7_75t_L g1394 ( 
.A(n_1316),
.B(n_1318),
.Y(n_1394)
);

INVxp67_ASAP7_75t_L g1395 ( 
.A(n_1248),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1292),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1332),
.B(n_1253),
.Y(n_1397)
);

NAND3xp33_ASAP7_75t_L g1398 ( 
.A(n_1342),
.B(n_1268),
.C(n_1242),
.Y(n_1398)
);

OAI22xp5_ASAP7_75t_L g1399 ( 
.A1(n_1387),
.A2(n_1310),
.B1(n_1253),
.B2(n_1236),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1342),
.A2(n_1232),
.B(n_1292),
.C(n_1318),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1355),
.B(n_1290),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1333),
.B(n_1265),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1388),
.B(n_1297),
.Y(n_1403)
);

INVx5_ASAP7_75t_L g1404 ( 
.A(n_1340),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1355),
.B(n_1311),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1388),
.B(n_1244),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1361),
.B(n_1307),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1365),
.A2(n_1338),
.B(n_1332),
.C(n_1346),
.Y(n_1408)
);

NAND2xp33_ASAP7_75t_R g1409 ( 
.A(n_1337),
.B(n_1224),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1371),
.B(n_1311),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1367),
.B(n_1239),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1367),
.B(n_1310),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1377),
.A2(n_1318),
.B(n_1245),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1353),
.B(n_1236),
.Y(n_1414)
);

O2A1O1Ixp33_ASAP7_75t_L g1415 ( 
.A1(n_1338),
.A2(n_1217),
.B(n_1323),
.C(n_1291),
.Y(n_1415)
);

AO32x2_ASAP7_75t_L g1416 ( 
.A1(n_1327),
.A2(n_1245),
.A3(n_1229),
.B1(n_1247),
.B2(n_1216),
.Y(n_1416)
);

AO32x2_ASAP7_75t_L g1417 ( 
.A1(n_1327),
.A2(n_1219),
.A3(n_1298),
.B1(n_1319),
.B2(n_1364),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1392),
.A2(n_1382),
.B1(n_1365),
.B2(n_1385),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1377),
.B(n_1372),
.Y(n_1419)
);

O2A1O1Ixp33_ASAP7_75t_L g1420 ( 
.A1(n_1363),
.A2(n_1347),
.B(n_1336),
.C(n_1368),
.Y(n_1420)
);

OAI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1363),
.A2(n_1327),
.B1(n_1385),
.B2(n_1336),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1359),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1340),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1331),
.A2(n_1347),
.B(n_1325),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1368),
.A2(n_1372),
.B(n_1346),
.C(n_1381),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1356),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_SL g1428 ( 
.A(n_1362),
.B(n_1340),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1390),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1430)
);

A2O1A1Ixp33_ASAP7_75t_L g1431 ( 
.A1(n_1391),
.A2(n_1356),
.B(n_1344),
.C(n_1393),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1356),
.A2(n_1344),
.B(n_1393),
.C(n_1366),
.Y(n_1432)
);

OAI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1382),
.A2(n_1327),
.B1(n_1384),
.B2(n_1389),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1330),
.A2(n_1345),
.B1(n_1384),
.B2(n_1348),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1373),
.B(n_1376),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1373),
.B(n_1379),
.Y(n_1436)
);

A2O1A1Ixp33_ASAP7_75t_L g1437 ( 
.A1(n_1393),
.A2(n_1374),
.B(n_1366),
.C(n_1370),
.Y(n_1437)
);

BUFx5_ASAP7_75t_L g1438 ( 
.A(n_1360),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1331),
.A2(n_1325),
.B(n_1341),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1425),
.B(n_1354),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1408),
.A2(n_1358),
.B1(n_1334),
.B2(n_1352),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1425),
.B(n_1354),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1430),
.B(n_1351),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1408),
.A2(n_1369),
.B1(n_1350),
.B2(n_1370),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1430),
.B(n_1357),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1425),
.B(n_1354),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1439),
.B(n_1354),
.Y(n_1447)
);

AOI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1418),
.A2(n_1419),
.B1(n_1421),
.B2(n_1409),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1439),
.B(n_1341),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1422),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1419),
.A2(n_1374),
.B1(n_1389),
.B2(n_1337),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1404),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1439),
.B(n_1341),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1431),
.B(n_1328),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1431),
.B(n_1329),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1435),
.B(n_1364),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1417),
.B(n_1364),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1436),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1438),
.Y(n_1459)
);

HB1xp67_ASAP7_75t_L g1460 ( 
.A(n_1409),
.Y(n_1460)
);

INVx4_ASAP7_75t_L g1461 ( 
.A(n_1452),
.Y(n_1461)
);

NAND3xp33_ASAP7_75t_L g1462 ( 
.A(n_1448),
.B(n_1420),
.C(n_1426),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1448),
.A2(n_1399),
.B1(n_1397),
.B2(n_1433),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1454),
.B(n_1455),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1449),
.B(n_1339),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1449),
.Y(n_1466)
);

HB1xp67_ASAP7_75t_L g1467 ( 
.A(n_1449),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1454),
.B(n_1417),
.Y(n_1468)
);

OAI221xp5_ASAP7_75t_L g1469 ( 
.A1(n_1448),
.A2(n_1398),
.B1(n_1432),
.B2(n_1415),
.C(n_1406),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1454),
.B(n_1417),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1453),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1442),
.B(n_1339),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1455),
.B(n_1428),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1455),
.B(n_1424),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1441),
.A2(n_1397),
.B1(n_1403),
.B2(n_1427),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1443),
.B(n_1335),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1453),
.B(n_1438),
.Y(n_1477)
);

NAND3x1_ASAP7_75t_SL g1478 ( 
.A(n_1457),
.B(n_1416),
.C(n_1411),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1447),
.B(n_1438),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1447),
.B(n_1438),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1442),
.B(n_1343),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1461),
.B(n_1459),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1471),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1465),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1476),
.B(n_1456),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1460),
.Y(n_1486)
);

NOR2x1_ASAP7_75t_L g1487 ( 
.A(n_1462),
.B(n_1441),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1465),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1465),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1469),
.B(n_1407),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1464),
.B(n_1460),
.Y(n_1491)
);

NAND4xp25_ASAP7_75t_L g1492 ( 
.A(n_1462),
.B(n_1444),
.C(n_1451),
.D(n_1457),
.Y(n_1492)
);

NOR2xp33_ASAP7_75t_L g1493 ( 
.A(n_1469),
.B(n_1405),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1465),
.B(n_1443),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1471),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1464),
.B(n_1456),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1472),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1476),
.B(n_1456),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1464),
.B(n_1458),
.Y(n_1499)
);

NOR2xp33_ASAP7_75t_L g1500 ( 
.A(n_1462),
.B(n_1423),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1472),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1472),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1461),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1473),
.B(n_1458),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1472),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1481),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1481),
.B(n_1445),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1463),
.B(n_1444),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1481),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1481),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1471),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1467),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1473),
.B(n_1458),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1467),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1476),
.B(n_1445),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1466),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1473),
.B(n_1450),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1514),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1514),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1486),
.B(n_1473),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1486),
.B(n_1468),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1483),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1483),
.Y(n_1523)
);

AOI32xp33_ASAP7_75t_L g1524 ( 
.A1(n_1487),
.A2(n_1468),
.A3(n_1470),
.B1(n_1451),
.B2(n_1457),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1499),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1468),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1491),
.B(n_1496),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1499),
.Y(n_1528)
);

OAI211xp5_ASAP7_75t_L g1529 ( 
.A1(n_1487),
.A2(n_1463),
.B(n_1475),
.C(n_1468),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1483),
.Y(n_1530)
);

INVxp67_ASAP7_75t_L g1531 ( 
.A(n_1500),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1493),
.B(n_1410),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1503),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1500),
.B(n_1470),
.Y(n_1534)
);

HB1xp67_ASAP7_75t_L g1535 ( 
.A(n_1512),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1512),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1503),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1515),
.B(n_1507),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1495),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1484),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1484),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1496),
.B(n_1470),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1490),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1488),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1488),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1489),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1489),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1515),
.B(n_1507),
.Y(n_1548)
);

AND2x4_ASAP7_75t_L g1549 ( 
.A(n_1503),
.B(n_1479),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1508),
.B(n_1470),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1495),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1497),
.Y(n_1553)
);

OAI22xp33_ASAP7_75t_SL g1554 ( 
.A1(n_1492),
.A2(n_1463),
.B1(n_1478),
.B2(n_1442),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1494),
.B(n_1466),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1492),
.B(n_1429),
.Y(n_1556)
);

NOR2x1p5_ASAP7_75t_SL g1557 ( 
.A(n_1495),
.B(n_1466),
.Y(n_1557)
);

NOR4xp25_ASAP7_75t_L g1558 ( 
.A(n_1497),
.B(n_1395),
.C(n_1457),
.D(n_1401),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1511),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1535),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1531),
.B(n_1543),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1538),
.B(n_1485),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1556),
.B(n_1513),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1527),
.B(n_1513),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1550),
.B(n_1485),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1538),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1558),
.B(n_1498),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1533),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1527),
.B(n_1503),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1548),
.B(n_1498),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1520),
.B(n_1517),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1529),
.B(n_1413),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1536),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1548),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1536),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1518),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1518),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1534),
.B(n_1517),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1554),
.B(n_1494),
.Y(n_1580)
);

OAI211xp5_ASAP7_75t_L g1581 ( 
.A1(n_1524),
.A2(n_1475),
.B(n_1432),
.C(n_1440),
.Y(n_1581)
);

NAND3xp33_ASAP7_75t_L g1582 ( 
.A(n_1524),
.B(n_1446),
.C(n_1440),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1519),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1520),
.B(n_1482),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1519),
.B(n_1501),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1522),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1554),
.B(n_1474),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1521),
.B(n_1482),
.Y(n_1588)
);

AOI221xp5_ASAP7_75t_L g1589 ( 
.A1(n_1532),
.A2(n_1501),
.B1(n_1502),
.B2(n_1505),
.C(n_1506),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1525),
.B(n_1502),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1540),
.Y(n_1591)
);

AOI21xp33_ASAP7_75t_SL g1592 ( 
.A1(n_1549),
.A2(n_1434),
.B(n_1478),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1525),
.B(n_1474),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1528),
.B(n_1521),
.Y(n_1594)
);

NAND3x1_ASAP7_75t_L g1595 ( 
.A(n_1533),
.B(n_1412),
.C(n_1478),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1540),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1567),
.B(n_1526),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1583),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1591),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1575),
.Y(n_1600)
);

NOR2x1_ASAP7_75t_L g1601 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1561),
.Y(n_1602)
);

AOI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1573),
.A2(n_1446),
.B1(n_1447),
.B2(n_1397),
.Y(n_1603)
);

AOI21xp33_ASAP7_75t_SL g1604 ( 
.A1(n_1573),
.A2(n_1478),
.B(n_1416),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1562),
.B(n_1528),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1573),
.A2(n_1478),
.B1(n_1397),
.B2(n_1437),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1564),
.B(n_1326),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1569),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1580),
.A2(n_1437),
.B(n_1400),
.Y(n_1609)
);

AOI32xp33_ASAP7_75t_L g1610 ( 
.A1(n_1568),
.A2(n_1526),
.A3(n_1549),
.B1(n_1542),
.B2(n_1480),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1582),
.A2(n_1446),
.B1(n_1447),
.B2(n_1549),
.Y(n_1611)
);

NAND3xp33_ASAP7_75t_L g1612 ( 
.A(n_1592),
.B(n_1544),
.C(n_1541),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1555),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1581),
.A2(n_1544),
.B(n_1541),
.Y(n_1614)
);

AOI31xp33_ASAP7_75t_L g1615 ( 
.A1(n_1587),
.A2(n_1589),
.A3(n_1578),
.B(n_1577),
.Y(n_1615)
);

AOI211x1_ASAP7_75t_L g1616 ( 
.A1(n_1566),
.A2(n_1542),
.B(n_1560),
.C(n_1551),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1569),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1563),
.B(n_1345),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1574),
.B(n_1545),
.Y(n_1619)
);

AOI222xp33_ASAP7_75t_L g1620 ( 
.A1(n_1594),
.A2(n_1557),
.B1(n_1446),
.B2(n_1402),
.C1(n_1480),
.C2(n_1479),
.Y(n_1620)
);

INVxp33_ASAP7_75t_L g1621 ( 
.A(n_1570),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_L g1622 ( 
.A(n_1563),
.B(n_1345),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1600),
.B(n_1565),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1618),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1602),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1597),
.B(n_1621),
.Y(n_1626)
);

OAI21xp5_ASAP7_75t_SL g1627 ( 
.A1(n_1615),
.A2(n_1570),
.B(n_1414),
.Y(n_1627)
);

INVxp67_ASAP7_75t_L g1628 ( 
.A(n_1622),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1598),
.B(n_1565),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1601),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1619),
.Y(n_1631)
);

AOI22xp33_ASAP7_75t_L g1632 ( 
.A1(n_1606),
.A2(n_1571),
.B1(n_1593),
.B2(n_1549),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1608),
.B(n_1617),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1619),
.Y(n_1634)
);

AOI221xp5_ASAP7_75t_L g1635 ( 
.A1(n_1604),
.A2(n_1612),
.B1(n_1610),
.B2(n_1614),
.C(n_1606),
.Y(n_1635)
);

INVx2_ASAP7_75t_SL g1636 ( 
.A(n_1605),
.Y(n_1636)
);

INVx1_ASAP7_75t_SL g1637 ( 
.A(n_1613),
.Y(n_1637)
);

AOI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1609),
.A2(n_1576),
.B1(n_1596),
.B2(n_1571),
.C(n_1585),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1609),
.A2(n_1595),
.B(n_1585),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1599),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1607),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1629),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1629),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1636),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1636),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1625),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1627),
.A2(n_1595),
.B1(n_1635),
.B2(n_1603),
.Y(n_1647)
);

O2A1O1Ixp33_ASAP7_75t_SL g1648 ( 
.A1(n_1630),
.A2(n_1611),
.B(n_1533),
.C(n_1537),
.Y(n_1648)
);

AOI222xp33_ASAP7_75t_L g1649 ( 
.A1(n_1638),
.A2(n_1557),
.B1(n_1616),
.B2(n_1588),
.C1(n_1572),
.C2(n_1620),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1623),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1633),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1639),
.A2(n_1637),
.B(n_1641),
.Y(n_1652)
);

INVx1_ASAP7_75t_SL g1653 ( 
.A(n_1644),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1642),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1651),
.Y(n_1655)
);

NOR2x1_ASAP7_75t_SL g1656 ( 
.A(n_1645),
.B(n_1633),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1651),
.B(n_1626),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1650),
.B(n_1641),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1643),
.B(n_1626),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_L g1660 ( 
.A(n_1652),
.B(n_1646),
.C(n_1628),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1648),
.Y(n_1661)
);

OAI22xp33_ASAP7_75t_L g1662 ( 
.A1(n_1647),
.A2(n_1624),
.B1(n_1631),
.B2(n_1634),
.Y(n_1662)
);

AOI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1662),
.A2(n_1640),
.B(n_1634),
.C(n_1649),
.Y(n_1663)
);

AOI311xp33_ASAP7_75t_L g1664 ( 
.A1(n_1660),
.A2(n_1632),
.A3(n_1547),
.B(n_1553),
.C(n_1546),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1661),
.B(n_1586),
.C(n_1590),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1658),
.B(n_1586),
.C(n_1588),
.D(n_1584),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1653),
.B(n_1656),
.Y(n_1667)
);

NAND4xp25_ASAP7_75t_L g1668 ( 
.A(n_1659),
.B(n_1584),
.C(n_1414),
.D(n_1590),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_SL g1669 ( 
.A(n_1657),
.B(n_1537),
.Y(n_1669)
);

NOR3xp33_ASAP7_75t_L g1670 ( 
.A(n_1667),
.B(n_1663),
.C(n_1654),
.Y(n_1670)
);

NAND4xp25_ASAP7_75t_L g1671 ( 
.A(n_1664),
.B(n_1655),
.C(n_1537),
.D(n_1572),
.Y(n_1671)
);

OAI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1666),
.A2(n_1655),
.B1(n_1537),
.B2(n_1545),
.C(n_1546),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1669),
.A2(n_1665),
.B(n_1668),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1667),
.A2(n_1553),
.B(n_1547),
.Y(n_1674)
);

AOI311xp33_ASAP7_75t_L g1675 ( 
.A1(n_1663),
.A2(n_1505),
.A3(n_1510),
.B(n_1506),
.C(n_1509),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1673),
.A2(n_1670),
.B1(n_1672),
.B2(n_1674),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1671),
.B(n_1555),
.Y(n_1677)
);

NAND4xp75_ASAP7_75t_L g1678 ( 
.A(n_1675),
.B(n_1416),
.C(n_1523),
.D(n_1530),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1670),
.B(n_1509),
.Y(n_1679)
);

NOR2x1_ASAP7_75t_L g1680 ( 
.A(n_1671),
.B(n_1522),
.Y(n_1680)
);

NOR3xp33_ASAP7_75t_SL g1681 ( 
.A(n_1676),
.B(n_1679),
.C(n_1678),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1680),
.B(n_1516),
.Y(n_1682)
);

A2O1A1Ixp33_ASAP7_75t_L g1683 ( 
.A1(n_1677),
.A2(n_1539),
.B(n_1559),
.C(n_1552),
.Y(n_1683)
);

AOI22xp5_ASAP7_75t_L g1684 ( 
.A1(n_1681),
.A2(n_1539),
.B1(n_1559),
.B2(n_1552),
.Y(n_1684)
);

OA22x2_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1682),
.B1(n_1683),
.B2(n_1552),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1685),
.B(n_1551),
.Y(n_1686)
);

OAI22xp33_ASAP7_75t_SL g1687 ( 
.A1(n_1685),
.A2(n_1559),
.B1(n_1539),
.B2(n_1530),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1686),
.A2(n_1530),
.B1(n_1523),
.B2(n_1522),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1687),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1689),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1688),
.A2(n_1523),
.B(n_1560),
.Y(n_1691)
);

OR2x6_ASAP7_75t_L g1692 ( 
.A(n_1690),
.B(n_1416),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1692),
.B(n_1691),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1693),
.Y(n_1694)
);

OAI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1694),
.A2(n_1394),
.B1(n_1383),
.B2(n_1375),
.C(n_1349),
.Y(n_1695)
);

AOI211xp5_ASAP7_75t_L g1696 ( 
.A1(n_1695),
.A2(n_1375),
.B(n_1383),
.C(n_1396),
.Y(n_1696)
);


endmodule