module fake_netlist_5_290_n_1687 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1687);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1687;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_2),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

BUFx8_ASAP7_75t_SL g157 ( 
.A(n_149),
.Y(n_157)
);

BUFx5_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_82),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_23),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_78),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_95),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_106),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_142),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_89),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_63),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_140),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_51),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_41),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_30),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_109),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_65),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_72),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_74),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_57),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_25),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_87),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_11),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_86),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_1),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_79),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_111),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_8),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_88),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_5),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_81),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_131),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_33),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_104),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_14),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_40),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_59),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_5),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_26),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_18),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_68),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_42),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_150),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_145),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_48),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_103),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_53),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_38),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_12),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_135),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_16),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_97),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_152),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_15),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_128),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_119),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_34),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_110),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_47),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_116),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_64),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_100),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_34),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_52),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_18),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_16),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_114),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_49),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_146),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_141),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_127),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_69),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_22),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_6),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_10),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_130),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_98),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_60),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_93),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_118),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_21),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_4),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_55),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_91),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_30),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_32),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_105),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_139),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_117),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_66),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_37),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_21),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_15),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_75),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_38),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_99),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_13),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_144),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_90),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_92),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_28),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_120),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_44),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_3),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_77),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_56),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_4),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_137),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_20),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_24),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_94),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_36),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_108),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_23),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_29),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_36),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_28),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_35),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_121),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_122),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_47),
.Y(n_296)
);

BUFx8_ASAP7_75t_SL g297 ( 
.A(n_22),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_71),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_148),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_83),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_39),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_43),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_7),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_96),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_3),
.Y(n_305)
);

HB1xp67_ASAP7_75t_SL g306 ( 
.A(n_24),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_277),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_277),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_299),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_157),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_297),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_194),
.Y(n_315)
);

INVxp33_ASAP7_75t_SL g316 ( 
.A(n_154),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_194),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_173),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_173),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_248),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g322 ( 
.A(n_274),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_186),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_186),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_160),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_192),
.Y(n_326)
);

BUFx2_ASAP7_75t_L g327 ( 
.A(n_154),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_158),
.Y(n_328)
);

INVxp67_ASAP7_75t_SL g329 ( 
.A(n_238),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_199),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_210),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_158),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_216),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_226),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_191),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_229),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_193),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_242),
.Y(n_338)
);

INVxp67_ASAP7_75t_SL g339 ( 
.A(n_238),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_252),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_265),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_176),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_289),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_200),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_305),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_204),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_292),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_175),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_211),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g351 ( 
.A(n_156),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g353 ( 
.A(n_237),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_253),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_158),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_306),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_212),
.Y(n_357)
);

INVxp33_ASAP7_75t_SL g358 ( 
.A(n_182),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_197),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_182),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_197),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_218),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_213),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_214),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_162),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_218),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_231),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_231),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_268),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_188),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_188),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_250),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_250),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_282),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_215),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_189),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_219),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_251),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_335),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_309),
.B(n_163),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_307),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_163),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_360),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_310),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_329),
.B(n_240),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

BUFx8_ASAP7_75t_L g393 ( 
.A(n_327),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_356),
.B(n_247),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_314),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_337),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_314),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_345),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_312),
.B(n_155),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_328),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_371),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_328),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_349),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_332),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_332),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_316),
.B(n_209),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_347),
.B(n_251),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_352),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_378),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_327),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_359),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_350),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_355),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_322),
.B(n_270),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_355),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_365),
.B(n_260),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_353),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_355),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_361),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

AND2x2_ASAP7_75t_SL g427 ( 
.A(n_370),
.B(n_260),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_357),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_262),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_362),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_364),
.B(n_375),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_362),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_320),
.A2(n_283),
.B1(n_303),
.B2(n_302),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_358),
.B(n_155),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_339),
.B(n_262),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_276),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_313),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_366),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

CKINVDCx6p67_ASAP7_75t_R g441 ( 
.A(n_342),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_318),
.B(n_280),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_311),
.B(n_159),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_400),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_380),
.Y(n_445)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_400),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_427),
.A2(n_376),
.B(n_276),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_379),
.Y(n_448)
);

INVx1_ASAP7_75t_SL g449 ( 
.A(n_441),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_376),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_400),
.Y(n_451)
);

OAI21xp33_ASAP7_75t_L g452 ( 
.A1(n_394),
.A2(n_331),
.B(n_321),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_391),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_379),
.B(n_367),
.Y(n_454)
);

BUFx4f_ASAP7_75t_L g455 ( 
.A(n_436),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_400),
.Y(n_456)
);

NOR3xp33_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_236),
.C(n_217),
.Y(n_457)
);

INVx6_ASAP7_75t_L g458 ( 
.A(n_382),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_436),
.B(n_382),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_390),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_441),
.Y(n_461)
);

BUFx3_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_382),
.B(n_367),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_429),
.B(n_331),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_380),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_392),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_392),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_391),
.B(n_318),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_395),
.Y(n_471)
);

AND2x6_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_222),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_386),
.B(n_368),
.Y(n_473)
);

INVxp67_ASAP7_75t_SL g474 ( 
.A(n_400),
.Y(n_474)
);

BUFx6f_ASAP7_75t_SL g475 ( 
.A(n_427),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_389),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_389),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_427),
.B(n_222),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_395),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_423),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_436),
.B(n_422),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_437),
.B(n_321),
.Y(n_482)
);

AND3x1_ASAP7_75t_L g483 ( 
.A(n_410),
.B(n_323),
.C(n_319),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_389),
.Y(n_484)
);

BUFx10_ASAP7_75t_L g485 ( 
.A(n_431),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_393),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_415),
.A2(n_254),
.B1(n_203),
.B2(n_205),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_397),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_419),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_435),
.B(n_319),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_385),
.B(n_442),
.Y(n_492)
);

INVx8_ASAP7_75t_L g493 ( 
.A(n_386),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_386),
.B(n_368),
.Y(n_494)
);

CKINVDCx11_ASAP7_75t_R g495 ( 
.A(n_423),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_323),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_404),
.Y(n_497)
);

CKINVDCx6p67_ASAP7_75t_R g498 ( 
.A(n_399),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_422),
.B(n_222),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_386),
.A2(n_422),
.B1(n_442),
.B2(n_421),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_388),
.B(n_381),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_422),
.B(n_372),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_383),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_405),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_396),
.B(n_222),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_405),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_401),
.B(n_324),
.C(n_206),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_402),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_398),
.B(n_222),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_409),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_417),
.B(n_168),
.Y(n_513)
);

BUFx6f_ASAP7_75t_SL g514 ( 
.A(n_409),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_411),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_408),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_384),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_428),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_408),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_439),
.B(n_171),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_411),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_408),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_R g523 ( 
.A(n_438),
.B(n_159),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_403),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_403),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_403),
.Y(n_526)
);

AO21x2_ASAP7_75t_L g527 ( 
.A1(n_418),
.A2(n_174),
.B(n_172),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_413),
.B(n_324),
.Y(n_528)
);

BUFx10_ASAP7_75t_L g529 ( 
.A(n_413),
.Y(n_529)
);

INVx1_ASAP7_75t_SL g530 ( 
.A(n_414),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_418),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_403),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_384),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_414),
.Y(n_534)
);

BUFx6f_ASAP7_75t_SL g535 ( 
.A(n_416),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_393),
.A2(n_207),
.B1(n_275),
.B2(n_245),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_418),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_416),
.Y(n_538)
);

AND2x6_ASAP7_75t_L g539 ( 
.A(n_403),
.B(n_178),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_403),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_L g542 ( 
.A(n_407),
.B(n_158),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_393),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_425),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_407),
.B(n_372),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_407),
.B(n_373),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_420),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_393),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_420),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_425),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_406),
.Y(n_551)
);

BUFx10_ASAP7_75t_L g552 ( 
.A(n_430),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_407),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_407),
.B(n_373),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_384),
.Y(n_555)
);

BUFx10_ASAP7_75t_L g556 ( 
.A(n_430),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_406),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_406),
.Y(n_558)
);

BUFx10_ASAP7_75t_L g559 ( 
.A(n_432),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_384),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_432),
.B(n_325),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_384),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_384),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_406),
.B(n_224),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_424),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_424),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_424),
.B(n_225),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_424),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_439),
.B(n_179),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_439),
.B(n_181),
.Y(n_571)
);

AND3x2_ASAP7_75t_L g572 ( 
.A(n_440),
.B(n_185),
.C(n_183),
.Y(n_572)
);

NOR3xp33_ASAP7_75t_L g573 ( 
.A(n_426),
.B(n_288),
.C(n_220),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_387),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_SL g575 ( 
.A1(n_440),
.A2(n_170),
.B1(n_369),
.B2(n_374),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_426),
.B(n_230),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_387),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_439),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_440),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_439),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_440),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_426),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_387),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_426),
.B(n_195),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_459),
.B(n_434),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_568),
.Y(n_586)
);

O2A1O1Ixp33_ASAP7_75t_L g587 ( 
.A1(n_478),
.A2(n_338),
.B(n_326),
.C(n_346),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_453),
.B(n_161),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_450),
.B(n_161),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_465),
.B(n_164),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_455),
.A2(n_434),
.B(n_196),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_458),
.A2(n_241),
.B1(n_198),
.B2(n_300),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_482),
.B(n_223),
.C(n_256),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_459),
.B(n_462),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_459),
.B(n_434),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_462),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_458),
.B(n_434),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_455),
.B(n_164),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_448),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_478),
.A2(n_221),
.B1(n_287),
.B2(n_285),
.Y(n_600)
);

NOR2xp67_ASAP7_75t_L g601 ( 
.A(n_579),
.B(n_348),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_568),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_481),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_492),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_458),
.B(n_202),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_481),
.B(n_325),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_447),
.B(n_266),
.C(n_201),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_452),
.B(n_165),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

INVxp67_ASAP7_75t_L g610 ( 
.A(n_496),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_208),
.Y(n_611)
);

A2O1A1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_500),
.A2(n_255),
.B(n_243),
.C(n_272),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_582),
.B(n_234),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_493),
.B(n_232),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_561),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_493),
.B(n_239),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_530),
.B(n_348),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

NAND2x1_ASAP7_75t_L g619 ( 
.A(n_444),
.B(n_446),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_527),
.A2(n_158),
.B1(n_293),
.B2(n_291),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_561),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_497),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_493),
.B(n_249),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_493),
.B(n_463),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_529),
.B(n_165),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_470),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_518),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_501),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_529),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_506),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_475),
.A2(n_257),
.B1(n_261),
.B2(n_263),
.Y(n_631)
);

BUFx12f_ASAP7_75t_SL g632 ( 
.A(n_495),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_508),
.Y(n_633)
);

NOR2x1p5_ASAP7_75t_L g634 ( 
.A(n_581),
.B(n_189),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_473),
.B(n_166),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_505),
.B(n_513),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_494),
.B(n_512),
.Y(n_637)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_488),
.B(n_326),
.Y(n_638)
);

O2A1O1Ixp5_ASAP7_75t_L g639 ( 
.A1(n_499),
.A2(n_346),
.B(n_344),
.C(n_343),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_515),
.B(n_166),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_521),
.B(n_167),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_551),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_534),
.B(n_167),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_538),
.B(n_169),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_541),
.B(n_169),
.Y(n_645)
);

BUFx5_ASAP7_75t_L g646 ( 
.A(n_539),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_544),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_551),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_491),
.B(n_513),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_557),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_529),
.B(n_177),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_552),
.B(n_177),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_550),
.B(n_180),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_507),
.B(n_330),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_504),
.B(n_180),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_527),
.A2(n_158),
.B1(n_291),
.B2(n_286),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_552),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_507),
.B(n_184),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_511),
.B(n_552),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_556),
.B(n_184),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_579),
.B(n_330),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_556),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_503),
.B(n_333),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_460),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_511),
.B(n_490),
.Y(n_665)
);

INVxp67_ASAP7_75t_L g666 ( 
.A(n_483),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_556),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_557),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_528),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_L g670 ( 
.A(n_509),
.B(n_573),
.C(n_457),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_464),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_559),
.B(n_187),
.Y(n_672)
);

A2O1A1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_467),
.A2(n_344),
.B(n_343),
.C(n_341),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_468),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_559),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_471),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_479),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_558),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_449),
.B(n_461),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_489),
.B(n_576),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_523),
.B(n_259),
.C(n_264),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_559),
.B(n_190),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_564),
.B(n_190),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_567),
.B(n_227),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_472),
.B(n_158),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_475),
.B(n_227),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_490),
.B(n_333),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_490),
.B(n_267),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_454),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_485),
.B(n_334),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_474),
.B(n_267),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_545),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_558),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_485),
.B(n_273),
.Y(n_694)
);

INVxp67_ASAP7_75t_L g695 ( 
.A(n_475),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_499),
.B(n_273),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_444),
.B(n_279),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_485),
.B(n_334),
.Y(n_698)
);

AO221x1_ASAP7_75t_L g699 ( 
.A1(n_444),
.A2(n_341),
.B1(n_340),
.B2(n_338),
.C(n_336),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_565),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_539),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_480),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_446),
.B(n_279),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_546),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_554),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_445),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_498),
.B(n_294),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_498),
.A2(n_294),
.B1(n_295),
.B2(n_298),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_518),
.B(n_336),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_446),
.B(n_295),
.Y(n_710)
);

NOR3x1_ASAP7_75t_L g711 ( 
.A(n_487),
.B(n_543),
.C(n_340),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_445),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_514),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_456),
.B(n_298),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_581),
.B(n_304),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_466),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_466),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_469),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_514),
.B(n_304),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_514),
.B(n_228),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_535),
.B(n_233),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_536),
.B(n_235),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_480),
.B(n_575),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_495),
.B(n_317),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_535),
.Y(n_725)
);

INVx2_ASAP7_75t_SL g726 ( 
.A(n_527),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_535),
.B(n_244),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_469),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_472),
.B(n_246),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_525),
.B(n_258),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_476),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_570),
.B(n_293),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_539),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_476),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_525),
.B(n_317),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_472),
.A2(n_286),
.B1(n_303),
.B2(n_302),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_566),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_477),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_472),
.A2(n_584),
.B1(n_539),
.B2(n_531),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_525),
.B(n_315),
.Y(n_740)
);

AO22x2_ASAP7_75t_L g741 ( 
.A1(n_584),
.A2(n_315),
.B1(n_1),
.B2(n_6),
.Y(n_741)
);

BUFx6f_ASAP7_75t_SL g742 ( 
.A(n_548),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_520),
.B(n_301),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_572),
.Y(n_744)
);

NOR2x1p5_ASAP7_75t_L g745 ( 
.A(n_548),
.B(n_296),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_539),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_609),
.B(n_517),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_649),
.A2(n_539),
.B1(n_477),
.B2(n_484),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_603),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_709),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_627),
.B(n_702),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_632),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_617),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_649),
.B(n_526),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_659),
.B(n_526),
.Y(n_755)
);

INVx2_ASAP7_75t_SL g756 ( 
.A(n_687),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_663),
.B(n_269),
.Y(n_757)
);

BUFx3_ASAP7_75t_L g758 ( 
.A(n_606),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_690),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_610),
.B(n_566),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_742),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_606),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_698),
.Y(n_763)
);

INVx5_ASAP7_75t_L g764 ( 
.A(n_701),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_589),
.A2(n_520),
.B1(n_569),
.B2(n_571),
.Y(n_765)
);

OR2x6_ASAP7_75t_L g766 ( 
.A(n_679),
.B(n_569),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_695),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_701),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_596),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_615),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_659),
.B(n_629),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_621),
.Y(n_772)
);

INVxp67_ASAP7_75t_SL g773 ( 
.A(n_594),
.Y(n_773)
);

INVx3_ASAP7_75t_L g774 ( 
.A(n_586),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_695),
.B(n_571),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_604),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_629),
.B(n_526),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_657),
.B(n_526),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_657),
.B(n_689),
.Y(n_779)
);

OR2x6_ASAP7_75t_L g780 ( 
.A(n_662),
.B(n_578),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_610),
.B(n_486),
.Y(n_781)
);

INVx5_ASAP7_75t_L g782 ( 
.A(n_701),
.Y(n_782)
);

HB1xp67_ASAP7_75t_L g783 ( 
.A(n_604),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_599),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_622),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_590),
.B(n_669),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_665),
.B(n_553),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_628),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_737),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_701),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_642),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_724),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_669),
.B(n_451),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_648),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_630),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_650),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_R g797 ( 
.A(n_667),
.B(n_269),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_626),
.B(n_271),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_733),
.Y(n_799)
);

INVx2_ASAP7_75t_SL g800 ( 
.A(n_654),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_741),
.A2(n_484),
.B1(n_271),
.B2(n_284),
.Y(n_801)
);

INVx5_ASAP7_75t_L g802 ( 
.A(n_733),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_733),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_680),
.B(n_486),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_633),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_636),
.B(n_553),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_611),
.Y(n_807)
);

BUFx6f_ASAP7_75t_L g808 ( 
.A(n_733),
.Y(n_808)
);

BUFx4f_ASAP7_75t_L g809 ( 
.A(n_661),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_637),
.B(n_502),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_732),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_647),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_746),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_664),
.Y(n_814)
);

AO22x1_ASAP7_75t_L g815 ( 
.A1(n_707),
.A2(n_278),
.B1(n_281),
.B2(n_284),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_671),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_607),
.B(n_553),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_674),
.Y(n_818)
);

BUFx6f_ASAP7_75t_L g819 ( 
.A(n_746),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_676),
.Y(n_820)
);

INVx2_ASAP7_75t_SL g821 ( 
.A(n_638),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_677),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_675),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_668),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_746),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_602),
.Y(n_826)
);

OR2x2_ASAP7_75t_SL g827 ( 
.A(n_681),
.B(n_593),
.Y(n_827)
);

BUFx4f_ASAP7_75t_L g828 ( 
.A(n_661),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_742),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_741),
.A2(n_620),
.B1(n_656),
.B2(n_600),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_735),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_666),
.A2(n_580),
.B1(n_578),
.B2(n_451),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_R g833 ( 
.A(n_686),
.B(n_278),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_678),
.Y(n_834)
);

NAND3xp33_ASAP7_75t_SL g835 ( 
.A(n_670),
.B(n_281),
.C(n_580),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_666),
.B(n_540),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_693),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_585),
.B(n_583),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_743),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_SL g840 ( 
.A1(n_741),
.A2(n_0),
.B1(n_9),
.B2(n_10),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_613),
.B(n_692),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_588),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_595),
.B(n_583),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_704),
.B(n_537),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_713),
.B(n_540),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_601),
.B(n_517),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_686),
.Y(n_847)
);

OAI22xp33_ASAP7_75t_L g848 ( 
.A1(n_661),
.A2(n_516),
.B1(n_510),
.B2(n_502),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_618),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_713),
.B(n_533),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_700),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_705),
.B(n_510),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_619),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_706),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_672),
.B(n_540),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_740),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_725),
.B(n_533),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_672),
.B(n_562),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_624),
.B(n_555),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_658),
.B(n_655),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_712),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_SL g862 ( 
.A1(n_707),
.A2(n_0),
.B1(n_9),
.B2(n_13),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_682),
.B(n_516),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_726),
.B(n_555),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_646),
.B(n_555),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_646),
.Y(n_866)
);

AND2x2_ASAP7_75t_SL g867 ( 
.A(n_620),
.B(n_542),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_716),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_646),
.B(n_682),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_717),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_658),
.B(n_547),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_718),
.Y(n_872)
);

AND2x4_ASAP7_75t_L g873 ( 
.A(n_725),
.B(n_562),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_728),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_730),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_731),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_635),
.B(n_547),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_734),
.Y(n_878)
);

AOI21xp33_ASAP7_75t_L g879 ( 
.A1(n_608),
.A2(n_542),
.B(n_522),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_744),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_646),
.B(n_555),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_670),
.B(n_519),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_738),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_608),
.B(n_537),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_646),
.B(n_560),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_688),
.B(n_519),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_640),
.Y(n_887)
);

INVx4_ASAP7_75t_L g888 ( 
.A(n_600),
.Y(n_888)
);

OAI22xp5_ASAP7_75t_SL g889 ( 
.A1(n_736),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_597),
.B(n_563),
.Y(n_890)
);

OAI22xp33_ASAP7_75t_L g891 ( 
.A1(n_708),
.A2(n_696),
.B1(n_722),
.B2(n_631),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_683),
.B(n_549),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_694),
.B(n_549),
.Y(n_893)
);

AO22x1_ASAP7_75t_L g894 ( 
.A1(n_719),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_894)
);

AND2x2_ASAP7_75t_SL g895 ( 
.A(n_656),
.B(n_560),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_723),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_720),
.B(n_25),
.Y(n_897)
);

BUFx2_ASAP7_75t_L g898 ( 
.A(n_600),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_736),
.A2(n_563),
.B1(n_560),
.B2(n_532),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_684),
.B(n_563),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_625),
.B(n_560),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_634),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_720),
.B(n_26),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_605),
.Y(n_904)
);

AO22x1_ASAP7_75t_L g905 ( 
.A1(n_721),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_641),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_587),
.B(n_563),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_721),
.B(n_27),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_639),
.Y(n_909)
);

BUFx8_ASAP7_75t_L g910 ( 
.A(n_711),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_697),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_703),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_651),
.B(n_31),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_587),
.B(n_532),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_727),
.Y(n_915)
);

NOR3xp33_ASAP7_75t_SL g916 ( 
.A(n_652),
.B(n_32),
.C(n_33),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_699),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_660),
.B(n_35),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_727),
.B(n_715),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_739),
.B(n_532),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_643),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_644),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_830),
.A2(n_612),
.B1(n_739),
.B2(n_653),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_919),
.B(n_645),
.C(n_598),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_786),
.B(n_616),
.Y(n_925)
);

A2O1A1Ixp33_ASAP7_75t_L g926 ( 
.A1(n_913),
.A2(n_591),
.B(n_714),
.C(n_710),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_750),
.B(n_614),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_841),
.B(n_691),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_785),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_807),
.B(n_623),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_764),
.B(n_532),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_788),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_753),
.B(n_592),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_860),
.B(n_673),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_911),
.B(n_729),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_807),
.B(n_685),
.Y(n_936)
);

AO22x1_ASAP7_75t_L g937 ( 
.A1(n_918),
.A2(n_745),
.B1(n_39),
.B2(n_40),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_759),
.B(n_37),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_795),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_854),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_896),
.A2(n_524),
.B1(n_574),
.B2(n_577),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_757),
.B(n_759),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_921),
.B(n_41),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_867),
.A2(n_577),
.B(n_574),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_922),
.B(n_42),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_781),
.B(n_44),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_756),
.B(n_763),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_805),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_773),
.B(n_45),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_868),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_880),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_830),
.A2(n_574),
.B1(n_46),
.B2(n_45),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_870),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_880),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_752),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_900),
.A2(n_574),
.B(n_50),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_776),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_758),
.B(n_84),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_821),
.B(n_46),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_839),
.B(n_776),
.Y(n_960)
);

O2A1O1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_835),
.A2(n_918),
.B(n_891),
.C(n_783),
.Y(n_961)
);

NOR2x1_ASAP7_75t_L g962 ( 
.A(n_823),
.B(n_54),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_887),
.B(n_574),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_751),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_814),
.Y(n_965)
);

NAND2x2_ASAP7_75t_L g966 ( 
.A(n_823),
.B(n_58),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_835),
.A2(n_61),
.B(n_62),
.C(n_70),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_768),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_847),
.B(n_73),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_768),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_768),
.Y(n_971)
);

AND2x4_ASAP7_75t_SL g972 ( 
.A(n_751),
.B(n_80),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_773),
.B(n_102),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_879),
.A2(n_107),
.B(n_112),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_891),
.A2(n_113),
.B(n_115),
.C(n_136),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_768),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_869),
.A2(n_855),
.B(n_817),
.C(n_771),
.Y(n_977)
);

CKINVDCx6p67_ASAP7_75t_R g978 ( 
.A(n_751),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_872),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_R g980 ( 
.A(n_915),
.B(n_761),
.Y(n_980)
);

A2O1A1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_867),
.A2(n_765),
.B(n_893),
.C(n_858),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_760),
.B(n_906),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_758),
.B(n_762),
.Y(n_983)
);

NAND2x1p5_ASAP7_75t_L g984 ( 
.A(n_764),
.B(n_782),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_798),
.B(n_800),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_863),
.B(n_858),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_875),
.B(n_836),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_762),
.B(n_784),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_883),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_784),
.B(n_812),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_882),
.B(n_904),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_818),
.Y(n_992)
);

A2O1A1Ixp33_ASAP7_75t_L g993 ( 
.A1(n_893),
.A2(n_842),
.B(n_882),
.C(n_836),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_799),
.Y(n_994)
);

INVx2_ASAP7_75t_SL g995 ( 
.A(n_792),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_820),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_801),
.A2(n_840),
.B1(n_895),
.B2(n_748),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_SL g998 ( 
.A(n_897),
.B(n_903),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_804),
.A2(n_810),
.B(n_754),
.Y(n_999)
);

AND2x4_ASAP7_75t_L g1000 ( 
.A(n_850),
.B(n_857),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_754),
.A2(n_884),
.B(n_869),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_812),
.B(n_816),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_871),
.A2(n_892),
.B(n_885),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_831),
.B(n_856),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_783),
.A2(n_771),
.B(n_779),
.C(n_908),
.Y(n_1005)
);

OR2x6_ASAP7_75t_SL g1006 ( 
.A(n_829),
.B(n_902),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_801),
.A2(n_840),
.B1(n_895),
.B2(n_748),
.Y(n_1007)
);

O2A1O1Ixp5_ASAP7_75t_L g1008 ( 
.A1(n_855),
.A2(n_817),
.B(n_917),
.C(n_787),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_816),
.B(n_809),
.Y(n_1009)
);

OAI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_889),
.A2(n_899),
.B1(n_888),
.B2(n_898),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_799),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_793),
.B(n_822),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_912),
.A2(n_901),
.B(n_770),
.C(n_772),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_767),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_809),
.B(n_828),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_865),
.A2(n_885),
.B(n_881),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_861),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_766),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_779),
.B(n_811),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_766),
.B(n_827),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_861),
.Y(n_1021)
);

INVxp67_ASAP7_75t_SL g1022 ( 
.A(n_799),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_766),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_899),
.A2(n_888),
.B1(n_828),
.B2(n_862),
.Y(n_1024)
);

AND2x6_ASAP7_75t_SL g1025 ( 
.A(n_775),
.B(n_845),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_833),
.B(n_912),
.Y(n_1026)
);

XOR2xp5_ASAP7_75t_L g1027 ( 
.A(n_886),
.B(n_850),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_799),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_775),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_749),
.A2(n_920),
.B1(n_916),
.B2(n_769),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_833),
.B(n_747),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_806),
.A2(n_916),
.B(n_848),
.C(n_787),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_838),
.A2(n_843),
.B(n_881),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_R g1034 ( 
.A(n_803),
.B(n_808),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_L g1035 ( 
.A(n_815),
.B(n_905),
.C(n_894),
.Y(n_1035)
);

O2A1O1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_806),
.A2(n_848),
.B(n_755),
.C(n_878),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_857),
.B(n_873),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_873),
.B(n_775),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_910),
.Y(n_1039)
);

BUFx3_ASAP7_75t_L g1040 ( 
.A(n_910),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_797),
.B(n_747),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_846),
.B(n_797),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_901),
.A2(n_877),
.B(n_876),
.C(n_874),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_L g1044 ( 
.A(n_777),
.B(n_778),
.C(n_755),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_791),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_832),
.A2(n_844),
.B(n_852),
.C(n_824),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_846),
.B(n_782),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_764),
.B(n_782),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_790),
.B(n_764),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_782),
.B(n_802),
.Y(n_1050)
);

BUFx6f_ASAP7_75t_L g1051 ( 
.A(n_803),
.Y(n_1051)
);

INVx5_ASAP7_75t_L g1052 ( 
.A(n_803),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_802),
.B(n_813),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_SL g1054 ( 
.A(n_802),
.B(n_813),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_774),
.B(n_849),
.Y(n_1055)
);

BUFx10_ASAP7_75t_L g1056 ( 
.A(n_845),
.Y(n_1056)
);

OAI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_920),
.A2(n_907),
.B1(n_813),
.B2(n_802),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_813),
.A2(n_909),
.B1(n_825),
.B2(n_819),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_780),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_865),
.A2(n_859),
.B(n_864),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_794),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_803),
.A2(n_825),
.B1(n_819),
.B2(n_808),
.Y(n_1062)
);

O2A1O1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_838),
.A2(n_843),
.B(n_859),
.C(n_777),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_929),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_1049),
.A2(n_999),
.B(n_926),
.Y(n_1065)
);

OAI22x1_ASAP7_75t_L g1066 ( 
.A1(n_1035),
.A2(n_1020),
.B1(n_1029),
.B2(n_1023),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_932),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_939),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_986),
.B(n_851),
.Y(n_1069)
);

OAI21xp33_ASAP7_75t_SL g1070 ( 
.A1(n_997),
.A2(n_890),
.B(n_914),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_995),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_942),
.B(n_834),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_961),
.A2(n_774),
.B(n_849),
.C(n_826),
.Y(n_1073)
);

NAND3x1_ASAP7_75t_L g1074 ( 
.A(n_969),
.B(n_826),
.C(n_780),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1004),
.B(n_837),
.Y(n_1075)
);

NOR4xp25_ASAP7_75t_L g1076 ( 
.A(n_997),
.B(n_796),
.C(n_789),
.D(n_845),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_954),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_1027),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1003),
.A2(n_808),
.B(n_819),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_928),
.A2(n_819),
.B(n_825),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1001),
.A2(n_825),
.B(n_853),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_948),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_1007),
.A2(n_1013),
.A3(n_1058),
.B(n_1057),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_930),
.B(n_853),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_965),
.Y(n_1085)
);

NOR2xp67_ASAP7_75t_L g1086 ( 
.A(n_991),
.B(n_853),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_992),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1000),
.B(n_853),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_977),
.A2(n_925),
.B(n_973),
.Y(n_1089)
);

BUFx10_ASAP7_75t_L g1090 ( 
.A(n_938),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_1063),
.A2(n_944),
.B(n_1058),
.Y(n_1091)
);

AO31x2_ASAP7_75t_L g1092 ( 
.A1(n_1057),
.A2(n_1043),
.A3(n_923),
.B(n_1030),
.Y(n_1092)
);

AO31x2_ASAP7_75t_L g1093 ( 
.A1(n_923),
.A2(n_1030),
.A3(n_1010),
.B(n_1046),
.Y(n_1093)
);

OAI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1008),
.A2(n_934),
.B(n_1036),
.Y(n_1094)
);

OAI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_934),
.A2(n_1032),
.B(n_993),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_996),
.Y(n_1096)
);

AOI21x1_ASAP7_75t_SL g1097 ( 
.A1(n_949),
.A2(n_935),
.B(n_946),
.Y(n_1097)
);

OAI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_974),
.A2(n_1005),
.B(n_944),
.Y(n_1098)
);

OA21x2_ASAP7_75t_L g1099 ( 
.A1(n_1044),
.A2(n_1012),
.B(n_956),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_968),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_985),
.B(n_1037),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_982),
.B(n_987),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_998),
.A2(n_1018),
.B1(n_924),
.B2(n_1024),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1010),
.A2(n_952),
.B1(n_1024),
.B2(n_991),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_940),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_984),
.A2(n_1052),
.B(n_936),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_980),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_950),
.Y(n_1108)
);

INVx4_ASAP7_75t_L g1109 ( 
.A(n_1052),
.Y(n_1109)
);

INVx4_ASAP7_75t_L g1110 ( 
.A(n_1052),
.Y(n_1110)
);

OAI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_959),
.A2(n_945),
.B(n_943),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1041),
.B(n_1000),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_953),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_947),
.B(n_957),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_979),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_989),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_936),
.B(n_1019),
.Y(n_1117)
);

O2A1O1Ixp5_ASAP7_75t_SL g1118 ( 
.A1(n_952),
.A2(n_927),
.B(n_1026),
.C(n_963),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1045),
.Y(n_1119)
);

AND2x4_ASAP7_75t_L g1120 ( 
.A(n_983),
.B(n_1009),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_968),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1061),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_1062),
.A2(n_1055),
.A3(n_1017),
.B(n_1021),
.Y(n_1123)
);

AO31x2_ASAP7_75t_L g1124 ( 
.A1(n_1038),
.A2(n_975),
.A3(n_967),
.B(n_1025),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1059),
.Y(n_1125)
);

CKINVDCx6p67_ASAP7_75t_R g1126 ( 
.A(n_1006),
.Y(n_1126)
);

AO21x2_ASAP7_75t_L g1127 ( 
.A1(n_933),
.A2(n_941),
.B(n_1034),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_966),
.A2(n_1056),
.A3(n_962),
.B(n_1054),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1011),
.B(n_1022),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_1031),
.A2(n_1042),
.B1(n_937),
.B2(n_1015),
.Y(n_1130)
);

OAI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_990),
.A2(n_1002),
.B(n_1047),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_931),
.A2(n_1053),
.B(n_1050),
.Y(n_1132)
);

AO21x2_ASAP7_75t_L g1133 ( 
.A1(n_1048),
.A2(n_988),
.B(n_958),
.Y(n_1133)
);

OA21x2_ASAP7_75t_L g1134 ( 
.A1(n_958),
.A2(n_960),
.B(n_983),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_968),
.Y(n_1135)
);

A2O1A1Ixp33_ASAP7_75t_L g1136 ( 
.A1(n_951),
.A2(n_972),
.B(n_964),
.C(n_1052),
.Y(n_1136)
);

OR2x2_ASAP7_75t_L g1137 ( 
.A(n_1014),
.B(n_978),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_931),
.A2(n_1028),
.B(n_970),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1056),
.A2(n_1051),
.A3(n_970),
.B(n_971),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1051),
.A2(n_994),
.B(n_970),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_955),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_971),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1039),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_971),
.B(n_976),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_976),
.A2(n_994),
.B(n_1028),
.Y(n_1145)
);

OA22x2_ASAP7_75t_L g1146 ( 
.A1(n_1040),
.A2(n_889),
.B1(n_862),
.B2(n_821),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1028),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_1051),
.Y(n_1148)
);

BUFx10_ASAP7_75t_L g1149 ( 
.A(n_969),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_981),
.A2(n_977),
.B(n_1008),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_968),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_986),
.B(n_1004),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_991),
.B(n_896),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_SL g1154 ( 
.A(n_997),
.B(n_1007),
.Y(n_1154)
);

AOI221xp5_ASAP7_75t_L g1155 ( 
.A1(n_961),
.A2(n_649),
.B1(n_589),
.B2(n_610),
.C(n_452),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1049),
.A2(n_455),
.B(n_866),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_986),
.B(n_786),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_997),
.A2(n_1007),
.B1(n_830),
.B2(n_649),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_929),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_986),
.B(n_1004),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_SL g1161 ( 
.A1(n_1005),
.A2(n_1032),
.B(n_975),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_930),
.B(n_847),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_986),
.B(n_786),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_929),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_930),
.B(n_786),
.Y(n_1165)
);

AO31x2_ASAP7_75t_L g1166 ( 
.A1(n_981),
.A2(n_1007),
.A3(n_997),
.B(n_1013),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_980),
.Y(n_1167)
);

NAND3x1_ASAP7_75t_L g1168 ( 
.A(n_969),
.B(n_723),
.C(n_913),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_968),
.Y(n_1169)
);

CKINVDCx16_ASAP7_75t_R g1170 ( 
.A(n_980),
.Y(n_1170)
);

A2O1A1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_961),
.A2(n_649),
.B(n_981),
.C(n_589),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_986),
.B(n_786),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_1052),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_986),
.B(n_786),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_986),
.B(n_786),
.Y(n_1175)
);

BUFx8_ASAP7_75t_L g1176 ( 
.A(n_1014),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_1014),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_981),
.A2(n_1001),
.B(n_1013),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1033),
.A2(n_1060),
.B(n_1016),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_986),
.B(n_786),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_929),
.Y(n_1181)
);

INVxp67_ASAP7_75t_L g1182 ( 
.A(n_960),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1049),
.A2(n_455),
.B(n_866),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_981),
.A2(n_1007),
.A3(n_997),
.B(n_1013),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1008),
.A2(n_977),
.B(n_1001),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_929),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_929),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_L g1188 ( 
.A(n_930),
.B(n_807),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_929),
.Y(n_1189)
);

AO32x2_ASAP7_75t_L g1190 ( 
.A1(n_997),
.A2(n_1007),
.A3(n_1010),
.B1(n_952),
.B2(n_1024),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_929),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1154),
.A2(n_1158),
.B1(n_1155),
.B2(n_1146),
.Y(n_1192)
);

NAND2x1p5_ASAP7_75t_L g1193 ( 
.A(n_1134),
.B(n_1109),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1156),
.A2(n_1183),
.B(n_1065),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1101),
.B(n_1072),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1085),
.Y(n_1196)
);

OR2x6_ASAP7_75t_L g1197 ( 
.A(n_1074),
.B(n_1168),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1165),
.B(n_1157),
.Y(n_1198)
);

INVx1_ASAP7_75t_SL g1199 ( 
.A(n_1114),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1158),
.A2(n_1154),
.B(n_1171),
.C(n_1070),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_SL g1201 ( 
.A1(n_1117),
.A2(n_1073),
.B(n_1095),
.C(n_1136),
.Y(n_1201)
);

OA21x2_ASAP7_75t_L g1202 ( 
.A1(n_1150),
.A2(n_1098),
.B(n_1094),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_1092),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_1170),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1091),
.A2(n_1089),
.B(n_1095),
.Y(n_1205)
);

OAI211xp5_ASAP7_75t_SL g1206 ( 
.A1(n_1070),
.A2(n_1162),
.B(n_1103),
.C(n_1111),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1147),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1163),
.A2(n_1172),
.B(n_1174),
.C(n_1180),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1175),
.B(n_1152),
.Y(n_1209)
);

BUFx8_ASAP7_75t_L g1210 ( 
.A(n_1078),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1186),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1179),
.A2(n_1081),
.B(n_1079),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1120),
.B(n_1088),
.Y(n_1213)
);

OA21x2_ASAP7_75t_L g1214 ( 
.A1(n_1161),
.A2(n_1111),
.B(n_1117),
.Y(n_1214)
);

NOR2xp33_ASAP7_75t_L g1215 ( 
.A(n_1152),
.B(n_1160),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1104),
.A2(n_1106),
.B(n_1080),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1187),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1189),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_SL g1219 ( 
.A1(n_1190),
.A2(n_1149),
.B1(n_1090),
.B2(n_1160),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1064),
.Y(n_1220)
);

NOR2xp67_ASAP7_75t_L g1221 ( 
.A(n_1107),
.B(n_1167),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1097),
.A2(n_1132),
.B(n_1118),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_SL g1223 ( 
.A(n_1127),
.B(n_1110),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1153),
.B(n_1104),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1084),
.A2(n_1188),
.B(n_1130),
.C(n_1102),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1067),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1082),
.Y(n_1227)
);

NOR2xp67_ASAP7_75t_SL g1228 ( 
.A(n_1110),
.B(n_1173),
.Y(n_1228)
);

BUFx8_ASAP7_75t_L g1229 ( 
.A(n_1177),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1176),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1087),
.Y(n_1231)
);

AND2x4_ASAP7_75t_SL g1232 ( 
.A(n_1120),
.B(n_1149),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_L g1233 ( 
.A1(n_1076),
.A2(n_1066),
.B1(n_1182),
.B2(n_1125),
.C(n_1069),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1185),
.A2(n_1099),
.B(n_1138),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1188),
.B(n_1075),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1185),
.A2(n_1099),
.B(n_1145),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1086),
.A2(n_1071),
.B1(n_1131),
.B2(n_1181),
.Y(n_1237)
);

INVx3_ASAP7_75t_L g1238 ( 
.A(n_1088),
.Y(n_1238)
);

INVxp67_ASAP7_75t_SL g1239 ( 
.A(n_1096),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1159),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1131),
.A2(n_1140),
.B(n_1129),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1164),
.Y(n_1242)
);

CKINVDCx20_ASAP7_75t_R g1243 ( 
.A(n_1176),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1191),
.Y(n_1244)
);

INVx2_ASAP7_75t_SL g1245 ( 
.A(n_1077),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1119),
.A2(n_1116),
.B(n_1115),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1105),
.A2(n_1108),
.B(n_1122),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1090),
.A2(n_1178),
.B1(n_1190),
.B2(n_1113),
.Y(n_1248)
);

BUFx8_ASAP7_75t_SL g1249 ( 
.A(n_1112),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1137),
.A2(n_1126),
.B1(n_1135),
.B2(n_1141),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1190),
.B(n_1148),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1123),
.Y(n_1252)
);

AO21x2_ASAP7_75t_L g1253 ( 
.A1(n_1133),
.A2(n_1142),
.B(n_1092),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1083),
.A2(n_1092),
.B(n_1093),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1166),
.B(n_1184),
.Y(n_1255)
);

AO21x2_ASAP7_75t_L g1256 ( 
.A1(n_1166),
.A2(n_1184),
.B(n_1124),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1166),
.A2(n_1184),
.B(n_1124),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1144),
.B(n_1100),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1143),
.B(n_1100),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1121),
.A2(n_1151),
.B1(n_1169),
.B2(n_1124),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1128),
.A2(n_1139),
.B(n_1121),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1128),
.Y(n_1262)
);

AO21x2_ASAP7_75t_L g1263 ( 
.A1(n_1065),
.A2(n_1098),
.B(n_1161),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_SL g1264 ( 
.A1(n_1161),
.A2(n_1005),
.B(n_1032),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1156),
.A2(n_1183),
.B(n_1065),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1171),
.A2(n_589),
.B(n_590),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1171),
.A2(n_589),
.B(n_649),
.C(n_786),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1101),
.B(n_1072),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1154),
.A2(n_1158),
.B1(n_889),
.B2(n_1155),
.Y(n_1269)
);

A2O1A1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1158),
.A2(n_649),
.B(n_1154),
.C(n_1007),
.Y(n_1270)
);

O2A1O1Ixp33_ASAP7_75t_SL g1271 ( 
.A1(n_1171),
.A2(n_981),
.B(n_1007),
.C(n_997),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1101),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1109),
.Y(n_1273)
);

AOI221xp5_ASAP7_75t_L g1274 ( 
.A1(n_1155),
.A2(n_649),
.B1(n_589),
.B2(n_1158),
.C(n_961),
.Y(n_1274)
);

NAND2x1p5_ASAP7_75t_L g1275 ( 
.A(n_1134),
.B(n_1054),
.Y(n_1275)
);

AOI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1168),
.A2(n_915),
.B1(n_847),
.B2(n_369),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1092),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1154),
.A2(n_1158),
.B1(n_889),
.B2(n_1155),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1065),
.A2(n_1098),
.B(n_1161),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1101),
.B(n_1072),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_L g1281 ( 
.A(n_1165),
.B(n_589),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1101),
.Y(n_1282)
);

NAND2x1p5_ASAP7_75t_L g1283 ( 
.A(n_1134),
.B(n_1054),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1158),
.A2(n_1171),
.A3(n_1089),
.B(n_1065),
.Y(n_1284)
);

BUFx2_ASAP7_75t_L g1285 ( 
.A(n_1147),
.Y(n_1285)
);

OAI22xp5_ASAP7_75t_L g1286 ( 
.A1(n_1168),
.A2(n_649),
.B1(n_847),
.B2(n_915),
.Y(n_1286)
);

OR2x2_ASAP7_75t_L g1287 ( 
.A(n_1153),
.B(n_1157),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1100),
.Y(n_1288)
);

NOR2xp33_ASAP7_75t_SL g1289 ( 
.A(n_1170),
.B(n_518),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1109),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_1158),
.A2(n_649),
.B(n_1154),
.C(n_1007),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1109),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1168),
.A2(n_649),
.B1(n_847),
.B2(n_915),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1068),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1154),
.A2(n_1158),
.B1(n_889),
.B2(n_1155),
.Y(n_1295)
);

BUFx10_ASAP7_75t_L g1296 ( 
.A(n_1107),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1215),
.B(n_1281),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1281),
.A2(n_1295),
.B1(n_1278),
.B2(n_1269),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1269),
.A2(n_1295),
.B1(n_1278),
.B2(n_1192),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1239),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1195),
.B(n_1268),
.Y(n_1301)
);

O2A1O1Ixp33_ASAP7_75t_L g1302 ( 
.A1(n_1266),
.A2(n_1267),
.B(n_1293),
.C(n_1286),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1215),
.B(n_1209),
.Y(n_1303)
);

O2A1O1Ixp33_ASAP7_75t_L g1304 ( 
.A1(n_1270),
.A2(n_1291),
.B(n_1274),
.C(n_1225),
.Y(n_1304)
);

BUFx4_ASAP7_75t_R g1305 ( 
.A(n_1249),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1280),
.B(n_1272),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1198),
.B(n_1287),
.Y(n_1307)
);

CKINVDCx6p67_ASAP7_75t_R g1308 ( 
.A(n_1230),
.Y(n_1308)
);

O2A1O1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1270),
.A2(n_1291),
.B(n_1225),
.C(n_1200),
.Y(n_1309)
);

BUFx8_ASAP7_75t_SL g1310 ( 
.A(n_1230),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1253),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1282),
.B(n_1199),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1200),
.A2(n_1206),
.B(n_1208),
.C(n_1271),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_L g1314 ( 
.A1(n_1206),
.A2(n_1271),
.B(n_1264),
.C(n_1201),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1224),
.B(n_1235),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1192),
.A2(n_1276),
.B1(n_1197),
.B2(n_1224),
.Y(n_1316)
);

NOR2xp67_ASAP7_75t_L g1317 ( 
.A(n_1221),
.B(n_1204),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1258),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1220),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1234),
.A2(n_1222),
.B(n_1236),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1252),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1201),
.A2(n_1237),
.B(n_1250),
.C(n_1233),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1204),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1197),
.A2(n_1263),
.B(n_1279),
.C(n_1260),
.Y(n_1324)
);

O2A1O1Ixp33_ASAP7_75t_L g1325 ( 
.A1(n_1197),
.A2(n_1279),
.B(n_1263),
.C(n_1242),
.Y(n_1325)
);

AOI21x1_ASAP7_75t_SL g1326 ( 
.A1(n_1255),
.A2(n_1277),
.B(n_1203),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1229),
.Y(n_1327)
);

AOI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1203),
.A2(n_1277),
.B(n_1251),
.Y(n_1328)
);

AOI21x1_ASAP7_75t_SL g1329 ( 
.A1(n_1213),
.A2(n_1223),
.B(n_1249),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1216),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1219),
.A2(n_1248),
.B1(n_1232),
.B2(n_1238),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1253),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1219),
.A2(n_1248),
.B1(n_1238),
.B2(n_1243),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1261),
.B(n_1211),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1205),
.A2(n_1216),
.B(n_1212),
.Y(n_1335)
);

NOR2xp67_ASAP7_75t_L g1336 ( 
.A(n_1245),
.B(n_1196),
.Y(n_1336)
);

AOI21x1_ASAP7_75t_SL g1337 ( 
.A1(n_1214),
.A2(n_1229),
.B(n_1243),
.Y(n_1337)
);

O2A1O1Ixp33_ASAP7_75t_L g1338 ( 
.A1(n_1226),
.A2(n_1240),
.B(n_1231),
.C(n_1227),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1289),
.Y(n_1339)
);

O2A1O1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1244),
.A2(n_1218),
.B(n_1294),
.C(n_1217),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_SL g1341 ( 
.A1(n_1228),
.A2(n_1241),
.B(n_1296),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1275),
.A2(n_1283),
.B(n_1205),
.Y(n_1342)
);

AOI22xp5_ASAP7_75t_L g1343 ( 
.A1(n_1207),
.A2(n_1285),
.B1(n_1210),
.B2(n_1259),
.Y(n_1343)
);

INVx3_ASAP7_75t_SL g1344 ( 
.A(n_1296),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1246),
.B(n_1247),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1258),
.B(n_1256),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1256),
.B(n_1288),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_1288),
.Y(n_1348)
);

O2A1O1Ixp33_ASAP7_75t_L g1349 ( 
.A1(n_1262),
.A2(n_1259),
.B(n_1193),
.C(n_1292),
.Y(n_1349)
);

BUFx2_ASAP7_75t_L g1350 ( 
.A(n_1288),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1257),
.B(n_1284),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1288),
.B(n_1257),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_R g1353 ( 
.A(n_1273),
.B(n_1290),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1284),
.B(n_1254),
.Y(n_1354)
);

O2A1O1Ixp5_ASAP7_75t_L g1355 ( 
.A1(n_1266),
.A2(n_1281),
.B(n_1200),
.C(n_1158),
.Y(n_1355)
);

AOI21x1_ASAP7_75t_SL g1356 ( 
.A1(n_1198),
.A2(n_786),
.B(n_897),
.Y(n_1356)
);

O2A1O1Ixp33_ASAP7_75t_L g1357 ( 
.A1(n_1281),
.A2(n_1266),
.B(n_1171),
.C(n_1267),
.Y(n_1357)
);

OAI211xp5_ASAP7_75t_L g1358 ( 
.A1(n_1281),
.A2(n_536),
.B(n_1192),
.C(n_589),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1270),
.A2(n_1291),
.B(n_1171),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1253),
.Y(n_1360)
);

O2A1O1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1281),
.A2(n_1266),
.B(n_1171),
.C(n_1267),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1287),
.B(n_1199),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1195),
.Y(n_1363)
);

O2A1O1Ixp5_ASAP7_75t_L g1364 ( 
.A1(n_1266),
.A2(n_1281),
.B(n_1200),
.C(n_1158),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1204),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1266),
.A2(n_1265),
.B(n_1194),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1195),
.B(n_1268),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1195),
.B(n_1268),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1207),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1239),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1195),
.B(n_1268),
.Y(n_1371)
);

A2O1A1Ixp33_ASAP7_75t_L g1372 ( 
.A1(n_1281),
.A2(n_1291),
.B(n_1270),
.C(n_1154),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_L g1373 ( 
.A1(n_1281),
.A2(n_1266),
.B(n_1171),
.C(n_1267),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1195),
.B(n_1268),
.Y(n_1374)
);

O2A1O1Ixp5_ASAP7_75t_L g1375 ( 
.A1(n_1266),
.A2(n_1281),
.B(n_1200),
.C(n_1158),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_SL g1376 ( 
.A1(n_1281),
.A2(n_862),
.B1(n_1276),
.B2(n_536),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1321),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1300),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1334),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1315),
.B(n_1303),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1351),
.B(n_1352),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1334),
.Y(n_1382)
);

AO21x2_ASAP7_75t_L g1383 ( 
.A1(n_1366),
.A2(n_1330),
.B(n_1335),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1334),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1370),
.B(n_1297),
.Y(n_1385)
);

INVxp67_ASAP7_75t_L g1386 ( 
.A(n_1319),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1320),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1298),
.A2(n_1299),
.B1(n_1376),
.B2(n_1316),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1354),
.Y(n_1389)
);

HB1xp67_ASAP7_75t_L g1390 ( 
.A(n_1311),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1332),
.B(n_1360),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1320),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1307),
.B(n_1372),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1320),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1345),
.Y(n_1395)
);

INVxp33_ASAP7_75t_L g1396 ( 
.A(n_1312),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1333),
.A2(n_1306),
.B1(n_1363),
.B2(n_1362),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1342),
.A2(n_1324),
.B(n_1325),
.Y(n_1398)
);

HB1xp67_ASAP7_75t_L g1399 ( 
.A(n_1347),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1338),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1369),
.A2(n_1358),
.B1(n_1374),
.B2(n_1301),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1357),
.A2(n_1373),
.B(n_1361),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1372),
.B(n_1313),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1346),
.B(n_1359),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1326),
.A2(n_1341),
.B(n_1342),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1355),
.A2(n_1375),
.B(n_1364),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1367),
.A2(n_1371),
.B1(n_1368),
.B2(n_1327),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1340),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1349),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1309),
.B(n_1304),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1314),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_1350),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1302),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1322),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1331),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1328),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1353),
.Y(n_1417)
);

HB1xp67_ASAP7_75t_L g1418 ( 
.A(n_1353),
.Y(n_1418)
);

AOI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1388),
.A2(n_1410),
.B1(n_1402),
.B2(n_1403),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1377),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1391),
.B(n_1343),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1381),
.B(n_1318),
.Y(n_1422)
);

OAI211xp5_ASAP7_75t_L g1423 ( 
.A1(n_1388),
.A2(n_1336),
.B(n_1339),
.C(n_1317),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1382),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1387),
.Y(n_1425)
);

HB1xp67_ASAP7_75t_L g1426 ( 
.A(n_1390),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1385),
.B(n_1344),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1395),
.B(n_1344),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1412),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1387),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1382),
.B(n_1308),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1405),
.B(n_1348),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1382),
.B(n_1308),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1387),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1385),
.B(n_1365),
.Y(n_1435)
);

BUFx2_ASAP7_75t_L g1436 ( 
.A(n_1382),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1378),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1410),
.A2(n_1327),
.B1(n_1310),
.B2(n_1323),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1382),
.B(n_1337),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1403),
.A2(n_1365),
.B1(n_1323),
.B2(n_1305),
.Y(n_1440)
);

INVx3_ASAP7_75t_SL g1441 ( 
.A(n_1391),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1391),
.B(n_1399),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1399),
.B(n_1356),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1384),
.B(n_1329),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1378),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1442),
.Y(n_1446)
);

OAI211xp5_ASAP7_75t_L g1447 ( 
.A1(n_1419),
.A2(n_1402),
.B(n_1410),
.C(n_1413),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1422),
.B(n_1379),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1425),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1419),
.A2(n_1401),
.B1(n_1414),
.B2(n_1413),
.Y(n_1450)
);

OAI211xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1427),
.A2(n_1413),
.B(n_1380),
.C(n_1407),
.Y(n_1451)
);

NOR5xp2_ASAP7_75t_SL g1452 ( 
.A(n_1440),
.B(n_1400),
.C(n_1414),
.D(n_1406),
.E(n_1310),
.Y(n_1452)
);

BUFx3_ASAP7_75t_L g1453 ( 
.A(n_1428),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_1435),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1421),
.A2(n_1415),
.B1(n_1404),
.B2(n_1414),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1425),
.Y(n_1456)
);

AOI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1423),
.A2(n_1400),
.B(n_1406),
.Y(n_1457)
);

AND2x4_ASAP7_75t_L g1458 ( 
.A(n_1424),
.B(n_1379),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1420),
.Y(n_1459)
);

OAI322xp33_ASAP7_75t_L g1460 ( 
.A1(n_1440),
.A2(n_1393),
.A3(n_1380),
.B1(n_1411),
.B2(n_1415),
.C1(n_1408),
.C2(n_1386),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1425),
.A2(n_1394),
.B(n_1392),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1430),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1428),
.Y(n_1463)
);

INVx2_ASAP7_75t_SL g1464 ( 
.A(n_1442),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1421),
.A2(n_1415),
.B1(n_1404),
.B2(n_1401),
.Y(n_1465)
);

NAND3xp33_ASAP7_75t_L g1466 ( 
.A(n_1423),
.B(n_1408),
.C(n_1411),
.Y(n_1466)
);

OAI211xp5_ASAP7_75t_L g1467 ( 
.A1(n_1427),
.A2(n_1397),
.B(n_1393),
.C(n_1407),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1422),
.B(n_1379),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_1429),
.Y(n_1469)
);

AOI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1435),
.A2(n_1408),
.B1(n_1411),
.B2(n_1396),
.C(n_1409),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1443),
.A2(n_1396),
.B1(n_1409),
.B2(n_1397),
.C(n_1386),
.Y(n_1471)
);

NAND3xp33_ASAP7_75t_L g1472 ( 
.A(n_1443),
.B(n_1406),
.C(n_1409),
.Y(n_1472)
);

OAI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1443),
.A2(n_1406),
.B(n_1405),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1384),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1429),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1421),
.A2(n_1418),
.B1(n_1417),
.B2(n_1406),
.Y(n_1476)
);

AOI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1430),
.A2(n_1394),
.B(n_1416),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1426),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1431),
.A2(n_1404),
.B1(n_1406),
.B2(n_1433),
.Y(n_1479)
);

INVxp67_ASAP7_75t_L g1480 ( 
.A(n_1428),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1441),
.B(n_1384),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1434),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1437),
.B(n_1389),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1431),
.A2(n_1433),
.B1(n_1439),
.B2(n_1444),
.Y(n_1484)
);

NOR3xp33_ASAP7_75t_SL g1485 ( 
.A(n_1447),
.B(n_1416),
.C(n_1438),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1459),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1453),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1478),
.Y(n_1488)
);

BUFx2_ASAP7_75t_L g1489 ( 
.A(n_1458),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1458),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1459),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1449),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1469),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1472),
.A2(n_1394),
.B(n_1383),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1483),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1451),
.B(n_1438),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1446),
.Y(n_1497)
);

BUFx3_ASAP7_75t_L g1498 ( 
.A(n_1453),
.Y(n_1498)
);

INVxp67_ASAP7_75t_L g1499 ( 
.A(n_1483),
.Y(n_1499)
);

OR2x6_ASAP7_75t_L g1500 ( 
.A(n_1457),
.B(n_1432),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1453),
.B(n_1436),
.Y(n_1501)
);

INVx4_ASAP7_75t_SL g1502 ( 
.A(n_1463),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1463),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1473),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1456),
.Y(n_1505)
);

INVx3_ASAP7_75t_L g1506 ( 
.A(n_1461),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1463),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1481),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1446),
.B(n_1437),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_SL g1510 ( 
.A(n_1470),
.B(n_1466),
.C(n_1471),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1477),
.A2(n_1456),
.B(n_1482),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1499),
.B(n_1464),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1502),
.B(n_1432),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1486),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1486),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1496),
.B(n_1475),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1488),
.B(n_1464),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1486),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1488),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1502),
.B(n_1480),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1499),
.B(n_1455),
.Y(n_1521)
);

BUFx3_ASAP7_75t_L g1522 ( 
.A(n_1507),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1493),
.B(n_1454),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1495),
.B(n_1462),
.Y(n_1524)
);

NOR3xp33_ASAP7_75t_SL g1525 ( 
.A(n_1510),
.B(n_1460),
.C(n_1467),
.Y(n_1525)
);

AND2x2_ASAP7_75t_SL g1526 ( 
.A(n_1504),
.B(n_1465),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1511),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1511),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1511),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_R g1530 ( 
.A(n_1493),
.B(n_1417),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1491),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1491),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1502),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1509),
.B(n_1474),
.Y(n_1534)
);

AND2x4_ASAP7_75t_SL g1535 ( 
.A(n_1485),
.B(n_1418),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1497),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1502),
.B(n_1432),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1502),
.B(n_1448),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1491),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1502),
.B(n_1448),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1497),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1507),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1495),
.B(n_1462),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1502),
.B(n_1468),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1509),
.B(n_1474),
.Y(n_1545)
);

AOI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1510),
.A2(n_1450),
.B1(n_1398),
.B2(n_1460),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1492),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1511),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1511),
.Y(n_1549)
);

NAND2xp67_ASAP7_75t_L g1550 ( 
.A(n_1501),
.B(n_1431),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1511),
.Y(n_1551)
);

OAI33xp33_ASAP7_75t_L g1552 ( 
.A1(n_1492),
.A2(n_1476),
.A3(n_1450),
.B1(n_1466),
.B2(n_1445),
.B3(n_1416),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1492),
.Y(n_1553)
);

NOR2xp67_ASAP7_75t_L g1554 ( 
.A(n_1538),
.B(n_1490),
.Y(n_1554)
);

OR2x6_ASAP7_75t_L g1555 ( 
.A(n_1533),
.B(n_1500),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_1530),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1525),
.B(n_1516),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1521),
.B(n_1519),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1533),
.B(n_1507),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1538),
.B(n_1487),
.Y(n_1560)
);

AND2x2_ASAP7_75t_SL g1561 ( 
.A(n_1526),
.B(n_1496),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1514),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1514),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1521),
.B(n_1503),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1522),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1526),
.B(n_1546),
.Y(n_1566)
);

NAND2xp33_ASAP7_75t_SL g1567 ( 
.A(n_1535),
.B(n_1485),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1526),
.B(n_1504),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1542),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1540),
.B(n_1487),
.Y(n_1570)
);

HB1xp67_ASAP7_75t_L g1571 ( 
.A(n_1536),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1515),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1535),
.B(n_1504),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1515),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1522),
.B(n_1487),
.Y(n_1575)
);

AOI32xp33_ASAP7_75t_L g1576 ( 
.A1(n_1535),
.A2(n_1503),
.A3(n_1487),
.B1(n_1498),
.B2(n_1489),
.Y(n_1576)
);

O2A1O1Ixp5_ASAP7_75t_L g1577 ( 
.A1(n_1552),
.A2(n_1501),
.B(n_1506),
.C(n_1505),
.Y(n_1577)
);

OAI21xp33_ASAP7_75t_L g1578 ( 
.A1(n_1550),
.A2(n_1500),
.B(n_1479),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1534),
.B(n_1508),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1550),
.B(n_1508),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1540),
.B(n_1498),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1523),
.B(n_1508),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1522),
.Y(n_1583)
);

AOI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1544),
.A2(n_1500),
.B1(n_1398),
.B2(n_1444),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1518),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1544),
.B(n_1498),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1541),
.B(n_1512),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1513),
.B(n_1498),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1561),
.A2(n_1500),
.B1(n_1513),
.B2(n_1537),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1561),
.A2(n_1557),
.B1(n_1566),
.B2(n_1567),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_L g1591 ( 
.A(n_1565),
.B(n_1517),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1556),
.B(n_1512),
.Y(n_1592)
);

INVxp67_ASAP7_75t_L g1593 ( 
.A(n_1571),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1558),
.B(n_1517),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1569),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1582),
.B(n_1520),
.Y(n_1596)
);

AND3x2_ASAP7_75t_L g1597 ( 
.A(n_1569),
.B(n_1520),
.C(n_1513),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1571),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1562),
.Y(n_1599)
);

INVx3_ASAP7_75t_L g1600 ( 
.A(n_1559),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1554),
.B(n_1513),
.Y(n_1601)
);

HB1xp67_ASAP7_75t_L g1602 ( 
.A(n_1583),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1581),
.B(n_1537),
.Y(n_1603)
);

AOI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1567),
.A2(n_1500),
.B1(n_1537),
.B2(n_1398),
.Y(n_1604)
);

AND3x1_ASAP7_75t_L g1605 ( 
.A(n_1568),
.B(n_1484),
.C(n_1501),
.Y(n_1605)
);

AOI22x1_ASAP7_75t_L g1606 ( 
.A1(n_1583),
.A2(n_1537),
.B1(n_1489),
.B2(n_1452),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1565),
.B(n_1587),
.Y(n_1607)
);

NAND2xp33_ASAP7_75t_L g1608 ( 
.A(n_1576),
.B(n_1433),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1581),
.B(n_1489),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_L g1610 ( 
.A(n_1564),
.B(n_1534),
.Y(n_1610)
);

AOI22xp33_ASAP7_75t_L g1611 ( 
.A1(n_1578),
.A2(n_1500),
.B1(n_1398),
.B2(n_1490),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1586),
.B(n_1490),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1559),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1594),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1605),
.A2(n_1577),
.B1(n_1573),
.B2(n_1580),
.C(n_1584),
.Y(n_1615)
);

AOI22xp33_ASAP7_75t_SL g1616 ( 
.A1(n_1606),
.A2(n_1586),
.B1(n_1560),
.B2(n_1570),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1590),
.A2(n_1575),
.B(n_1559),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1595),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1594),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1600),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1595),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1597),
.Y(n_1622)
);

OAI31xp33_ASAP7_75t_L g1623 ( 
.A1(n_1604),
.A2(n_1588),
.A3(n_1575),
.B(n_1579),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1607),
.B(n_1545),
.Y(n_1624)
);

AOI32xp33_ASAP7_75t_L g1625 ( 
.A1(n_1605),
.A2(n_1588),
.A3(n_1575),
.B1(n_1585),
.B2(n_1574),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1606),
.A2(n_1500),
.B(n_1555),
.Y(n_1626)
);

AOI21xp33_ASAP7_75t_L g1627 ( 
.A1(n_1593),
.A2(n_1572),
.B(n_1563),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1518),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1591),
.Y(n_1629)
);

INVx2_ASAP7_75t_SL g1630 ( 
.A(n_1600),
.Y(n_1630)
);

AND3x2_ASAP7_75t_L g1631 ( 
.A(n_1602),
.B(n_1532),
.C(n_1531),
.Y(n_1631)
);

AOI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1608),
.A2(n_1524),
.B1(n_1543),
.B2(n_1494),
.C(n_1532),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1614),
.B(n_1619),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1629),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_1630),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1622),
.B(n_1613),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_SL g1637 ( 
.A(n_1624),
.B(n_1613),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1617),
.B(n_1592),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1620),
.B(n_1598),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1625),
.B(n_1600),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1618),
.B(n_1600),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1621),
.B(n_1596),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1628),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1638),
.A2(n_1616),
.B1(n_1615),
.B2(n_1611),
.Y(n_1644)
);

NOR3xp33_ASAP7_75t_L g1645 ( 
.A(n_1633),
.B(n_1627),
.C(n_1626),
.Y(n_1645)
);

OAI31xp33_ASAP7_75t_L g1646 ( 
.A1(n_1637),
.A2(n_1623),
.A3(n_1627),
.B(n_1610),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1640),
.A2(n_1591),
.B(n_1632),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_L g1648 ( 
.A(n_1636),
.B(n_1628),
.C(n_1599),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_SL g1649 ( 
.A1(n_1634),
.A2(n_1601),
.B1(n_1555),
.B2(n_1599),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1641),
.Y(n_1650)
);

NOR5xp2_ASAP7_75t_L g1651 ( 
.A(n_1643),
.B(n_1631),
.C(n_1539),
.D(n_1531),
.E(n_1547),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1635),
.A2(n_1603),
.B1(n_1589),
.B2(n_1612),
.Y(n_1652)
);

AOI211xp5_ASAP7_75t_SL g1653 ( 
.A1(n_1639),
.A2(n_1603),
.B(n_1612),
.C(n_1609),
.Y(n_1653)
);

OAI21xp33_ASAP7_75t_L g1654 ( 
.A1(n_1642),
.A2(n_1609),
.B(n_1601),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1650),
.Y(n_1655)
);

OAI22xp5_ASAP7_75t_L g1656 ( 
.A1(n_1644),
.A2(n_1555),
.B1(n_1601),
.B2(n_1490),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1649),
.B(n_1601),
.Y(n_1657)
);

AOI22x1_ASAP7_75t_L g1658 ( 
.A1(n_1647),
.A2(n_1529),
.B1(n_1551),
.B2(n_1549),
.Y(n_1658)
);

A2O1A1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1646),
.A2(n_1527),
.B(n_1551),
.C(n_1549),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1657),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1655),
.B(n_1653),
.Y(n_1661)
);

AOI21xp5_ASAP7_75t_L g1662 ( 
.A1(n_1659),
.A2(n_1645),
.B(n_1648),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1658),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1656),
.B(n_1654),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1657),
.Y(n_1665)
);

NOR2x1_ASAP7_75t_L g1666 ( 
.A(n_1660),
.B(n_1651),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1665),
.B(n_1652),
.Y(n_1667)
);

AO22x2_ASAP7_75t_L g1668 ( 
.A1(n_1662),
.A2(n_1539),
.B1(n_1553),
.B2(n_1547),
.Y(n_1668)
);

CKINVDCx14_ASAP7_75t_R g1669 ( 
.A(n_1661),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1663),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_L g1671 ( 
.A(n_1666),
.B(n_1664),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1670),
.Y(n_1672)
);

INVxp33_ASAP7_75t_L g1673 ( 
.A(n_1667),
.Y(n_1673)
);

NOR3xp33_ASAP7_75t_L g1674 ( 
.A(n_1671),
.B(n_1669),
.C(n_1672),
.Y(n_1674)
);

NOR2x1_ASAP7_75t_L g1675 ( 
.A(n_1674),
.B(n_1662),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1675),
.Y(n_1676)
);

AO22x1_ASAP7_75t_L g1677 ( 
.A1(n_1676),
.A2(n_1673),
.B1(n_1668),
.B2(n_1490),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1677),
.Y(n_1678)
);

OAI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1528),
.B(n_1551),
.Y(n_1679)
);

OA21x2_ASAP7_75t_L g1680 ( 
.A1(n_1678),
.A2(n_1528),
.B(n_1549),
.Y(n_1680)
);

AOI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1548),
.B(n_1529),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1679),
.Y(n_1682)
);

NOR2xp67_ASAP7_75t_L g1683 ( 
.A(n_1682),
.B(n_1553),
.Y(n_1683)
);

OA21x2_ASAP7_75t_L g1684 ( 
.A1(n_1681),
.A2(n_1548),
.B(n_1529),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1548),
.B1(n_1528),
.B2(n_1527),
.Y(n_1685)
);

AOI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1685),
.A2(n_1684),
.B1(n_1527),
.B2(n_1543),
.Y(n_1686)
);

AOI211xp5_ASAP7_75t_L g1687 ( 
.A1(n_1686),
.A2(n_1524),
.B(n_1545),
.C(n_1505),
.Y(n_1687)
);


endmodule