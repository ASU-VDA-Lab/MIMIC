module real_jpeg_6934_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_131;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_120;
wire n_113;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_148;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_9;
wire n_137;
wire n_129;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_74;
wire n_70;
wire n_32;
wire n_20;
wire n_80;
wire n_30;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_1),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_2),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_2),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_2),
.A2(n_45),
.B1(n_51),
.B2(n_54),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_2),
.B(n_65),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_2),
.A2(n_45),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

O2A1O1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_2),
.A2(n_104),
.B(n_106),
.C(n_107),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_2),
.B(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_2),
.B(n_132),
.C(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_2),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_2),
.B(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_4),
.Y(n_145)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_7),
.Y(n_92)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_7),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_117),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_115),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_110),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_11),
.B(n_110),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_73),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_14),
.B1(n_46),
.B2(n_47),
.Y(n_12)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_13),
.A2(n_75),
.B(n_111),
.C(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_13),
.B(n_75),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_13),
.A2(n_14),
.B1(n_74),
.B2(n_75),
.Y(n_123)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

AO21x2_ASAP7_75t_SL g14 ( 
.A1(n_15),
.A2(n_29),
.B(n_41),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_29),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_16)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

OA22x2_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_35),
.B2(n_38),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_30),
.A2(n_33),
.B(n_45),
.Y(n_106)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_63),
.B2(n_64),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_48),
.A2(n_49),
.B1(n_103),
.B2(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_48),
.B(n_74),
.C(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_48),
.B(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_48),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_49),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_49),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_56),
.Y(n_49)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AO22x1_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_101),
.B2(n_102),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_74),
.A2(n_75),
.B1(n_120),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_74),
.A2(n_75),
.B1(n_129),
.B2(n_130),
.Y(n_150)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_129),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_82),
.Y(n_75)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_78),
.Y(n_134)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_93),
.Y(n_82)
);

NAND2x1_ASAP7_75t_SL g93 ( 
.A(n_83),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_83),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B1(n_88),
.B2(n_92),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_84),
.B(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_100),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_103),
.Y(n_112)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_111),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_126),
.B(n_152),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_138),
.B(n_151),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_135),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_135),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_131),
.B(n_134),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_149),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);


endmodule