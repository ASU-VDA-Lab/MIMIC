module real_jpeg_11328_n_12 (n_5, n_4, n_8, n_0, n_251, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_251;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_244;
wire n_167;
wire n_179;
wire n_128;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_9),
.B(n_25),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g82 ( 
.A(n_3),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_58),
.Y(n_53)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_5),
.A2(n_40),
.B(n_53),
.C(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_40),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_5),
.A2(n_9),
.B(n_55),
.Y(n_134)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_11),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_8),
.A2(n_20),
.B1(n_40),
.B2(n_42),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_8),
.A2(n_20),
.B1(n_54),
.B2(n_55),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_11),
.B1(n_21),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_29),
.B1(n_40),
.B2(n_42),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_9),
.A2(n_29),
.B1(n_54),
.B2(n_55),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_9),
.B(n_73),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_9),
.A2(n_24),
.B(n_39),
.C(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_9),
.B(n_22),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_10),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_10),
.A2(n_37),
.B1(n_54),
.B2(n_55),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_11),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_23),
.B(n_26),
.C(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_26),
.Y(n_31)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_26),
.B(n_29),
.C(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_115),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_113),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_92),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_15),
.B(n_92),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_74),
.B1(n_75),
.B2(n_91),
.Y(n_15)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_16),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_65),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_32),
.B1(n_33),
.B2(n_64),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_18),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_18),
.A2(n_64),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_18),
.B(n_106),
.C(n_185),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_18),
.A2(n_64),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_18),
.B(n_216),
.C(n_218),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_22),
.B(n_27),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_19),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_23),
.B(n_30),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_23),
.A2(n_28),
.B1(n_30),
.B2(n_105),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_24),
.A2(n_38),
.B(n_39),
.C(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_24),
.B(n_39),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_28),
.Y(n_89)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_29),
.A2(n_42),
.B(n_58),
.C(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_29),
.B(n_81),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_29),
.B(n_53),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_SL g163 ( 
.A1(n_29),
.A2(n_40),
.B(n_43),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_49),
.B1(n_50),
.B2(n_63),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_34),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_38),
.B(n_44),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_39),
.Y(n_43)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_45),
.A2(n_70),
.B(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_47),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_46),
.B(n_220),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_61),
.Y(n_50)
);

INVxp33_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_52),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_59),
.B1(n_61),
.B2(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_67),
.B(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_59),
.B1(n_87),
.B2(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_54),
.B(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_65),
.A2(n_66),
.B(n_68),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_68),
.A2(n_69),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_68),
.A2(n_69),
.B1(n_103),
.B2(n_104),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_69),
.B(n_123),
.C(n_174),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_69),
.B(n_103),
.C(n_208),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_71),
.B(n_73),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_83),
.B(n_88),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_76),
.A2(n_88),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_76),
.A2(n_84),
.B1(n_111),
.B2(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_78),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_78),
.B(n_127),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_82),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_80),
.A2(n_81),
.B1(n_125),
.B2(n_127),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_81),
.A2(n_203),
.B(n_204),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_82),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_83),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_84),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_86),
.A2(n_130),
.B(n_131),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_87),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_107),
.C(n_108),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_93),
.A2(n_94),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_103),
.C(n_106),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_95),
.A2(n_96),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_97),
.A2(n_100),
.B1(n_101),
.B2(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_97),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_98),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_100),
.A2(n_101),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_100),
.A2(n_101),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_143),
.C(n_151),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_101),
.B(n_170),
.C(n_177),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_103),
.A2(n_104),
.B1(n_106),
.B2(n_160),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_106),
.A2(n_129),
.B1(n_135),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_106),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_106),
.B(n_129),
.C(n_165),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_106),
.A2(n_160),
.B1(n_185),
.B2(n_187),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_107),
.A2(n_108),
.B1(n_109),
.B2(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_107),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AOI321xp33_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_225),
.A3(n_238),
.B1(n_244),
.B2(n_249),
.C(n_251),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_197),
.C(n_222),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_179),
.B(n_196),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_167),
.B(n_178),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_155),
.B(n_166),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_146),
.B(n_154),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_136),
.B(n_145),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_128),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_138),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_133),
.B2(n_135),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_129),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_129),
.B(n_133),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_129),
.A2(n_135),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_135),
.B(n_202),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_141),
.B(n_144),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_142),
.B(n_143),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_143),
.A2(n_149),
.B1(n_150),
.B2(n_153),
.Y(n_148)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_143),
.A2(n_153),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_143),
.B(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_147),
.B(n_148),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_156),
.B(n_157),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_161),
.B2(n_165),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_161),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_164),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_168),
.B(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_176),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_181),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_189),
.C(n_195),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_189),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_193),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_198),
.A2(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_209),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_199),
.B(n_209),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_205),
.CI(n_206),
.CON(n_199),
.SN(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_221),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_215),
.C(n_221),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_224),
.Y(n_246)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_226),
.A2(n_245),
.B(n_248),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_228),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_235),
.C(n_237),
.Y(n_239)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);


endmodule