module fake_jpeg_30821_n_104 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx8_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_43),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_38),
.B1(n_44),
.B2(n_39),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_14),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_52),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_53),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_36),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_0),
.Y(n_69)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_35),
.B1(n_40),
.B2(n_3),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

NAND3xp33_ASAP7_75t_L g67 ( 
.A(n_58),
.B(n_16),
.C(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_61),
.A2(n_35),
.B1(n_2),
.B2(n_4),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_54),
.B1(n_64),
.B2(n_7),
.Y(n_83)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_4),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_72),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_35),
.C(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

OR2x4_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_5),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

NOR2x1_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_6),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_77),
.B(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_67),
.Y(n_78)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_82),
.B(n_84),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_75),
.A2(n_8),
.B(n_54),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_77),
.C(n_66),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_91),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_25),
.C(n_9),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_84),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_96),
.C(n_86),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_88),
.B(n_86),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_90),
.B(n_68),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_83),
.B(n_8),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_10),
.B(n_11),
.Y(n_102)
);

OAI321xp33_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_13),
.A3(n_17),
.B1(n_22),
.B2(n_27),
.C(n_29),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_30),
.Y(n_104)
);


endmodule