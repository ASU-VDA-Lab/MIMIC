module fake_jpeg_30770_n_103 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_103);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_27),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_45),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_2),
.Y(n_60)
);

AOI21xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_0),
.B(n_1),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_53),
.B1(n_3),
.B2(n_4),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_38),
.B1(n_34),
.B2(n_42),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_54),
.B(n_60),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_47),
.A2(n_39),
.B(n_3),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_59),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_41),
.C(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_62),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_44),
.Y(n_62)
);

AOI32xp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_32),
.A3(n_39),
.B1(n_17),
.B2(n_19),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_7),
.B(n_11),
.C(n_12),
.Y(n_85)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

NOR2x1_ASAP7_75t_L g65 ( 
.A(n_58),
.B(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_65),
.B(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_4),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_71),
.B(n_73),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_6),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_18),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_58),
.A2(n_20),
.B1(n_30),
.B2(n_9),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_70),
.B(n_6),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_84),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_23),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_85),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_69),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_24),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_86),
.A2(n_68),
.B1(n_77),
.B2(n_65),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_92),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_88),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_87),
.C(n_83),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_98),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_81),
.C(n_79),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_95),
.B(n_97),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_91),
.B(n_94),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_85),
.B1(n_89),
.B2(n_15),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_26),
.Y(n_103)
);


endmodule