module real_aes_5761_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_153;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_150;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_649;
wire n_193;
wire n_293;
wire n_162;
wire n_397;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_646;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g287 ( .A(n_0), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_1), .B(n_302), .Y(n_420) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_2), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g421 ( .A(n_2), .B(n_422), .Y(n_421) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_3), .A2(n_28), .B1(n_301), .B2(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g174 ( .A1(n_4), .A2(n_8), .B1(n_175), .B2(n_177), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g341 ( .A1(n_5), .A2(n_31), .B1(n_276), .B2(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_6), .A2(n_49), .B1(n_250), .B2(n_253), .Y(n_266) );
HB1xp67_ASAP7_75t_L g651 ( .A(n_6), .Y(n_651) );
INVx1_ASAP7_75t_L g282 ( .A(n_7), .Y(n_282) );
INVx1_ASAP7_75t_L g107 ( .A(n_9), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_9), .B(n_58), .Y(n_126) );
INVxp67_ASAP7_75t_L g146 ( .A(n_9), .Y(n_146) );
INVx1_ASAP7_75t_L g285 ( .A(n_10), .Y(n_285) );
AOI21xp33_ASAP7_75t_SL g110 ( .A1(n_11), .A2(n_111), .B(n_117), .Y(n_110) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_12), .A2(n_53), .B(n_246), .Y(n_245) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_12), .A2(n_53), .B(n_246), .Y(n_261) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_13), .B(n_92), .Y(n_103) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_14), .A2(n_51), .B1(n_250), .B2(n_253), .Y(n_249) );
INVx1_ASAP7_75t_L g275 ( .A(n_15), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_16), .A2(n_60), .B1(n_136), .B2(n_138), .Y(n_135) );
BUFx3_ASAP7_75t_L g205 ( .A(n_17), .Y(n_205) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_18), .Y(n_80) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_19), .Y(n_92) );
AO22x1_ASAP7_75t_L g415 ( .A1(n_20), .A2(n_62), .B1(n_288), .B2(n_416), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_21), .Y(n_305) );
AND2x2_ASAP7_75t_L g319 ( .A(n_22), .B(n_276), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_23), .B(n_288), .Y(n_311) );
AOI22x1_ASAP7_75t_L g348 ( .A1(n_24), .A2(n_75), .B1(n_250), .B2(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_25), .B(n_57), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_26), .B(n_351), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g164 ( .A1(n_27), .A2(n_29), .B1(n_165), .B2(n_170), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_30), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_32), .B(n_385), .Y(n_384) );
HB1xp67_ASAP7_75t_L g197 ( .A(n_33), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_34), .B(n_280), .Y(n_310) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_35), .A2(n_37), .B1(n_158), .B2(n_162), .Y(n_157) );
INVx1_ASAP7_75t_L g246 ( .A(n_36), .Y(n_246) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_38), .Y(n_216) );
AND2x4_ASAP7_75t_L g230 ( .A(n_38), .B(n_214), .Y(n_230) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_39), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_40), .A2(n_42), .B1(n_149), .B2(n_152), .Y(n_148) );
INVx2_ASAP7_75t_L g257 ( .A(n_41), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g84 ( .A(n_43), .B(n_85), .Y(n_84) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_44), .A2(n_59), .B1(n_301), .B2(n_349), .Y(n_362) );
CKINVDCx14_ASAP7_75t_R g424 ( .A(n_45), .Y(n_424) );
AND2x2_ASAP7_75t_L g325 ( .A(n_46), .B(n_288), .Y(n_325) );
OA22x2_ASAP7_75t_L g97 ( .A1(n_47), .A2(n_58), .B1(n_92), .B2(n_96), .Y(n_97) );
INVx1_ASAP7_75t_L g133 ( .A(n_47), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_48), .B(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_50), .B(n_378), .Y(n_377) );
NAND2x1p5_ASAP7_75t_L g329 ( .A(n_52), .B(n_259), .Y(n_329) );
INVx1_ASAP7_75t_L g118 ( .A(n_54), .Y(n_118) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_55), .A2(n_67), .B1(n_182), .B2(n_185), .Y(n_181) );
CKINVDCx14_ASAP7_75t_R g354 ( .A(n_56), .Y(n_354) );
INVx1_ASAP7_75t_L g109 ( .A(n_57), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_57), .B(n_130), .Y(n_129) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_57), .Y(n_208) );
OAI21xp33_ASAP7_75t_L g155 ( .A1(n_58), .A2(n_63), .B(n_147), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_61), .B(n_302), .Y(n_382) );
INVx1_ASAP7_75t_L g95 ( .A(n_63), .Y(n_95) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_63), .B(n_74), .Y(n_127) );
INVx1_ASAP7_75t_L g192 ( .A(n_64), .Y(n_192) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_65), .Y(n_193) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_66), .Y(n_224) );
BUFx5_ASAP7_75t_L g252 ( .A(n_66), .Y(n_252) );
INVx1_ASAP7_75t_L g345 ( .A(n_66), .Y(n_345) );
INVx2_ASAP7_75t_L g290 ( .A(n_68), .Y(n_290) );
NAND2xp33_ASAP7_75t_L g321 ( .A(n_69), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_SL g214 ( .A(n_70), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_71), .A2(n_81), .B1(n_188), .B2(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_71), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_72), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_73), .B(n_328), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_74), .B(n_102), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_76), .B(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_200), .B1(n_217), .B2(n_231), .C(n_649), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_189), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_187), .B2(n_188), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_80), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_81), .Y(n_188) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_81), .A2(n_188), .B1(n_651), .B2(n_652), .Y(n_650) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NOR4xp75_ASAP7_75t_L g82 ( .A(n_83), .B(n_134), .C(n_156), .D(n_173), .Y(n_82) );
NAND2xp5_ASAP7_75t_L g83 ( .A(n_84), .B(n_110), .Y(n_83) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_98), .Y(n_88) );
AND2x2_ASAP7_75t_L g137 ( .A(n_89), .B(n_116), .Y(n_137) );
AND2x2_ASAP7_75t_L g166 ( .A(n_89), .B(n_167), .Y(n_166) );
AND2x4_ASAP7_75t_L g183 ( .A(n_89), .B(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_97), .Y(n_89) );
INVx1_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g90 ( .A(n_91), .B(n_94), .Y(n_90) );
NAND2xp33_ASAP7_75t_L g91 ( .A(n_92), .B(n_93), .Y(n_91) );
INVx2_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx3_ASAP7_75t_L g102 ( .A(n_92), .Y(n_102) );
NAND2xp33_ASAP7_75t_L g108 ( .A(n_92), .B(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
INVx1_ASAP7_75t_L g147 ( .A(n_92), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_93), .B(n_133), .Y(n_132) );
INVxp67_ASAP7_75t_L g209 ( .A(n_93), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g94 ( .A(n_95), .B(n_96), .Y(n_94) );
OAI21xp5_ASAP7_75t_L g145 ( .A1(n_95), .A2(n_146), .B(n_147), .Y(n_145) );
AND2x2_ASAP7_75t_L g114 ( .A(n_97), .B(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g144 ( .A(n_97), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g161 ( .A(n_97), .Y(n_161) );
AND2x4_ASAP7_75t_L g151 ( .A(n_98), .B(n_114), .Y(n_151) );
AND2x4_ASAP7_75t_L g153 ( .A(n_98), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g163 ( .A(n_98), .B(n_160), .Y(n_163) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_104), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
AND2x4_ASAP7_75t_L g116 ( .A(n_100), .B(n_104), .Y(n_116) );
AND2x2_ASAP7_75t_L g141 ( .A(n_100), .B(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g167 ( .A(n_100), .B(n_168), .Y(n_167) );
OR2x2_ASAP7_75t_L g180 ( .A(n_100), .B(n_169), .Y(n_180) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_103), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_102), .B(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g130 ( .A(n_102), .Y(n_130) );
NAND3xp33_ASAP7_75t_L g128 ( .A(n_103), .B(n_129), .C(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g169 ( .A(n_105), .Y(n_169) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_116), .Y(n_113) );
AND2x4_ASAP7_75t_L g160 ( .A(n_115), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g159 ( .A(n_116), .B(n_160), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g117 ( .A(n_118), .B(n_119), .Y(n_117) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AO21x2_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_125), .B(n_128), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_124), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_130), .B(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g154 ( .A(n_131), .B(n_155), .Y(n_154) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_133), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_148), .Y(n_134) );
BUFx3_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx5_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_144), .Y(n_140) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_143), .Y(n_206) );
INVx2_ASAP7_75t_SL g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g172 ( .A(n_154), .B(n_167), .Y(n_172) );
AND2x4_ASAP7_75t_L g186 ( .A(n_154), .B(n_179), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g156 ( .A(n_157), .B(n_164), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x4_ASAP7_75t_L g176 ( .A(n_160), .B(n_167), .Y(n_176) );
AND2x4_ASAP7_75t_L g178 ( .A(n_160), .B(n_179), .Y(n_178) );
BUFx5_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx8_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_174), .B(n_181), .Y(n_173) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g184 ( .A(n_180), .Y(n_184) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
BUFx12f_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_191), .B1(n_194), .B2(n_199), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g190 ( .A(n_191), .Y(n_190) );
XNOR2xp5_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
INVx1_ASAP7_75t_L g199 ( .A(n_194), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B1(n_197), .B2(n_198), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_195), .Y(n_198) );
INVx1_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_202), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_203), .B(n_211), .Y(n_202) );
INVxp67_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g654 ( .A(n_204), .B(n_211), .Y(n_654) );
AOI211xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_206), .B(n_207), .C(n_210), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_212), .B(n_215), .Y(n_211) );
OR2x2_ASAP7_75t_L g658 ( .A(n_212), .B(n_216), .Y(n_658) );
INVx1_ASAP7_75t_L g661 ( .A(n_212), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_212), .B(n_215), .Y(n_662) );
HB1xp67_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
HB1xp67_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_229), .Y(n_218) );
OA21x2_ASAP7_75t_L g660 ( .A1(n_219), .A2(n_661), .B(n_662), .Y(n_660) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_225), .Y(n_219) );
CKINVDCx16_ASAP7_75t_R g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g280 ( .A(n_223), .Y(n_280) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx3_ASAP7_75t_L g255 ( .A(n_224), .Y(n_255) );
INVx6_ASAP7_75t_L g278 ( .A(n_224), .Y(n_278) );
INVx2_ASAP7_75t_L g308 ( .A(n_224), .Y(n_308) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_226), .B(n_304), .Y(n_303) );
OAI22x1_ASAP7_75t_L g340 ( .A1(n_226), .A2(n_341), .B1(n_346), .B2(n_348), .Y(n_340) );
INVx4_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_227), .A2(n_301), .B1(n_303), .B2(n_306), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_227), .B(n_360), .Y(n_359) );
AOI21xp5_ASAP7_75t_L g380 ( .A1(n_227), .A2(n_381), .B(n_382), .Y(n_380) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx4_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
INVx3_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_228), .B(n_275), .Y(n_274) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_228), .B(n_282), .Y(n_281) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_228), .Y(n_313) );
INVxp67_ASAP7_75t_L g323 ( .A(n_228), .Y(n_323) );
INVx1_ASAP7_75t_L g347 ( .A(n_228), .Y(n_347) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_229), .A2(n_300), .B(n_309), .Y(n_299) );
AO31x2_ASAP7_75t_L g339 ( .A1(n_229), .A2(n_340), .A3(n_350), .B(n_353), .Y(n_339) );
AO31x2_ASAP7_75t_L g394 ( .A1(n_229), .A2(n_340), .A3(n_350), .B(n_353), .Y(n_394) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx3_ASAP7_75t_L g248 ( .A(n_230), .Y(n_248) );
INVx1_ASAP7_75t_L g271 ( .A(n_230), .Y(n_271) );
INVx3_ASAP7_75t_L g361 ( .A(n_230), .Y(n_361) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_235), .B(n_523), .Y(n_234) );
NOR4xp75_ASAP7_75t_L g235 ( .A(n_236), .B(n_436), .C(n_454), .D(n_480), .Y(n_235) );
AO21x1_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_292), .B(n_400), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
HB1xp67_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_239), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g444 ( .A(n_239), .B(n_410), .Y(n_444) );
INVx2_ASAP7_75t_L g506 ( .A(n_239), .Y(n_506) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_267), .Y(n_239) );
INVx1_ASAP7_75t_L g371 ( .A(n_240), .Y(n_371) );
INVx1_ASAP7_75t_L g399 ( .A(n_240), .Y(n_399) );
AND2x2_ASAP7_75t_L g426 ( .A(n_240), .B(n_268), .Y(n_426) );
INVx1_ASAP7_75t_L g457 ( .A(n_240), .Y(n_457) );
INVx2_ASAP7_75t_L g489 ( .A(n_240), .Y(n_489) );
NOR2x1_ASAP7_75t_L g531 ( .A(n_240), .B(n_532), .Y(n_531) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_240), .Y(n_546) );
AND2x2_ASAP7_75t_L g595 ( .A(n_240), .B(n_375), .Y(n_595) );
OR2x6_ASAP7_75t_L g240 ( .A(n_241), .B(n_262), .Y(n_240) );
OAI21x1_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_249), .B(n_256), .Y(n_241) );
NAND3xp33_ASAP7_75t_SL g242 ( .A(n_243), .B(n_244), .C(n_247), .Y(n_242) );
NOR2xp33_ASAP7_75t_SL g284 ( .A(n_243), .B(n_285), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_243), .B(n_287), .Y(n_286) );
NAND3xp33_ASAP7_75t_L g263 ( .A(n_244), .B(n_247), .C(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g270 ( .A(n_244), .Y(n_270) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g352 ( .A(n_245), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_245), .B(n_361), .Y(n_360) );
AOI21xp33_ASAP7_75t_SL g332 ( .A1(n_247), .A2(n_333), .B(n_335), .Y(n_332) );
INVx2_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_248), .B(n_378), .Y(n_389) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g288 ( .A(n_252), .Y(n_288) );
INVx2_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
INVx2_ASAP7_75t_L g387 ( .A(n_252), .Y(n_387) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g366 ( .A(n_254), .Y(n_366) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g385 ( .A(n_255), .Y(n_385) );
INVx1_ASAP7_75t_L g422 ( .A(n_255), .Y(n_422) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g316 ( .A(n_258), .Y(n_316) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g334 ( .A(n_260), .Y(n_334) );
INVx4_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g291 ( .A(n_261), .Y(n_291) );
BUFx3_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx3_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g488 ( .A(n_267), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
OR2x2_ASAP7_75t_L g493 ( .A(n_268), .B(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g513 ( .A(n_268), .Y(n_513) );
INVx1_ASAP7_75t_L g532 ( .A(n_268), .Y(n_532) );
AND2x2_ASAP7_75t_L g594 ( .A(n_268), .B(n_459), .Y(n_594) );
INVxp67_ASAP7_75t_L g624 ( .A(n_268), .Y(n_624) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_289), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_270), .B(n_271), .Y(n_269) );
OR2x2_ASAP7_75t_L g412 ( .A(n_271), .B(n_316), .Y(n_412) );
NAND3xp33_ASAP7_75t_SL g272 ( .A(n_273), .B(n_279), .C(n_283), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g322 ( .A(n_278), .Y(n_322) );
INVx1_ASAP7_75t_L g328 ( .A(n_278), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AOI22xp5_ASAP7_75t_L g283 ( .A1(n_280), .A2(n_284), .B1(n_286), .B2(n_288), .Y(n_283) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx3_ASAP7_75t_L g378 ( .A(n_291), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_368), .B1(n_390), .B2(n_397), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_336), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g565 ( .A(n_296), .Y(n_565) );
OR2x2_ASAP7_75t_L g647 ( .A(n_296), .B(n_479), .Y(n_647) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g478 ( .A(n_297), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_317), .Y(n_297) );
AND2x2_ASAP7_75t_L g391 ( .A(n_298), .B(n_392), .Y(n_391) );
NAND2x1_ASAP7_75t_L g440 ( .A(n_298), .B(n_338), .Y(n_440) );
AND2x2_ASAP7_75t_L g575 ( .A(n_298), .B(n_357), .Y(n_575) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_314), .B(n_315), .Y(n_298) );
OA21x2_ASAP7_75t_L g406 ( .A1(n_299), .A2(n_314), .B(n_315), .Y(n_406) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_312), .Y(n_309) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_SL g331 ( .A(n_313), .Y(n_331) );
INVx1_ASAP7_75t_L g388 ( .A(n_313), .Y(n_388) );
INVx1_ASAP7_75t_L g414 ( .A(n_313), .Y(n_414) );
INVx3_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
AND2x2_ASAP7_75t_L g401 ( .A(n_317), .B(n_394), .Y(n_401) );
AND2x4_ASAP7_75t_L g429 ( .A(n_317), .B(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g548 ( .A(n_317), .B(n_394), .Y(n_548) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_324), .B(n_332), .Y(n_317) );
AO21x2_ASAP7_75t_L g396 ( .A1(n_318), .A2(n_324), .B(n_332), .Y(n_396) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_320), .B(n_323), .Y(n_318) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
OAI21x1_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_326), .B(n_330), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_329), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_329), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g335 ( .A(n_329), .Y(n_335) );
AOI21x1_ASAP7_75t_L g419 ( .A1(n_331), .A2(n_420), .B(n_421), .Y(n_419) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_356), .Y(n_336) );
INVx2_ASAP7_75t_L g431 ( .A(n_337), .Y(n_431) );
INVx1_ASAP7_75t_L g463 ( .A(n_337), .Y(n_463) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g453 ( .A(n_338), .B(n_396), .Y(n_453) );
INVx1_ASAP7_75t_L g467 ( .A(n_338), .Y(n_467) );
AND2x2_ASAP7_75t_L g607 ( .A(n_338), .B(n_407), .Y(n_607) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g418 ( .A(n_345), .Y(n_418) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_347), .B(n_360), .Y(n_364) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2xp67_ASAP7_75t_SL g353 ( .A(n_354), .B(n_355), .Y(n_353) );
OR2x2_ASAP7_75t_L g423 ( .A(n_355), .B(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g479 ( .A(n_356), .Y(n_479) );
OR2x2_ASAP7_75t_L g591 ( .A(n_356), .B(n_440), .Y(n_591) );
INVx2_ASAP7_75t_L g599 ( .A(n_356), .Y(n_599) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_363), .Y(n_357) );
NAND2x1p5_ASAP7_75t_L g392 ( .A(n_358), .B(n_363), .Y(n_392) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_367), .Y(n_363) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g514 ( .A(n_371), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g539 ( .A(n_373), .B(n_499), .Y(n_539) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g473 ( .A(n_374), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g410 ( .A(n_375), .B(n_411), .Y(n_410) );
INVx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g435 ( .A(n_376), .Y(n_435) );
AND2x2_ASAP7_75t_L g458 ( .A(n_376), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g470 ( .A(n_376), .B(n_411), .Y(n_470) );
AND2x4_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .Y(n_376) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_383), .B(n_389), .Y(n_379) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .B(n_388), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AND2x2_ASAP7_75t_L g495 ( .A(n_391), .B(n_439), .Y(n_495) );
INVx1_ASAP7_75t_L g608 ( .A(n_391), .Y(n_608) );
AND2x2_ASAP7_75t_L g640 ( .A(n_391), .B(n_467), .Y(n_640) );
INVx2_ASAP7_75t_L g407 ( .A(n_392), .Y(n_407) );
AND2x2_ASAP7_75t_L g450 ( .A(n_392), .B(n_405), .Y(n_450) );
INVx1_ASAP7_75t_L g500 ( .A(n_392), .Y(n_500) );
INVx1_ASAP7_75t_L g552 ( .A(n_392), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_392), .B(n_519), .Y(n_560) );
BUFx3_ASAP7_75t_L g447 ( .A(n_393), .Y(n_447) );
NOR2xp67_ASAP7_75t_L g567 ( .A(n_393), .B(n_449), .Y(n_567) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx1_ASAP7_75t_L g477 ( .A(n_394), .Y(n_477) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVxp67_ASAP7_75t_L g439 ( .A(n_396), .Y(n_439) );
INVx1_ASAP7_75t_L g519 ( .A(n_396), .Y(n_519) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g469 ( .A(n_398), .B(n_470), .Y(n_469) );
OR2x2_ASAP7_75t_L g472 ( .A(n_398), .B(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_398), .Y(n_501) );
OR2x2_ASAP7_75t_L g628 ( .A(n_398), .B(n_505), .Y(n_628) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AND2x2_ASAP7_75t_L g491 ( .A(n_399), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_399), .B(n_557), .Y(n_556) );
OAI32xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .A3(n_408), .B1(n_427), .B2(n_432), .Y(n_400) );
INVx2_ASAP7_75t_L g563 ( .A(n_401), .Y(n_563) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g590 ( .A(n_403), .Y(n_590) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g510 ( .A(n_404), .Y(n_510) );
OR2x2_ASAP7_75t_L g517 ( .A(n_404), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .Y(n_404) );
INVx1_ASAP7_75t_L g602 ( .A(n_405), .Y(n_602) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g430 ( .A(n_406), .Y(n_430) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_406), .Y(n_558) );
INVx1_ASAP7_75t_L g452 ( .A(n_407), .Y(n_452) );
INVx2_ASAP7_75t_L g442 ( .A(n_408), .Y(n_442) );
OR2x2_ASAP7_75t_L g408 ( .A(n_409), .B(n_425), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x4_ASAP7_75t_L g530 ( .A(n_410), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g617 ( .A(n_410), .B(n_488), .Y(n_617) );
INVx2_ASAP7_75t_SL g459 ( .A(n_411), .Y(n_459) );
OAI21x1_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B(n_423), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g494 ( .A1(n_412), .A2(n_413), .B(n_423), .Y(n_494) );
AOI21x1_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B(n_419), .Y(n_413) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g566 ( .A(n_426), .B(n_470), .Y(n_566) );
NAND2x1_ASAP7_75t_SL g588 ( .A(n_426), .B(n_458), .Y(n_588) );
AND2x2_ASAP7_75t_L g597 ( .A(n_426), .B(n_486), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_426), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x2_ASAP7_75t_L g641 ( .A(n_428), .B(n_499), .Y(n_641) );
AND2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_431), .Y(n_428) );
AND2x4_ASAP7_75t_SL g466 ( .A(n_429), .B(n_467), .Y(n_466) );
BUFx3_ASAP7_75t_L g542 ( .A(n_429), .Y(n_542) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_430), .Y(n_535) );
INVx1_ASAP7_75t_L g568 ( .A(n_432), .Y(n_568) );
AOI211xp5_ASAP7_75t_SL g555 ( .A1(n_433), .A2(n_467), .B(n_556), .C(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
AND2x2_ASAP7_75t_L g512 ( .A(n_434), .B(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g570 ( .A(n_434), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g637 ( .A(n_434), .B(n_488), .Y(n_637) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g521 ( .A(n_435), .B(n_457), .Y(n_521) );
OR2x2_ASAP7_75t_L g536 ( .A(n_435), .B(n_493), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_435), .B(n_624), .Y(n_623) );
OAI22xp5_ASAP7_75t_SL g436 ( .A1(n_437), .A2(n_441), .B1(n_443), .B2(n_445), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_439), .Y(n_534) );
AND3x2_ASAP7_75t_L g614 ( .A(n_439), .B(n_599), .C(n_602), .Y(n_614) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_446), .A2(n_448), .B(n_451), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g633 ( .A(n_448), .Y(n_633) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g464 ( .A(n_450), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
BUFx3_ASAP7_75t_L g528 ( .A(n_453), .Y(n_528) );
AND2x2_ASAP7_75t_L g598 ( .A(n_453), .B(n_599), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_460), .B(n_468), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
AND2x2_ASAP7_75t_L g578 ( .A(n_458), .B(n_488), .Y(n_578) );
INVx2_ASAP7_75t_L g586 ( .A(n_458), .Y(n_586) );
INVx1_ASAP7_75t_L g474 ( .A(n_459), .Y(n_474) );
INVx1_ASAP7_75t_L g503 ( .A(n_459), .Y(n_503) );
INVxp67_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_462), .B(n_465), .Y(n_461) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_462), .A2(n_483), .B1(n_498), .B2(n_504), .Y(n_497) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
OR2x2_ASAP7_75t_L g573 ( .A(n_463), .B(n_574), .Y(n_573) );
INVx2_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g483 ( .A(n_466), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_471), .B(n_475), .Y(n_468) );
INVx2_ASAP7_75t_L g505 ( .A(n_470), .Y(n_505) );
AND2x2_ASAP7_75t_L g550 ( .A(n_470), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g600 ( .A1(n_472), .A2(n_573), .B1(n_601), .B2(n_603), .Y(n_600) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_474), .Y(n_486) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_476), .B(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_476), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND3x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_496), .C(n_507), .Y(n_480) );
AOI21x1_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B(n_490), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_485), .A2(n_570), .B1(n_647), .B2(n_648), .Y(n_646) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_487), .Y(n_485) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .Y(n_490) );
INVx1_ASAP7_75t_L g540 ( .A(n_492), .Y(n_540) );
AND2x2_ASAP7_75t_L g620 ( .A(n_492), .B(n_546), .Y(n_620) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g522 ( .A(n_493), .Y(n_522) );
BUFx2_ASAP7_75t_L g515 ( .A(n_494), .Y(n_515) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND3xp33_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .C(n_502), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g554 ( .A(n_503), .B(n_513), .Y(n_554) );
OR2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVxp67_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_511), .B1(n_516), .B2(n_520), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND3xp33_ASAP7_75t_SL g562 ( .A(n_509), .B(n_563), .C(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
AND2x2_ASAP7_75t_L g622 ( .A(n_514), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_514), .B(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g557 ( .A(n_515), .Y(n_557) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_518), .B(n_552), .Y(n_648) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_519), .A2(n_544), .B1(n_545), .B2(n_547), .Y(n_543) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
NAND2x2_ASAP7_75t_L g631 ( .A(n_521), .B(n_632), .Y(n_631) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_609), .Y(n_523) );
NAND4xp25_ASAP7_75t_L g524 ( .A(n_525), .B(n_561), .C(n_576), .D(n_596), .Y(n_524) );
NOR2xp67_ASAP7_75t_L g525 ( .A(n_526), .B(n_537), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_529), .B1(n_533), .B2(n_536), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_529), .A2(n_541), .B(n_619), .Y(n_618) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g571 ( .A(n_531), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
OAI211xp5_ASAP7_75t_SL g553 ( .A1(n_535), .A2(n_554), .B(n_555), .C(n_559), .Y(n_553) );
INVx1_ASAP7_75t_L g580 ( .A(n_535), .Y(n_580) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_536), .A2(n_606), .B(n_608), .Y(n_605) );
OAI321xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_540), .A3(n_541), .B1(n_543), .B2(n_549), .C(n_553), .Y(n_537) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g603 ( .A(n_540), .B(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_542), .B(n_583), .Y(n_582) );
NOR2x1_ASAP7_75t_R g625 ( .A(n_542), .B(n_606), .Y(n_625) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g626 ( .A(n_547), .B(n_575), .Y(n_626) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g601 ( .A(n_548), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g613 ( .A(n_548), .Y(n_613) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g583 ( .A(n_552), .Y(n_583) );
INVxp67_ASAP7_75t_L g639 ( .A(n_557), .Y(n_639) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI222xp33_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_566), .B1(n_567), .B2(n_568), .C1(n_569), .C2(n_572), .Y(n_561) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g630 ( .A(n_565), .Y(n_630) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g585 ( .A(n_571), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI221x1_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_579), .B1(n_581), .B2(n_584), .C(n_587), .Y(n_576) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
OAI22xp33_ASAP7_75t_SL g587 ( .A1(n_588), .A2(n_589), .B1(n_591), .B2(n_592), .Y(n_587) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
BUFx3_ASAP7_75t_L g632 ( .A(n_594), .Y(n_632) );
INVx2_ASAP7_75t_L g604 ( .A(n_595), .Y(n_604) );
AOI211xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_600), .C(n_605), .Y(n_596) );
NAND2x1_ASAP7_75t_L g612 ( .A(n_599), .B(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_SL g629 ( .A1(n_603), .A2(n_630), .B1(n_631), .B2(n_633), .Y(n_629) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND3xp33_ASAP7_75t_SL g609 ( .A(n_610), .B(n_621), .C(n_634), .Y(n_609) );
O2A1O1Ixp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_614), .B(n_615), .C(n_618), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_625), .B1(n_626), .B2(n_627), .C(n_629), .Y(n_621) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_624), .Y(n_645) );
INVxp67_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_640), .B1(n_641), .B2(n_642), .C(n_646), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI222xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_653), .B2(n_655), .C1(n_657), .C2(n_659), .Y(n_649) );
CKINVDCx5p33_ASAP7_75t_R g652 ( .A(n_651), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
BUFx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
endmodule