module fake_ariane_1241_n_1795 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1795);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1795;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_131),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_158),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_59),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_148),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_89),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_94),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_19),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_97),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_117),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_86),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_26),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_112),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_3),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_92),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_121),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_35),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_22),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_65),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_75),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_118),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_80),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_27),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_143),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_141),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_77),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_52),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_129),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_14),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_103),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_38),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_21),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_30),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_22),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_23),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_38),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_18),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_64),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_98),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_50),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_144),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_57),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_76),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_145),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_165),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_113),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_35),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_29),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_49),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_54),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_43),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_26),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_160),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_4),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_14),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_47),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_154),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_9),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_153),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_58),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_107),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_56),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_11),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_72),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_87),
.Y(n_241)
);

BUFx8_ASAP7_75t_SL g242 ( 
.A(n_17),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_136),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_19),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_69),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_104),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_119),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_130),
.Y(n_248)
);

BUFx2_ASAP7_75t_SL g249 ( 
.A(n_50),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_101),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_102),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_78),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_41),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_91),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_166),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_11),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_120),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_73),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_114),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_62),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_25),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_128),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_138),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_68),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_29),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_108),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_5),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_55),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_15),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_132),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_8),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_23),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_55),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_0),
.Y(n_278)
);

INVx2_ASAP7_75t_SL g279 ( 
.A(n_74),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_4),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_99),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_150),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_36),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_134),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g285 ( 
.A(n_25),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_18),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_13),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_51),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_95),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_81),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_147),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_36),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_116),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_0),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_51),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_24),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_111),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_96),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_17),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_164),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_60),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_133),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_39),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_67),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_28),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_46),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_110),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_70),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_31),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_32),
.Y(n_310)
);

INVx2_ASAP7_75t_SL g311 ( 
.A(n_20),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_84),
.Y(n_312)
);

INVxp67_ASAP7_75t_R g313 ( 
.A(n_15),
.Y(n_313)
);

BUFx2_ASAP7_75t_L g314 ( 
.A(n_32),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_168),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_10),
.Y(n_316)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_149),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_151),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_20),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_7),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_13),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_21),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_125),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_127),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_46),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_71),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_126),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_82),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_163),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_33),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_159),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_52),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_135),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_42),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_31),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_1),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_224),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_242),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_260),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_314),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_172),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_209),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_209),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_203),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_216),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_299),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_299),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_336),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_238),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_336),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_203),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_183),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_187),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_212),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_232),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_203),
.Y(n_357)
);

INVxp67_ASAP7_75t_SL g358 ( 
.A(n_203),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_238),
.Y(n_359)
);

BUFx6f_ASAP7_75t_SL g360 ( 
.A(n_238),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_208),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_186),
.B(n_1),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_235),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_281),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_289),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_215),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_223),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_300),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_226),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_281),
.Y(n_370)
);

INVxp67_ASAP7_75t_SL g371 ( 
.A(n_203),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_230),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_281),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_239),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_181),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_177),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_169),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_250),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_263),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_270),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_169),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_271),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_204),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_323),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_274),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_275),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_170),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_249),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_280),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_170),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_187),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_331),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_181),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_171),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_208),
.Y(n_396)
);

NOR2xp67_ASAP7_75t_L g397 ( 
.A(n_311),
.B(n_199),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_171),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_283),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_295),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_173),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_173),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_176),
.B(n_180),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_217),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_174),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_208),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_174),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_175),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_310),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_175),
.Y(n_410)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_210),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_210),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_199),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_210),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_254),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_254),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_345),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_391),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_404),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_345),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_352),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_352),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_393),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_393),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_417),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_375),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_360),
.B(n_229),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_190),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_418),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_388),
.B(n_324),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_375),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_403),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_353),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_355),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_361),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_348),
.B(n_193),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_367),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_369),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_372),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_374),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_286),
.Y(n_450)
);

AND2x2_ASAP7_75t_SL g451 ( 
.A(n_362),
.B(n_246),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_379),
.Y(n_453)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_360),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_382),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_343),
.B(n_286),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_385),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_386),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_389),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_341),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_377),
.B(n_198),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_399),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_400),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_344),
.B(n_195),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_409),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_413),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_377),
.B(n_198),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_347),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_349),
.B(n_246),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_351),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_397),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_395),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_381),
.B(n_279),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_337),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_360),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_354),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_350),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_387),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_387),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_350),
.B(n_197),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_411),
.B(n_296),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_390),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_390),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_359),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_359),
.B(n_296),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_416),
.B(n_335),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_440),
.B(n_364),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_479),
.B(n_340),
.Y(n_494)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_480),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_419),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_451),
.A2(n_433),
.B1(n_468),
.B2(n_462),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_419),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_419),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_398),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_454),
.Y(n_502)
);

NAND2xp33_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_401),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_423),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_423),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_480),
.B(n_401),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_480),
.B(n_402),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_SL g508 ( 
.A1(n_433),
.A2(n_451),
.B1(n_338),
.B2(n_406),
.Y(n_508)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_451),
.B(n_405),
.C(n_402),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_423),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_427),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_421),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_440),
.B(n_462),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_364),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_468),
.B(n_370),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_445),
.B(n_396),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_475),
.B(n_370),
.Y(n_517)
);

CKINVDCx6p67_ASAP7_75t_R g518 ( 
.A(n_443),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

INVxp67_ASAP7_75t_SL g520 ( 
.A(n_435),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_422),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_445),
.B(n_373),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_427),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_451),
.A2(n_335),
.B1(n_373),
.B2(n_326),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_476),
.A2(n_285),
.B1(n_412),
.B2(n_408),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_480),
.B(n_405),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_424),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_475),
.B(n_407),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_480),
.B(n_407),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_422),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_479),
.B(n_340),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_424),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_434),
.B(n_477),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_427),
.Y(n_535)
);

OR2x6_ASAP7_75t_L g536 ( 
.A(n_479),
.B(n_279),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_476),
.A2(n_410),
.B1(n_408),
.B2(n_306),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_427),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_434),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_426),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_439),
.A2(n_410),
.B1(n_322),
.B2(n_321),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_434),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_435),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_454),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_480),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_477),
.B(n_184),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_488),
.A2(n_188),
.B1(n_207),
.B2(n_206),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_420),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_426),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_422),
.Y(n_550)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_487),
.Y(n_551)
);

OR2x6_ASAP7_75t_L g552 ( 
.A(n_479),
.B(n_485),
.Y(n_552)
);

BUFx4f_ASAP7_75t_L g553 ( 
.A(n_487),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_485),
.B(n_188),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_422),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_485),
.B(n_189),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_426),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_485),
.B(n_342),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_427),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_430),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_428),
.Y(n_562)
);

AO22x1_ASAP7_75t_L g563 ( 
.A1(n_476),
.A2(n_332),
.B1(n_294),
.B2(n_194),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_477),
.B(n_220),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_428),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_428),
.Y(n_566)
);

AND3x1_ASAP7_75t_L g567 ( 
.A(n_478),
.B(n_313),
.C(n_244),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_487),
.B(n_178),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_428),
.Y(n_569)
);

NOR2x1p5_ASAP7_75t_L g570 ( 
.A(n_490),
.B(n_339),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_428),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_445),
.B(n_229),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_430),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_430),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_430),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_472),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_487),
.B(n_178),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_487),
.B(n_179),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_472),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_428),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_428),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_428),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_470),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_484),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_472),
.Y(n_585)
);

INVx3_ASAP7_75t_L g586 ( 
.A(n_429),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_429),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_472),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_477),
.B(n_319),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_429),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g591 ( 
.A(n_461),
.B(n_339),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_429),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_487),
.B(n_179),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_470),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_429),
.Y(n_595)
);

NOR3xp33_ASAP7_75t_L g596 ( 
.A(n_439),
.B(n_482),
.C(n_481),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_461),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_486),
.B(n_491),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_487),
.B(n_443),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_476),
.B(n_486),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_429),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_487),
.B(n_182),
.Y(n_602)
);

AND2x6_ASAP7_75t_L g603 ( 
.A(n_484),
.B(n_332),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_486),
.B(n_182),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_429),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_429),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_486),
.B(n_346),
.Y(n_607)
);

NAND3xp33_ASAP7_75t_L g608 ( 
.A(n_458),
.B(n_211),
.C(n_202),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_445),
.B(n_229),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_445),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_453),
.B(n_244),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_453),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_458),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_425),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_453),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_453),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_453),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_458),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_458),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_491),
.B(n_185),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_443),
.B(n_185),
.Y(n_621)
);

AO21x2_ASAP7_75t_L g622 ( 
.A1(n_483),
.A2(n_241),
.B(n_233),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_458),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_458),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_490),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_458),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_491),
.B(n_191),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_425),
.Y(n_628)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_478),
.B(n_189),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_491),
.B(n_356),
.Y(n_630)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_454),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_425),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_483),
.B(n_191),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_478),
.A2(n_244),
.B1(n_306),
.B2(n_258),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_425),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_458),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_481),
.B(n_363),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_460),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_488),
.A2(n_489),
.B1(n_482),
.B2(n_481),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_478),
.A2(n_306),
.B1(n_269),
.B2(n_292),
.Y(n_640)
);

NAND2xp33_ASAP7_75t_L g641 ( 
.A(n_513),
.B(n_482),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_521),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_548),
.B(n_488),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_521),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_584),
.B(n_490),
.Y(n_645)
);

O2A1O1Ixp5_ASAP7_75t_L g646 ( 
.A1(n_568),
.A2(n_489),
.B(n_437),
.C(n_456),
.Y(n_646)
);

INVxp33_ASAP7_75t_L g647 ( 
.A(n_548),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_530),
.Y(n_648)
);

NOR2xp67_ASAP7_75t_L g649 ( 
.A(n_597),
.B(n_443),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_497),
.B(n_490),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_497),
.B(n_489),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_520),
.B(n_443),
.Y(n_652)
);

BUFx5_ASAP7_75t_L g653 ( 
.A(n_545),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_583),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_493),
.B(n_443),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_563),
.B(n_437),
.C(n_421),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_594),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_591),
.B(n_474),
.Y(n_658)
);

BUFx3_ASAP7_75t_L g659 ( 
.A(n_594),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_570),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_495),
.A2(n_444),
.B(n_442),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_516),
.B(n_474),
.Y(n_662)
);

NOR2xp67_ASAP7_75t_L g663 ( 
.A(n_509),
.B(n_443),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_495),
.B(n_443),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_516),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_530),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_514),
.B(n_443),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_550),
.Y(n_668)
);

NOR3xp33_ASAP7_75t_L g669 ( 
.A(n_563),
.B(n_201),
.C(n_194),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_550),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_495),
.B(n_460),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_543),
.B(n_444),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_559),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_572),
.B(n_454),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_572),
.B(n_454),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_555),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_609),
.B(n_454),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_555),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_551),
.B(n_460),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_609),
.B(n_450),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_558),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_551),
.B(n_460),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_611),
.B(n_450),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_610),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_509),
.A2(n_492),
.B1(n_442),
.B2(n_441),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_528),
.B(n_450),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_611),
.B(n_474),
.Y(n_687)
);

OAI221xp5_ASAP7_75t_L g688 ( 
.A1(n_524),
.A2(n_470),
.B1(n_466),
.B2(n_464),
.C(n_446),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_515),
.B(n_474),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_598),
.B(n_522),
.Y(n_690)
);

INVx4_ASAP7_75t_L g691 ( 
.A(n_518),
.Y(n_691)
);

OAI22x1_ASAP7_75t_SL g692 ( 
.A1(n_512),
.A2(n_383),
.B1(n_384),
.B2(n_376),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_584),
.B(n_492),
.Y(n_693)
);

NOR2xp67_ASAP7_75t_L g694 ( 
.A(n_517),
.B(n_464),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_494),
.B(n_492),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_552),
.A2(n_492),
.B1(n_441),
.B2(n_456),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_539),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_522),
.B(n_492),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_610),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_612),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_531),
.B(n_492),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_600),
.B(n_441),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_512),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_554),
.B(n_442),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_625),
.B(n_466),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_612),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_551),
.B(n_460),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_559),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_615),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_553),
.B(n_460),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_554),
.B(n_556),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_554),
.B(n_446),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_496),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_554),
.B(n_446),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_556),
.B(n_447),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_556),
.B(n_447),
.Y(n_716)
);

NOR2xp67_ASAP7_75t_L g717 ( 
.A(n_591),
.B(n_447),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_496),
.Y(n_718)
);

INVx1_ASAP7_75t_SL g719 ( 
.A(n_629),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_603),
.A2(n_449),
.B1(n_452),
.B2(n_467),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_498),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_615),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_552),
.A2(n_456),
.B1(n_448),
.B2(n_459),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_556),
.B(n_448),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_639),
.B(n_448),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_553),
.B(n_460),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_639),
.B(n_459),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_616),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_633),
.B(n_459),
.Y(n_729)
);

OR2x2_ASAP7_75t_L g730 ( 
.A(n_629),
.B(n_473),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_607),
.B(n_365),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_616),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_539),
.B(n_463),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_559),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_542),
.B(n_463),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_604),
.B(n_463),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_603),
.A2(n_449),
.B1(n_452),
.B2(n_455),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_559),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_620),
.B(n_460),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_596),
.B(n_469),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_542),
.B(n_431),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_617),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_603),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_498),
.Y(n_744)
);

INVxp67_ASAP7_75t_SL g745 ( 
.A(n_559),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_630),
.B(n_368),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_603),
.B(n_431),
.Y(n_747)
);

BUFx6f_ASAP7_75t_L g748 ( 
.A(n_518),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_637),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_603),
.B(n_431),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_552),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_617),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_603),
.B(n_431),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_547),
.B(n_525),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_570),
.B(n_552),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_499),
.Y(n_756)
);

INVx2_ASAP7_75t_SL g757 ( 
.A(n_546),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_567),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_603),
.B(n_431),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_552),
.B(n_469),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_499),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_564),
.B(n_432),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_547),
.B(n_457),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_589),
.B(n_469),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_537),
.B(n_469),
.C(n_207),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_504),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_567),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_622),
.B(n_432),
.Y(n_768)
);

NOR2xp33_ASAP7_75t_L g769 ( 
.A(n_534),
.B(n_469),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_504),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_553),
.B(n_469),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_L g772 ( 
.A(n_506),
.B(n_469),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_541),
.B(n_457),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_505),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_622),
.B(n_432),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_505),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_613),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_507),
.B(n_469),
.Y(n_778)
);

OR2x6_ASAP7_75t_L g779 ( 
.A(n_536),
.B(n_457),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_622),
.B(n_432),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_510),
.Y(n_781)
);

INVx8_ASAP7_75t_L g782 ( 
.A(n_536),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_536),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_510),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_536),
.B(n_560),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_545),
.B(n_449),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_519),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_519),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_L g789 ( 
.A(n_526),
.B(n_471),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_599),
.A2(n_465),
.B(n_452),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_529),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_508),
.B(n_473),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_536),
.B(n_465),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_560),
.B(n_432),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_627),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_573),
.B(n_449),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_527),
.B(n_452),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_527),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_573),
.B(n_455),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_574),
.B(n_455),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_532),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_532),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_540),
.B(n_549),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_540),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_576),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_574),
.B(n_455),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_500),
.A2(n_467),
.B1(n_325),
.B2(n_192),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_545),
.B(n_467),
.Y(n_808)
);

NOR2x2_ASAP7_75t_L g809 ( 
.A(n_779),
.B(n_392),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_690),
.A2(n_503),
.B(n_577),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_681),
.B(n_749),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_686),
.B(n_634),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_652),
.A2(n_593),
.B(n_578),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_713),
.Y(n_814)
);

OAI321xp33_ASAP7_75t_L g815 ( 
.A1(n_651),
.A2(n_640),
.A3(n_473),
.B1(n_608),
.B2(n_436),
.C(n_579),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_671),
.A2(n_602),
.B(n_621),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_671),
.A2(n_544),
.B(n_502),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_718),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_721),
.Y(n_819)
);

NAND3xp33_ASAP7_75t_L g820 ( 
.A(n_651),
.B(n_557),
.C(n_549),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_643),
.B(n_436),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_658),
.Y(n_822)
);

O2A1O1Ixp5_ASAP7_75t_L g823 ( 
.A1(n_650),
.A2(n_557),
.B(n_575),
.C(n_588),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_744),
.B(n_502),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_719),
.B(n_436),
.Y(n_825)
);

AOI22x1_ASAP7_75t_L g826 ( 
.A1(n_766),
.A2(n_575),
.B1(n_636),
.B2(n_613),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_661),
.A2(n_619),
.B(n_618),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_686),
.B(n_579),
.Y(n_828)
);

OAI21xp5_ASAP7_75t_L g829 ( 
.A1(n_790),
.A2(n_803),
.B(n_769),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_679),
.A2(n_544),
.B(n_502),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_695),
.B(n_585),
.Y(n_831)
);

OR2x2_ASAP7_75t_L g832 ( 
.A(n_731),
.B(n_438),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_695),
.B(n_585),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_781),
.Y(n_834)
);

INVx5_ASAP7_75t_L g835 ( 
.A(n_748),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_679),
.A2(n_631),
.B(n_544),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_755),
.B(n_438),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_682),
.A2(n_631),
.B(n_619),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_701),
.B(n_588),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_701),
.B(n_438),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_665),
.B(n_757),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_689),
.B(n_438),
.Y(n_842)
);

OAI21xp5_ASAP7_75t_L g843 ( 
.A1(n_803),
.A2(n_769),
.B(n_739),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_744),
.B(n_751),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_689),
.B(n_501),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_682),
.A2(n_710),
.B(n_707),
.Y(n_846)
);

INVx3_ASAP7_75t_L g847 ( 
.A(n_751),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_672),
.B(n_501),
.Y(n_848)
);

CKINVDCx8_ASAP7_75t_R g849 ( 
.A(n_703),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_662),
.B(n_501),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_754),
.B(n_511),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_751),
.B(n_631),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_650),
.A2(n_638),
.B(n_618),
.C(n_623),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_801),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_680),
.B(n_511),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_729),
.A2(n_638),
.B(n_623),
.C(n_624),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_802),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_756),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_751),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_805),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_656),
.B(n_225),
.C(n_222),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_683),
.B(n_729),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_739),
.A2(n_626),
.B(n_624),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_687),
.B(n_511),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_707),
.A2(n_626),
.B(n_605),
.Y(n_865)
);

AOI21x1_ASAP7_75t_L g866 ( 
.A1(n_710),
.A2(n_605),
.B(n_562),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_726),
.A2(n_636),
.B(n_613),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_726),
.A2(n_562),
.B(n_561),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_771),
.A2(n_675),
.B(n_674),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_642),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_705),
.B(n_523),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_771),
.A2(n_636),
.B(n_533),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_761),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_770),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_677),
.A2(n_533),
.B(n_523),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_705),
.B(n_523),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_653),
.B(n_743),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_653),
.B(n_533),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_736),
.A2(n_565),
.B(n_561),
.Y(n_879)
);

BUFx2_ASAP7_75t_L g880 ( 
.A(n_746),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_702),
.A2(n_538),
.B(n_535),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_645),
.A2(n_538),
.B1(n_535),
.B2(n_586),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_655),
.A2(n_538),
.B(n_535),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_642),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_655),
.A2(n_586),
.B(n_566),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_698),
.B(n_566),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_774),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_667),
.A2(n_808),
.B(n_786),
.Y(n_888)
);

BUFx6f_ASAP7_75t_L g889 ( 
.A(n_748),
.Y(n_889)
);

AO21x1_ASAP7_75t_L g890 ( 
.A1(n_768),
.A2(n_569),
.B(n_565),
.Y(n_890)
);

NOR2xp33_ASAP7_75t_L g891 ( 
.A(n_758),
.B(n_586),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_676),
.Y(n_892)
);

AO21x2_ASAP7_75t_L g893 ( 
.A1(n_775),
.A2(n_608),
.B(n_571),
.Y(n_893)
);

AOI21x1_ASAP7_75t_L g894 ( 
.A1(n_786),
.A2(n_571),
.B(n_569),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_676),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_793),
.B(n_580),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_793),
.B(n_580),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_767),
.B(n_581),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_664),
.A2(n_582),
.B(n_581),
.Y(n_899)
);

AOI21x1_ASAP7_75t_L g900 ( 
.A1(n_808),
.A2(n_587),
.B(n_582),
.Y(n_900)
);

INVx4_ASAP7_75t_L g901 ( 
.A(n_782),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_725),
.B(n_587),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_667),
.A2(n_606),
.B(n_592),
.Y(n_903)
);

NOR2x1_ASAP7_75t_L g904 ( 
.A(n_717),
.B(n_590),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_763),
.B(n_206),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_647),
.B(n_294),
.Y(n_906)
);

AO21x1_ASAP7_75t_L g907 ( 
.A1(n_780),
.A2(n_590),
.B(n_592),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_653),
.B(n_595),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_727),
.B(n_595),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_693),
.B(n_601),
.Y(n_910)
);

AO21x1_ASAP7_75t_L g911 ( 
.A1(n_764),
.A2(n_601),
.B(n_606),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_647),
.B(n_614),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_644),
.Y(n_913)
);

OAI321xp33_ASAP7_75t_L g914 ( 
.A1(n_765),
.A2(n_290),
.A3(n_248),
.B1(n_253),
.B2(n_256),
.C(n_312),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_776),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_648),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_745),
.A2(n_635),
.B(n_632),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_664),
.A2(n_635),
.B(n_632),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_641),
.A2(n_736),
.B(n_794),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_748),
.Y(n_920)
);

AO21x1_ASAP7_75t_L g921 ( 
.A1(n_764),
.A2(n_264),
.B(n_259),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_697),
.B(n_628),
.Y(n_922)
);

INVx6_ASAP7_75t_L g923 ( 
.A(n_660),
.Y(n_923)
);

INVx11_ASAP7_75t_L g924 ( 
.A(n_692),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_773),
.B(n_303),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_653),
.B(n_628),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_741),
.A2(n_205),
.B(n_200),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_694),
.B(n_704),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_712),
.B(n_303),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_714),
.B(n_305),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_762),
.A2(n_205),
.B(n_200),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_715),
.B(n_305),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_716),
.B(n_309),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_733),
.A2(n_328),
.B(n_315),
.C(n_297),
.Y(n_934)
);

NOR2x1_ASAP7_75t_R g935 ( 
.A(n_660),
.B(n_309),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_691),
.Y(n_936)
);

OAI21xp33_ASAP7_75t_L g937 ( 
.A1(n_685),
.A2(n_320),
.B(n_321),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_784),
.Y(n_938)
);

INVx2_ASAP7_75t_L g939 ( 
.A(n_666),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_724),
.B(n_320),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_796),
.A2(n_196),
.B(n_251),
.Y(n_941)
);

O2A1O1Ixp33_ASAP7_75t_SL g942 ( 
.A1(n_787),
.A2(n_329),
.B(n_3),
.C(n_5),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_711),
.B(n_322),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_799),
.A2(n_196),
.B(n_251),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_800),
.A2(n_252),
.B(n_298),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_806),
.A2(n_252),
.B(n_298),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_668),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_735),
.B(n_227),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_691),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_646),
.A2(n_471),
.B(n_334),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_670),
.Y(n_951)
);

OAI21xp33_ASAP7_75t_L g952 ( 
.A1(n_788),
.A2(n_231),
.B(n_234),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_659),
.B(n_255),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_797),
.A2(n_301),
.B(n_302),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_778),
.A2(n_471),
.B(n_425),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_792),
.B(n_267),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_678),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_797),
.A2(n_772),
.B(n_699),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_659),
.B(n_276),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_653),
.B(n_301),
.Y(n_960)
);

AOI21xp33_ASAP7_75t_L g961 ( 
.A1(n_730),
.A2(n_288),
.B(n_277),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_696),
.B(n_278),
.Y(n_962)
);

INVx2_ASAP7_75t_SL g963 ( 
.A(n_660),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_798),
.Y(n_964)
);

OAI21xp5_ASAP7_75t_L g965 ( 
.A1(n_684),
.A2(n_471),
.B(n_325),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_700),
.A2(n_471),
.B(n_318),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_804),
.A2(n_287),
.B(n_6),
.C(n_7),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_706),
.A2(n_302),
.B(n_304),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_709),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_722),
.A2(n_471),
.B(n_304),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_728),
.A2(n_307),
.B(n_308),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_755),
.B(n_471),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_782),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_723),
.A2(n_307),
.B(n_334),
.C(n_330),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_732),
.Y(n_975)
);

INVx6_ASAP7_75t_L g976 ( 
.A(n_777),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_743),
.B(n_425),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_742),
.A2(n_308),
.B(n_318),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_752),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_653),
.B(n_327),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_748),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_740),
.A2(n_330),
.B(n_213),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_778),
.A2(n_261),
.B(n_218),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_669),
.A2(n_425),
.B(n_262),
.C(n_293),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_654),
.B(n_471),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_657),
.B(n_471),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_777),
.B(n_425),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_688),
.B(n_214),
.C(n_219),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_777),
.A2(n_257),
.B(n_291),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_795),
.B(n_471),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_791),
.B(n_2),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_783),
.B(n_284),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_880),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_811),
.B(n_782),
.Y(n_994)
);

BUFx3_ASAP7_75t_L g995 ( 
.A(n_849),
.Y(n_995)
);

BUFx6f_ASAP7_75t_L g996 ( 
.A(n_889),
.Y(n_996)
);

BUFx8_ASAP7_75t_L g997 ( 
.A(n_963),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_862),
.A2(n_737),
.B1(n_720),
.B2(n_779),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_812),
.A2(n_760),
.B(n_663),
.C(n_785),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_814),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_L g1001 ( 
.A1(n_956),
.A2(n_737),
.B1(n_720),
.B2(n_760),
.Y(n_1001)
);

AOI21xp33_ASAP7_75t_L g1002 ( 
.A1(n_956),
.A2(n_747),
.B(n_750),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_843),
.A2(n_738),
.B(n_673),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_811),
.B(n_649),
.Y(n_1004)
);

INVx8_ASAP7_75t_L g1005 ( 
.A(n_835),
.Y(n_1005)
);

NAND3xp33_ASAP7_75t_SL g1006 ( 
.A(n_861),
.B(n_967),
.C(n_988),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_988),
.A2(n_753),
.B(n_759),
.C(n_807),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_822),
.B(n_777),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_831),
.B(n_673),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_833),
.A2(n_738),
.B(n_734),
.Y(n_1010)
);

BUFx2_ASAP7_75t_L g1011 ( 
.A(n_822),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_961),
.A2(n_789),
.B(n_8),
.C(n_12),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_851),
.A2(n_738),
.B(n_734),
.C(n_708),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_905),
.B(n_738),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_925),
.B(n_734),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_906),
.B(n_734),
.Y(n_1016)
);

AOI22xp33_ASAP7_75t_L g1017 ( 
.A1(n_937),
.A2(n_991),
.B1(n_825),
.B2(n_819),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_818),
.Y(n_1018)
);

A2O1A1Ixp33_ASAP7_75t_L g1019 ( 
.A1(n_851),
.A2(n_708),
.B(n_673),
.C(n_282),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_835),
.B(n_708),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_834),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_820),
.A2(n_673),
.B(n_273),
.C(n_272),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_839),
.A2(n_243),
.B1(n_266),
.B2(n_265),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_991),
.B(n_2),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_SL g1025 ( 
.A1(n_824),
.A2(n_12),
.B(n_16),
.C(n_24),
.Y(n_1025)
);

OAI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_828),
.A2(n_268),
.B1(n_247),
.B2(n_245),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_898),
.A2(n_240),
.B(n_237),
.C(n_236),
.Y(n_1027)
);

NAND2xp33_ASAP7_75t_L g1028 ( 
.A(n_889),
.B(n_228),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_889),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_821),
.B(n_27),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_840),
.A2(n_221),
.B(n_79),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_841),
.B(n_30),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_858),
.B(n_33),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_889),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_845),
.A2(n_83),
.B(n_162),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_832),
.B(n_34),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_920),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_861),
.A2(n_34),
.B(n_37),
.C(n_39),
.Y(n_1038)
);

NAND2x1_ASAP7_75t_L g1039 ( 
.A(n_976),
.B(n_920),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_829),
.A2(n_85),
.B(n_156),
.Y(n_1040)
);

OAI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_873),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_1041)
);

AOI21x1_ASAP7_75t_L g1042 ( 
.A1(n_868),
.A2(n_88),
.B(n_152),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_920),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_837),
.B(n_40),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_837),
.B(n_42),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_874),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_919),
.A2(n_93),
.B(n_140),
.Y(n_1047)
);

CKINVDCx8_ASAP7_75t_R g1048 ( 
.A(n_835),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_958),
.A2(n_90),
.B(n_139),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_869),
.A2(n_842),
.B(n_848),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_848),
.A2(n_66),
.B(n_124),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_887),
.B(n_45),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_854),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_915),
.B(n_47),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_923),
.Y(n_1055)
);

O2A1O1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_974),
.A2(n_48),
.B(n_49),
.C(n_53),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_920),
.B(n_48),
.Y(n_1057)
);

OR2x6_ASAP7_75t_SL g1058 ( 
.A(n_953),
.B(n_53),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_894),
.A2(n_900),
.B(n_866),
.Y(n_1059)
);

NOR2xp67_ASAP7_75t_R g1060 ( 
.A(n_901),
.B(n_54),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_888),
.A2(n_61),
.B(n_63),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_938),
.B(n_100),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_964),
.A2(n_105),
.B1(n_106),
.B2(n_109),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_929),
.B(n_115),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_912),
.A2(n_167),
.B1(n_844),
.B2(n_898),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_857),
.A2(n_916),
.B1(n_913),
.B2(n_939),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_859),
.B(n_959),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_859),
.B(n_847),
.Y(n_1068)
);

O2A1O1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_974),
.A2(n_948),
.B(n_942),
.C(n_932),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_908),
.A2(n_926),
.B(n_885),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_942),
.A2(n_930),
.B(n_933),
.C(n_940),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_975),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_969),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_912),
.B(n_943),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_935),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_908),
.A2(n_926),
.B(n_883),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_847),
.B(n_891),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_SL g1078 ( 
.A(n_901),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_863),
.A2(n_846),
.B(n_903),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_960),
.A2(n_980),
.B(n_911),
.C(n_810),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_973),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_947),
.A2(n_951),
.B1(n_957),
.B2(n_979),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_879),
.A2(n_878),
.B(n_875),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_891),
.B(n_972),
.Y(n_1084)
);

OR2x6_ASAP7_75t_SL g1085 ( 
.A(n_962),
.B(n_924),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_934),
.A2(n_815),
.B(n_823),
.C(n_928),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_952),
.B(n_844),
.Y(n_1087)
);

AND2x6_ASAP7_75t_L g1088 ( 
.A(n_981),
.B(n_936),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_878),
.A2(n_830),
.B(n_836),
.Y(n_1089)
);

O2A1O1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_984),
.A2(n_856),
.B(n_871),
.C(n_876),
.Y(n_1090)
);

NOR3xp33_ASAP7_75t_SL g1091 ( 
.A(n_968),
.B(n_971),
.C(n_978),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_817),
.A2(n_824),
.B(n_881),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_992),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_864),
.A2(n_838),
.B(n_813),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_SL g1095 ( 
.A1(n_809),
.A2(n_936),
.B1(n_949),
.B2(n_981),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_981),
.Y(n_1096)
);

AOI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_949),
.A2(n_852),
.B1(n_877),
.B2(n_960),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_860),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_SL g1099 ( 
.A1(n_827),
.A2(n_950),
.B(n_931),
.C(n_927),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_976),
.B(n_990),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_SL g1101 ( 
.A(n_896),
.B(n_897),
.Y(n_1101)
);

CKINVDCx16_ASAP7_75t_R g1102 ( 
.A(n_809),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_870),
.Y(n_1103)
);

O2A1O1Ixp5_ASAP7_75t_L g1104 ( 
.A1(n_980),
.A2(n_921),
.B(n_816),
.C(n_856),
.Y(n_1104)
);

O2A1O1Ixp5_ASAP7_75t_L g1105 ( 
.A1(n_823),
.A2(n_955),
.B(n_984),
.C(n_852),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_914),
.A2(n_853),
.B(n_970),
.C(n_966),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_902),
.B(n_909),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_976),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_850),
.A2(n_855),
.B1(n_910),
.B2(n_886),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_954),
.B(n_884),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_892),
.B(n_895),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_SL g1112 ( 
.A(n_941),
.B(n_945),
.C(n_946),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_SL g1113 ( 
.A(n_982),
.B(n_983),
.C(n_944),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_882),
.B(n_977),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_918),
.A2(n_872),
.B(n_867),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_853),
.B(n_922),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_965),
.A2(n_826),
.B1(n_977),
.B2(n_904),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_985),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_893),
.B(n_989),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_893),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_865),
.A2(n_917),
.B(n_877),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_987),
.B(n_986),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_987),
.B(n_907),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_890),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_899),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_862),
.A2(n_651),
.B1(n_497),
.B2(n_831),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_811),
.B(n_681),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_843),
.A2(n_551),
.B(n_495),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_811),
.B(n_749),
.Y(n_1129)
);

HB1xp67_ASAP7_75t_L g1130 ( 
.A(n_822),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_R g1131 ( 
.A(n_849),
.B(n_703),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_814),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_889),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_822),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_862),
.B(n_651),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_814),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_880),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_812),
.A2(n_651),
.B(n_497),
.C(n_695),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_1131),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1121),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1141)
);

O2A1O1Ixp5_ASAP7_75t_L g1142 ( 
.A1(n_1104),
.A2(n_1106),
.B(n_1126),
.C(n_1080),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1126),
.A2(n_1135),
.B(n_1127),
.C(n_1138),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_1069),
.A2(n_1032),
.B(n_1071),
.C(n_1087),
.Y(n_1144)
);

OAI21xp5_ASAP7_75t_SL g1145 ( 
.A1(n_1024),
.A2(n_1046),
.B(n_1041),
.Y(n_1145)
);

BUFx12f_ASAP7_75t_L g1146 ( 
.A(n_997),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_998),
.A2(n_1006),
.B1(n_1084),
.B2(n_1001),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1128),
.A2(n_1050),
.B(n_1009),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1092),
.A2(n_1115),
.B(n_1094),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1048),
.Y(n_1150)
);

INVx3_ASAP7_75t_SL g1151 ( 
.A(n_995),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_993),
.Y(n_1152)
);

AO32x2_ASAP7_75t_L g1153 ( 
.A1(n_1109),
.A2(n_1046),
.A3(n_1041),
.B1(n_1095),
.B2(n_998),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1056),
.A2(n_1038),
.B1(n_1134),
.B2(n_1023),
.C(n_1026),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1120),
.A2(n_1124),
.A3(n_1109),
.B(n_1083),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1079),
.A2(n_1086),
.A3(n_1117),
.B(n_1013),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1070),
.A2(n_1076),
.B(n_1042),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1017),
.A2(n_1102),
.B1(n_1137),
.B2(n_1074),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_1003),
.A2(n_1010),
.B(n_1049),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1107),
.A2(n_1090),
.B(n_1101),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1005),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1011),
.B(n_1130),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1072),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_L g1164 ( 
.A(n_1096),
.B(n_1081),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1023),
.A2(n_1026),
.B(n_1099),
.C(n_1027),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1117),
.A2(n_1116),
.B(n_1007),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1137),
.B(n_1044),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_994),
.B(n_1067),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1105),
.A2(n_1123),
.B(n_1061),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_999),
.A2(n_1110),
.A3(n_1019),
.B(n_1062),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_SL g1171 ( 
.A1(n_1033),
.A2(n_1052),
.B(n_1097),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1008),
.B(n_1093),
.Y(n_1172)
);

INVx8_ASAP7_75t_L g1173 ( 
.A(n_1005),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_1075),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1000),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1018),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1047),
.A2(n_1031),
.B(n_1113),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1065),
.A2(n_1012),
.B(n_1002),
.C(n_1077),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1040),
.A2(n_1119),
.B(n_1035),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1021),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_1064),
.A2(n_1125),
.B(n_1051),
.Y(n_1181)
);

O2A1O1Ixp33_ASAP7_75t_L g1182 ( 
.A1(n_1004),
.A2(n_1025),
.B(n_1030),
.C(n_1033),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1114),
.A2(n_1062),
.B(n_1020),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_997),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1053),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1122),
.A2(n_1022),
.A3(n_1103),
.B(n_1111),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1132),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1014),
.A2(n_1063),
.B(n_1100),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1015),
.A2(n_1091),
.B(n_1052),
.C(n_1054),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1063),
.A2(n_1028),
.B(n_1020),
.Y(n_1190)
);

INVx1_ASAP7_75t_SL g1191 ( 
.A(n_1016),
.Y(n_1191)
);

BUFx10_ASAP7_75t_L g1192 ( 
.A(n_1078),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1136),
.Y(n_1193)
);

NOR2xp67_ASAP7_75t_SL g1194 ( 
.A(n_996),
.B(n_1133),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1045),
.B(n_1036),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1055),
.B(n_1068),
.Y(n_1196)
);

BUFx4_ASAP7_75t_SL g1197 ( 
.A(n_1108),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1098),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1096),
.A2(n_1112),
.A3(n_1118),
.B(n_1066),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1005),
.A2(n_1057),
.B(n_1039),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1060),
.A2(n_1088),
.B(n_1058),
.C(n_1034),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_SL g1202 ( 
.A1(n_1082),
.A2(n_1088),
.B(n_1078),
.Y(n_1202)
);

HB1xp67_ASAP7_75t_L g1203 ( 
.A(n_996),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_SL g1204 ( 
.A(n_1088),
.B(n_996),
.Y(n_1204)
);

NAND2xp33_ASAP7_75t_L g1205 ( 
.A(n_1088),
.B(n_1029),
.Y(n_1205)
);

OAI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1029),
.A2(n_1034),
.B(n_1037),
.Y(n_1206)
);

OAI22x1_ASAP7_75t_L g1207 ( 
.A1(n_1085),
.A2(n_1029),
.B1(n_1034),
.B2(n_1037),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1037),
.A2(n_1043),
.B(n_1133),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1043),
.A2(n_651),
.B(n_1135),
.C(n_497),
.Y(n_1209)
);

BUFx2_ASAP7_75t_R g1210 ( 
.A(n_1085),
.Y(n_1210)
);

AOI22x1_ASAP7_75t_L g1211 ( 
.A1(n_1050),
.A2(n_479),
.B1(n_486),
.B2(n_485),
.Y(n_1211)
);

AOI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1092),
.A2(n_1050),
.B(n_1079),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1121),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1072),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1073),
.Y(n_1218)
);

INVx2_ASAP7_75t_L g1219 ( 
.A(n_1073),
.Y(n_1219)
);

AOI31xp67_ASAP7_75t_L g1220 ( 
.A1(n_1123),
.A2(n_1065),
.A3(n_1101),
.B(n_1097),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1131),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1073),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1005),
.Y(n_1225)
);

NAND3x1_ASAP7_75t_L g1226 ( 
.A(n_1024),
.B(n_1032),
.C(n_656),
.Y(n_1226)
);

O2A1O1Ixp5_ASAP7_75t_L g1227 ( 
.A1(n_1104),
.A2(n_651),
.B(n_1106),
.C(n_1126),
.Y(n_1227)
);

AOI221xp5_ASAP7_75t_L g1228 ( 
.A1(n_1126),
.A2(n_754),
.B1(n_749),
.B2(n_637),
.C(n_651),
.Y(n_1228)
);

CKINVDCx6p67_ASAP7_75t_R g1229 ( 
.A(n_995),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1079),
.A2(n_1050),
.B(n_1115),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1121),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1232)
);

OAI21xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1024),
.A2(n_497),
.B(n_651),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1048),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1120),
.A2(n_890),
.A3(n_907),
.B(n_911),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_1135),
.B(n_1129),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1137),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1126),
.A2(n_651),
.B1(n_754),
.B2(n_1129),
.Y(n_1243)
);

AO32x2_ASAP7_75t_L g1244 ( 
.A1(n_1109),
.A2(n_1126),
.A3(n_1046),
.B1(n_1041),
.B2(n_1095),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1245)
);

OAI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1121),
.Y(n_1246)
);

OR2x2_ASAP7_75t_L g1247 ( 
.A(n_1127),
.B(n_1137),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1131),
.Y(n_1248)
);

CKINVDCx14_ASAP7_75t_R g1249 ( 
.A(n_1131),
.Y(n_1249)
);

AO31x2_ASAP7_75t_L g1250 ( 
.A1(n_1120),
.A2(n_890),
.A3(n_907),
.B(n_911),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1121),
.Y(n_1251)
);

AND2x6_ASAP7_75t_SL g1252 ( 
.A(n_1129),
.B(n_637),
.Y(n_1252)
);

AOI21xp33_ASAP7_75t_L g1253 ( 
.A1(n_1069),
.A2(n_749),
.B(n_956),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_993),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1085),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1073),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1120),
.A2(n_890),
.A3(n_907),
.B(n_911),
.Y(n_1261)
);

AO31x2_ASAP7_75t_L g1262 ( 
.A1(n_1120),
.A2(n_890),
.A3(n_907),
.B(n_911),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1072),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1024),
.A2(n_956),
.B1(n_342),
.B2(n_356),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1072),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1267)
);

AO21x1_ASAP7_75t_L g1268 ( 
.A1(n_1126),
.A2(n_651),
.B(n_1109),
.Y(n_1268)
);

CKINVDCx16_ASAP7_75t_R g1269 ( 
.A(n_1131),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1138),
.A2(n_1126),
.B(n_651),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1271)
);

NOR2xp67_ASAP7_75t_L g1272 ( 
.A(n_1096),
.B(n_835),
.Y(n_1272)
);

INVx2_ASAP7_75t_SL g1273 ( 
.A(n_997),
.Y(n_1273)
);

OA21x2_ASAP7_75t_L g1274 ( 
.A1(n_1079),
.A2(n_1050),
.B(n_1115),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1275)
);

AOI31xp67_ASAP7_75t_L g1276 ( 
.A1(n_1123),
.A2(n_1065),
.A3(n_1101),
.B(n_1097),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1135),
.A2(n_651),
.B(n_497),
.C(n_1138),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1072),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1121),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1129),
.B(n_811),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1089),
.A2(n_1059),
.B(n_1121),
.Y(n_1281)
);

OAI22x1_ASAP7_75t_L g1282 ( 
.A1(n_1024),
.A2(n_754),
.B1(n_512),
.B2(n_749),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1072),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1072),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1073),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1135),
.A2(n_1126),
.B1(n_497),
.B2(n_651),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_1073),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1129),
.B(n_1135),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1135),
.A2(n_551),
.B(n_495),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1146),
.Y(n_1292)
);

NAND2x1p5_ASAP7_75t_L g1293 ( 
.A(n_1242),
.B(n_1194),
.Y(n_1293)
);

INVx4_ASAP7_75t_L g1294 ( 
.A(n_1151),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1173),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1163),
.Y(n_1296)
);

INVx8_ASAP7_75t_L g1297 ( 
.A(n_1173),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1216),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1249),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1287),
.A2(n_1270),
.B1(n_1280),
.B2(n_1243),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1243),
.A2(n_1228),
.B1(n_1145),
.B2(n_1233),
.Y(n_1301)
);

INVxp67_ASAP7_75t_SL g1302 ( 
.A(n_1230),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1167),
.B(n_1141),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1263),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1139),
.Y(n_1305)
);

INVx6_ASAP7_75t_L g1306 ( 
.A(n_1173),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_SL g1307 ( 
.A1(n_1265),
.A2(n_1269),
.B1(n_1282),
.B2(n_1270),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1155),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1150),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1218),
.Y(n_1310)
);

CKINVDCx20_ASAP7_75t_R g1311 ( 
.A(n_1221),
.Y(n_1311)
);

CKINVDCx11_ASAP7_75t_R g1312 ( 
.A(n_1256),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1248),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1233),
.A2(n_1254),
.B1(n_1223),
.B2(n_1238),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1266),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1145),
.A2(n_1147),
.B1(n_1277),
.B2(n_1226),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_1229),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1225),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1278),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1283),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1219),
.Y(n_1321)
);

AO22x1_ASAP7_75t_L g1322 ( 
.A1(n_1215),
.A2(n_1240),
.B1(n_1257),
.B2(n_1236),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1222),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1285),
.Y(n_1324)
);

AOI22x1_ASAP7_75t_SL g1325 ( 
.A1(n_1184),
.A2(n_1152),
.B1(n_1210),
.B2(n_1234),
.Y(n_1325)
);

OAI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1147),
.A2(n_1290),
.B1(n_1284),
.B2(n_1289),
.Y(n_1326)
);

BUFx8_ASAP7_75t_L g1327 ( 
.A(n_1255),
.Y(n_1327)
);

OR2x2_ASAP7_75t_L g1328 ( 
.A(n_1247),
.B(n_1242),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_SL g1329 ( 
.A1(n_1195),
.A2(n_1244),
.B1(n_1153),
.B2(n_1252),
.Y(n_1329)
);

OAI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1144),
.A2(n_1154),
.B1(n_1143),
.B2(n_1209),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1207),
.A2(n_1172),
.B1(n_1252),
.B2(n_1168),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1225),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1174),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_SL g1334 ( 
.A1(n_1244),
.A2(n_1153),
.B1(n_1158),
.B2(n_1171),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1239),
.A2(n_1253),
.B1(n_1162),
.B2(n_1166),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1268),
.A2(n_1193),
.B1(n_1175),
.B2(n_1176),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1180),
.A2(n_1185),
.B1(n_1288),
.B2(n_1286),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1244),
.A2(n_1153),
.B1(n_1227),
.B2(n_1211),
.Y(n_1338)
);

INVx6_ASAP7_75t_L g1339 ( 
.A(n_1192),
.Y(n_1339)
);

INVx4_ASAP7_75t_L g1340 ( 
.A(n_1161),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1160),
.A2(n_1204),
.B1(n_1196),
.B2(n_1191),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1260),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1234),
.B(n_1198),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1203),
.Y(n_1344)
);

CKINVDCx6p67_ASAP7_75t_R g1345 ( 
.A(n_1192),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1155),
.Y(n_1346)
);

BUFx12f_ASAP7_75t_L g1347 ( 
.A(n_1174),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_1273),
.Y(n_1348)
);

BUFx8_ASAP7_75t_SL g1349 ( 
.A(n_1197),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1201),
.B(n_1206),
.Y(n_1350)
);

BUFx6f_ASAP7_75t_L g1351 ( 
.A(n_1208),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1186),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1199),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1186),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1204),
.A2(n_1190),
.B1(n_1188),
.B2(n_1164),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1202),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1186),
.Y(n_1357)
);

BUFx8_ASAP7_75t_L g1358 ( 
.A(n_1205),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1199),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1155),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1183),
.A2(n_1169),
.B1(n_1179),
.B2(n_1181),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1177),
.A2(n_1142),
.B1(n_1291),
.B2(n_1258),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1178),
.A2(n_1165),
.B(n_1189),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1182),
.B(n_1164),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1213),
.A2(n_1271),
.B1(n_1241),
.B2(n_1259),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1272),
.B(n_1156),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1200),
.A2(n_1232),
.B1(n_1275),
.B2(n_1245),
.Y(n_1367)
);

CKINVDCx11_ASAP7_75t_R g1368 ( 
.A(n_1220),
.Y(n_1368)
);

CKINVDCx9p33_ASAP7_75t_R g1369 ( 
.A(n_1276),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1156),
.B(n_1170),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_1212),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1217),
.A2(n_1267),
.B(n_1264),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1224),
.A2(n_1235),
.B1(n_1230),
.B2(n_1274),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1148),
.A2(n_1274),
.B1(n_1170),
.B2(n_1157),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1140),
.Y(n_1375)
);

BUFx8_ASAP7_75t_L g1376 ( 
.A(n_1237),
.Y(n_1376)
);

OAI22xp5_ASAP7_75t_L g1377 ( 
.A1(n_1149),
.A2(n_1159),
.B1(n_1214),
.B2(n_1231),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1250),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1261),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_SL g1380 ( 
.A1(n_1246),
.A2(n_1251),
.B1(n_1279),
.B2(n_1281),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1262),
.A2(n_1243),
.B1(n_1135),
.B2(n_497),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1262),
.A2(n_1228),
.B1(n_1243),
.B2(n_956),
.Y(n_1382)
);

CKINVDCx20_ASAP7_75t_R g1383 ( 
.A(n_1139),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_956),
.B2(n_1270),
.Y(n_1384)
);

CKINVDCx11_ASAP7_75t_R g1385 ( 
.A(n_1139),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1249),
.Y(n_1386)
);

CKINVDCx6p67_ASAP7_75t_R g1387 ( 
.A(n_1146),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1187),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_956),
.B2(n_1270),
.Y(n_1389)
);

INVx4_ASAP7_75t_L g1390 ( 
.A(n_1151),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1287),
.A2(n_1270),
.B1(n_754),
.B2(n_956),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1187),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_1139),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1139),
.Y(n_1394)
);

BUFx10_ASAP7_75t_L g1395 ( 
.A(n_1221),
.Y(n_1395)
);

INVx6_ASAP7_75t_L g1396 ( 
.A(n_1173),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1280),
.B(n_1167),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1287),
.A2(n_1270),
.B1(n_754),
.B2(n_956),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1280),
.B(n_1167),
.Y(n_1399)
);

BUFx12f_ASAP7_75t_L g1400 ( 
.A(n_1221),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_956),
.B2(n_1270),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_956),
.B2(n_1270),
.Y(n_1402)
);

INVx6_ASAP7_75t_L g1403 ( 
.A(n_1173),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1218),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_956),
.B2(n_1270),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_956),
.B2(n_1270),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1151),
.Y(n_1407)
);

OAI21xp33_ASAP7_75t_L g1408 ( 
.A1(n_1144),
.A2(n_1145),
.B(n_497),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1243),
.A2(n_1135),
.B1(n_497),
.B2(n_1228),
.Y(n_1409)
);

INVx1_ASAP7_75t_SL g1410 ( 
.A(n_1151),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1218),
.Y(n_1411)
);

INVx3_ASAP7_75t_L g1412 ( 
.A(n_1173),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1228),
.A2(n_1243),
.B1(n_956),
.B2(n_1270),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1287),
.A2(n_1270),
.B1(n_754),
.B2(n_956),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1322),
.B(n_1326),
.Y(n_1415)
);

BUFx2_ASAP7_75t_L g1416 ( 
.A(n_1366),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1378),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1379),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1372),
.A2(n_1377),
.B(n_1373),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1360),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1300),
.B(n_1296),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1354),
.Y(n_1422)
);

OA21x2_ASAP7_75t_L g1423 ( 
.A1(n_1373),
.A2(n_1362),
.B(n_1370),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1300),
.B(n_1298),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1328),
.B(n_1301),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1361),
.A2(n_1365),
.B(n_1362),
.Y(n_1426)
);

INVx4_ASAP7_75t_L g1427 ( 
.A(n_1350),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1304),
.B(n_1315),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1319),
.B(n_1320),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1361),
.A2(n_1365),
.B(n_1302),
.Y(n_1430)
);

OAI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1384),
.A2(n_1406),
.B1(n_1405),
.B2(n_1413),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1308),
.Y(n_1432)
);

OA21x2_ASAP7_75t_L g1433 ( 
.A1(n_1302),
.A2(n_1363),
.B(n_1359),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1391),
.A2(n_1398),
.B1(n_1414),
.B2(n_1389),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1344),
.Y(n_1435)
);

BUFx4f_ASAP7_75t_L g1436 ( 
.A(n_1297),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1352),
.A2(n_1357),
.B(n_1336),
.Y(n_1437)
);

INVx3_ASAP7_75t_SL g1438 ( 
.A(n_1339),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1324),
.B(n_1397),
.Y(n_1439)
);

HB1xp67_ASAP7_75t_L g1440 ( 
.A(n_1343),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1399),
.B(n_1303),
.Y(n_1441)
);

INVx2_ASAP7_75t_SL g1442 ( 
.A(n_1351),
.Y(n_1442)
);

OR2x2_ASAP7_75t_L g1443 ( 
.A(n_1381),
.B(n_1316),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1349),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1346),
.Y(n_1445)
);

AOI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1364),
.A2(n_1330),
.B(n_1409),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1329),
.B(n_1314),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1391),
.A2(n_1414),
.B1(n_1398),
.B2(n_1406),
.Y(n_1448)
);

AOI222xp33_ASAP7_75t_L g1449 ( 
.A1(n_1307),
.A2(n_1413),
.B1(n_1384),
.B2(n_1389),
.C1(n_1405),
.C2(n_1402),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1346),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1401),
.A2(n_1402),
.B1(n_1326),
.B2(n_1314),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1371),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1376),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1310),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1329),
.B(n_1334),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1376),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1334),
.B(n_1338),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1351),
.Y(n_1458)
);

AOI222xp33_ASAP7_75t_L g1459 ( 
.A1(n_1401),
.A2(n_1408),
.B1(n_1382),
.B2(n_1368),
.C1(n_1335),
.C2(n_1341),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1321),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1353),
.A2(n_1382),
.B(n_1375),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1305),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1371),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1367),
.A2(n_1355),
.B(n_1392),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1388),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1338),
.B(n_1337),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1337),
.B(n_1374),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1371),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1323),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1293),
.B(n_1331),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1342),
.Y(n_1471)
);

AO31x2_ASAP7_75t_L g1472 ( 
.A1(n_1404),
.A2(n_1411),
.A3(n_1369),
.B(n_1374),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1369),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1355),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1356),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1380),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1380),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1340),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1318),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1309),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1318),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1332),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1358),
.A2(n_1325),
.B1(n_1339),
.B2(n_1347),
.Y(n_1483)
);

INVxp33_ASAP7_75t_L g1484 ( 
.A(n_1385),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1412),
.B(n_1407),
.Y(n_1485)
);

OAI211xp5_ASAP7_75t_L g1486 ( 
.A1(n_1410),
.A2(n_1390),
.B(n_1294),
.C(n_1312),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1348),
.A2(n_1317),
.B1(n_1394),
.B2(n_1393),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1295),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1295),
.Y(n_1489)
);

OAI21x1_ASAP7_75t_L g1490 ( 
.A1(n_1306),
.A2(n_1403),
.B(n_1396),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1333),
.B(n_1345),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1403),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1396),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_L g1494 ( 
.A1(n_1327),
.A2(n_1387),
.B1(n_1292),
.B2(n_1396),
.Y(n_1494)
);

BUFx2_ASAP7_75t_L g1495 ( 
.A(n_1327),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1451),
.A2(n_1383),
.B(n_1311),
.Y(n_1496)
);

INVx3_ASAP7_75t_L g1497 ( 
.A(n_1427),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1451),
.A2(n_1386),
.B(n_1299),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1440),
.B(n_1292),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1441),
.B(n_1395),
.Y(n_1500)
);

AO32x2_ASAP7_75t_L g1501 ( 
.A1(n_1427),
.A2(n_1313),
.A3(n_1400),
.B1(n_1431),
.B2(n_1442),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1416),
.B(n_1439),
.Y(n_1502)
);

NAND4xp25_ASAP7_75t_L g1503 ( 
.A(n_1449),
.B(n_1459),
.C(n_1415),
.D(n_1448),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1439),
.B(n_1441),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1416),
.B(n_1476),
.Y(n_1505)
);

OAI21xp5_ASAP7_75t_L g1506 ( 
.A1(n_1446),
.A2(n_1443),
.B(n_1434),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1476),
.B(n_1477),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1477),
.B(n_1428),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1428),
.B(n_1429),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1453),
.B(n_1456),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1419),
.A2(n_1426),
.B(n_1430),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1425),
.B(n_1435),
.Y(n_1512)
);

AO32x2_ASAP7_75t_L g1513 ( 
.A1(n_1442),
.A2(n_1458),
.A3(n_1455),
.B1(n_1421),
.B2(n_1424),
.Y(n_1513)
);

OAI211xp5_ASAP7_75t_L g1514 ( 
.A1(n_1447),
.A2(n_1457),
.B(n_1425),
.C(n_1455),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1423),
.B(n_1433),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1447),
.A2(n_1457),
.B(n_1466),
.C(n_1474),
.Y(n_1516)
);

NAND3xp33_ASAP7_75t_L g1517 ( 
.A(n_1474),
.B(n_1482),
.C(n_1481),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1433),
.Y(n_1518)
);

AND2x4_ASAP7_75t_L g1519 ( 
.A(n_1490),
.B(n_1475),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1423),
.B(n_1433),
.Y(n_1520)
);

INVx3_ASAP7_75t_L g1521 ( 
.A(n_1475),
.Y(n_1521)
);

OAI211xp5_ASAP7_75t_L g1522 ( 
.A1(n_1470),
.A2(n_1467),
.B(n_1486),
.C(n_1479),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1423),
.B(n_1433),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1432),
.A2(n_1450),
.B(n_1445),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1464),
.A2(n_1423),
.B(n_1473),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1465),
.B(n_1480),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1468),
.A2(n_1420),
.B(n_1417),
.Y(n_1527)
);

AOI211xp5_ASAP7_75t_L g1528 ( 
.A1(n_1488),
.A2(n_1489),
.B(n_1493),
.C(n_1492),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1436),
.A2(n_1494),
.B1(n_1487),
.B2(n_1483),
.Y(n_1529)
);

AO32x2_ASAP7_75t_L g1530 ( 
.A1(n_1458),
.A2(n_1454),
.A3(n_1460),
.B1(n_1469),
.B2(n_1471),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1512),
.B(n_1472),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1503),
.A2(n_1461),
.B1(n_1437),
.B2(n_1422),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1506),
.A2(n_1461),
.B1(n_1437),
.B2(n_1418),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1509),
.B(n_1502),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1509),
.B(n_1472),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1527),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1502),
.B(n_1472),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1528),
.B(n_1478),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1504),
.B(n_1461),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1524),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1519),
.B(n_1463),
.Y(n_1541)
);

INVx3_ASAP7_75t_L g1542 ( 
.A(n_1521),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1501),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1527),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1522),
.B(n_1438),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1526),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1530),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1501),
.Y(n_1548)
);

NOR2xp33_ASAP7_75t_L g1549 ( 
.A(n_1499),
.B(n_1485),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1530),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1530),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1511),
.B(n_1463),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1511),
.B(n_1452),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1518),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1515),
.B(n_1452),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1515),
.B(n_1452),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1536),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1535),
.B(n_1520),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1543),
.B(n_1520),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1544),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1532),
.A2(n_1496),
.B1(n_1507),
.B2(n_1523),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1544),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1535),
.B(n_1523),
.Y(n_1563)
);

INVxp67_ASAP7_75t_L g1564 ( 
.A(n_1543),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1532),
.A2(n_1514),
.B1(n_1516),
.B2(n_1498),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1535),
.B(n_1513),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1540),
.Y(n_1567)
);

NOR2x1_ASAP7_75t_SL g1568 ( 
.A(n_1538),
.B(n_1517),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1554),
.B(n_1525),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1543),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1555),
.B(n_1513),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1554),
.B(n_1508),
.Y(n_1572)
);

INVx5_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1519),
.Y(n_1574)
);

AOI22xp33_ASAP7_75t_L g1575 ( 
.A1(n_1533),
.A2(n_1507),
.B1(n_1505),
.B2(n_1510),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1555),
.B(n_1513),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1555),
.B(n_1556),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1552),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1556),
.B(n_1513),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1541),
.B(n_1519),
.Y(n_1580)
);

NAND2x1p5_ASAP7_75t_L g1581 ( 
.A(n_1538),
.B(n_1497),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1548),
.Y(n_1582)
);

INVxp67_ASAP7_75t_L g1583 ( 
.A(n_1548),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1581),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1581),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1571),
.B(n_1548),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1560),
.Y(n_1587)
);

INVx2_ASAP7_75t_L g1588 ( 
.A(n_1557),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1568),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1571),
.B(n_1534),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1571),
.B(n_1534),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1564),
.B(n_1546),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1557),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1568),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1559),
.B(n_1539),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1571),
.B(n_1534),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1559),
.B(n_1564),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1576),
.B(n_1553),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1576),
.B(n_1553),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1576),
.B(n_1553),
.Y(n_1600)
);

NAND2xp33_ASAP7_75t_R g1601 ( 
.A(n_1566),
.B(n_1495),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1573),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1562),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1581),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1567),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1579),
.B(n_1537),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1559),
.B(n_1539),
.Y(n_1607)
);

BUFx3_ASAP7_75t_L g1608 ( 
.A(n_1581),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1568),
.B(n_1484),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1579),
.B(n_1537),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1579),
.B(n_1577),
.Y(n_1611)
);

BUFx2_ASAP7_75t_L g1612 ( 
.A(n_1581),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1579),
.B(n_1537),
.Y(n_1613)
);

AND2x4_ASAP7_75t_SL g1614 ( 
.A(n_1574),
.B(n_1580),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1559),
.B(n_1539),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1594),
.B(n_1570),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1603),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1594),
.B(n_1570),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1590),
.B(n_1570),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1590),
.B(n_1570),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1611),
.B(n_1570),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1587),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1588),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1588),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1611),
.B(n_1582),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1592),
.B(n_1583),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1592),
.B(n_1583),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1587),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1597),
.B(n_1582),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1611),
.B(n_1582),
.Y(n_1630)
);

AOI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1601),
.A2(n_1565),
.B1(n_1516),
.B2(n_1561),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1590),
.B(n_1582),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1597),
.B(n_1582),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1597),
.B(n_1572),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1588),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_1609),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1586),
.B(n_1572),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1588),
.Y(n_1638)
);

AND3x2_ASAP7_75t_L g1639 ( 
.A(n_1589),
.B(n_1495),
.C(n_1545),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1586),
.B(n_1558),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1593),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1603),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1591),
.B(n_1578),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1586),
.B(n_1572),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1593),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1606),
.B(n_1558),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1609),
.B(n_1444),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1593),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1591),
.B(n_1574),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1605),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1652)
);

OAI31xp33_ASAP7_75t_L g1653 ( 
.A1(n_1589),
.A2(n_1561),
.A3(n_1566),
.B(n_1545),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1587),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1591),
.B(n_1578),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1584),
.B(n_1462),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1596),
.B(n_1578),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1595),
.B(n_1569),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1621),
.B(n_1614),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1636),
.B(n_1558),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1636),
.B(n_1558),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1622),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1595),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1631),
.B(n_1563),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1631),
.B(n_1563),
.Y(n_1665)
);

AND2x4_ASAP7_75t_L g1666 ( 
.A(n_1621),
.B(n_1614),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1626),
.B(n_1563),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1648),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1639),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1656),
.Y(n_1670)
);

AOI211x1_ASAP7_75t_SL g1671 ( 
.A1(n_1626),
.A2(n_1529),
.B(n_1569),
.C(n_1593),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1634),
.B(n_1607),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1640),
.B(n_1607),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1616),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1621),
.B(n_1614),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1625),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1627),
.B(n_1563),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1639),
.B(n_1491),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1640),
.B(n_1607),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1627),
.B(n_1606),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1629),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1622),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1616),
.B(n_1606),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1616),
.B(n_1610),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1637),
.B(n_1615),
.Y(n_1685)
);

BUFx2_ASAP7_75t_L g1686 ( 
.A(n_1618),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1625),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1618),
.B(n_1610),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1628),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1625),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1637),
.B(n_1615),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1629),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1644),
.B(n_1615),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1630),
.B(n_1614),
.Y(n_1694)
);

AND2x4_ASAP7_75t_SL g1695 ( 
.A(n_1666),
.B(n_1500),
.Y(n_1695)
);

CKINVDCx14_ASAP7_75t_R g1696 ( 
.A(n_1686),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1668),
.B(n_1630),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1664),
.A2(n_1565),
.B1(n_1633),
.B2(n_1630),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1665),
.A2(n_1653),
.B(n_1565),
.C(n_1566),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1674),
.A2(n_1653),
.B(n_1633),
.Y(n_1700)
);

OAI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1669),
.A2(n_1601),
.B1(n_1531),
.B2(n_1647),
.Y(n_1701)
);

OAI21xp33_ASAP7_75t_SL g1702 ( 
.A1(n_1659),
.A2(n_1655),
.B(n_1643),
.Y(n_1702)
);

OAI211xp5_ASAP7_75t_SL g1703 ( 
.A1(n_1671),
.A2(n_1658),
.B(n_1652),
.C(n_1628),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1662),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1678),
.A2(n_1566),
.B1(n_1533),
.B2(n_1613),
.Y(n_1705)
);

INVxp67_ASAP7_75t_L g1706 ( 
.A(n_1681),
.Y(n_1706)
);

AOI21xp33_ASAP7_75t_SL g1707 ( 
.A1(n_1692),
.A2(n_1632),
.B(n_1620),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1671),
.B(n_1619),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1663),
.B(n_1644),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1662),
.Y(n_1710)
);

OAI31xp33_ASAP7_75t_L g1711 ( 
.A1(n_1660),
.A2(n_1613),
.A3(n_1610),
.B(n_1632),
.Y(n_1711)
);

AOI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1661),
.A2(n_1674),
.B(n_1686),
.C(n_1680),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1676),
.B(n_1619),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1676),
.B(n_1620),
.Y(n_1714)
);

OAI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1670),
.A2(n_1632),
.B(n_1652),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1663),
.B(n_1647),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1687),
.B(n_1643),
.Y(n_1717)
);

OAI221xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1683),
.A2(n_1658),
.B1(n_1575),
.B2(n_1613),
.C(n_1655),
.Y(n_1718)
);

OR2x2_ASAP7_75t_L g1719 ( 
.A(n_1672),
.B(n_1643),
.Y(n_1719)
);

NOR4xp25_ASAP7_75t_L g1720 ( 
.A(n_1682),
.B(n_1654),
.C(n_1657),
.D(n_1655),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1699),
.A2(n_1666),
.B1(n_1684),
.B2(n_1688),
.Y(n_1721)
);

OAI21xp33_ASAP7_75t_L g1722 ( 
.A1(n_1720),
.A2(n_1690),
.B(n_1687),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1697),
.B(n_1690),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1704),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1719),
.B(n_1672),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1710),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1709),
.B(n_1716),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1706),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1717),
.B(n_1685),
.Y(n_1729)
);

AOI21xp33_ASAP7_75t_SL g1730 ( 
.A1(n_1708),
.A2(n_1666),
.B(n_1685),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1713),
.Y(n_1731)
);

INVx1_ASAP7_75t_SL g1732 ( 
.A(n_1695),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1696),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1714),
.B(n_1691),
.Y(n_1734)
);

AND2x2_ASAP7_75t_SL g1735 ( 
.A(n_1703),
.B(n_1666),
.Y(n_1735)
);

OAI22xp5_ASAP7_75t_L g1736 ( 
.A1(n_1700),
.A2(n_1694),
.B1(n_1675),
.B2(n_1659),
.Y(n_1736)
);

NAND3xp33_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1712),
.C(n_1698),
.Y(n_1737)
);

AOI222xp33_ASAP7_75t_L g1738 ( 
.A1(n_1698),
.A2(n_1547),
.B1(n_1551),
.B2(n_1550),
.C1(n_1677),
.C2(n_1667),
.Y(n_1738)
);

NOR3xp33_ASAP7_75t_L g1739 ( 
.A(n_1715),
.B(n_1689),
.C(n_1682),
.Y(n_1739)
);

NOR4xp25_ASAP7_75t_SL g1740 ( 
.A(n_1718),
.B(n_1689),
.C(n_1612),
.D(n_1654),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1725),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1727),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1734),
.B(n_1691),
.Y(n_1743)
);

XNOR2xp5_ASAP7_75t_L g1744 ( 
.A(n_1733),
.B(n_1705),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1729),
.Y(n_1745)
);

NOR2xp33_ASAP7_75t_L g1746 ( 
.A(n_1732),
.B(n_1707),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1737),
.B(n_1693),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1723),
.B(n_1711),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1728),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1737),
.A2(n_1701),
.B1(n_1702),
.B2(n_1694),
.Y(n_1750)
);

NOR3xp33_ASAP7_75t_L g1751 ( 
.A(n_1730),
.B(n_1693),
.C(n_1679),
.Y(n_1751)
);

OAI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1738),
.A2(n_1679),
.B1(n_1673),
.B2(n_1641),
.C(n_1635),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1745),
.B(n_1731),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1747),
.A2(n_1740),
.B1(n_1735),
.B2(n_1721),
.Y(n_1754)
);

OAI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1747),
.A2(n_1752),
.B1(n_1750),
.B2(n_1722),
.C(n_1744),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1743),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1742),
.B(n_1739),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1741),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1751),
.B(n_1675),
.Y(n_1759)
);

NOR3x1_ASAP7_75t_L g1760 ( 
.A(n_1748),
.B(n_1736),
.C(n_1726),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1749),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1746),
.B(n_1724),
.Y(n_1762)
);

NAND3xp33_ASAP7_75t_L g1763 ( 
.A(n_1747),
.B(n_1740),
.C(n_1624),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1754),
.A2(n_1638),
.B1(n_1624),
.B2(n_1641),
.C(n_1623),
.Y(n_1764)
);

NOR3x1_ASAP7_75t_L g1765 ( 
.A(n_1755),
.B(n_1491),
.C(n_1673),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_L g1766 ( 
.A(n_1756),
.B(n_1617),
.Y(n_1766)
);

AOI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1763),
.A2(n_1638),
.B1(n_1624),
.B2(n_1635),
.C(n_1649),
.Y(n_1767)
);

AOI221x1_ASAP7_75t_L g1768 ( 
.A1(n_1763),
.A2(n_1617),
.B1(n_1651),
.B2(n_1642),
.C(n_1646),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1764),
.A2(n_1757),
.B1(n_1761),
.B2(n_1762),
.C(n_1758),
.Y(n_1769)
);

O2A1O1Ixp5_ASAP7_75t_SL g1770 ( 
.A1(n_1768),
.A2(n_1753),
.B(n_1760),
.C(n_1765),
.Y(n_1770)
);

AOI322xp5_ASAP7_75t_L g1771 ( 
.A1(n_1766),
.A2(n_1759),
.A3(n_1767),
.B1(n_1635),
.B2(n_1623),
.C1(n_1649),
.C2(n_1638),
.Y(n_1771)
);

AOI31xp33_ASAP7_75t_L g1772 ( 
.A1(n_1766),
.A2(n_1657),
.A3(n_1604),
.B(n_1650),
.Y(n_1772)
);

AOI211xp5_ASAP7_75t_SL g1773 ( 
.A1(n_1764),
.A2(n_1602),
.B(n_1657),
.C(n_1650),
.Y(n_1773)
);

OAI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1768),
.A2(n_1641),
.B1(n_1649),
.B2(n_1623),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1769),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_L g1776 ( 
.A(n_1770),
.B(n_1642),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1774),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1773),
.B(n_1596),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1772),
.B(n_1646),
.Y(n_1779)
);

OAI22xp33_ASAP7_75t_L g1780 ( 
.A1(n_1777),
.A2(n_1645),
.B1(n_1771),
.B2(n_1584),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1779),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1775),
.B(n_1651),
.Y(n_1782)
);

AOI22x1_ASAP7_75t_L g1783 ( 
.A1(n_1781),
.A2(n_1778),
.B1(n_1776),
.B2(n_1612),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1783),
.A2(n_1776),
.B1(n_1780),
.B2(n_1782),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1784),
.B(n_1645),
.Y(n_1785)
);

NAND3x1_ASAP7_75t_L g1786 ( 
.A(n_1784),
.B(n_1602),
.C(n_1596),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1785),
.A2(n_1786),
.B1(n_1645),
.B2(n_1599),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1785),
.Y(n_1788)
);

OAI21xp33_ASAP7_75t_L g1789 ( 
.A1(n_1788),
.A2(n_1585),
.B(n_1584),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1787),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1598),
.B1(n_1599),
.B2(n_1600),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1791),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1792),
.Y(n_1793)
);

OAI221xp5_ASAP7_75t_R g1794 ( 
.A1(n_1793),
.A2(n_1789),
.B1(n_1612),
.B2(n_1585),
.C(n_1584),
.Y(n_1794)
);

AOI211xp5_ASAP7_75t_L g1795 ( 
.A1(n_1794),
.A2(n_1604),
.B(n_1549),
.C(n_1608),
.Y(n_1795)
);


endmodule