module fake_jpeg_2173_n_207 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_207);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_207;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_93;
wire n_91;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_18),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_41),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_48),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_33),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_12),
.Y(n_66)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx16f_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_22),
.B(n_24),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_53),
.Y(n_80)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_64),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_93),
.Y(n_105)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_81),
.Y(n_96)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_78),
.A2(n_71),
.B1(n_59),
.B2(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_89),
.B1(n_63),
.B2(n_67),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_71),
.B1(n_62),
.B2(n_61),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_88),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_66),
.B1(n_56),
.B2(n_49),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_87),
.A2(n_91),
.B1(n_57),
.B2(n_65),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g88 ( 
.A(n_79),
.B(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_67),
.B1(n_58),
.B2(n_56),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_72),
.A2(n_49),
.B1(n_58),
.B2(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_SL g99 ( 
.A1(n_88),
.A2(n_63),
.B(n_54),
.C(n_60),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_82),
.A3(n_54),
.B1(n_55),
.B2(n_52),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_94),
.Y(n_100)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_102),
.B(n_108),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_84),
.B1(n_83),
.B2(n_54),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_2),
.B(n_3),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_107),
.Y(n_120)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_106),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_60),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_114),
.B(n_119),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_95),
.A2(n_86),
.B1(n_84),
.B2(n_83),
.Y(n_115)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_118),
.B(n_25),
.C(n_46),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_84),
.B1(n_83),
.B2(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_57),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_84),
.B1(n_83),
.B2(n_54),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_124),
.B1(n_128),
.B2(n_26),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_122),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_70),
.B1(n_1),
.B2(n_2),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_0),
.B(n_1),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_110),
.B(n_5),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_132),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_3),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_4),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_134),
.B(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_5),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_110),
.C(n_23),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_149),
.C(n_17),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_6),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_140),
.B(n_141),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_6),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_147),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_7),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_7),
.Y(n_144)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_8),
.Y(n_145)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_8),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_11),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_12),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_150),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_30),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_47),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_151),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_13),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_154),
.Y(n_171)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_113),
.B(n_121),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_45),
.B(n_43),
.Y(n_157)
);

OAI21xp33_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_153),
.B(n_38),
.Y(n_184)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_166),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_165),
.A2(n_150),
.B1(n_153),
.B2(n_142),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_173),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_18),
.B(n_19),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_37),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_142),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_161),
.B1(n_164),
.B2(n_152),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_179),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_153),
.C(n_139),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_182),
.C(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_184),
.A2(n_186),
.B(n_157),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_180),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_160),
.B1(n_171),
.B2(n_158),
.C(n_163),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_187),
.A2(n_188),
.B(n_192),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_176),
.B(n_177),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_191),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_169),
.B(n_165),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_185),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_168),
.C(n_36),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_193),
.B(n_167),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_178),
.B1(n_163),
.B2(n_172),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_198),
.A2(n_170),
.B1(n_162),
.B2(n_174),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_195),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_197),
.B(n_200),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_204),
.A2(n_203),
.B1(n_194),
.B2(n_39),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_40),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_20),
.Y(n_207)
);


endmodule