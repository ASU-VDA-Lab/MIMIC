module fake_netlist_5_1959_n_160 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_160);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;

output n_160;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_136;
wire n_86;
wire n_124;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_53;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_64;
wire n_77;
wire n_106;
wire n_102;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_141;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_28),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVxp67_ASAP7_75t_SL g51 ( 
.A(n_15),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_1),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_37),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_45),
.B(n_6),
.Y(n_65)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_33),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_48),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_7),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_46),
.B(n_43),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_46),
.B(n_43),
.Y(n_75)
);

NAND2x1p5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_38),
.B(n_33),
.C(n_10),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_23),
.Y(n_80)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_8),
.B(n_9),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_9),
.B(n_10),
.C(n_11),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_60),
.B(n_21),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_11),
.C(n_12),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_22),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_12),
.B(n_13),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_73),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_77),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_71),
.Y(n_94)
);

O2A1O1Ixp5_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_71),
.B(n_58),
.C(n_63),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_62),
.B(n_72),
.Y(n_96)
);

AND2x4_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_70),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_68),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_62),
.B(n_72),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_79),
.A2(n_64),
.B1(n_70),
.B2(n_67),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_83),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_75),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_66),
.Y(n_109)
);

OAI221xp5_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_100),
.B1(n_76),
.B2(n_90),
.C(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_104),
.A2(n_97),
.B1(n_76),
.B2(n_74),
.Y(n_111)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_90),
.C(n_100),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_103),
.A2(n_66),
.B1(n_85),
.B2(n_88),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_105),
.B(n_84),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_82),
.B1(n_93),
.B2(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_108),
.B1(n_105),
.B2(n_106),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_117),
.B(n_106),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_113),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_102),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_127),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_108),
.Y(n_129)
);

NAND3x1_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_89),
.C(n_63),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_98),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_120),
.B(n_122),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_126),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NAND4xp75_ASAP7_75t_SL g137 ( 
.A(n_130),
.B(n_122),
.C(n_132),
.D(n_95),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_SL g138 ( 
.A(n_130),
.B(n_55),
.C(n_56),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_133),
.B(n_124),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_134),
.B(n_124),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_129),
.B1(n_57),
.B2(n_56),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_129),
.B1(n_114),
.B2(n_68),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_123),
.Y(n_147)
);

AND3x4_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_123),
.C(n_14),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_13),
.B1(n_15),
.B2(n_68),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_148),
.A2(n_145),
.B1(n_107),
.B2(n_101),
.Y(n_153)
);

AOI211x1_ASAP7_75t_L g154 ( 
.A1(n_150),
.A2(n_96),
.B(n_101),
.C(n_98),
.Y(n_154)
);

A2O1A1Ixp33_ASAP7_75t_L g155 ( 
.A1(n_149),
.A2(n_96),
.B(n_107),
.C(n_83),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_153),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_155),
.A2(n_149),
.B1(n_152),
.B2(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_154),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g159 ( 
.A(n_157),
.B(n_155),
.C(n_146),
.Y(n_159)
);

OAI221xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_156),
.B1(n_158),
.B2(n_151),
.C(n_146),
.Y(n_160)
);


endmodule