module fake_netlist_1_3614_n_543 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_543);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_543;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_67), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_17), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_23), .Y(n_80) );
INVxp67_ASAP7_75t_SL g81 ( .A(n_25), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_1), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_22), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_62), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_16), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_49), .Y(n_86) );
INVx2_ASAP7_75t_SL g87 ( .A(n_60), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_20), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_32), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_66), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_35), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_71), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_34), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_4), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_15), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_75), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_4), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_59), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_69), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_42), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_65), .Y(n_102) );
INVx2_ASAP7_75t_L g103 ( .A(n_55), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_26), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_77), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_46), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_64), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_2), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_53), .Y(n_110) );
INVxp67_ASAP7_75t_L g111 ( .A(n_74), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_10), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_68), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_58), .Y(n_114) );
INVx5_ASAP7_75t_L g115 ( .A(n_106), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_109), .B(n_0), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_106), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_78), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_106), .Y(n_119) );
INVx2_ASAP7_75t_SL g120 ( .A(n_113), .Y(n_120) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_106), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
AND2x4_ASAP7_75t_L g123 ( .A(n_82), .B(n_94), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_85), .Y(n_125) );
HB1xp67_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_87), .B(n_0), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_106), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
OAI22xp5_ASAP7_75t_SL g131 ( .A1(n_112), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_89), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_91), .Y(n_133) );
BUFx8_ASAP7_75t_L g134 ( .A(n_87), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_96), .Y(n_136) );
BUFx3_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_135), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_120), .B(n_111), .Y(n_139) );
INVx8_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
OAI22xp33_ASAP7_75t_L g142 ( .A1(n_126), .A2(n_108), .B1(n_82), .B2(n_95), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_120), .B(n_93), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_135), .Y(n_145) );
INVx3_ASAP7_75t_L g146 ( .A(n_123), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_123), .B(n_94), .Y(n_147) );
OR2x2_ASAP7_75t_SL g148 ( .A(n_116), .B(n_95), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_134), .B(n_90), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_135), .Y(n_150) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_123), .B(n_114), .Y(n_151) );
INVx5_ASAP7_75t_L g152 ( .A(n_115), .Y(n_152) );
INVx4_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_134), .B(n_100), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_135), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_118), .B(n_97), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_122), .B(n_114), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_119), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_125), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_125), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_122), .B(n_110), .Y(n_162) );
OR2x2_ASAP7_75t_L g163 ( .A(n_157), .B(n_131), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_153), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_155), .B(n_134), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_140), .B(n_134), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_140), .Y(n_167) );
AND2x4_ASAP7_75t_L g168 ( .A(n_147), .B(n_124), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_147), .B(n_124), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_140), .B(n_132), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_139), .B(n_132), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_140), .B(n_133), .Y(n_172) );
AND2x6_ASAP7_75t_SL g173 ( .A(n_157), .B(n_127), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_153), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_153), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_140), .B(n_146), .Y(n_177) );
NAND2x1p5_ASAP7_75t_L g178 ( .A(n_151), .B(n_125), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_146), .B(n_133), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_151), .B(n_79), .Y(n_180) );
INVx2_ASAP7_75t_SL g181 ( .A(n_151), .Y(n_181) );
NOR2xp67_ASAP7_75t_L g182 ( .A(n_144), .B(n_129), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_160), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_146), .A2(n_129), .B1(n_137), .B2(n_130), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_162), .B(n_129), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
BUFx2_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_161), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_149), .B(n_80), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_148), .B(n_129), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_158), .B(n_137), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_158), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_154), .B(n_137), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_142), .B(n_84), .Y(n_195) );
OAI22x1_ASAP7_75t_L g196 ( .A1(n_187), .A2(n_81), .B1(n_86), .B2(n_98), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_165), .A2(n_161), .B(n_156), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_173), .B(n_88), .Y(n_198) );
INVx4_ASAP7_75t_L g199 ( .A(n_167), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_178), .A2(n_136), .B1(n_130), .B2(n_98), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_193), .B(n_130), .Y(n_201) );
NAND2x1p5_ASAP7_75t_L g202 ( .A(n_167), .B(n_136), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_181), .A2(n_136), .B1(n_91), .B2(n_92), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_193), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_164), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_191), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_183), .A2(n_141), .B(n_156), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_179), .Y(n_209) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_178), .A2(n_92), .B1(n_99), .B2(n_104), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_183), .A2(n_141), .B(n_150), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_186), .A2(n_143), .B(n_150), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_195), .A2(n_99), .B(n_101), .C(n_104), .Y(n_213) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_178), .A2(n_101), .B1(n_100), .B2(n_103), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g215 ( .A1(n_171), .A2(n_103), .B(n_107), .C(n_117), .Y(n_215) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_167), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_186), .A2(n_145), .B(n_143), .Y(n_217) );
AOI222xp33_ASAP7_75t_L g218 ( .A1(n_187), .A2(n_107), .B1(n_105), .B2(n_102), .C1(n_128), .C2(n_117), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_168), .B(n_3), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_191), .Y(n_220) );
OR2x6_ASAP7_75t_L g221 ( .A(n_181), .B(n_117), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_191), .Y(n_222) );
OAI21xp33_ASAP7_75t_L g223 ( .A1(n_170), .A2(n_145), .B(n_128), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_188), .A2(n_138), .B(n_128), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_188), .A2(n_152), .B(n_115), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_168), .B(n_152), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_174), .A2(n_152), .B(n_115), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_168), .B(n_5), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_197), .A2(n_194), .B(n_185), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_209), .B(n_169), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_220), .B(n_169), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_199), .B(n_166), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_202), .A2(n_169), .B1(n_172), .B2(n_190), .Y(n_233) );
AO31x2_ASAP7_75t_L g234 ( .A1(n_215), .A2(n_174), .A3(n_175), .B(n_176), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_205), .B(n_163), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_199), .B(n_163), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_219), .Y(n_237) );
AO32x2_ASAP7_75t_L g238 ( .A1(n_214), .A2(n_184), .A3(n_182), .B1(n_180), .B2(n_121), .Y(n_238) );
AO32x2_ASAP7_75t_L g239 ( .A1(n_214), .A2(n_119), .A3(n_121), .B1(n_189), .B2(n_8), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_198), .Y(n_240) );
INVxp33_ASAP7_75t_SL g241 ( .A(n_216), .Y(n_241) );
NOR2xp67_ASAP7_75t_L g242 ( .A(n_196), .B(n_5), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_L g243 ( .A1(n_210), .A2(n_177), .B(n_175), .C(n_176), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_210), .A2(n_6), .B(n_7), .C(n_8), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_207), .B(n_6), .Y(n_245) );
OAI21x1_ASAP7_75t_L g246 ( .A1(n_208), .A2(n_192), .B(n_121), .Y(n_246) );
CKINVDCx11_ASAP7_75t_R g247 ( .A(n_222), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_218), .A2(n_192), .B1(n_115), .B2(n_121), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_211), .A2(n_192), .B(n_159), .Y(n_249) );
INVx2_ASAP7_75t_L g250 ( .A(n_204), .Y(n_250) );
OAI21x1_ASAP7_75t_L g251 ( .A1(n_212), .A2(n_192), .B(n_121), .Y(n_251) );
INVx5_ASAP7_75t_L g252 ( .A(n_221), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_SL g253 ( .A1(n_228), .A2(n_41), .B(n_54), .C(n_76), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_226), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_217), .A2(n_192), .B(n_121), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_252), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_250), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_230), .Y(n_258) );
INVx2_ASAP7_75t_SL g259 ( .A(n_252), .Y(n_259) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_246), .A2(n_224), .B(n_200), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_235), .B(n_218), .Y(n_261) );
INVx8_ASAP7_75t_L g262 ( .A(n_252), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_229), .A2(n_221), .B(n_201), .Y(n_263) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_251), .A2(n_202), .B(n_225), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_230), .Y(n_265) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_229), .A2(n_223), .B(n_213), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_249), .A2(n_221), .B(n_206), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_237), .B(n_226), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_235), .B(n_203), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_255), .A2(n_227), .B(n_159), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_232), .A2(n_159), .B(n_119), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_253), .A2(n_159), .B(n_119), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_236), .B(n_7), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_236), .A2(n_119), .B1(n_115), .B2(n_11), .Y(n_275) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_242), .A2(n_119), .B(n_115), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_234), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_274), .Y(n_278) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_272), .A2(n_244), .B(n_233), .Y(n_279) );
AND2x4_ASAP7_75t_L g280 ( .A(n_256), .B(n_252), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_274), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g282 ( .A1(n_262), .A2(n_241), .B1(n_254), .B2(n_245), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_256), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_274), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_270), .A2(n_243), .B(n_248), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_257), .B(n_239), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_277), .Y(n_287) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_268), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_257), .B(n_239), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_277), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_261), .B(n_231), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_277), .Y(n_292) );
OA21x2_ASAP7_75t_L g293 ( .A1(n_263), .A2(n_239), .B(n_238), .Y(n_293) );
INVxp67_ASAP7_75t_L g294 ( .A(n_268), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_258), .B(n_234), .Y(n_296) );
OR2x6_ASAP7_75t_L g297 ( .A(n_262), .B(n_231), .Y(n_297) );
INVx5_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_258), .B(n_238), .Y(n_299) );
HB1xp67_ASAP7_75t_L g300 ( .A(n_288), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_296), .B(n_265), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_296), .B(n_276), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_278), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_273), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
BUFx3_ASAP7_75t_L g306 ( .A(n_298), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_281), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_298), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_299), .B(n_265), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_281), .B(n_273), .Y(n_311) );
OAI211xp5_ASAP7_75t_L g312 ( .A1(n_282), .A2(n_247), .B(n_275), .C(n_240), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_299), .B(n_238), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_286), .B(n_276), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_283), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_284), .B(n_256), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_286), .B(n_276), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_289), .B(n_256), .Y(n_318) );
BUFx2_ASAP7_75t_L g319 ( .A(n_283), .Y(n_319) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_297), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_284), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_289), .B(n_266), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_284), .B(n_266), .Y(n_323) );
INVx3_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_287), .B(n_259), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_287), .B(n_259), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_290), .Y(n_327) );
INVxp67_ASAP7_75t_L g328 ( .A(n_295), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_290), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_305), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_302), .B(n_290), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_301), .B(n_292), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_318), .B(n_292), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_300), .B(n_291), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_307), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_318), .B(n_292), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_303), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_303), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_314), .B(n_293), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_324), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_314), .B(n_293), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_324), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_317), .B(n_293), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_308), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_310), .B(n_294), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_317), .B(n_293), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_301), .B(n_297), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_321), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_322), .B(n_279), .Y(n_353) );
INVx4_ASAP7_75t_L g354 ( .A(n_306), .Y(n_354) );
AND2x4_ASAP7_75t_SL g355 ( .A(n_309), .B(n_280), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_326), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_310), .B(n_280), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_328), .B(n_280), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_302), .B(n_298), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_322), .B(n_279), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_324), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_313), .B(n_279), .Y(n_363) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_312), .B(n_295), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_285), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_319), .B(n_297), .Y(n_366) );
OR2x6_ASAP7_75t_L g367 ( .A(n_319), .B(n_262), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_304), .B(n_280), .Y(n_368) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_315), .A2(n_275), .B1(n_269), .B2(n_295), .C(n_271), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g370 ( .A1(n_302), .A2(n_297), .B1(n_298), .B2(n_266), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_327), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_326), .Y(n_372) );
OAI21xp33_ASAP7_75t_SL g373 ( .A1(n_309), .A2(n_297), .B(n_285), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_342), .B(n_302), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_356), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_372), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_351), .B(n_304), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_337), .B(n_320), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_342), .B(n_323), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_330), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_330), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_333), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_349), .B(n_311), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_353), .B(n_311), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_351), .B(n_316), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_335), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_344), .B(n_323), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_353), .B(n_325), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_344), .B(n_324), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_361), .B(n_325), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_333), .Y(n_391) );
NOR2x1p5_ASAP7_75t_SL g392 ( .A(n_366), .B(n_316), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_334), .B(n_325), .Y(n_393) );
OR2x6_ASAP7_75t_L g394 ( .A(n_367), .B(n_306), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_358), .B(n_327), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_336), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_346), .B(n_329), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_361), .B(n_325), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_364), .B(n_306), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_346), .B(n_329), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_335), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_350), .B(n_298), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_336), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_350), .B(n_298), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_334), .B(n_9), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_340), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_363), .B(n_9), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_338), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_338), .Y(n_409) );
NAND2x1_ASAP7_75t_L g410 ( .A(n_354), .B(n_267), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_347), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_340), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_347), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_348), .Y(n_414) );
INVx1_ASAP7_75t_SL g415 ( .A(n_355), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_348), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_354), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_352), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_341), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_352), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g421 ( .A(n_354), .B(n_264), .Y(n_421) );
INVxp67_ASAP7_75t_L g422 ( .A(n_366), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_332), .B(n_10), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_357), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_357), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g426 ( .A1(n_402), .A2(n_355), .B1(n_360), .B2(n_367), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_376), .B(n_363), .Y(n_428) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_394), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_380), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_397), .B(n_365), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_381), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_401), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_382), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_391), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_386), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_417), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_374), .B(n_339), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_396), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_386), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g441 ( .A1(n_394), .A2(n_367), .B1(n_373), .B2(n_370), .C(n_368), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g442 ( .A1(n_399), .A2(n_359), .B1(n_365), .B2(n_367), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_417), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_415), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_374), .B(n_379), .Y(n_445) );
INVx1_ASAP7_75t_SL g446 ( .A(n_402), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_403), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_379), .B(n_339), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_397), .B(n_332), .Y(n_449) );
INVx1_ASAP7_75t_SL g450 ( .A(n_404), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_408), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_409), .Y(n_452) );
NOR2x1_ASAP7_75t_L g453 ( .A(n_394), .B(n_360), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_400), .B(n_422), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_411), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_400), .B(n_371), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_413), .Y(n_457) );
AND2x4_ASAP7_75t_SL g458 ( .A(n_404), .B(n_360), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_422), .B(n_371), .Y(n_459) );
INVx2_ASAP7_75t_SL g460 ( .A(n_393), .Y(n_460) );
AOI33xp33_ASAP7_75t_L g461 ( .A1(n_405), .A2(n_331), .A3(n_360), .B1(n_369), .B2(n_345), .B3(n_343), .Y(n_461) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_378), .B(n_331), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_407), .B(n_331), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_387), .B(n_331), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_389), .Y(n_465) );
OR2x2_ASAP7_75t_L g466 ( .A(n_387), .B(n_341), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_414), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_384), .B(n_362), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_395), .B(n_362), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_423), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_445), .B(n_389), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_459), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_456), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_430), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_470), .B(n_398), .Y(n_476) );
NOR4xp25_ASAP7_75t_L g477 ( .A(n_441), .B(n_399), .C(n_383), .D(n_424), .Y(n_477) );
NOR2xp67_ASAP7_75t_L g478 ( .A(n_440), .B(n_390), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
INVxp33_ASAP7_75t_L g481 ( .A(n_453), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_470), .B(n_388), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_435), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_436), .Y(n_484) );
AOI32xp33_ASAP7_75t_L g485 ( .A1(n_426), .A2(n_392), .A3(n_385), .B1(n_377), .B2(n_420), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_461), .B(n_425), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_436), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_461), .B(n_416), .Y(n_488) );
OAI221xp5_ASAP7_75t_L g489 ( .A1(n_441), .A2(n_410), .B1(n_421), .B2(n_418), .C(n_412), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_426), .B(n_401), .C(n_419), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
AOI21xp33_ASAP7_75t_L g492 ( .A1(n_427), .A2(n_421), .B(n_419), .Y(n_492) );
OAI22xp5_ASAP7_75t_SL g493 ( .A1(n_429), .A2(n_406), .B1(n_412), .B2(n_345), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_428), .B(n_406), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_438), .B(n_343), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_433), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_437), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_466), .B(n_11), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_447), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_475), .Y(n_501) );
NAND2xp33_ASAP7_75t_SL g502 ( .A(n_481), .B(n_443), .Y(n_502) );
OAI21x1_ASAP7_75t_SL g503 ( .A1(n_472), .A2(n_460), .B(n_454), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_477), .A2(n_462), .B1(n_463), .B2(n_450), .C(n_446), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_486), .A2(n_463), .B1(n_442), .B2(n_462), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_489), .A2(n_458), .B1(n_465), .B2(n_449), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_488), .A2(n_458), .B1(n_464), .B2(n_431), .Y(n_507) );
AOI32xp33_ASAP7_75t_L g508 ( .A1(n_481), .A2(n_448), .A3(n_469), .B1(n_467), .B2(n_457), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_491), .A2(n_455), .B(n_452), .C(n_451), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_485), .A2(n_468), .B1(n_433), .B2(n_14), .C(n_15), .Y(n_510) );
AOI322xp5_ASAP7_75t_L g511 ( .A1(n_476), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_260), .C1(n_264), .C2(n_21), .Y(n_511) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_499), .Y(n_512) );
AOI221xp5_ASAP7_75t_L g513 ( .A1(n_490), .A2(n_12), .B1(n_13), .B2(n_159), .C(n_19), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_473), .A2(n_18), .B1(n_24), .B2(n_27), .C(n_28), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_474), .B(n_260), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_482), .B(n_29), .Y(n_516) );
OAI22xp33_ASAP7_75t_SL g517 ( .A1(n_499), .A2(n_30), .B1(n_31), .B2(n_33), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_478), .A2(n_36), .B1(n_37), .B2(n_38), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_504), .A2(n_500), .B1(n_498), .B2(n_480), .C(n_483), .Y(n_519) );
BUFx8_ASAP7_75t_L g520 ( .A(n_501), .Y(n_520) );
AOI21xp33_ASAP7_75t_L g521 ( .A1(n_510), .A2(n_484), .B(n_487), .Y(n_521) );
OR3x1_ASAP7_75t_L g522 ( .A(n_506), .B(n_492), .C(n_479), .Y(n_522) );
AOI22xp5_ASAP7_75t_SL g523 ( .A1(n_512), .A2(n_497), .B1(n_484), .B2(n_487), .Y(n_523) );
AOI211xp5_ASAP7_75t_L g524 ( .A1(n_517), .A2(n_493), .B(n_472), .C(n_494), .Y(n_524) );
O2A1O1Ixp5_ASAP7_75t_L g525 ( .A1(n_502), .A2(n_496), .B(n_471), .C(n_495), .Y(n_525) );
OAI22xp5_ASAP7_75t_L g526 ( .A1(n_507), .A2(n_471), .B1(n_495), .B2(n_496), .Y(n_526) );
OAI21xp5_ASAP7_75t_SL g527 ( .A1(n_508), .A2(n_39), .B(n_43), .Y(n_527) );
OAI211xp5_ASAP7_75t_L g528 ( .A1(n_524), .A2(n_513), .B(n_505), .C(n_511), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_519), .B(n_509), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_527), .A2(n_503), .B(n_515), .Y(n_530) );
NAND4xp25_ASAP7_75t_L g531 ( .A(n_525), .B(n_518), .C(n_514), .D(n_516), .Y(n_531) );
OAI211xp5_ASAP7_75t_SL g532 ( .A1(n_521), .A2(n_44), .B(n_45), .C(n_47), .Y(n_532) );
INVx3_ASAP7_75t_SL g533 ( .A(n_528), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_529), .B(n_523), .Y(n_534) );
NOR5xp2_ASAP7_75t_L g535 ( .A(n_532), .B(n_522), .C(n_520), .D(n_526), .E(n_52), .Y(n_535) );
OR3x1_ASAP7_75t_L g536 ( .A(n_533), .B(n_531), .C(n_530), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_534), .Y(n_537) );
OAI22xp5_ASAP7_75t_SL g538 ( .A1(n_536), .A2(n_535), .B1(n_50), .B2(n_51), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_538), .A2(n_537), .B1(n_152), .B2(n_57), .Y(n_539) );
XOR2xp5_ASAP7_75t_L g540 ( .A(n_539), .B(n_48), .Y(n_540) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_540), .A2(n_56), .B(n_61), .Y(n_541) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_541), .A2(n_70), .B(n_72), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g543 ( .A1(n_542), .A2(n_73), .B1(n_152), .B2(n_537), .Y(n_543) );
endmodule