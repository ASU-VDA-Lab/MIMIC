module fake_jpeg_20843_n_354 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_354);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_354;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_15),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_7),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_19),
.B(n_16),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_48),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g92 ( 
.A(n_46),
.Y(n_92)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_22),
.B(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_62),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_21),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g55 ( 
.A(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_60),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_23),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g61 ( 
.A(n_36),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_63),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_0),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_28),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_71),
.B(n_84),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_31),
.C(n_30),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_86),
.C(n_31),
.Y(n_136)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVxp67_ASAP7_75t_SL g122 ( 
.A(n_75),
.Y(n_122)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_90),
.Y(n_124)
);

CKINVDCx9p33_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_82),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_83),
.B(n_89),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_28),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_31),
.C(n_30),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_37),
.Y(n_89)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_93),
.B(n_100),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_44),
.A2(n_28),
.B1(n_24),
.B2(n_40),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_101),
.B1(n_107),
.B2(n_20),
.Y(n_144)
);

CKINVDCx12_ASAP7_75t_R g97 ( 
.A(n_61),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_98),
.B(n_102),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_53),
.A2(n_24),
.B1(n_35),
.B2(n_40),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_22),
.Y(n_102)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_117),
.Y(n_127)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_105),
.Y(n_151)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_24),
.B(n_39),
.C(n_37),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_65),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_66),
.B(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_116),
.Y(n_152)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_59),
.B(n_25),
.Y(n_117)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_82),
.B(n_31),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_139),
.Y(n_187)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_67),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_126),
.A2(n_132),
.B(n_110),
.Y(n_179)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_96),
.A2(n_25),
.B1(n_26),
.B2(n_34),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_144),
.B1(n_99),
.B2(n_113),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_27),
.B1(n_34),
.B2(n_20),
.Y(n_132)
);

AO22x2_ASAP7_75t_L g133 ( 
.A1(n_86),
.A2(n_27),
.B1(n_18),
.B2(n_20),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_92),
.B1(n_105),
.B2(n_75),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_138),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_72),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_149),
.Y(n_161)
);

OR2x4_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_35),
.Y(n_138)
);

NOR2x1_ASAP7_75t_L g139 ( 
.A(n_107),
.B(n_20),
.Y(n_139)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_145),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_85),
.Y(n_146)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_110),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_101),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_95),
.B(n_20),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_133),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_81),
.A2(n_18),
.B1(n_8),
.B2(n_15),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_94),
.C(n_71),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_156),
.B(n_159),
.C(n_162),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_125),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_168),
.C(n_189),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_158),
.A2(n_148),
.B1(n_140),
.B2(n_141),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_150),
.B(n_84),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_111),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_69),
.Y(n_162)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_167),
.Y(n_219)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_10),
.B(n_12),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_78),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_169),
.B(n_176),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_149),
.A2(n_80),
.B1(n_77),
.B2(n_81),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_147),
.B1(n_146),
.B2(n_140),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_171),
.A2(n_179),
.B(n_120),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_142),
.B(n_88),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_172),
.B(n_174),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_137),
.B(n_135),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_88),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_122),
.Y(n_177)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_100),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_181),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_124),
.B(n_100),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_144),
.B(n_18),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_184),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_127),
.B(n_5),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_191),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_85),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_115),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_18),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_134),
.B(n_139),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_133),
.B(n_115),
.Y(n_192)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_193),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g194 ( 
.A(n_131),
.Y(n_194)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_195),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_196),
.A2(n_203),
.B(n_206),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_198),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_202),
.Y(n_243)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_132),
.B(n_133),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_176),
.A2(n_133),
.B1(n_132),
.B2(n_129),
.Y(n_205)
);

A2O1A1O1Ixp25_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_132),
.B(n_155),
.C(n_18),
.D(n_123),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_213),
.B(n_166),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_129),
.B1(n_123),
.B2(n_77),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_106),
.B1(n_114),
.B2(n_92),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_155),
.B(n_114),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_207),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_186),
.A2(n_79),
.B1(n_73),
.B2(n_93),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_216),
.B(n_218),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g217 ( 
.A(n_185),
.Y(n_217)
);

BUFx4f_ASAP7_75t_SL g249 ( 
.A(n_217),
.Y(n_249)
);

AND2x6_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_120),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_187),
.A2(n_73),
.B1(n_119),
.B2(n_70),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_161),
.A2(n_27),
.B1(n_119),
.B2(n_2),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_170),
.A2(n_6),
.B1(n_14),
.B2(n_13),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_178),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_226),
.B(n_228),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_6),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_156),
.C(n_159),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_233),
.C(n_238),
.Y(n_262)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_201),
.A2(n_169),
.A3(n_179),
.B1(n_187),
.B2(n_160),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_247),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_157),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_236),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_162),
.C(n_160),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_160),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_234),
.B(n_241),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_199),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_163),
.C(n_164),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_239),
.A2(n_215),
.B(n_221),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_163),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_242),
.A2(n_204),
.B(n_203),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_225),
.B(n_164),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_250),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g245 ( 
.A1(n_210),
.A2(n_207),
.B1(n_203),
.B2(n_206),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_245),
.A2(n_204),
.B1(n_210),
.B2(n_205),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_193),
.C(n_175),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_255),
.C(n_257),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_189),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_200),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_254),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_199),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_229),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_175),
.C(n_165),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_194),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_211),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_201),
.B(n_213),
.Y(n_257)
);

NAND3xp33_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_197),
.C(n_228),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_259),
.B(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_260),
.Y(n_292)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_269),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_264),
.A2(n_266),
.B(n_248),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_265),
.A2(n_252),
.B(n_231),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_257),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_271),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_222),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_224),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_245),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_280),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_237),
.A2(n_196),
.B1(n_209),
.B2(n_208),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_277),
.A2(n_242),
.B1(n_237),
.B2(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

BUFx12_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_233),
.B(n_165),
.Y(n_280)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_277),
.A2(n_258),
.B1(n_275),
.B2(n_274),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_284),
.B1(n_295),
.B2(n_276),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_272),
.B1(n_266),
.B2(n_273),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_279),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_173),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_230),
.C(n_241),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_296),
.C(n_297),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_240),
.Y(n_304)
);

BUFx12_ASAP7_75t_L g291 ( 
.A(n_260),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_291),
.B(n_198),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_273),
.A2(n_269),
.B1(n_252),
.B2(n_264),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_262),
.B(n_234),
.C(n_253),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_240),
.C(n_239),
.Y(n_297)
);

AO21x1_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_268),
.B(n_267),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_263),
.C(n_270),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_307),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_263),
.C(n_295),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_302),
.B(n_303),
.C(n_308),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_265),
.C(n_261),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_306),
.Y(n_328)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_270),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_267),
.C(n_268),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_311),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_278),
.B(n_271),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_292),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_281),
.C(n_293),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_281),
.B(n_229),
.C(n_202),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_313),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_287),
.A2(n_197),
.B1(n_198),
.B2(n_249),
.Y(n_313)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_314),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_301),
.A2(n_289),
.B(n_293),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_317),
.A2(n_320),
.B(n_322),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_307),
.B(n_290),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_318),
.B(n_327),
.Y(n_333)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_308),
.B(n_290),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_303),
.A2(n_302),
.B1(n_315),
.B2(n_292),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_282),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_315),
.B(n_283),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_331),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_317),
.A2(n_291),
.B(n_290),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_305),
.C(n_288),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_291),
.Y(n_332)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_319),
.A2(n_288),
.B(n_285),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_334),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_325),
.B(n_288),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_335),
.B(n_336),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_321),
.B(n_249),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_326),
.B(n_151),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_338),
.A2(n_217),
.B(n_211),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_333),
.A2(n_316),
.B(n_328),
.Y(n_340)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_340),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_343),
.Y(n_348)
);

OAI211xp5_ASAP7_75t_L g344 ( 
.A1(n_332),
.A2(n_324),
.B(n_328),
.C(n_8),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_344),
.A2(n_345),
.B(n_13),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_337),
.A2(n_330),
.B1(n_151),
.B2(n_4),
.Y(n_345)
);

NOR2xp67_ASAP7_75t_SL g347 ( 
.A(n_341),
.B(n_10),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_347),
.A2(n_349),
.B(n_350),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_0),
.C(n_1),
.Y(n_350)
);

AOI322xp5_ASAP7_75t_L g351 ( 
.A1(n_348),
.A2(n_346),
.A3(n_342),
.B1(n_340),
.B2(n_345),
.C1(n_350),
.C2(n_3),
.Y(n_351)
);

O2A1O1Ixp33_ASAP7_75t_L g353 ( 
.A1(n_351),
.A2(n_2),
.B(n_3),
.C(n_352),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_353),
.B(n_3),
.Y(n_354)
);


endmodule