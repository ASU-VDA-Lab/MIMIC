module fake_jpeg_18662_n_128 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_128);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_128;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_14),
.B(n_0),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_30),
.Y(n_42)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_14),
.B(n_1),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_6),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_12),
.B(n_10),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_2),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_35),
.A2(n_15),
.B1(n_20),
.B2(n_26),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_17),
.B(n_3),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_3),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_3),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_18),
.B1(n_24),
.B2(n_21),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_62),
.B1(n_35),
.B2(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_53),
.Y(n_67)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_28),
.A2(n_24),
.B1(n_18),
.B2(n_21),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_48),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_75)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_30),
.B(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_55),
.Y(n_66)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_26),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_57),
.B(n_61),
.Y(n_77)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_15),
.B1(n_19),
.B2(n_22),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_70),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_4),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_42),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_71),
.B(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_46),
.B1(n_55),
.B2(n_59),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_58),
.B(n_41),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_76),
.B(n_77),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_43),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_78),
.A2(n_52),
.B(n_47),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_52),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_86),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_51),
.B(n_49),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_89),
.Y(n_102)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_56),
.Y(n_85)
);

BUFx12_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_87),
.A2(n_90),
.B1(n_63),
.B2(n_69),
.Y(n_101)
);

AO22x2_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_49),
.B1(n_79),
.B2(n_75),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_94),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_100),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_93),
.B(n_79),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_84),
.B1(n_90),
.B2(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_90),
.B(n_65),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_108),
.Y(n_114)
);

AO21x1_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_89),
.B(n_84),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_91),
.C(n_92),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_96),
.C(n_97),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_90),
.B1(n_83),
.B2(n_65),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_102),
.B(n_104),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_105),
.Y(n_119)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_97),
.B(n_102),
.Y(n_115)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_97),
.C(n_106),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_109),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_114),
.C(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_122),
.B(n_69),
.C(n_95),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_120),
.A2(n_108),
.B(n_103),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_123),
.B(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_124),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_126),
.A2(n_125),
.B(n_68),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_127),
.B(n_74),
.Y(n_128)
);


endmodule