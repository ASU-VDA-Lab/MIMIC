module fake_jpeg_13211_n_154 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_154);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_154;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_0),
.B(n_29),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_7),
.B(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_32),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_1),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_74),
.Y(n_86)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_72),
.B(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_2),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_66),
.Y(n_84)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_77),
.Y(n_80)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_71),
.A2(n_63),
.B1(n_47),
.B2(n_58),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_78),
.A2(n_83),
.B1(n_91),
.B2(n_92),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_67),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_87),
.C(n_50),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_68),
.A2(n_63),
.B1(n_65),
.B2(n_59),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_60),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_49),
.B1(n_56),
.B2(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_90),
.A2(n_50),
.B1(n_3),
.B2(n_4),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_76),
.A2(n_62),
.B1(n_61),
.B2(n_48),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_76),
.A2(n_54),
.B1(n_46),
.B2(n_45),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_57),
.B1(n_52),
.B2(n_4),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_7),
.B(n_8),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_21),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_96),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_89),
.B1(n_82),
.B2(n_88),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_100),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_88),
.B(n_5),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_9),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_10),
.Y(n_104)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_81),
.B(n_10),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g119 ( 
.A(n_106),
.B(n_24),
.Y(n_119)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_12),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_13),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_30),
.Y(n_129)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_97),
.A2(n_50),
.B(n_16),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_115),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_14),
.B(n_19),
.Y(n_115)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_22),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_129),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_120),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_111),
.B(n_27),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_40),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_110),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_114),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_131),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_128),
.A2(n_105),
.B1(n_95),
.B2(n_36),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_123),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_137),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_141),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_122),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_138),
.C(n_134),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_143),
.A2(n_127),
.A3(n_137),
.B1(n_133),
.B2(n_118),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_147),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_149),
.A2(n_146),
.B(n_145),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_150),
.B(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_151),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_148),
.C(n_142),
.Y(n_153)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);


endmodule