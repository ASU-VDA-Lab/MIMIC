module fake_jpeg_1113_n_589 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_589);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_589;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx24_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

CKINVDCx5p33_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_8),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_5),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_15),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_58),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_59),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_62),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_63),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_46),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_64),
.B(n_79),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_66),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_67),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_68),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_69),
.Y(n_129)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_22),
.Y(n_70)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx8_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_17),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_72),
.B(n_4),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_73),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_77),
.Y(n_134)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g154 ( 
.A(n_78),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_33),
.B(n_1),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_80),
.Y(n_132)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_86),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

BUFx4f_ASAP7_75t_SL g188 ( 
.A(n_88),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_33),
.B(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_91),
.B(n_99),
.Y(n_164)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_34),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_97),
.Y(n_151)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_33),
.B(n_2),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_45),
.Y(n_101)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_102),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_51),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_103),
.B(n_25),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_32),
.Y(n_105)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_106),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_109),
.Y(n_173)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_53),
.Y(n_110)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_37),
.Y(n_113)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_21),
.Y(n_114)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_114),
.Y(n_177)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_21),
.Y(n_115)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_37),
.Y(n_116)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_52),
.Y(n_120)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_121),
.B(n_125),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_36),
.B(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_122),
.B(n_127),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_124),
.Y(n_182)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_41),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_52),
.Y(n_126)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_36),
.B(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_64),
.B(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_128),
.B(n_157),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_40),
.B1(n_52),
.B2(n_57),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_152),
.A2(n_155),
.B1(n_162),
.B2(n_178),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_79),
.A2(n_40),
.B1(n_57),
.B2(n_35),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_91),
.B(n_27),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_99),
.A2(n_27),
.B1(n_50),
.B2(n_49),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_168),
.B(n_7),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_107),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_176),
.B(n_7),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_60),
.A2(n_54),
.B1(n_48),
.B2(n_44),
.Y(n_178)
);

OA22x2_ASAP7_75t_L g179 ( 
.A1(n_71),
.A2(n_54),
.B1(n_48),
.B2(n_38),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_SL g230 ( 
.A1(n_179),
.A2(n_42),
.B(n_9),
.C(n_10),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_69),
.A2(n_44),
.B1(n_43),
.B2(n_55),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_181),
.A2(n_199),
.B(n_201),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_185),
.B(n_202),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_61),
.A2(n_20),
.B1(n_50),
.B2(n_49),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_187),
.A2(n_193),
.B1(n_200),
.B2(n_7),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_126),
.A2(n_43),
.B1(n_20),
.B2(n_35),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_70),
.B(n_55),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_206),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_97),
.A2(n_119),
.B1(n_30),
.B2(n_25),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_124),
.A2(n_30),
.B1(n_23),
.B2(n_41),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_63),
.A2(n_23),
.B1(n_47),
.B2(n_41),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_65),
.B(n_4),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_67),
.Y(n_203)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_120),
.B(n_47),
.C(n_42),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_7),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_68),
.B(n_73),
.Y(n_206)
);

INVx6_ASAP7_75t_SL g207 ( 
.A(n_76),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_209),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_82),
.B(n_5),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_212),
.B(n_214),
.Y(n_252)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_88),
.B(n_5),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_93),
.A2(n_117),
.B1(n_112),
.B2(n_111),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_216),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g219 ( 
.A1(n_216),
.A2(n_101),
.B1(n_96),
.B2(n_95),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_219),
.A2(n_256),
.B1(n_259),
.B2(n_270),
.Y(n_298)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_220),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_221),
.B(n_235),
.Y(n_314)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_150),
.Y(n_222)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_222),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g317 ( 
.A(n_223),
.Y(n_317)
);

CKINVDCx6p67_ASAP7_75t_R g224 ( 
.A(n_180),
.Y(n_224)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_224),
.Y(n_299)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_129),
.Y(n_225)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_130),
.A2(n_47),
.B(n_42),
.C(n_10),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_226),
.B(n_227),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_210),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_229),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_230),
.A2(n_278),
.B1(n_288),
.B2(n_290),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_231),
.Y(n_309)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_140),
.Y(n_232)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_232),
.Y(n_304)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_131),
.Y(n_233)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_233),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_234),
.B(n_236),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_147),
.Y(n_237)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_197),
.Y(n_238)
);

INVx4_ASAP7_75t_L g344 ( 
.A(n_238),
.Y(n_344)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_158),
.Y(n_239)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_239),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_136),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_240),
.B(n_246),
.Y(n_345)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_129),
.Y(n_242)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_242),
.Y(n_301)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_165),
.Y(n_243)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_151),
.Y(n_245)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_245),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_183),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_132),
.Y(n_247)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_197),
.Y(n_249)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_9),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_250),
.B(n_264),
.Y(n_312)
);

AND2x2_ASAP7_75t_SL g254 ( 
.A(n_194),
.B(n_9),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_254),
.B(n_153),
.C(n_161),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_134),
.Y(n_255)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_255),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_184),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_133),
.Y(n_257)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_257),
.Y(n_305)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_138),
.Y(n_258)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_171),
.Y(n_260)
);

BUFx2_ASAP7_75t_SL g351 ( 
.A(n_260),
.Y(n_351)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_177),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_261),
.Y(n_337)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_198),
.Y(n_263)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_263),
.Y(n_327)
);

AOI32xp33_ASAP7_75t_L g264 ( 
.A1(n_130),
.A2(n_13),
.A3(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_264)
);

INVx4_ASAP7_75t_SL g266 ( 
.A(n_173),
.Y(n_266)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_186),
.Y(n_267)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

BUFx12_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_268),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_164),
.B(n_16),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_269),
.B(n_271),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_164),
.A2(n_13),
.B1(n_14),
.B2(n_214),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_160),
.B(n_14),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

INVx6_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_139),
.Y(n_275)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_144),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_276),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_212),
.B(n_208),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_277),
.B(n_279),
.Y(n_332)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_178),
.A2(n_14),
.B1(n_201),
.B2(n_181),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_179),
.B(n_154),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_141),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_283),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_134),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_281),
.Y(n_333)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_137),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_282),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_149),
.B(n_166),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_285),
.Y(n_341)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_135),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_179),
.B(n_154),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_286),
.A2(n_191),
.B1(n_189),
.B2(n_146),
.Y(n_313)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_142),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_188),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_174),
.B(n_172),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_289),
.Y(n_324)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_148),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_143),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_156),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_175),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_182),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_294),
.A2(n_145),
.B1(n_148),
.B2(n_204),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_145),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_295),
.A2(n_211),
.B1(n_224),
.B2(n_223),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_252),
.A2(n_253),
.B1(n_244),
.B2(n_228),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_300),
.A2(n_321),
.B1(n_328),
.B2(n_346),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_313),
.B(n_281),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_SL g318 ( 
.A(n_250),
.B(n_199),
.C(n_192),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_318),
.B(n_326),
.C(n_251),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_319),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_259),
.A2(n_215),
.B1(n_196),
.B2(n_163),
.Y(n_321)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_262),
.B(n_137),
.C(n_217),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_219),
.A2(n_204),
.B1(n_143),
.B2(n_159),
.Y(n_328)
);

AOI32xp33_ASAP7_75t_L g336 ( 
.A1(n_226),
.A2(n_153),
.A3(n_159),
.B1(n_161),
.B2(n_190),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_238),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_340),
.B(n_268),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_230),
.A2(n_217),
.B1(n_190),
.B2(n_211),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_347),
.Y(n_387)
);

OA21x2_ASAP7_75t_L g352 ( 
.A1(n_339),
.A2(n_300),
.B(n_328),
.Y(n_352)
);

AO21x2_ASAP7_75t_L g399 ( 
.A1(n_352),
.A2(n_354),
.B(n_331),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_254),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_364),
.Y(n_397)
);

OA22x2_ASAP7_75t_L g354 ( 
.A1(n_338),
.A2(n_278),
.B1(n_261),
.B2(n_241),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_393),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_345),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_361),
.Y(n_408)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_297),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_358),
.Y(n_417)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_298),
.A2(n_343),
.B1(n_309),
.B2(n_338),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_360),
.A2(n_367),
.B(n_373),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_348),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_320),
.Y(n_362)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_363),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_221),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_302),
.Y(n_365)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_348),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_369),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_299),
.A2(n_249),
.B1(n_239),
.B2(n_284),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_248),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_372),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_343),
.A2(n_275),
.B(n_260),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_389),
.B1(n_392),
.B2(n_394),
.Y(n_398)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_310),
.Y(n_375)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_310),
.Y(n_376)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_322),
.Y(n_377)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_377),
.Y(n_425)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_322),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_378),
.B(n_383),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_334),
.B(n_233),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_390),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_321),
.A2(n_265),
.B1(n_273),
.B2(n_272),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_380),
.A2(n_385),
.B1(n_299),
.B2(n_349),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_381),
.A2(n_382),
.B1(n_384),
.B2(n_351),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_L g382 ( 
.A1(n_350),
.A2(n_267),
.B1(n_290),
.B2(n_243),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_296),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g384 ( 
.A1(n_333),
.A2(n_311),
.B1(n_297),
.B2(n_330),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_340),
.A2(n_266),
.B1(n_255),
.B2(n_242),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_296),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_386),
.B(n_388),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_341),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_312),
.A2(n_282),
.B1(n_225),
.B2(n_263),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_318),
.A2(n_224),
.B(n_292),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_303),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_391),
.B(n_349),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_312),
.A2(n_274),
.B1(n_293),
.B2(n_245),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_314),
.A2(n_268),
.B1(n_325),
.B2(n_308),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_396),
.B(n_370),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_399),
.A2(n_355),
.B1(n_354),
.B2(n_389),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_364),
.C(n_357),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_411),
.C(n_412),
.Y(n_445)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_404),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_353),
.B(n_369),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g447 ( 
.A(n_406),
.B(n_410),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_393),
.B(n_324),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_360),
.B(n_305),
.C(n_327),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_352),
.B(n_342),
.C(n_323),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_352),
.A2(n_311),
.B1(n_337),
.B2(n_315),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_416),
.A2(n_355),
.B1(n_385),
.B2(n_380),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g418 ( 
.A(n_352),
.B(n_303),
.C(n_337),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_418),
.B(n_423),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_315),
.C(n_335),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_379),
.Y(n_424)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_427),
.C(n_316),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_316),
.Y(n_427)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_428),
.Y(n_453)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_354),
.A2(n_374),
.B1(n_381),
.B2(n_371),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_429),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_419),
.Y(n_430)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_431),
.A2(n_440),
.B1(n_407),
.B2(n_400),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_392),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_432),
.B(n_448),
.C(n_418),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_420),
.A2(n_390),
.B(n_387),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_433),
.A2(n_438),
.B(n_450),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_408),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_434),
.B(n_446),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_410),
.B(n_359),
.Y(n_435)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_406),
.C(n_411),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_437),
.B1(n_439),
.B2(n_443),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_420),
.A2(n_354),
.B(n_394),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_398),
.A2(n_354),
.B1(n_366),
.B2(n_361),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_399),
.A2(n_362),
.B1(n_358),
.B2(n_383),
.Y(n_440)
);

AOI22x1_ASAP7_75t_L g443 ( 
.A1(n_399),
.A2(n_368),
.B1(n_386),
.B2(n_378),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_402),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_428),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_449),
.B(n_452),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_395),
.A2(n_413),
.B(n_398),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_395),
.A2(n_306),
.B(n_377),
.Y(n_451)
);

AO21x1_ASAP7_75t_L g484 ( 
.A1(n_451),
.A2(n_461),
.B(n_407),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_422),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_421),
.Y(n_454)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_454),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_396),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_457),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_397),
.B(n_391),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_425),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_403),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_403),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_405),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_423),
.Y(n_460)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_460),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_412),
.B(n_376),
.Y(n_461)
);

XOR2x2_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_397),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_462),
.B(n_463),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_464),
.B(n_473),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_439),
.A2(n_399),
.B1(n_416),
.B2(n_401),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_467),
.A2(n_431),
.B1(n_440),
.B2(n_442),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g470 ( 
.A(n_434),
.B(n_400),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_470),
.A2(n_485),
.B1(n_443),
.B2(n_454),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_445),
.B(n_426),
.C(n_425),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_472),
.B(n_477),
.C(n_478),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_399),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_487),
.Y(n_504)
);

OA21x2_ASAP7_75t_L g476 ( 
.A1(n_437),
.A2(n_405),
.B(n_414),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_476),
.A2(n_484),
.B(n_489),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_445),
.B(n_414),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_409),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_409),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_482),
.B(n_488),
.C(n_490),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_446),
.Y(n_486)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_486),
.Y(n_491)
);

INVxp33_ASAP7_75t_SL g487 ( 
.A(n_450),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_456),
.B(n_375),
.Y(n_488)
);

FAx1_ASAP7_75t_L g489 ( 
.A(n_438),
.B(n_417),
.CI(n_372),
.CON(n_489),
.SN(n_489)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_365),
.C(n_306),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_489),
.A2(n_441),
.B1(n_455),
.B2(n_453),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_493),
.A2(n_497),
.B1(n_499),
.B2(n_508),
.Y(n_520)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_474),
.Y(n_494)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_494),
.Y(n_527)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_474),
.Y(n_495)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_495),
.Y(n_530)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_481),
.Y(n_496)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_496),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_489),
.A2(n_441),
.B1(n_485),
.B2(n_481),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_465),
.A2(n_453),
.B1(n_461),
.B2(n_442),
.Y(n_499)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_480),
.Y(n_502)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_502),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_477),
.B(n_444),
.C(n_433),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_513),
.C(n_462),
.Y(n_516)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_483),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_505),
.B(n_506),
.Y(n_521)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_507),
.A2(n_510),
.B1(n_512),
.B2(n_514),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_469),
.A2(n_444),
.B1(n_457),
.B2(n_451),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_476),
.Y(n_509)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_509),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_476),
.A2(n_443),
.B1(n_458),
.B2(n_459),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_472),
.B(n_344),
.C(n_417),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_466),
.A2(n_401),
.B1(n_363),
.B2(n_344),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_516),
.B(n_519),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_496),
.A2(n_469),
.B1(n_471),
.B2(n_484),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_517),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_498),
.B(n_464),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g522 ( 
.A(n_504),
.B(n_468),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_523),
.C(n_525),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_513),
.B(n_490),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_499),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_524),
.B(n_497),
.Y(n_545)
);

NAND2xp33_ASAP7_75t_R g525 ( 
.A(n_501),
.B(n_478),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_507),
.A2(n_473),
.B1(n_482),
.B2(n_475),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_526),
.A2(n_508),
.B1(n_517),
.B2(n_504),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_500),
.B(n_471),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_528),
.B(n_529),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_498),
.B(n_488),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_528),
.B(n_503),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_533),
.B(n_540),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_521),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_534),
.B(n_535),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_492),
.C(n_529),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_520),
.A2(n_495),
.B1(n_494),
.B2(n_491),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_537),
.B(n_538),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_492),
.C(n_500),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_SL g542 ( 
.A1(n_515),
.A2(n_511),
.B(n_531),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_542),
.A2(n_493),
.B(n_510),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_SL g543 ( 
.A(n_520),
.B(n_511),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_543),
.B(n_545),
.Y(n_550)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_521),
.Y(n_544)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_544),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g546 ( 
.A1(n_531),
.A2(n_509),
.B1(n_491),
.B2(n_514),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_527),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_536),
.A2(n_542),
.B(n_533),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_549),
.B(n_552),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_R g551 ( 
.A(n_543),
.B(n_530),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_551),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_518),
.C(n_515),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_539),
.B(n_530),
.C(n_527),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_546),
.C(n_541),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_556),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_538),
.B(n_522),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_559),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_547),
.B(n_532),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_552),
.B(n_539),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_562),
.B(n_568),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_565),
.B(n_548),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g566 ( 
.A1(n_560),
.A2(n_532),
.B1(n_505),
.B2(n_502),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_566),
.B(n_570),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_555),
.B(n_541),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_557),
.B(n_506),
.Y(n_569)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_569),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_467),
.C(n_363),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_565),
.B(n_550),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_571),
.B(n_572),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_564),
.B(n_550),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_575),
.B(n_576),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_561),
.B(n_548),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_SL g578 ( 
.A1(n_575),
.A2(n_563),
.B(n_556),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g582 ( 
.A1(n_578),
.A2(n_579),
.B(n_573),
.Y(n_582)
);

NOR3xp33_ASAP7_75t_L g579 ( 
.A(n_577),
.B(n_563),
.C(n_567),
.Y(n_579)
);

OAI31xp33_ASAP7_75t_SL g584 ( 
.A1(n_582),
.A2(n_583),
.A3(n_581),
.B(n_551),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_L g583 ( 
.A1(n_580),
.A2(n_574),
.B(n_567),
.Y(n_583)
);

MAJx2_ASAP7_75t_L g586 ( 
.A(n_584),
.B(n_585),
.C(n_329),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_582),
.A2(n_570),
.B(n_329),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_586),
.A2(n_317),
.B(n_320),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_587),
.B(n_307),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g589 ( 
.A(n_588),
.B(n_307),
.Y(n_589)
);


endmodule