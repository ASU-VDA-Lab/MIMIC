module real_jpeg_11917_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_313, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_313;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g85 ( 
.A(n_0),
.Y(n_85)
);

BUFx16f_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_45),
.B1(n_50),
.B2(n_55),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_55),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_5),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_5),
.B(n_45),
.C(n_49),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g134 ( 
.A(n_5),
.B(n_31),
.Y(n_134)
);

OAI21xp33_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_141),
.B(n_144),
.Y(n_161)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_5),
.A2(n_27),
.B(n_30),
.C(n_172),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_126),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_5),
.B(n_60),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_6),
.A2(n_45),
.B1(n_50),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_6),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_143),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_143),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_6),
.A2(n_60),
.B1(n_61),
.B2(n_143),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_7),
.A2(n_40),
.B1(n_45),
.B2(n_50),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_9),
.A2(n_60),
.B1(n_61),
.B2(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_69),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_9),
.A2(n_45),
.B1(n_50),
.B2(n_69),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_69),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_10),
.A2(n_45),
.B1(n_50),
.B2(n_138),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_138),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_10),
.A2(n_60),
.B1(n_61),
.B2(n_138),
.Y(n_245)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_12),
.A2(n_60),
.B1(n_61),
.B2(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_12),
.A2(n_45),
.B1(n_50),
.B2(n_62),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_62),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_12),
.A2(n_28),
.B1(n_30),
.B2(n_62),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_13),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_14),
.A2(n_60),
.B1(n_61),
.B2(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_14),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_14),
.A2(n_32),
.B1(n_33),
.B2(n_97),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_45),
.B1(n_50),
.B2(n_97),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_97),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_28),
.B1(n_30),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_15),
.A2(n_37),
.B1(n_60),
.B2(n_61),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_15),
.A2(n_37),
.B1(n_45),
.B2(n_50),
.Y(n_235)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_111),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_109),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_20),
.B(n_98),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_71),
.C(n_79),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_21),
.B(n_71),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_57),
.B1(n_58),
.B2(n_70),
.Y(n_21)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_23),
.B(n_42),
.C(n_58),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_24),
.B(n_179),
.Y(n_193)
);

NOR2x1_ASAP7_75t_R g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_26),
.A2(n_32),
.B(n_126),
.Y(n_172)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_28),
.A2(n_30),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g231 ( 
.A(n_28),
.B(n_65),
.Y(n_231)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_30),
.A2(n_61),
.A3(n_66),
.B1(n_218),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_31),
.B(n_179),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_32),
.A2(n_33),
.B1(n_48),
.B2(n_49),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_33),
.B(n_130),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_36),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_72)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_39),
.A2(n_73),
.B1(n_75),
.B2(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_41),
.A2(n_42),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_51),
.B(n_53),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_43),
.A2(n_51),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_43),
.B(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_43),
.A2(n_51),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_43),
.A2(n_51),
.B1(n_224),
.B2(n_252),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_43),
.A2(n_51),
.B1(n_90),
.B2(n_252),
.Y(n_258)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_54),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_44),
.A2(n_137),
.B(n_139),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_44),
.B(n_126),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_44),
.A2(n_139),
.B(n_223),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_44)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_50),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_50),
.B(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_51),
.B(n_128),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_57),
.A2(n_58),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_64),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_60),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_67)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

O2A1O1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_61),
.A2(n_63),
.B(n_126),
.C(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_63),
.A2(n_64),
.B1(n_245),
.B2(n_265),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_63),
.A2(n_265),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_64),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_64),
.B(n_96),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_64),
.A2(n_93),
.B(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_71),
.A2(n_72),
.B(n_76),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_73),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_73),
.A2(n_75),
.B1(n_192),
.B2(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_73),
.A2(n_178),
.B(n_221),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_267),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_75),
.A2(n_192),
.B(n_193),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_75),
.A2(n_193),
.B(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_77),
.A2(n_125),
.B(n_127),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_77),
.A2(n_127),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_79),
.B(n_309),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B(n_92),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_80),
.A2(n_81),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_82),
.A2(n_83),
.B1(n_92),
.B2(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_84),
.A2(n_85),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_84),
.B(n_145),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_84),
.A2(n_85),
.B1(n_235),
.B2(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_85),
.B(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_85),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_87),
.A2(n_141),
.B1(n_158),
.B2(n_261),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_92),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_108),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_307),
.B(n_311),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_294),
.B(n_306),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_277),
.B(n_293),
.Y(n_115)
);

OAI321xp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_237),
.A3(n_270),
.B1(n_275),
.B2(n_276),
.C(n_313),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_209),
.B(n_236),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_186),
.B(n_208),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_167),
.B(n_185),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_146),
.B(n_166),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_131),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_122),
.B(n_131),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_129),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_123),
.A2(n_124),
.B1(n_129),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_126),
.B(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_140),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_136),
.C(n_140),
.Y(n_168)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_137),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B(n_144),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_141),
.A2(n_158),
.B1(n_174),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_141),
.A2(n_158),
.B1(n_200),
.B2(n_234),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_154),
.B(n_165),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_148),
.B(n_152),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_150),
.A2(n_158),
.B(n_159),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_160),
.B(n_164),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_156),
.B(n_157),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_159),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_168),
.B(n_169),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_175),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_180),
.C(n_184),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_173),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_175)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_187),
.B(n_188),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_201),
.B2(n_202),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_204),
.C(n_206),
.Y(n_210)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_195),
.C(n_199),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_198),
.B2(n_199),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_203),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_204),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_210),
.B(n_211),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_226),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_227),
.C(n_228),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_219),
.B2(n_225),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_220),
.C(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_219),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_228),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_233),
.Y(n_247)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_254),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_254),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_248),
.C(n_253),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_239),
.A2(n_240),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_247),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_246),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_246),
.C(n_247),
.Y(n_269)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_248),
.B(n_253),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_251),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_250),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_269),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_262),
.C(n_269),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_260),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_266),
.C(n_268),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_271),
.B(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_292),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_292),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_282),
.C(n_283),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_290),
.B2(n_291),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.C(n_291),
.Y(n_305)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_296),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_305),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_300),
.C(n_305),
.Y(n_310)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_310),
.Y(n_311)
);


endmodule