module real_jpeg_4006_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_1),
.Y(n_174)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_2),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_2),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_2),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_3),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_3),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_3),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_3),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_3),
.B(n_88),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_273),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_4),
.B(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_4),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_4),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_4),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_4),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_4),
.B(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_6),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_6),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_6),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_6),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_6),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_6),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_7),
.B(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_7),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_7),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_7),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_7),
.B(n_46),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_7),
.B(n_88),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_7),
.B(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_9),
.Y(n_74)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_9),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_9),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g282 ( 
.A(n_9),
.Y(n_282)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_10),
.B(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_10),
.B(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_10),
.B(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_12),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_71),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_12),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g137 ( 
.A(n_12),
.B(n_138),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_12),
.B(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_13),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_14),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_14),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g157 ( 
.A(n_14),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_14),
.B(n_166),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_15),
.Y(n_98)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_15),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_195),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_193),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_144),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_19),
.B(n_144),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_92),
.C(n_129),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_20),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_62),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_21),
.B(n_63),
.C(n_78),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_41),
.C(n_52),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_22),
.B(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_28),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_23),
.B(n_29),
.C(n_40),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_27),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_34),
.B2(n_40),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_31),
.B(n_66),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_33),
.Y(n_139)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_33),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_33),
.Y(n_237)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g142 ( 
.A(n_39),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_39),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_39),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_41),
.A2(n_52),
.B1(n_53),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_41),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.C(n_49),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_42),
.A2(n_49),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_42),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_45),
.B(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_49),
.Y(n_205)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_50),
.Y(n_217)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_51),
.Y(n_153)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_57),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_54),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_54),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_54),
.A2(n_57),
.B1(n_58),
.B2(n_156),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_55),
.Y(n_247)
);

INVx8_ASAP7_75t_L g271 ( 
.A(n_55),
.Y(n_271)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_56),
.Y(n_280)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_78),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_65),
.B(n_69),
.C(n_76),
.Y(n_192)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_69),
.A2(n_70),
.B1(n_119),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_70),
.B(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_74),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_86),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_81),
.B(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_79),
.B(n_87),
.C(n_89),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_83),
.Y(n_81)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_92),
.B(n_129),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_111),
.C(n_116),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_93),
.B(n_111),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_107),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_100),
.B2(n_106),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_95),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_100),
.C(n_107),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_105),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_113),
.B(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_116),
.B(n_200),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_123),
.C(n_126),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_117),
.A2(n_118),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_119),
.Y(n_298)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_123),
.A2(n_124),
.B1(n_126),
.B2(n_127),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_143),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_132),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_136),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_162),
.C(n_163),
.Y(n_161)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_140),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_137),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_177),
.C(n_178),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_175),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_160),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_157),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_157),
.A2(n_159),
.B1(n_254),
.B2(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_157),
.B(n_256),
.Y(n_299)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_158),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.Y(n_164)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_173),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_172),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_192),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_186),
.B1(n_190),
.B2(n_191),
.Y(n_182)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_183),
.Y(n_190)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_189),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_225),
.B(n_323),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_223),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_198),
.B(n_223),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.C(n_220),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_199),
.B(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_201),
.B(n_220),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.C(n_218),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_202),
.B(n_314),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_206),
.A2(n_218),
.B1(n_219),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_206),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.C(n_214),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_207),
.A2(n_208),
.B1(n_214),
.B2(n_215),
.Y(n_303)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_211),
.B(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_318),
.B(n_322),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_305),
.B(n_317),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_291),
.B(n_304),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_265),
.B(n_290),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_257),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_231),
.B(n_257),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_243),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_232),
.B(n_244),
.C(n_253),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_233),
.B(n_239),
.C(n_240),
.Y(n_301)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_248),
.Y(n_258)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.C(n_263),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_258),
.B(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_259),
.A2(n_263),
.B1(n_264),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_259),
.Y(n_288)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_284),
.B(n_289),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_276),
.B(n_283),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_268),
.B(n_275),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_275),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_272),
.Y(n_285)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_SL g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_281),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_285),
.B(n_286),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_300),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_301),
.C(n_302),
.Y(n_316)
);

FAx1_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_297),
.CI(n_299),
.CON(n_294),
.SN(n_294)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_316),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_316),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_313),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_310),
.C(n_313),
.Y(n_319)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_311),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_320),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);


endmodule