module fake_jpeg_28421_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx4f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_21),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g58 ( 
.A(n_19),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_1),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_68),
.Y(n_72)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_2),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_2),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g70 ( 
.A(n_56),
.Y(n_70)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_57),
.B1(n_42),
.B2(n_45),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_52),
.B1(n_55),
.B2(n_54),
.Y(n_99)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_61),
.B(n_60),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_82),
.B(n_51),
.C(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_81),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_50),
.B1(n_61),
.B2(n_60),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_86),
.A2(n_99),
.B1(n_58),
.B2(n_47),
.Y(n_100)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_46),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_3),
.Y(n_107)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_95),
.Y(n_105)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_100),
.B(n_102),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_3),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_87),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_85),
.Y(n_114)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_33),
.C(n_40),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_113),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_91),
.B1(n_88),
.B2(n_96),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_111),
.A2(n_112),
.B1(n_105),
.B2(n_109),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_96),
.B1(n_85),
.B2(n_62),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_5),
.Y(n_128)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_39),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_123),
.B1(n_127),
.B2(n_122),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_120),
.Y(n_131)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_44),
.B1(n_48),
.B2(n_6),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_25),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_126),
.B(n_129),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_115),
.A2(n_29),
.B(n_38),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_115),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_132),
.B(n_135),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_119),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_131),
.C(n_134),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_137),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_136),
.B(n_130),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_125),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_140),
.A2(n_15),
.B1(n_16),
.B2(n_22),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_24),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_142),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_30),
.B(n_31),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_36),
.Y(n_145)
);


endmodule