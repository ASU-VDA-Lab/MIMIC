module real_jpeg_15914_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AND2x2_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_0),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_0),
.B(n_120),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_0),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_0),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_0),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_0),
.B(n_137),
.Y(n_410)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_1),
.Y(n_416)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_2),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_2),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_2),
.Y(n_344)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_2),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_3),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_3),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_36),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_4),
.B(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_4),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_4),
.B(n_418),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_5),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_5),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_6),
.B(n_61),
.Y(n_60)
);

AND2x4_ASAP7_75t_SL g76 ( 
.A(n_6),
.B(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_6),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_6),
.B(n_134),
.Y(n_146)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_6),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_6),
.B(n_393),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_7),
.Y(n_135)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_7),
.Y(n_202)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_7),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_8),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_8),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_8),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_8),
.B(n_69),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_8),
.B(n_41),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_8),
.B(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_8),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_9),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_9),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_9),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_9),
.B(n_199),
.Y(n_325)
);

BUFx2_ASAP7_75t_R g345 ( 
.A(n_9),
.Y(n_345)
);

NAND2x1_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_28),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_10),
.B(n_79),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_10),
.B(n_72),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_10),
.B(n_220),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_10),
.B(n_298),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_11),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g228 ( 
.A(n_11),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_12),
.B(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_12),
.A2(n_15),
.B1(n_41),
.B2(n_45),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_12),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_12),
.B(n_123),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_12),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_12),
.B(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_13),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_14),
.Y(n_99)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_15),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_15),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_15),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_15),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_15),
.B(n_67),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_15),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_15),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_15),
.B(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_16),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_381),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_210),
.B(n_380),
.Y(n_18)
);

AND2x2_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_166),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_20),
.B(n_166),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_89),
.Y(n_20)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_21),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_64),
.C(n_81),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_23),
.B(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.C(n_50),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_24),
.B(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_27),
.B(n_32),
.C(n_35),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_27),
.B(n_160),
.Y(n_425)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_34),
.Y(n_352)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_38),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_39),
.A2(n_40),
.B1(n_50),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_40),
.A2(n_231),
.B(n_235),
.Y(n_230)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_49),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_49),
.Y(n_399)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_50),
.Y(n_264)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_56),
.C(n_60),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_51),
.A2(n_52),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_51),
.A2(n_52),
.B1(n_60),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

MAJx2_ASAP7_75t_L g426 ( 
.A(n_52),
.B(n_94),
.C(n_101),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_56),
.B(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_58),
.Y(n_121)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_59),
.Y(n_144)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_60),
.Y(n_181)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_63),
.Y(n_221)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_63),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_64),
.A2(n_81),
.B1(n_82),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_75),
.C(n_77),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_65),
.B(n_205),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_68),
.C(n_71),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_66),
.A2(n_71),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_66),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_66),
.B(n_278),
.Y(n_277)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_67),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_68),
.B(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_71),
.Y(n_243)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_73),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_77),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_80),
.Y(n_234)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_80),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2x1_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_88),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_84),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_84),
.B(n_218),
.C(n_224),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_84),
.A2(n_156),
.B1(n_224),
.B2(n_225),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_88),
.B(n_155),
.C(n_156),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_125),
.B1(n_164),
.B2(n_165),
.Y(n_89)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_90),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_106),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_91),
.B(n_107),
.C(n_113),
.Y(n_431)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_94),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g400 ( 
.A1(n_94),
.A2(n_105),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_95),
.B(n_403),
.Y(n_402)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_99),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_101),
.B1(n_112),
.B2(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_108),
.C(n_112),
.Y(n_107)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_114),
.B(n_119),
.C(n_122),
.Y(n_408)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_122),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_125),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_153),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_126),
.B(n_154),
.C(n_157),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.C(n_145),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_130),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.C(n_141),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_136),
.A2(n_141),
.B1(n_142),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_141),
.B(n_251),
.C(n_254),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_141),
.A2(n_142),
.B1(n_251),
.B2(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_143),
.Y(n_281)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_148),
.C(n_152),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.Y(n_153)
);

XNOR2x1_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_158),
.B(n_163),
.C(n_430),
.Y(n_429)
);

XNOR2x1_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_160),
.Y(n_430)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_164),
.B(n_385),
.C(n_386),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.C(n_175),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_168),
.A2(n_169),
.B1(n_172),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_172),
.Y(n_271)
);

XOR2x2_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_176),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_203),
.C(n_207),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_177),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_182),
.C(n_192),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2x1_ASAP7_75t_L g257 ( 
.A(n_179),
.B(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_182),
.B(n_192),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_183),
.B(n_189),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.C(n_198),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_193),
.A2(n_197),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_193),
.Y(n_247)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_197),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_197),
.B(n_322),
.C(n_324),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_197),
.A2(n_248),
.B1(n_324),
.B2(n_325),
.Y(n_335)
);

XOR2x1_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_204),
.B(n_207),
.Y(n_266)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_376),
.Y(n_212)
);

NAND3xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_267),
.C(n_272),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_259),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_215),
.B(n_259),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_244),
.C(n_257),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_216),
.B(n_374),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_229),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_230),
.C(n_240),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g365 ( 
.A(n_218),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_SL g311 ( 
.A(n_219),
.B(n_222),
.Y(n_311)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_219),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_219),
.A2(n_329),
.B1(n_330),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_240),
.Y(n_229)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_242),
.B(n_279),
.C(n_282),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_244),
.B(n_257),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.C(n_255),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_245),
.B(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_250),
.B(n_256),
.Y(n_361)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2x2_ASAP7_75t_SL g305 ( 
.A(n_254),
.B(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_262),
.C(n_265),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_268),
.Y(n_378)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_269),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_371),
.B(n_375),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_357),
.B(n_370),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_316),
.B(n_356),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_302),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_276),
.B(n_302),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_286),
.C(n_293),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_277),
.B(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_282),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_286),
.A2(n_287),
.B1(n_293),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_292),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_288),
.B(n_292),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

AO22x1_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_297),
.B1(n_300),
.B2(n_301),
.Y(n_293)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_297),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_300),
.Y(n_309)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_301),
.B(n_349),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_308),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_304),
.B(n_305),
.C(n_308),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g368 ( 
.A(n_309),
.B(n_311),
.C(n_312),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_326),
.B(n_355),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_321),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_322),
.A2(n_323),
.B1(n_334),
.B2(n_335),
.Y(n_333)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_327),
.A2(n_336),
.B(n_354),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_333),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_328),
.B(n_333),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_330),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_348),
.B(n_353),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_346),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_346),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_345),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_345),
.B(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_358),
.B(n_369),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_369),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_362),
.B2(n_363),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_359),
.B(n_364),
.C(n_368),
.Y(n_372)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_367),
.B2(n_368),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_372),
.B(n_373),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.C(n_379),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_432),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_387),
.Y(n_383)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_384),
.B(n_387),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_422),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_407),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_400),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_409),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_417),
.Y(n_411)
);

INVx8_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx6_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx5_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_431),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_429),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_424)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_425),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_426),
.Y(n_428)
);


endmodule