module fake_jpeg_29522_n_104 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_32),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_1),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_3),
.Y(n_58)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_44),
.B(n_45),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_37),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_4),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_34),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_35),
.B1(n_36),
.B2(n_30),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_63),
.B1(n_68),
.B2(n_73),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_67),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_35),
.B1(n_5),
.B2(n_6),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_66),
.B(n_70),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_50),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_53),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_75),
.B(n_29),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_28),
.B1(n_38),
.B2(n_29),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_18),
.B1(n_19),
.B2(n_23),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_71),
.B1(n_62),
.B2(n_60),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_89),
.B1(n_88),
.B2(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_79),
.B(n_80),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_9),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_10),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_89),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_13),
.B(n_14),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_87),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_15),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_92),
.B(n_85),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_93),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_90),
.B(n_83),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_94),
.C(n_77),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_94),
.B1(n_91),
.B2(n_86),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_98),
.B(n_99),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_95),
.B(n_24),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_101),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_96),
.B1(n_81),
.B2(n_76),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_86),
.Y(n_104)
);


endmodule