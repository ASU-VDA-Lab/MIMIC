module real_jpeg_4986_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_1),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_1),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_1),
.B(n_148),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g195 ( 
.A(n_1),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_2),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_2),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_2),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_2),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_2),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_3),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_3),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_3),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_3),
.B(n_76),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_3),
.B(n_286),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_3),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_3),
.B(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_4),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_5),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_5),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_5),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_175),
.Y(n_174)
);

AND2x2_ASAP7_75t_SL g245 ( 
.A(n_5),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_5),
.B(n_329),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_5),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_6),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_6),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_6),
.B(n_196),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_6),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_6),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_6),
.B(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_6),
.B(n_109),
.Y(n_362)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_8),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_8),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_8),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_8),
.B(n_249),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_8),
.B(n_196),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_8),
.B(n_332),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_8),
.B(n_198),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_9),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_9),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_10),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_10),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_10),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_10),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_10),
.B(n_193),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_10),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_10),
.B(n_329),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_11),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_11),
.B(n_39),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_11),
.B(n_266),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_11),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_11),
.B(n_100),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_11),
.B(n_348),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_11),
.B(n_359),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_12),
.Y(n_123)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g99 ( 
.A(n_14),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_14),
.B(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_15),
.Y(n_93)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_15),
.Y(n_144)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_15),
.Y(n_190)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_15),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_16),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_16),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_16),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_16),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_16),
.B(n_105),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_16),
.B(n_340),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_16),
.B(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_17),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_17),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_204),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_203),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_160),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_22),
.B(n_160),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_94),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_67),
.C(n_80),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_24),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.C(n_48),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_25),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_31),
.C(n_36),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_41),
.C(n_45),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_30),
.A2(n_31),
.B1(n_101),
.B2(n_107),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_31),
.B(n_101),
.C(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_35),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_40),
.B(n_48),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_41),
.B(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_45),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_47),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g266 ( 
.A(n_47),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_47),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_54),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_49),
.B(n_55),
.C(n_60),
.Y(n_158)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_53),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_57),
.Y(n_180)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_57),
.Y(n_314)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_64),
.Y(n_371)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_66),
.Y(n_87)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_66),
.Y(n_296)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_66),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_67),
.B(n_80),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_74),
.C(n_79),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_74),
.B1(n_75),
.B2(n_79),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_74),
.A2(n_75),
.B1(n_91),
.B2(n_92),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_81),
.C(n_91),
.Y(n_80)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_77),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_77),
.Y(n_228)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g346 ( 
.A(n_78),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_82),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.C(n_88),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_83),
.B(n_88),
.Y(n_168)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_86),
.B(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_90),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_134),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_113),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_108),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_101),
.B2(n_107),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_106),
.Y(n_246)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_106),
.Y(n_292)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_112),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_115),
.B(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.C(n_128),
.Y(n_120)
);

FAx1_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_124),
.CI(n_128),
.CON(n_159),
.SN(n_159)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_127),
.Y(n_249)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_132),
.Y(n_368)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_133),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_155),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_154),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_151),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_159),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g448 ( 
.A(n_159),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_163),
.C(n_165),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_161),
.B(n_163),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_208),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_184),
.C(n_186),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_169),
.C(n_181),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_167),
.B(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_169),
.A2(n_170),
.B1(n_181),
.B2(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_174),
.C(n_178),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_171),
.B(n_178),
.Y(n_422)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_174),
.B(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_181),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_186),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_197),
.C(n_200),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_238),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.C(n_195),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_188),
.B(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_192),
.B(n_195),
.Y(n_221)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_197),
.B(n_200),
.Y(n_238)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_254),
.B(n_446),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_207),
.B(n_209),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_213),
.C(n_216),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_211),
.B(n_214),
.Y(n_442)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_216),
.B(n_442),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_236),
.C(n_239),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_218),
.B(n_435),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.C(n_229),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_219),
.A2(n_220),
.B1(n_413),
.B2(n_414),
.Y(n_412)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_222),
.A2(n_223),
.B(n_225),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_222),
.B(n_229),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_224),
.Y(n_269)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.C(n_234),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_390)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_234),
.B(n_390),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_235),
.B(n_326),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_236),
.A2(n_237),
.B1(n_239),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_239),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_250),
.C(n_253),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_241),
.B(n_424),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_247),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_242),
.B(n_402),
.Y(n_401)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_403),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g403 ( 
.A(n_245),
.Y(n_403)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_250),
.B(n_253),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_252),
.Y(n_326)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_440),
.B(n_445),
.Y(n_254)
);

OAI21x1_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_427),
.B(n_439),
.Y(n_255)
);

AOI21x1_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_409),
.B(n_426),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_383),
.B(n_408),
.Y(n_257)
);

AOI21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_353),
.B(n_382),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_318),
.B(n_352),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_298),
.B(n_317),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_275),
.B(n_297),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_272),
.B(n_274),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_270),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_264),
.B(n_270),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_267),
.Y(n_276)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_277),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_288),
.B2(n_289),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_278),
.B(n_291),
.C(n_293),
.Y(n_316)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_285),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_285),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_293),
.B2(n_294),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_316),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_316),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_308),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_307),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_307),
.C(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_306),
.Y(n_323)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_308),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_336),
.C(n_337),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_315),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_321),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_334),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_322),
.B(n_335),
.C(n_338),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_325),
.C(n_327),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_327),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_330),
.B1(n_331),
.B2(n_333),
.Y(n_327)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_333),
.Y(n_363)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_SL g377 ( 
.A(n_332),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_343),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_339),
.B(n_347),
.C(n_350),
.Y(n_380)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_347),
.B1(n_350),
.B2(n_351),
.Y(n_343)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_344),
.Y(n_350)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_347),
.Y(n_351)
);

INVx6_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_354),
.B(n_381),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_381),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g354 ( 
.A(n_355),
.B(n_365),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_364),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_356),
.B(n_364),
.C(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_363),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_358),
.Y(n_397)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_363),
.B(n_397),
.C(n_398),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_372),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_374),
.C(n_379),
.Y(n_386)
);

BUFx24_ASAP7_75t_SL g449 ( 
.A(n_366),
.Y(n_449)
);

FAx1_ASAP7_75t_SL g366 ( 
.A(n_367),
.B(n_369),
.CI(n_370),
.CON(n_366),
.SN(n_366)
);

MAJx2_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_369),
.C(n_370),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_373),
.A2(n_374),
.B1(n_379),
.B2(n_380),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_378),
.Y(n_393)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_406),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_384),
.B(n_406),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_395),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_387),
.C(n_395),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_391),
.B2(n_392),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_418),
.C(n_419),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_393),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_399),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_396),
.B(n_400),
.C(n_405),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B1(n_404),
.B2(n_405),
.Y(n_399)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_400),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_401),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_425),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_410),
.B(n_425),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_416),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_412),
.B(n_415),
.C(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_413),
.Y(n_414)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_420),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_421),
.C(n_423),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_437),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_428),
.B(n_437),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_434),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_431),
.B(n_434),
.C(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_441),
.B(n_443),
.Y(n_445)
);


endmodule