module fake_ariane_816_n_27 (n_8, n_3, n_2, n_7, n_5, n_1, n_0, n_6, n_9, n_4, n_27);

input n_8;
input n_3;
input n_2;
input n_7;
input n_5;
input n_1;
input n_0;
input n_6;
input n_9;
input n_4;

output n_27;

wire n_24;
wire n_22;
wire n_13;
wire n_20;
wire n_17;
wire n_18;
wire n_11;
wire n_26;
wire n_14;
wire n_19;
wire n_16;
wire n_12;
wire n_15;
wire n_21;
wire n_23;
wire n_10;
wire n_25;

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_5),
.B(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_1),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_2),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx4_ASAP7_75t_SL g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

AO31x2_ASAP7_75t_L g18 ( 
.A1(n_13),
.A2(n_0),
.A3(n_2),
.B(n_3),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_10),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_20),
.A2(n_12),
.B1(n_17),
.B2(n_14),
.Y(n_22)
);

AOI221xp5_ASAP7_75t_L g23 ( 
.A1(n_21),
.A2(n_14),
.B1(n_18),
.B2(n_6),
.C(n_3),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g24 ( 
.A1(n_22),
.A2(n_18),
.B(n_6),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_18),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g26 ( 
.A1(n_25),
.A2(n_23),
.B1(n_16),
.B2(n_20),
.Y(n_26)
);

AO21x1_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_4),
.B(n_9),
.Y(n_27)
);


endmodule