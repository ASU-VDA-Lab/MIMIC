module fake_jpeg_18389_n_253 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_253);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_253;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_10),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_17),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_26),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_29),
.B1(n_19),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_47),
.B1(n_37),
.B2(n_36),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_29),
.B1(n_19),
.B2(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_36),
.A2(n_29),
.B1(n_30),
.B2(n_24),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_23),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_18),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_23),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_58),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_36),
.A2(n_29),
.B1(n_19),
.B2(n_24),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_23),
.B1(n_27),
.B2(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_72),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_68),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_100)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_47),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_57),
.A2(n_37),
.B1(n_36),
.B2(n_33),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_77),
.B(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_57),
.A2(n_37),
.B1(n_20),
.B2(n_33),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_87),
.C(n_34),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_37),
.B1(n_31),
.B2(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_31),
.B1(n_25),
.B2(n_32),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_85),
.Y(n_98)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_86),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_59),
.A2(n_18),
.B1(n_21),
.B2(n_27),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_88),
.B(n_102),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_111),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_101),
.B1(n_83),
.B2(n_62),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_52),
.B1(n_47),
.B2(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_71),
.B(n_56),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_58),
.B(n_34),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_67),
.B(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_106),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_65),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_51),
.B1(n_76),
.B2(n_69),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_112),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_34),
.B(n_23),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_70),
.B(n_41),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_63),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_86),
.B1(n_74),
.B2(n_68),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_98),
.B1(n_60),
.B2(n_85),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_117),
.A2(n_101),
.B1(n_112),
.B2(n_98),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_124),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_63),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_125),
.Y(n_140)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_109),
.B(n_18),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_39),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_129),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_39),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_18),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_95),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_133),
.B(n_105),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_90),
.C(n_102),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_132),
.C(n_96),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_34),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_39),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_90),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_134),
.B(n_64),
.Y(n_162)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_94),
.B(n_39),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_92),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_139),
.B(n_154),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_99),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_159),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_128),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_142),
.A2(n_145),
.B(n_149),
.Y(n_185)
);

MAJx2_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_88),
.C(n_107),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_148),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_115),
.B(n_100),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_149),
.A2(n_133),
.B(n_21),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_160),
.B1(n_163),
.B2(n_152),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_156),
.B1(n_136),
.B2(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_79),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_108),
.B1(n_79),
.B2(n_60),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_34),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_117),
.A2(n_108),
.B1(n_60),
.B2(n_41),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_161),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_162),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_122),
.A2(n_41),
.B1(n_32),
.B2(n_25),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_41),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_120),
.C(n_125),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_166),
.C(n_172),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_120),
.C(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_155),
.B(n_114),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_175),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_130),
.C(n_126),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_144),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_164),
.Y(n_176)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_176),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_184),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_150),
.B1(n_160),
.B2(n_176),
.Y(n_201)
);

OAI322xp33_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_127),
.A3(n_130),
.B1(n_122),
.B2(n_133),
.C1(n_28),
.C2(n_22),
.Y(n_179)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_179),
.B(n_186),
.C(n_22),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_180),
.A2(n_185),
.B1(n_156),
.B2(n_153),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_182),
.A2(n_177),
.B(n_152),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_28),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_163),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_147),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_145),
.B(n_14),
.C(n_13),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_190),
.Y(n_208)
);

OAI21x1_ASAP7_75t_L g216 ( 
.A1(n_189),
.A2(n_32),
.B(n_25),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_140),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_203),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_197),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_170),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_173),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_142),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_198),
.B(n_14),
.Y(n_215)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_168),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_169),
.C(n_165),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_172),
.C(n_183),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_204),
.B1(n_191),
.B2(n_196),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_202),
.Y(n_212)
);

OAI21x1_ASAP7_75t_L g203 ( 
.A1(n_185),
.A2(n_151),
.B(n_22),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_169),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_209),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_174),
.C(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_213),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_214),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_215),
.B(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_216),
.B(n_3),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_217),
.A2(n_201),
.B1(n_204),
.B2(n_202),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_219),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_222),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_212),
.A2(n_189),
.B1(n_193),
.B2(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_227),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_228),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_208),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_206),
.B(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_236),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_190),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_234),
.B(n_3),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_209),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_231),
.A2(n_223),
.B1(n_225),
.B2(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_239),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_227),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_242),
.B(n_5),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_4),
.C(n_5),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_241),
.A2(n_233),
.B(n_7),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_4),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_246),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_238),
.A2(n_229),
.B(n_7),
.Y(n_245)
);

AOI321xp33_ASAP7_75t_SL g247 ( 
.A1(n_245),
.A2(n_241),
.A3(n_240),
.B1(n_9),
.B2(n_10),
.C(n_7),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_247),
.A2(n_248),
.B(n_8),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_243),
.A2(n_229),
.B(n_9),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_251),
.B(n_8),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_249),
.A2(n_8),
.B(n_11),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_11),
.Y(n_253)
);


endmodule