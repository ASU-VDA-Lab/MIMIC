module fake_jpeg_28049_n_55 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_55);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_51;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_17;
wire n_25;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_32;

BUFx4f_ASAP7_75t_SL g16 ( 
.A(n_14),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_2),
.B(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_30),
.C(n_31),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_37),
.B(n_39),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_47),
.B1(n_41),
.B2(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_42),
.B1(n_38),
.B2(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_16),
.C(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_20),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_53),
.A2(n_50),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_25),
.Y(n_55)
);


endmodule