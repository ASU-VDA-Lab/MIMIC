module fake_jpeg_21730_n_238 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_15),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_35),
.B(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

CKINVDCx9p33_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_49),
.Y(n_82)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_40),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_50),
.A2(n_57),
.B1(n_63),
.B2(n_71),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_34),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_51),
.A2(n_0),
.B(n_1),
.Y(n_98)
);

BUFx4f_ASAP7_75t_SL g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_32),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_19),
.B1(n_28),
.B2(n_17),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_59),
.B(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_31),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_40),
.A2(n_19),
.B1(n_28),
.B2(n_17),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_24),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_68),
.Y(n_84)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_21),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_42),
.A2(n_17),
.B1(n_23),
.B2(n_21),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_70),
.A2(n_77),
.B1(n_44),
.B2(n_18),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_26),
.B1(n_22),
.B2(n_20),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_37),
.B(n_26),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_73),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_37),
.A2(n_22),
.B(n_18),
.C(n_29),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_38),
.B(n_43),
.C(n_44),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_36),
.B(n_29),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_75),
.Y(n_104)
);

OA22x2_ASAP7_75t_L g76 ( 
.A1(n_37),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_76)
);

OA22x2_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_42),
.A2(n_27),
.B1(n_18),
.B2(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_38),
.C(n_44),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_95),
.C(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_79),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_87),
.Y(n_134)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_100),
.B1(n_78),
.B2(n_54),
.Y(n_120)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_93),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_SL g136 ( 
.A(n_94),
.B(n_103),
.C(n_52),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_27),
.C(n_16),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_16),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_108),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_60),
.B1(n_47),
.B2(n_49),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_9),
.B1(n_3),
.B2(n_4),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_0),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_61),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_74),
.A2(n_0),
.B(n_4),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_105),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_53),
.B(n_14),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_125),
.Y(n_139)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_53),
.A3(n_76),
.B1(n_70),
.B2(n_77),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_123),
.Y(n_147)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_116),
.B(n_119),
.Y(n_148)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_106),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_129),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_121),
.B1(n_127),
.B2(n_96),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_67),
.B1(n_58),
.B2(n_47),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_102),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_128),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_46),
.Y(n_125)
);

NAND2xp33_ASAP7_75t_R g126 ( 
.A(n_99),
.B(n_52),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_94),
.B(n_109),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_61),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_135),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_46),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_60),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_66),
.C(n_46),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_136),
.A2(n_103),
.B(n_96),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_98),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_105),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_145),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_160),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_86),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_138),
.Y(n_144)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_144),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_SL g151 ( 
.A(n_137),
.B(n_92),
.C(n_99),
.Y(n_151)
);

NOR4xp25_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_155),
.C(n_143),
.D(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_153),
.A2(n_135),
.B1(n_122),
.B2(n_124),
.Y(n_175)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_157),
.B(n_148),
.Y(n_177)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_158),
.B(n_162),
.Y(n_170)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_80),
.B(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_108),
.Y(n_161)
);

AO22x1_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_110),
.B1(n_118),
.B2(n_114),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_80),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_116),
.B(n_88),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_133),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_149),
.A2(n_119),
.B1(n_113),
.B2(n_124),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_168),
.B1(n_175),
.B2(n_147),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_119),
.B1(n_124),
.B2(n_127),
.Y(n_168)
);

XNOR2x2_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_122),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_169),
.A2(n_177),
.B(n_148),
.Y(n_190)
);

XNOR2x2_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_110),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_178),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_115),
.Y(n_179)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_182),
.A2(n_194),
.B1(n_178),
.B2(n_177),
.Y(n_201)
);

OAI321xp33_ASAP7_75t_L g183 ( 
.A1(n_171),
.A2(n_147),
.A3(n_150),
.B1(n_161),
.B2(n_151),
.C(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_183),
.B(n_184),
.Y(n_199)
);

OAI321xp33_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_169),
.A3(n_168),
.B1(n_150),
.B2(n_166),
.C(n_175),
.Y(n_184)
);

OA21x2_ASAP7_75t_SL g204 ( 
.A1(n_186),
.A2(n_189),
.B(n_191),
.Y(n_204)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_181),
.B(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_169),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_190),
.A2(n_192),
.B(n_193),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_153),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_180),
.B(n_159),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_163),
.C(n_144),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_180),
.B(n_158),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_196),
.A2(n_156),
.B(n_140),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_195),
.A2(n_172),
.B1(n_164),
.B2(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_197),
.A2(n_202),
.B1(n_205),
.B2(n_207),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_177),
.B(n_172),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_129),
.B(n_66),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_201),
.B(n_194),
.C(n_189),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_195),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_146),
.B1(n_154),
.B2(n_152),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_192),
.B(n_185),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_141),
.B1(n_162),
.B2(n_93),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_212),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_198),
.A2(n_186),
.B(n_187),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_211),
.A2(n_215),
.B(n_217),
.Y(n_220)
);

NOR3xp33_ASAP7_75t_SL g212 ( 
.A(n_199),
.B(n_141),
.C(n_12),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_208),
.A2(n_81),
.B1(n_89),
.B2(n_83),
.Y(n_214)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_214),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_208),
.A2(n_87),
.B(n_114),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_202),
.B(n_203),
.Y(n_222)
);

OA21x2_ASAP7_75t_SL g217 ( 
.A1(n_204),
.A2(n_10),
.B(n_13),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_201),
.C(n_204),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_223),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_222),
.B(n_211),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_216),
.B(n_203),
.C(n_207),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_225),
.A2(n_220),
.B(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_213),
.B1(n_200),
.B2(n_212),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_228),
.B(n_229),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_218),
.B(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_227),
.A2(n_221),
.B(n_223),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_232),
.A2(n_226),
.B(n_14),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_231),
.B(n_226),
.C(n_14),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_235),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_13),
.C(n_60),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_236),
.Y(n_238)
);


endmodule