module fake_jpeg_653_n_530 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_530);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_530;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_352;
wire n_350;
wire n_150;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_133;
wire n_132;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

NAND2x1_ASAP7_75t_SL g46 ( 
.A(n_27),
.B(n_12),
.Y(n_46)
);

OR2x4_ASAP7_75t_L g141 ( 
.A(n_46),
.B(n_33),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_47),
.B(n_55),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_13),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_60),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_64),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_32),
.B(n_11),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_65),
.B(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_66),
.Y(n_119)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx12f_ASAP7_75t_SL g70 ( 
.A(n_37),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_80),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_77),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_11),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_78),
.B(n_92),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVxp67_ASAP7_75t_SL g80 ( 
.A(n_33),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx11_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_88),
.Y(n_150)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_35),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_22),
.B(n_11),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_15),
.Y(n_95)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_57),
.B(n_22),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_98),
.B(n_100),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_101),
.B(n_128),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_31),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_103),
.B(n_108),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_31),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_31),
.B1(n_30),
.B2(n_40),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_41),
.B1(n_16),
.B2(n_34),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_80),
.A2(n_17),
.B1(n_30),
.B2(n_40),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_118),
.A2(n_122),
.B1(n_138),
.B2(n_140),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_46),
.A2(n_17),
.B1(n_30),
.B2(n_40),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_38),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_124),
.B(n_137),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_69),
.A2(n_39),
.B(n_15),
.C(n_28),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_39),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_60),
.A2(n_17),
.B1(n_39),
.B2(n_28),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_17),
.B1(n_28),
.B2(n_38),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_141),
.B(n_24),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_62),
.A2(n_74),
.B1(n_63),
.B2(n_87),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_148),
.A2(n_29),
.B1(n_41),
.B2(n_34),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_91),
.B(n_36),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_149),
.B(n_29),
.Y(n_201)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_156),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_160),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

BUFx2_ASAP7_75t_SL g218 ( 
.A(n_161),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_99),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_162),
.B(n_172),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_102),
.A2(n_36),
.B(n_38),
.Y(n_163)
);

NAND2x1_ASAP7_75t_L g231 ( 
.A(n_163),
.B(n_186),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_164),
.A2(n_165),
.B1(n_187),
.B2(n_26),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_L g165 ( 
.A1(n_122),
.A2(n_68),
.B1(n_86),
.B2(n_79),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_166),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_106),
.B(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_167),
.B(n_175),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_109),
.A2(n_59),
.B1(n_61),
.B2(n_48),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_168),
.A2(n_183),
.B1(n_140),
.B2(n_157),
.Y(n_232)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_102),
.Y(n_170)
);

INVx5_ASAP7_75t_SL g225 ( 
.A(n_170),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_156),
.Y(n_171)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_97),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_110),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_178),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_128),
.B(n_90),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_141),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_200),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_129),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_180),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_117),
.A2(n_36),
.B1(n_41),
.B2(n_24),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_107),
.Y(n_182)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_182),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_138),
.A2(n_56),
.B1(n_53),
.B2(n_75),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_130),
.C(n_112),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_191),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_117),
.B(n_16),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_105),
.A2(n_71),
.B1(n_16),
.B2(n_20),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_189),
.B(n_195),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_190),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_107),
.B(n_34),
.Y(n_191)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_139),
.Y(n_193)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_97),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_196),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_135),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_197),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_204),
.B1(n_26),
.B2(n_24),
.Y(n_210)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_151),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_199),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_113),
.B(n_29),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_202),
.Y(n_228)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_175),
.A2(n_118),
.B1(n_157),
.B2(n_155),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_209),
.A2(n_232),
.B1(n_233),
.B2(n_182),
.Y(n_267)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

OR2x2_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_123),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_211),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_164),
.A2(n_111),
.B1(n_155),
.B2(n_144),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_216),
.A2(n_168),
.B1(n_158),
.B2(n_200),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_187),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_167),
.B(n_152),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_178),
.C(n_207),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_120),
.B1(n_144),
.B2(n_142),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_206),
.A2(n_178),
.B(n_179),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_241),
.A2(n_253),
.B(n_163),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g299 ( 
.A(n_243),
.B(n_263),
.C(n_266),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_244),
.A2(n_219),
.B1(n_236),
.B2(n_234),
.Y(n_280)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_214),
.Y(n_245)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_246),
.B(n_248),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_213),
.B(n_188),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_247),
.B(n_269),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_184),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_205),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_262),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_159),
.B1(n_183),
.B2(n_165),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_250),
.A2(n_261),
.B1(n_267),
.B2(n_225),
.Y(n_283)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_229),
.Y(n_251)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_251),
.Y(n_271)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_231),
.B(n_221),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_209),
.A2(n_170),
.B(n_172),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_254),
.A2(n_221),
.B(n_231),
.Y(n_277)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_214),
.Y(n_255)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_255),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_228),
.B(n_203),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_258),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g257 ( 
.A(n_208),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_257),
.A2(n_222),
.B1(n_174),
.B2(n_199),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_228),
.B(n_186),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_186),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_268),
.Y(n_285)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_214),
.Y(n_260)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_207),
.B(n_185),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_226),
.B(n_173),
.C(n_177),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_191),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_162),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_234),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_272),
.B(n_295),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_273),
.Y(n_324)
);

AO22x1_ASAP7_75t_SL g275 ( 
.A1(n_261),
.A2(n_227),
.B1(n_233),
.B2(n_221),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_281),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_277),
.A2(n_265),
.B(n_253),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_279),
.B(n_290),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_280),
.A2(n_283),
.B1(n_292),
.B2(n_298),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_269),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_264),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_286),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_264),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_252),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_287),
.B(n_235),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_248),
.B(n_211),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_267),
.A2(n_261),
.B1(n_254),
.B2(n_246),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_291),
.A2(n_241),
.B1(n_258),
.B2(n_244),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_250),
.A2(n_237),
.B1(n_222),
.B2(n_215),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_219),
.Y(n_293)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

OA21x2_ASAP7_75t_SL g295 ( 
.A1(n_247),
.A2(n_225),
.B(n_236),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_261),
.A2(n_237),
.B1(n_215),
.B2(n_225),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_263),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_304),
.C(n_310),
.Y(n_334)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_263),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_303),
.B(n_313),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_243),
.C(n_259),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_305),
.A2(n_315),
.B(n_326),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_270),
.B(n_262),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_307),
.B(n_314),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_309),
.A2(n_311),
.B1(n_318),
.B2(n_320),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_268),
.C(n_265),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_242),
.B1(n_251),
.B2(n_266),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_272),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_312),
.B(n_301),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_189),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_270),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_277),
.A2(n_242),
.B(n_212),
.Y(n_315)
);

NAND4xp25_ASAP7_75t_SL g317 ( 
.A(n_285),
.B(n_33),
.C(n_151),
.D(n_192),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_317),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_245),
.B1(n_255),
.B2(n_260),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_195),
.C(n_166),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_319),
.B(n_321),
.C(n_190),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_255),
.B1(n_245),
.B2(n_240),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_276),
.B(n_235),
.C(n_196),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_280),
.A2(n_274),
.B1(n_276),
.B2(n_293),
.Y(n_322)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_322),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_279),
.B(n_191),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_323),
.B(n_289),
.Y(n_349)
);

A2O1A1O1Ixp25_ASAP7_75t_L g326 ( 
.A1(n_279),
.A2(n_290),
.B(n_281),
.C(n_295),
.D(n_274),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_292),
.A2(n_240),
.B1(n_238),
.B2(n_212),
.Y(n_327)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_275),
.A2(n_287),
.B1(n_284),
.B2(n_271),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_328),
.A2(n_298),
.B1(n_275),
.B2(n_289),
.Y(n_338)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_329),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_275),
.A2(n_238),
.B1(n_224),
.B2(n_190),
.Y(n_330)
);

OAI22x1_ASAP7_75t_L g357 ( 
.A1(n_330),
.A2(n_297),
.B1(n_294),
.B2(n_160),
.Y(n_357)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_271),
.Y(n_332)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_332),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_338),
.A2(n_357),
.B1(n_360),
.B2(n_127),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_326),
.A2(n_273),
.B(n_275),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_339),
.A2(n_330),
.B(n_318),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_340),
.B(n_352),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_306),
.A2(n_282),
.B1(n_286),
.B2(n_288),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_341),
.A2(n_358),
.B1(n_332),
.B2(n_325),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_315),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_363),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_346),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_331),
.B(n_288),
.Y(n_348)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_348),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g388 ( 
.A(n_349),
.B(n_154),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_296),
.Y(n_350)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_350),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_223),
.C(n_180),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_359),
.C(n_323),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_303),
.B(n_180),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_355),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_296),
.Y(n_354)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_304),
.B(n_176),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_316),
.A2(n_294),
.B1(n_297),
.B2(n_257),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_310),
.B(n_223),
.C(n_123),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_328),
.A2(n_208),
.B1(n_160),
.B2(n_171),
.Y(n_360)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_302),
.Y(n_362)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_362),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_321),
.B(n_220),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_305),
.A2(n_324),
.B(n_311),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_364),
.A2(n_324),
.B(n_309),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_365),
.B(n_370),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_367),
.A2(n_368),
.B(n_378),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_319),
.C(n_308),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_369),
.B(n_375),
.C(n_379),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g413 ( 
.A(n_372),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_334),
.B(n_308),
.C(n_317),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_337),
.B(n_220),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_376),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_193),
.Y(n_377)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_377),
.Y(n_402)
);

FAx1_ASAP7_75t_L g378 ( 
.A(n_353),
.B(n_218),
.CI(n_143),
.CON(n_378),
.SN(n_378)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_171),
.C(n_150),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_204),
.Y(n_380)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_388),
.C(n_335),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_361),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_383),
.A2(n_394),
.B1(n_335),
.B2(n_363),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_344),
.B(n_202),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_384),
.B(n_350),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_143),
.C(n_127),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_390),
.C(n_340),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_347),
.B(n_111),
.C(n_142),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_336),
.B(n_26),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_391),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_348),
.B(n_354),
.Y(n_393)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_356),
.A2(n_136),
.B1(n_120),
.B2(n_134),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_374),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_395),
.B(n_407),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_396),
.A2(n_404),
.B1(n_409),
.B2(n_383),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_374),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_398),
.B(n_10),
.Y(n_440)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_399),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_367),
.A2(n_364),
.B1(n_339),
.B2(n_345),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_401),
.A2(n_386),
.B1(n_134),
.B2(n_132),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_368),
.A2(n_343),
.B1(n_338),
.B2(n_341),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_370),
.B(n_353),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_410),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_393),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_349),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_387),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_382),
.A2(n_357),
.B1(n_358),
.B2(n_360),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_365),
.B(n_371),
.C(n_375),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_412),
.B(n_415),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_362),
.Y(n_414)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_414),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_371),
.B(n_359),
.C(n_333),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_416),
.B(n_387),
.Y(n_436)
);

OAI211xp5_ASAP7_75t_SL g418 ( 
.A1(n_382),
.A2(n_342),
.B(n_333),
.C(n_136),
.Y(n_418)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_418),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_378),
.A2(n_342),
.B(n_20),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_419),
.A2(n_392),
.B(n_377),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_422),
.B(n_440),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_420),
.A2(n_378),
.B(n_413),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g457 ( 
.A1(n_425),
.A2(n_445),
.B(n_20),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_380),
.C(n_379),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_426),
.B(n_427),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_389),
.C(n_390),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_385),
.C(n_388),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_114),
.C(n_104),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_429),
.A2(n_404),
.B1(n_409),
.B2(n_398),
.Y(n_449)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_430),
.Y(n_447)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g463 ( 
.A(n_435),
.B(n_442),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_121),
.Y(n_458)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_414),
.Y(n_437)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_438),
.A2(n_153),
.B1(n_42),
.B2(n_10),
.Y(n_465)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_397),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_441),
.B(n_443),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_413),
.B(n_132),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_402),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_406),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_416),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_420),
.A2(n_419),
.B(n_401),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_411),
.B(n_417),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_125),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_449),
.A2(n_450),
.B1(n_452),
.B2(n_454),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_432),
.A2(n_405),
.B1(n_403),
.B2(n_410),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_451),
.B(n_456),
.Y(n_467)
);

INVx11_ASAP7_75t_L g452 ( 
.A(n_441),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_423),
.A2(n_403),
.B1(n_415),
.B2(n_408),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_121),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_457),
.B(n_440),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_458),
.B(n_424),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_423),
.A2(n_114),
.B1(n_104),
.B2(n_125),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_438),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_SL g470 ( 
.A(n_461),
.B(n_462),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_10),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_10),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_465),
.A2(n_431),
.B1(n_455),
.B2(n_430),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_460),
.B(n_434),
.Y(n_468)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_468),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_469),
.B(n_471),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_472),
.B(n_475),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_454),
.B(n_428),
.C(n_434),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_474),
.B(n_480),
.Y(n_484)
);

NOR2xp67_ASAP7_75t_SL g476 ( 
.A(n_450),
.B(n_427),
.Y(n_476)
);

AOI21x1_ASAP7_75t_L g493 ( 
.A1(n_476),
.A2(n_424),
.B(n_452),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_453),
.A2(n_437),
.B1(n_444),
.B2(n_443),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_477),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_0),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_449),
.B(n_426),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_479),
.B(n_459),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_445),
.C(n_425),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_436),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_481),
.B(n_457),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_447),
.B(n_455),
.Y(n_483)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_483),
.A2(n_448),
.B(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_485),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_479),
.B(n_466),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_486),
.B(n_0),
.Y(n_503)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_488),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_490),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_458),
.C(n_447),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_497),
.B(n_1),
.Y(n_507)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_495),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_467),
.B(n_465),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_496),
.B(n_498),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_483),
.A2(n_153),
.B(n_42),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_484),
.B(n_470),
.Y(n_499)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_487),
.A2(n_472),
.B(n_475),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_500),
.A2(n_494),
.B(n_491),
.Y(n_511)
);

OAI21x1_ASAP7_75t_SL g518 ( 
.A1(n_503),
.A2(n_506),
.B(n_507),
.Y(n_518)
);

A2O1A1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_492),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_490),
.B(n_494),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_508),
.A2(n_491),
.B(n_3),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_495),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_4),
.B(n_5),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_511),
.A2(n_512),
.B(n_513),
.Y(n_523)
);

A2O1A1O1Ixp25_ASAP7_75t_L g513 ( 
.A1(n_501),
.A2(n_1),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_3),
.C(n_4),
.Y(n_515)
);

MAJx2_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_516),
.C(n_517),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_504),
.A2(n_505),
.B(n_509),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_514),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_521),
.C(n_522),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_518),
.B(n_506),
.C(n_6),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_506),
.C(n_6),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_519),
.B(n_5),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_524),
.A2(n_525),
.B(n_7),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_5),
.C(n_6),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_6),
.B(n_7),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_527),
.A2(n_528),
.B1(n_6),
.B2(n_9),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_529),
.B(n_9),
.Y(n_530)
);


endmodule