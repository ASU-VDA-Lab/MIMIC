module fake_jpeg_11624_n_639 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_639);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_639;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_519;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_1),
.B(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_11),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_18),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

INVxp33_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_4),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_0),
.Y(n_53)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_60),
.Y(n_150)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_61),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_62),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_65),
.B(n_73),
.Y(n_182)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_66),
.B(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_24),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_69),
.B(n_119),
.Y(n_133)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_71),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_72),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_43),
.B(n_11),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_75),
.Y(n_141)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_76),
.B(n_89),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_77),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_78),
.Y(n_191)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_24),
.Y(n_79)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_79),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_80),
.Y(n_179)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_81),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_82),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_83),
.Y(n_185)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_85),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_87),
.Y(n_202)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_59),
.Y(n_88)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_25),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_90),
.B(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_91),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_39),
.B(n_11),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_92),
.B(n_124),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_25),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_94),
.B(n_99),
.Y(n_156)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_30),
.A2(n_9),
.B1(n_17),
.B2(n_3),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_97),
.A2(n_46),
.B1(n_44),
.B2(n_27),
.Y(n_176)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_100),
.Y(n_187)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_33),
.Y(n_102)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_25),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_106),
.Y(n_162)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_39),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_107),
.B(n_116),
.Y(n_166)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_33),
.Y(n_108)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_109),
.Y(n_213)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_41),
.Y(n_110)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_23),
.Y(n_111)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_23),
.Y(n_112)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_34),
.Y(n_113)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_26),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_52),
.B(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_122),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_52),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_118),
.B(n_123),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_120),
.B(n_121),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_34),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_52),
.B(n_9),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_22),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_32),
.Y(n_125)
);

NOR2x1_ASAP7_75t_R g196 ( 
.A(n_125),
.B(n_127),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_22),
.B(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_126),
.B(n_128),
.Y(n_180)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_35),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_32),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_130),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_35),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_58),
.B1(n_35),
.B2(n_38),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_131),
.A2(n_154),
.B1(n_167),
.B2(n_176),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_105),
.A2(n_28),
.B1(n_57),
.B2(n_31),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_134),
.A2(n_157),
.B1(n_165),
.B2(n_175),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_69),
.A2(n_53),
.B1(n_54),
.B2(n_58),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_139),
.A2(n_153),
.B1(n_173),
.B2(n_181),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_28),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_145),
.B(n_198),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_70),
.A2(n_53),
.B1(n_58),
.B2(n_50),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_122),
.A2(n_38),
.B1(n_45),
.B2(n_50),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_61),
.A2(n_38),
.B1(n_45),
.B2(n_50),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_85),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_158),
.B(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_129),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_161),
.B(n_163),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_60),
.B(n_27),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_100),
.A2(n_57),
.B1(n_31),
.B2(n_37),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_84),
.A2(n_45),
.B1(n_55),
.B2(n_40),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_70),
.A2(n_55),
.B1(n_46),
.B2(n_44),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_113),
.A2(n_130),
.B1(n_128),
.B2(n_124),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_63),
.A2(n_40),
.B1(n_37),
.B2(n_3),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_104),
.A2(n_13),
.B1(n_17),
.B2(n_3),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_183),
.A2(n_203),
.B1(n_219),
.B2(n_222),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_SL g186 ( 
.A(n_64),
.Y(n_186)
);

INVx13_ASAP7_75t_L g261 ( 
.A(n_186),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_114),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_190),
.B(n_194),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_110),
.A2(n_14),
.B1(n_17),
.B2(n_4),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_200),
.C(n_133),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_111),
.B(n_112),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_95),
.A2(n_8),
.B1(n_16),
.B2(n_4),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_195),
.A2(n_211),
.B1(n_176),
.B2(n_154),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_96),
.B(n_8),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_98),
.A2(n_8),
.B1(n_16),
.B2(n_4),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_199),
.A2(n_206),
.B1(n_216),
.B2(n_197),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_101),
.B(n_6),
.C(n_15),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_81),
.A2(n_6),
.B1(n_16),
.B2(n_18),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_79),
.A2(n_6),
.B(n_18),
.C(n_0),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g270 ( 
.A1(n_204),
.A2(n_192),
.B(n_205),
.C(n_218),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g206 ( 
.A1(n_121),
.A2(n_86),
.B1(n_62),
.B2(n_83),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_120),
.B(n_2),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_208),
.B(n_209),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_102),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_108),
.B(n_2),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_210),
.B(n_217),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_80),
.A2(n_2),
.B1(n_91),
.B2(n_109),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_78),
.B(n_2),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_215),
.B(n_148),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_88),
.A2(n_68),
.B1(n_87),
.B2(n_127),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_82),
.B(n_119),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_71),
.A2(n_118),
.B1(n_69),
.B2(n_53),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_72),
.A2(n_118),
.B1(n_69),
.B2(n_53),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_150),
.Y(n_223)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_150),
.Y(n_228)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_230),
.Y(n_329)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_231),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_133),
.B(n_77),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_232),
.B(n_241),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_235),
.B(n_240),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_236),
.A2(n_239),
.B1(n_287),
.B2(n_290),
.Y(n_301)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_169),
.Y(n_237)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_237),
.Y(n_308)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_174),
.Y(n_238)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_206),
.B1(n_207),
.B2(n_201),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_148),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_133),
.B(n_161),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_163),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_246),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_138),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_152),
.Y(n_247)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_247),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_193),
.A2(n_196),
.B1(n_152),
.B2(n_220),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_248),
.Y(n_316)
);

AOI21xp33_ASAP7_75t_L g249 ( 
.A1(n_145),
.A2(n_135),
.B(n_182),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_249),
.B(n_252),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_250),
.B(n_288),
.Y(n_327)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_174),
.Y(n_251)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_251),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_171),
.B(n_135),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_168),
.C(n_178),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_269),
.C(n_272),
.Y(n_334)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_254),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_162),
.B(n_166),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_255),
.B(n_263),
.Y(n_312)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_168),
.B(n_178),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_281),
.Y(n_324)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_160),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_257),
.Y(n_328)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_179),
.Y(n_258)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_258),
.Y(n_333)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_191),
.Y(n_259)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_259),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_160),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_180),
.B(n_200),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_262),
.B(n_270),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_156),
.B(n_141),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_193),
.A2(n_196),
.B1(n_220),
.B2(n_158),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_264),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_198),
.B(n_205),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_265),
.B(n_266),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_144),
.B(n_147),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_179),
.Y(n_267)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_268),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_132),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_151),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_132),
.B(n_142),
.Y(n_272)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_273),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_157),
.A2(n_199),
.B1(n_216),
.B2(n_204),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_274),
.A2(n_285),
.B1(n_296),
.B2(n_234),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_151),
.A2(n_214),
.B1(n_140),
.B2(n_169),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_191),
.Y(n_276)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_276),
.Y(n_356)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_149),
.Y(n_277)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_277),
.Y(n_358)
);

OR2x2_ASAP7_75t_SL g278 ( 
.A(n_190),
.B(n_137),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g303 ( 
.A(n_278),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_218),
.A2(n_214),
.B1(n_201),
.B2(n_187),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_279),
.A2(n_232),
.B(n_281),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_137),
.B(n_142),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_280),
.B(n_272),
.C(n_282),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_177),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g282 ( 
.A(n_149),
.B(n_164),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_282),
.B(n_292),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_189),
.B(n_209),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_283),
.B(n_284),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_140),
.B(n_170),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_187),
.A2(n_159),
.B1(n_172),
.B2(n_143),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_155),
.B(n_164),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_289),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_136),
.A2(n_202),
.B1(n_177),
.B2(n_170),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_185),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_155),
.B(n_159),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_136),
.A2(n_202),
.B1(n_177),
.B2(n_212),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_188),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_294),
.Y(n_348)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_218),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_212),
.A2(n_197),
.B1(n_188),
.B2(n_221),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_293),
.A2(n_224),
.B1(n_226),
.B2(n_279),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_146),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_172),
.B(n_221),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_295),
.B(n_297),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_146),
.B(n_161),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_146),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_298),
.B(n_300),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_171),
.B(n_118),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_299),
.B(n_243),
.Y(n_349)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_213),
.Y(n_300)
);

AND2x2_ASAP7_75t_SL g302 ( 
.A(n_242),
.B(n_253),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_302),
.B(n_323),
.Y(n_365)
);

OAI32xp33_ASAP7_75t_L g304 ( 
.A1(n_225),
.A2(n_270),
.A3(n_242),
.B1(n_262),
.B2(n_252),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_304),
.B(n_321),
.Y(n_400)
);

NAND2xp67_ASAP7_75t_L g309 ( 
.A(n_225),
.B(n_233),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_309),
.B(n_255),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_236),
.A2(n_229),
.B1(n_265),
.B2(n_230),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_311),
.A2(n_303),
.B1(n_305),
.B2(n_347),
.Y(n_390)
);

OAI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_317),
.A2(n_300),
.B1(n_254),
.B2(n_231),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_227),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_326),
.B(n_259),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_256),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_330),
.B(n_341),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_296),
.A2(n_234),
.B1(n_229),
.B2(n_241),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_332),
.A2(n_346),
.B1(n_317),
.B2(n_334),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_256),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_286),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_330),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_241),
.A2(n_269),
.B1(n_292),
.B2(n_235),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_297),
.B(n_244),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_347),
.B(n_350),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_349),
.B(n_359),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_L g350 ( 
.A1(n_269),
.A2(n_278),
.B(n_243),
.C(n_232),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_223),
.B(n_228),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_351),
.B(n_295),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_282),
.B(n_280),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_354),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_276),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_299),
.B(n_246),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_351),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_360),
.B(n_373),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_302),
.B(n_289),
.C(n_272),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_364),
.C(n_379),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_280),
.C(n_277),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_377),
.B1(n_406),
.B2(n_354),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_240),
.B(n_247),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_367),
.A2(n_374),
.B(n_386),
.Y(n_425)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_370),
.B(n_390),
.Y(n_436)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_372),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_353),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_322),
.A2(n_237),
.B(n_268),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_375),
.B(n_383),
.Y(n_422)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_332),
.A2(n_268),
.B1(n_251),
.B2(n_258),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_325),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_378),
.B(n_382),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_308),
.Y(n_380)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_380),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_381),
.A2(n_356),
.B(n_335),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_353),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_342),
.B(n_238),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_340),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_384),
.B(n_388),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_356),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_385),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_316),
.A2(n_298),
.B(n_294),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_306),
.B(n_266),
.C(n_267),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_389),
.C(n_335),
.Y(n_444)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_305),
.B(n_271),
.Y(n_389)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_319),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_391),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_316),
.A2(n_261),
.B(n_273),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_396),
.B(n_320),
.Y(n_429)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_393),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_301),
.A2(n_288),
.B1(n_291),
.B2(n_261),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_394),
.A2(n_339),
.B1(n_333),
.B2(n_343),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_331),
.B(n_309),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_395),
.B(n_402),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_326),
.A2(n_336),
.B(n_350),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_353),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_397),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_321),
.B(n_307),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_398),
.B(n_399),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_348),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_310),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_405),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_354),
.B(n_357),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_404),
.B(n_344),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_310),
.B(n_304),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_396),
.A2(n_336),
.B(n_341),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_SL g466 ( 
.A1(n_407),
.A2(n_433),
.B(n_381),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_390),
.A2(n_346),
.B1(n_334),
.B2(n_338),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_408),
.A2(n_417),
.B1(n_441),
.B2(n_360),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_369),
.B(n_318),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_413),
.B(n_370),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_414),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_406),
.A2(n_306),
.B1(n_344),
.B2(n_324),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_415),
.A2(n_427),
.B1(n_428),
.B2(n_438),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_383),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_421),
.B(n_426),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_442),
.C(n_364),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_375),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_377),
.A2(n_306),
.B1(n_344),
.B2(n_324),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_365),
.A2(n_324),
.B1(n_329),
.B2(n_314),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_429),
.A2(n_432),
.B(n_367),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_365),
.A2(n_386),
.B(n_363),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_365),
.A2(n_329),
.B1(n_314),
.B2(n_352),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_363),
.B(n_312),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_444),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_405),
.A2(n_327),
.B1(n_343),
.B2(n_333),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_379),
.B(n_358),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_401),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_445),
.B(n_399),
.Y(n_451)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_418),
.Y(n_446)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_446),
.Y(n_483)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_449),
.A2(n_455),
.B1(n_458),
.B2(n_459),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_450),
.B(n_463),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_451),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_409),
.B(n_395),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_460),
.C(n_474),
.Y(n_482)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_434),
.Y(n_453)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_453),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_441),
.A2(n_403),
.B1(n_362),
.B2(n_404),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_421),
.A2(n_362),
.B1(n_404),
.B2(n_387),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_445),
.A2(n_381),
.B1(n_371),
.B2(n_368),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_409),
.B(n_389),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_440),
.Y(n_461)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_461),
.Y(n_511)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_440),
.Y(n_462)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_462),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_431),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_429),
.B(n_425),
.Y(n_486)
);

MAJx2_ASAP7_75t_L g509 ( 
.A(n_465),
.B(n_416),
.C(n_313),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_466),
.A2(n_425),
.B(n_420),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_426),
.B(n_378),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_469),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_414),
.A2(n_400),
.B1(n_394),
.B2(n_361),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_468),
.A2(n_408),
.B1(n_422),
.B2(n_407),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_437),
.B(n_376),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_423),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_470),
.B(n_472),
.Y(n_496)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_423),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_471),
.B(n_478),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_413),
.B(n_328),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g485 ( 
.A1(n_473),
.A2(n_475),
.B1(n_476),
.B2(n_478),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_443),
.B(n_374),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_435),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_431),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_442),
.B(n_373),
.C(n_382),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_477),
.B(n_479),
.C(n_430),
.Y(n_507)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_420),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_358),
.C(n_388),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_437),
.B(n_384),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_480),
.A2(n_481),
.B1(n_410),
.B2(n_419),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_422),
.B(n_393),
.Y(n_481)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_485),
.Y(n_516)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_486),
.A2(n_501),
.B(n_504),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_443),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_490),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_489),
.A2(n_510),
.B(n_513),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_465),
.B(n_415),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_491),
.B(n_372),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_424),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_492),
.B(n_498),
.Y(n_533)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_493),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_457),
.B(n_424),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_456),
.A2(n_436),
.B1(n_438),
.B2(n_428),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_499),
.A2(n_446),
.B1(n_391),
.B2(n_418),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_456),
.A2(n_417),
.B1(n_433),
.B2(n_411),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_500),
.A2(n_503),
.B1(n_501),
.B2(n_510),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_454),
.A2(n_468),
.B1(n_462),
.B2(n_461),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_454),
.A2(n_411),
.B1(n_436),
.B2(n_410),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_464),
.B(n_432),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_457),
.B(n_439),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_506),
.B(n_508),
.C(n_509),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_507),
.B(n_447),
.C(n_471),
.Y(n_528)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_479),
.B(n_427),
.C(n_416),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_474),
.A2(n_392),
.B(n_419),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_466),
.A2(n_412),
.B(n_320),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_458),
.B(n_412),
.C(n_308),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_514),
.B(n_339),
.C(n_337),
.Y(n_543)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_502),
.Y(n_518)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_518),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_484),
.B(n_448),
.Y(n_519)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_519),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_494),
.B(n_467),
.Y(n_520)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_484),
.B(n_481),
.Y(n_521)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_521),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_499),
.A2(n_477),
.B1(n_469),
.B2(n_480),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_523),
.A2(n_535),
.B1(n_541),
.B2(n_508),
.Y(n_561)
);

FAx1_ASAP7_75t_SL g524 ( 
.A(n_482),
.B(n_455),
.CI(n_449),
.CON(n_524),
.SN(n_524)
);

A2O1A1Ixp33_ASAP7_75t_L g548 ( 
.A1(n_524),
.A2(n_489),
.B(n_482),
.C(n_491),
.Y(n_548)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_502),
.Y(n_525)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_497),
.B(n_453),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_526),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_528),
.B(n_507),
.C(n_509),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_512),
.Y(n_529)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_529),
.Y(n_554)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_503),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_530),
.B(n_536),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_495),
.B(n_505),
.Y(n_531)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_531),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_532),
.A2(n_530),
.B1(n_517),
.B2(n_541),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_514),
.Y(n_534)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_534),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_496),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_483),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_537),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_539),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_513),
.B(n_380),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_540),
.B(n_504),
.Y(n_559)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_488),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_486),
.A2(n_355),
.B(n_345),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_542),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_487),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_548),
.A2(n_538),
.B(n_515),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_549),
.B(n_561),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_SL g552 ( 
.A(n_533),
.B(n_498),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_565),
.Y(n_578)
);

BUFx12_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_557),
.Y(n_567)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_558),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_559),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_563),
.B(n_527),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_532),
.A2(n_504),
.B1(n_490),
.B2(n_492),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_564),
.B(n_524),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_527),
.B(n_506),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_568),
.B(n_581),
.Y(n_600)
);

BUFx24_ASAP7_75t_SL g569 ( 
.A(n_546),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g590 ( 
.A(n_569),
.B(n_576),
.Y(n_590)
);

FAx1_ASAP7_75t_SL g570 ( 
.A(n_563),
.B(n_519),
.CI(n_522),
.CON(n_570),
.SN(n_570)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_570),
.B(n_579),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_550),
.B(n_536),
.Y(n_571)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_571),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_549),
.B(n_528),
.C(n_527),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_574),
.B(n_580),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_575),
.B(n_515),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_520),
.Y(n_576)
);

BUFx24_ASAP7_75t_SL g579 ( 
.A(n_560),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_565),
.B(n_522),
.C(n_534),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_558),
.B(n_522),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_560),
.B(n_526),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_582),
.B(n_584),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_550),
.B(n_531),
.Y(n_583)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_583),
.Y(n_601)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_556),
.A2(n_538),
.B(n_523),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g593 ( 
.A1(n_585),
.A2(n_540),
.B(n_539),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_552),
.C(n_564),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_586),
.B(n_588),
.C(n_589),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_543),
.C(n_533),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_543),
.C(n_533),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_591),
.B(n_597),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_593),
.B(n_594),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_572),
.A2(n_548),
.B1(n_517),
.B2(n_547),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_SL g595 ( 
.A1(n_572),
.A2(n_566),
.B1(n_544),
.B2(n_516),
.Y(n_595)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_595),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_570),
.B(n_516),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_581),
.B(n_551),
.C(n_535),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_599),
.B(n_589),
.C(n_588),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_596),
.B(n_553),
.Y(n_602)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_602),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_601),
.B(n_553),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_603),
.B(n_608),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_590),
.B(n_573),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_605),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_587),
.B(n_580),
.Y(n_605)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_595),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_599),
.B(n_524),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_609),
.B(n_613),
.Y(n_618)
);

INVx11_ASAP7_75t_L g610 ( 
.A(n_594),
.Y(n_610)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_610),
.B(n_611),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_600),
.B(n_524),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_606),
.B(n_592),
.C(n_598),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_617),
.B(n_620),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_606),
.B(n_611),
.Y(n_619)
);

INVxp33_ASAP7_75t_L g628 ( 
.A(n_619),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_602),
.B(n_554),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_612),
.B(n_600),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_621),
.B(n_603),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_607),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_622),
.A2(n_578),
.B1(n_554),
.B2(n_555),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_615),
.B(n_607),
.C(n_586),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_626),
.B(n_630),
.Y(n_634)
);

AOI321xp33_ASAP7_75t_SL g627 ( 
.A1(n_618),
.A2(n_610),
.A3(n_608),
.B1(n_614),
.B2(n_567),
.C(n_593),
.Y(n_627)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_627),
.A2(n_629),
.B(n_623),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g635 ( 
.A(n_631),
.B(n_632),
.C(n_633),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_628),
.A2(n_625),
.B(n_627),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_625),
.A2(n_624),
.B(n_616),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_634),
.B(n_616),
.C(n_555),
.Y(n_636)
);

AOI221xp5_ASAP7_75t_L g637 ( 
.A1(n_636),
.A2(n_562),
.B1(n_525),
.B2(n_518),
.C(n_529),
.Y(n_637)
);

XNOR2xp5_ASAP7_75t_L g638 ( 
.A(n_637),
.B(n_635),
.Y(n_638)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_578),
.Y(n_639)
);


endmodule