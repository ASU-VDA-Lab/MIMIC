module fake_jpeg_30031_n_100 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_21),
.B(n_2),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_38),
.B(n_42),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_45),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_62)
);

AOI21xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_1),
.B(n_3),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_49),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_1),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_57),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_62),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_37),
.B1(n_33),
.B2(n_43),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_3),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_5),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_58),
.A2(n_47),
.B1(n_50),
.B2(n_48),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_56),
.B(n_4),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_18),
.Y(n_84)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_62),
.B(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_8),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_72),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_20),
.B(n_24),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_74),
.Y(n_83)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_75),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_72),
.A2(n_53),
.B1(n_13),
.B2(n_15),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_76),
.A2(n_79),
.B1(n_86),
.B2(n_75),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_12),
.B1(n_16),
.B2(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_25),
.C(n_26),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_67),
.B(n_63),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_80),
.Y(n_89)
);

AO221x1_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_91),
.B1(n_76),
.B2(n_77),
.C(n_31),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_77),
.C(n_85),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_93),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_95),
.B(n_83),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_87),
.B1(n_85),
.B2(n_89),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_68),
.B1(n_78),
.B2(n_32),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_78),
.C(n_27),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_30),
.Y(n_100)
);


endmodule