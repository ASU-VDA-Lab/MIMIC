module fake_netlist_5_1122_n_2077 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2077);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2077;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_877;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2038;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_2034;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_199),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_114),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_32),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_97),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_72),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_138),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_145),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_99),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_16),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_28),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_72),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_105),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_121),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_64),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_176),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_19),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_47),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_21),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_164),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_78),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_17),
.Y(n_227)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_26),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_60),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_54),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_104),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_40),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_184),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_81),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_103),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_34),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_155),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_160),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_163),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_192),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_14),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_142),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_113),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_165),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_17),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_70),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_133),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_139),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_124),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_2),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_93),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_85),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_28),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_200),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_62),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_53),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_51),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_64),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_175),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_151),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_125),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_158),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_117),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_156),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_187),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_152),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_193),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_35),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_179),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_67),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_146),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_53),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_70),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_58),
.Y(n_275)
);

BUFx8_ASAP7_75t_SL g276 ( 
.A(n_106),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_13),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_118),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_161),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_111),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_132),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_141),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_95),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_162),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_68),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_21),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_98),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_25),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_14),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_122),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_108),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_54),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_196),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_171),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_166),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_35),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_79),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_1),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_40),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_13),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_22),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_6),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_60),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_195),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_110),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_185),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_4),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_16),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_144),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_129),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_63),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_19),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_68),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_120),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_7),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_88),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_157),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_194),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_119),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_127),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_148),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_169),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_12),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_96),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_23),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_23),
.Y(n_330)
);

BUFx10_ASAP7_75t_L g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_130),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_173),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_198),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_65),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_143),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_46),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_0),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_123),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_190),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_91),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_76),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_67),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_57),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_48),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_89),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_82),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_4),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_137),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_167),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_59),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_8),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_149),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_61),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_62),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_58),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_38),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_134),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_112),
.Y(n_359)
);

CKINVDCx11_ASAP7_75t_R g360 ( 
.A(n_10),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_43),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_22),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_27),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_135),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_92),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_46),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_94),
.Y(n_367)
);

BUFx5_ASAP7_75t_L g368 ( 
.A(n_15),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_27),
.Y(n_369)
);

INVx1_ASAP7_75t_SL g370 ( 
.A(n_15),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_38),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_33),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_153),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_1),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_71),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_197),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_12),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_186),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_56),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_31),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_11),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_5),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_51),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_80),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_31),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_90),
.Y(n_386)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_150),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_25),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_87),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_10),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_42),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_29),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_178),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_180),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_43),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_188),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_84),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_74),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_52),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_75),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_244),
.B(n_0),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_276),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_368),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_230),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_368),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_368),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_368),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_241),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_226),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_2),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_260),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_R g412 ( 
.A(n_201),
.B(n_204),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_284),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_360),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_294),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_243),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_245),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_237),
.B(n_3),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_248),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_368),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_319),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_368),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_329),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_271),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_250),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_271),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_323),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_271),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_271),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_314),
.B(n_3),
.Y(n_432)
);

BUFx6f_ASAP7_75t_SL g433 ( 
.A(n_249),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_271),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_295),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_345),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_253),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_255),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_295),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_228),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_206),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_262),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_263),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_387),
.B(n_5),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_396),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_295),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_295),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_278),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_295),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_264),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_324),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_265),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_267),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_268),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_272),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_312),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_324),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_279),
.Y(n_458)
);

BUFx6f_ASAP7_75t_SL g459 ( 
.A(n_249),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_280),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_282),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_324),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g463 ( 
.A(n_226),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_324),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_206),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g466 ( 
.A(n_214),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_292),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_297),
.Y(n_468)
);

INVxp33_ASAP7_75t_SL g469 ( 
.A(n_214),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_215),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_329),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_324),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_332),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_387),
.B(n_6),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_299),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g476 ( 
.A(n_203),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_249),
.Y(n_477)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_281),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_307),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_308),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_361),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_361),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_347),
.B(n_9),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_361),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_361),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_361),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_313),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_322),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_325),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_326),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_328),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_329),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_258),
.Y(n_493)
);

NOR2xp67_ASAP7_75t_L g494 ( 
.A(n_390),
.B(n_9),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_258),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_343),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_333),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_334),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_336),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_386),
.B(n_11),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_340),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_406),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_441),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_425),
.B(n_211),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_465),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_471),
.B(n_211),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_406),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_426),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_423),
.Y(n_509)
);

CKINVDCx6p67_ASAP7_75t_R g510 ( 
.A(n_473),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_426),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_428),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_430),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_430),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_423),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_403),
.Y(n_517)
);

INVx6_ASAP7_75t_L g518 ( 
.A(n_463),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_L g519 ( 
.A(n_432),
.B(n_390),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_492),
.B(n_219),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_410),
.B(n_281),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_440),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_403),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_444),
.B(n_201),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_474),
.B(n_204),
.Y(n_526)
);

AND2x2_ASAP7_75t_SL g527 ( 
.A(n_432),
.B(n_219),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_405),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_431),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_407),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_463),
.B(n_252),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_407),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_431),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_492),
.B(n_252),
.Y(n_535)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_416),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_448),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_434),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_421),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_421),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_424),
.Y(n_542)
);

CKINVDCx11_ASAP7_75t_R g543 ( 
.A(n_404),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g544 ( 
.A(n_401),
.B(n_266),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_434),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_435),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_435),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_439),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_439),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_463),
.B(n_266),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_446),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_447),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_449),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_449),
.Y(n_557)
);

OR2x6_ASAP7_75t_L g558 ( 
.A(n_494),
.B(n_296),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_477),
.A2(n_330),
.B1(n_285),
.B2(n_257),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_451),
.Y(n_560)
);

NOR2x1_ASAP7_75t_L g561 ( 
.A(n_451),
.B(n_296),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_466),
.B(n_317),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_457),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_457),
.B(n_462),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_462),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_409),
.B(n_378),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_470),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_494),
.B(n_228),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_409),
.B(n_378),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_472),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_481),
.B(n_482),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_481),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_482),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_484),
.B(n_240),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_484),
.B(n_209),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_485),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_456),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_558),
.B(n_522),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_504),
.B(n_496),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_518),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_509),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_577),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_518),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_518),
.Y(n_588)
);

BUFx4f_ASAP7_75t_L g589 ( 
.A(n_527),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_577),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_502),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_SL g592 ( 
.A(n_522),
.B(n_433),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_523),
.B(n_433),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g594 ( 
.A(n_562),
.B(n_417),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_527),
.B(n_418),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_570),
.B(n_477),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_518),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_509),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_523),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_544),
.A2(n_500),
.B1(n_483),
.B2(n_343),
.Y(n_600)
);

BUFx6f_ASAP7_75t_SL g601 ( 
.A(n_544),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

AND2x2_ASAP7_75t_SL g603 ( 
.A(n_527),
.B(n_544),
.Y(n_603)
);

BUFx6f_ASAP7_75t_SL g604 ( 
.A(n_544),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_509),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_502),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_505),
.B(n_436),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_577),
.Y(n_608)
);

XOR2x2_ASAP7_75t_L g609 ( 
.A(n_562),
.B(n_419),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_570),
.B(n_478),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_L g611 ( 
.A1(n_544),
.A2(n_475),
.B1(n_501),
.B2(n_490),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_527),
.B(n_420),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_577),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g614 ( 
.A(n_581),
.Y(n_614)
);

INVxp33_ASAP7_75t_SL g615 ( 
.A(n_570),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_574),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_527),
.B(n_478),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_574),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_518),
.Y(n_620)
);

INVxp33_ASAP7_75t_SL g621 ( 
.A(n_538),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_574),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_518),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_518),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_525),
.B(n_427),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_577),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_574),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_547),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_574),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_577),
.Y(n_630)
);

AND3x2_ASAP7_75t_L g631 ( 
.A(n_523),
.B(n_289),
.C(n_251),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_SL g632 ( 
.A(n_559),
.B(n_419),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_531),
.Y(n_633)
);

AO21x2_ASAP7_75t_L g634 ( 
.A1(n_525),
.A2(n_205),
.B(n_202),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_531),
.Y(n_635)
);

OR2x6_ASAP7_75t_L g636 ( 
.A(n_558),
.B(n_207),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_502),
.Y(n_637)
);

XNOR2x2_ASAP7_75t_L g638 ( 
.A(n_538),
.B(n_300),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_502),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_504),
.B(n_506),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_505),
.B(n_436),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_504),
.B(n_506),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_504),
.B(n_240),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_574),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_578),
.B(n_437),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_502),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_503),
.A2(n_242),
.B1(n_567),
.B2(n_370),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_506),
.B(n_493),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_543),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_531),
.Y(n_650)
);

BUFx2_ASAP7_75t_L g651 ( 
.A(n_503),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_506),
.B(n_438),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_578),
.B(n_442),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_548),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_548),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_502),
.Y(n_656)
);

AND3x2_ASAP7_75t_L g657 ( 
.A(n_567),
.B(n_374),
.C(n_352),
.Y(n_657)
);

BUFx6f_ASAP7_75t_L g658 ( 
.A(n_502),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_531),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_526),
.B(n_443),
.Y(n_660)
);

OR2x6_ASAP7_75t_L g661 ( 
.A(n_558),
.B(n_235),
.Y(n_661)
);

BUFx10_ASAP7_75t_L g662 ( 
.A(n_558),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_526),
.B(n_450),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_548),
.Y(n_664)
);

AOI22xp33_ASAP7_75t_L g665 ( 
.A1(n_558),
.A2(n_374),
.B1(n_377),
.B2(n_352),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_558),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_548),
.Y(n_667)
);

CKINVDCx16_ASAP7_75t_R g668 ( 
.A(n_581),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_531),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_553),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_532),
.B(n_452),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_553),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_532),
.B(n_453),
.Y(n_673)
);

NAND3xp33_ASAP7_75t_L g674 ( 
.A(n_519),
.B(n_486),
.C(n_412),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_553),
.Y(n_675)
);

INVx4_ASAP7_75t_SL g676 ( 
.A(n_558),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_559),
.B(n_454),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_532),
.B(n_455),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_502),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_531),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_553),
.Y(n_681)
);

INVx8_ASAP7_75t_L g682 ( 
.A(n_558),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_536),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_532),
.B(n_458),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_519),
.B(n_486),
.C(n_261),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_507),
.Y(n_686)
);

NAND3xp33_ASAP7_75t_L g687 ( 
.A(n_551),
.B(n_270),
.C(n_236),
.Y(n_687)
);

INVx3_ASAP7_75t_L g688 ( 
.A(n_507),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_536),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_566),
.B(n_283),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_507),
.Y(n_691)
);

BUFx4f_ASAP7_75t_L g692 ( 
.A(n_528),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_510),
.A2(n_298),
.B1(n_246),
.B2(n_247),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_554),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_554),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_554),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_551),
.B(n_460),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_551),
.B(n_461),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_554),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_556),
.Y(n_700)
);

BUFx3_ASAP7_75t_L g701 ( 
.A(n_547),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_507),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_536),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_536),
.Y(n_704)
);

INVxp33_ASAP7_75t_L g705 ( 
.A(n_543),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_536),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_507),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_536),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_542),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_556),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_542),
.Y(n_711)
);

BUFx6f_ASAP7_75t_L g712 ( 
.A(n_507),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_566),
.B(n_467),
.Y(n_713)
);

AND2x2_ASAP7_75t_SL g714 ( 
.A(n_551),
.B(n_240),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_542),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_507),
.Y(n_716)
);

NAND3xp33_ASAP7_75t_L g717 ( 
.A(n_566),
.B(n_288),
.C(n_287),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_566),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_521),
.A2(n_377),
.B1(n_348),
.B2(n_314),
.Y(n_719)
);

INVx4_ASAP7_75t_SL g720 ( 
.A(n_528),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_571),
.B(n_493),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_556),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_542),
.B(n_468),
.Y(n_723)
);

BUFx3_ASAP7_75t_L g724 ( 
.A(n_547),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_571),
.B(n_479),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_571),
.B(n_480),
.Y(n_726)
);

AO22x2_ASAP7_75t_L g727 ( 
.A1(n_571),
.A2(n_383),
.B1(n_305),
.B2(n_304),
.Y(n_727)
);

INVx5_ASAP7_75t_L g728 ( 
.A(n_528),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_521),
.B(n_487),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_556),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_547),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_542),
.Y(n_732)
);

BUFx6f_ASAP7_75t_L g733 ( 
.A(n_507),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_581),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_625),
.B(n_488),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_585),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_586),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_586),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_663),
.B(n_489),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_585),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_642),
.B(n_491),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_628),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_598),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_598),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_642),
.B(n_603),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_594),
.B(n_497),
.Y(n_746)
);

NOR2x1p5_ASAP7_75t_L g747 ( 
.A(n_607),
.B(n_510),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_603),
.B(n_498),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_590),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_603),
.B(n_499),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_718),
.B(n_542),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_718),
.B(n_546),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_589),
.B(n_714),
.Y(n_753)
);

A2O1A1Ixp33_ASAP7_75t_L g754 ( 
.A1(n_589),
.A2(n_640),
.B(n_600),
.C(n_583),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_714),
.B(n_546),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_714),
.B(n_546),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_660),
.B(n_595),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_602),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_612),
.B(n_546),
.Y(n_759)
);

NAND3xp33_ASAP7_75t_L g760 ( 
.A(n_674),
.B(n_402),
.C(n_256),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_590),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_608),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_608),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_721),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_589),
.B(n_528),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_613),
.Y(n_766)
);

OR2x2_ASAP7_75t_L g767 ( 
.A(n_599),
.B(n_510),
.Y(n_767)
);

AND2x4_ASAP7_75t_L g768 ( 
.A(n_721),
.B(n_552),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_583),
.B(n_546),
.Y(n_769)
);

O2A1O1Ixp33_ASAP7_75t_L g770 ( 
.A1(n_617),
.A2(n_546),
.B(n_524),
.C(n_529),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_652),
.B(n_552),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_725),
.B(n_552),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_648),
.B(n_552),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_601),
.A2(n_535),
.B1(n_521),
.B2(n_524),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_648),
.B(n_555),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_613),
.Y(n_776)
);

AND2x6_ASAP7_75t_SL g777 ( 
.A(n_632),
.B(n_208),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_602),
.Y(n_778)
);

INVxp33_ASAP7_75t_L g779 ( 
.A(n_607),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_601),
.A2(n_411),
.B1(n_413),
.B2(n_408),
.Y(n_780)
);

BUFx5_ASAP7_75t_L g781 ( 
.A(n_633),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_601),
.A2(n_535),
.B1(n_521),
.B2(n_524),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_615),
.B(n_645),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_676),
.B(n_528),
.Y(n_784)
);

O2A1O1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_671),
.A2(n_524),
.B(n_529),
.C(n_517),
.Y(n_785)
);

INVxp67_ASAP7_75t_L g786 ( 
.A(n_651),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_676),
.B(n_528),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_621),
.Y(n_788)
);

NOR3xp33_ASAP7_75t_L g789 ( 
.A(n_611),
.B(n_414),
.C(n_269),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_615),
.B(n_469),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_676),
.B(n_528),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_682),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_599),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_626),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_676),
.B(n_555),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_SL g796 ( 
.A(n_604),
.B(n_433),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_666),
.B(n_528),
.Y(n_797)
);

BUFx8_ASAP7_75t_L g798 ( 
.A(n_651),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_645),
.B(n_415),
.Y(n_799)
);

INVx4_ASAP7_75t_L g800 ( 
.A(n_682),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_596),
.B(n_273),
.C(n_254),
.Y(n_801)
);

NAND3xp33_ASAP7_75t_L g802 ( 
.A(n_674),
.B(n_275),
.C(n_274),
.Y(n_802)
);

AND2x6_ASAP7_75t_SL g803 ( 
.A(n_632),
.B(n_213),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_723),
.B(n_555),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_666),
.B(n_616),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_626),
.B(n_630),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_616),
.B(n_528),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_618),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_630),
.Y(n_809)
);

AOI22xp33_ASAP7_75t_L g810 ( 
.A1(n_604),
.A2(n_521),
.B1(n_535),
.B2(n_517),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_605),
.Y(n_811)
);

NAND2xp33_ASAP7_75t_L g812 ( 
.A(n_682),
.B(n_643),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_628),
.B(n_555),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_618),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_673),
.B(n_517),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_622),
.B(n_240),
.Y(n_816)
);

A2O1A1Ixp33_ASAP7_75t_L g817 ( 
.A1(n_665),
.A2(n_521),
.B(n_535),
.C(n_259),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_678),
.B(n_517),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_605),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_604),
.A2(n_422),
.B1(n_429),
.B2(n_445),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_622),
.B(n_240),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_684),
.B(n_529),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_634),
.A2(n_535),
.B1(n_529),
.B2(n_541),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_SL g824 ( 
.A(n_647),
.B(n_222),
.C(n_215),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_641),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_697),
.B(n_533),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_627),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_627),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_629),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_653),
.B(n_698),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_629),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_653),
.B(n_476),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_644),
.B(n_533),
.Y(n_833)
);

HB1xp67_ASAP7_75t_L g834 ( 
.A(n_734),
.Y(n_834)
);

BUFx4_ASAP7_75t_L g835 ( 
.A(n_621),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_641),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_644),
.B(n_309),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_633),
.B(n_533),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_635),
.B(n_533),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_635),
.B(n_537),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_650),
.B(n_537),
.Y(n_841)
);

INVx2_ASAP7_75t_SL g842 ( 
.A(n_713),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_619),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_734),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_726),
.Y(n_845)
);

NOR2xp67_ASAP7_75t_L g846 ( 
.A(n_685),
.B(n_520),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_650),
.B(n_537),
.Y(n_847)
);

INVx4_ASAP7_75t_L g848 ( 
.A(n_682),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_654),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_662),
.B(n_659),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_654),
.Y(n_851)
);

NAND2x1_ASAP7_75t_L g852 ( 
.A(n_584),
.B(n_520),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_662),
.B(n_309),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_655),
.Y(n_854)
);

NAND2x1_ASAP7_75t_L g855 ( 
.A(n_584),
.B(n_520),
.Y(n_855)
);

OR2x2_ASAP7_75t_L g856 ( 
.A(n_614),
.B(n_510),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_655),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_662),
.B(n_309),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_662),
.B(n_309),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_659),
.B(n_537),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_664),
.Y(n_861)
);

AND3x1_ASAP7_75t_L g862 ( 
.A(n_647),
.B(n_227),
.C(n_218),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_582),
.A2(n_306),
.B1(n_320),
.B2(n_321),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_620),
.A2(n_564),
.B(n_541),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_669),
.B(n_680),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_634),
.A2(n_535),
.B1(n_540),
.B2(n_541),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_669),
.B(n_540),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_680),
.B(n_309),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_631),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_683),
.B(n_540),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_664),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_610),
.B(n_433),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_683),
.B(n_540),
.Y(n_873)
);

OR2x6_ASAP7_75t_L g874 ( 
.A(n_682),
.B(n_348),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_643),
.B(n_339),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_634),
.A2(n_541),
.B1(n_520),
.B2(n_561),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_689),
.B(n_520),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_689),
.B(n_520),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_717),
.A2(n_355),
.B(n_277),
.C(n_302),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_677),
.B(n_459),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_703),
.B(n_339),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_667),
.Y(n_882)
);

OAI21xp33_ASAP7_75t_L g883 ( 
.A1(n_719),
.A2(n_327),
.B(n_303),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_703),
.B(n_339),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_667),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_670),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_638),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_614),
.B(n_228),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_701),
.Y(n_889)
);

NAND2xp33_ASAP7_75t_L g890 ( 
.A(n_643),
.B(n_342),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_704),
.B(n_339),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_704),
.B(n_507),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_706),
.B(n_516),
.Y(n_893)
);

NOR3xp33_ASAP7_75t_L g894 ( 
.A(n_668),
.B(n_693),
.C(n_729),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_706),
.B(n_516),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_708),
.B(n_516),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_708),
.B(n_516),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_709),
.B(n_516),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_582),
.A2(n_690),
.B1(n_592),
.B2(n_593),
.Y(n_899)
);

OAI22xp33_ASAP7_75t_L g900 ( 
.A1(n_582),
.A2(n_353),
.B1(n_359),
.B2(n_341),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_657),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_670),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_709),
.B(n_516),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_701),
.Y(n_904)
);

A2O1A1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_717),
.A2(n_362),
.B(n_344),
.C(n_351),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_711),
.B(n_508),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_844),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_757),
.B(n_582),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_765),
.A2(n_692),
.B(n_623),
.Y(n_909)
);

BUFx5_ASAP7_75t_L g910 ( 
.A(n_795),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_765),
.A2(n_692),
.B(n_623),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_830),
.B(n_582),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_746),
.B(n_724),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_815),
.A2(n_692),
.B(n_620),
.Y(n_914)
);

INVxp67_ASAP7_75t_L g915 ( 
.A(n_834),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_783),
.B(n_668),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_745),
.A2(n_685),
.B(n_687),
.C(n_724),
.Y(n_917)
);

A2O1A1Ixp33_ASAP7_75t_L g918 ( 
.A1(n_754),
.A2(n_687),
.B(n_731),
.C(n_715),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_735),
.B(n_731),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_818),
.A2(n_588),
.B(n_587),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_792),
.B(n_587),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_792),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_739),
.B(n_711),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_822),
.A2(n_826),
.B(n_812),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_808),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_843),
.A2(n_597),
.B(n_588),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_769),
.A2(n_624),
.B(n_597),
.Y(n_927)
);

AO21x1_ASAP7_75t_L g928 ( 
.A1(n_863),
.A2(n_389),
.B(n_384),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_792),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_793),
.Y(n_930)
);

O2A1O1Ixp5_ASAP7_75t_L g931 ( 
.A1(n_771),
.A2(n_715),
.B(n_732),
.C(n_730),
.Y(n_931)
);

NOR2x1_ASAP7_75t_SL g932 ( 
.A(n_800),
.B(n_636),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_764),
.B(n_742),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_804),
.A2(n_624),
.B(n_646),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_754),
.A2(n_802),
.B(n_748),
.C(n_750),
.Y(n_935)
);

INVxp67_ASAP7_75t_L g936 ( 
.A(n_832),
.Y(n_936)
);

AOI22xp5_ASAP7_75t_L g937 ( 
.A1(n_753),
.A2(n_690),
.B1(n_661),
.B2(n_636),
.Y(n_937)
);

AOI33xp33_ASAP7_75t_L g938 ( 
.A1(n_825),
.A2(n_398),
.A3(n_372),
.B1(n_366),
.B2(n_380),
.B3(n_363),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_753),
.A2(n_690),
.B1(n_661),
.B2(n_636),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_800),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_741),
.B(n_790),
.Y(n_941)
);

NAND3xp33_ASAP7_75t_L g942 ( 
.A(n_786),
.B(n_690),
.C(n_290),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_808),
.Y(n_943)
);

O2A1O1Ixp5_ASAP7_75t_L g944 ( 
.A1(n_759),
.A2(n_732),
.B(n_700),
.C(n_730),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_788),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_833),
.A2(n_656),
.B(n_646),
.Y(n_946)
);

O2A1O1Ixp33_ASAP7_75t_SL g947 ( 
.A1(n_900),
.A2(n_394),
.B(n_397),
.C(n_688),
.Y(n_947)
);

OAI22x1_ASAP7_75t_L g948 ( 
.A1(n_887),
.A2(n_780),
.B1(n_799),
.B2(n_836),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_755),
.A2(n_606),
.B(n_591),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_768),
.A2(n_845),
.B1(n_842),
.B2(n_805),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_813),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_773),
.A2(n_775),
.B(n_752),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_767),
.B(n_609),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_779),
.B(n_609),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_751),
.A2(n_656),
.B(n_646),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_808),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_756),
.A2(n_679),
.B(n_656),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_807),
.A2(n_702),
.B(n_679),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_807),
.A2(n_702),
.B(n_679),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_888),
.B(n_727),
.Y(n_960)
);

INVx3_ASAP7_75t_L g961 ( 
.A(n_813),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_779),
.B(n_638),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_805),
.A2(n_702),
.B(n_639),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_824),
.B(n_690),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_768),
.B(n_727),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_781),
.B(n_619),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_797),
.A2(n_639),
.B(n_619),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_770),
.A2(n_606),
.B(n_591),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_879),
.A2(n_636),
.B(n_661),
.C(n_382),
.Y(n_969)
);

A2O1A1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_880),
.A2(n_691),
.B(n_606),
.C(n_716),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_797),
.A2(n_639),
.B(n_619),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_828),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_813),
.Y(n_973)
);

NAND2x1p5_ASAP7_75t_L g974 ( 
.A(n_800),
.B(n_591),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_768),
.B(n_643),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_760),
.B(n_637),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_877),
.A2(n_639),
.B(n_619),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_781),
.B(n_639),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_878),
.A2(n_712),
.B(n_658),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_852),
.A2(n_712),
.B(n_658),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_772),
.A2(n_661),
.B1(n_636),
.B2(n_643),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_855),
.A2(n_712),
.B(n_658),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_742),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_781),
.B(n_658),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_814),
.B(n_827),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_829),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_795),
.Y(n_987)
);

OAI21xp33_ASAP7_75t_L g988 ( 
.A1(n_883),
.A2(n_727),
.B(n_223),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_829),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_850),
.A2(n_712),
.B(n_658),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_894),
.B(n_727),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_904),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_850),
.A2(n_733),
.B(n_712),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_795),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_831),
.Y(n_995)
);

AOI21xp33_ASAP7_75t_L g996 ( 
.A1(n_872),
.A2(n_661),
.B(n_705),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_879),
.A2(n_388),
.B(n_391),
.C(n_371),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_737),
.B(n_643),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_SL g999 ( 
.A(n_899),
.B(n_904),
.Y(n_999)
);

OAI21xp33_ASAP7_75t_L g1000 ( 
.A1(n_789),
.A2(n_223),
.B(n_222),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_738),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_798),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_806),
.A2(n_733),
.B(n_686),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_848),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_781),
.B(n_733),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_853),
.A2(n_733),
.B(n_686),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_781),
.B(n_733),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_749),
.B(n_643),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_848),
.B(n_649),
.Y(n_1009)
);

INVxp67_ASAP7_75t_R g1010 ( 
.A(n_820),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_761),
.B(n_637),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_853),
.A2(n_686),
.B(n_637),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_858),
.A2(n_691),
.B(n_688),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_905),
.A2(n_392),
.B(n_722),
.C(n_672),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_762),
.B(n_688),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_848),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_763),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_889),
.B(n_691),
.Y(n_1018)
);

AO21x1_ASAP7_75t_L g1019 ( 
.A1(n_858),
.A2(n_675),
.B(n_672),
.Y(n_1019)
);

NOR2x1p5_ASAP7_75t_L g1020 ( 
.A(n_856),
.B(n_224),
.Y(n_1020)
);

INVx3_ASAP7_75t_L g1021 ( 
.A(n_766),
.Y(n_1021)
);

OAI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_862),
.A2(n_229),
.B(n_224),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_776),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_849),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_794),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_859),
.A2(n_716),
.B(n_707),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_809),
.B(n_774),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_859),
.A2(n_716),
.B(n_707),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_865),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_782),
.A2(n_707),
.B1(n_225),
.B2(n_393),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_869),
.B(n_459),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_784),
.A2(n_728),
.B(n_681),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_784),
.A2(n_728),
.B(n_681),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_865),
.A2(n_694),
.B(n_675),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_781),
.B(n_720),
.Y(n_1035)
);

O2A1O1Ixp5_ASAP7_75t_L g1036 ( 
.A1(n_816),
.A2(n_694),
.B(n_722),
.C(n_695),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_785),
.A2(n_810),
.B(n_801),
.C(n_817),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_864),
.A2(n_696),
.B(n_695),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_798),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_781),
.B(n_696),
.Y(n_1040)
);

AND2x4_ASAP7_75t_L g1041 ( 
.A(n_901),
.B(n_649),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_787),
.A2(n_791),
.B(n_892),
.Y(n_1042)
);

HB1xp67_ASAP7_75t_L g1043 ( 
.A(n_874),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_874),
.A2(n_866),
.B1(n_823),
.B2(n_791),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_849),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_874),
.A2(n_212),
.B1(n_210),
.B2(n_239),
.Y(n_1046)
);

O2A1O1Ixp5_ASAP7_75t_L g1047 ( 
.A1(n_816),
.A2(n_699),
.B(n_700),
.C(n_710),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_851),
.B(n_699),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_906),
.B(n_459),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_851),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_R g1051 ( 
.A(n_835),
.B(n_229),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_787),
.A2(n_728),
.B(n_710),
.Y(n_1052)
);

AO21x1_ASAP7_75t_L g1053 ( 
.A1(n_821),
.A2(n_511),
.B(n_508),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_854),
.B(n_720),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_854),
.B(n_857),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_857),
.B(n_720),
.Y(n_1056)
);

O2A1O1Ixp5_ASAP7_75t_L g1057 ( 
.A1(n_821),
.A2(n_508),
.B(n_513),
.C(n_580),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_861),
.B(n_720),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_861),
.Y(n_1059)
);

BUFx2_ASAP7_75t_L g1060 ( 
.A(n_798),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_871),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_871),
.B(n_511),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_882),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_838),
.A2(n_728),
.B(n_564),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_882),
.B(n_511),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_885),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_885),
.B(n_512),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_839),
.A2(n_728),
.B(n_561),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_840),
.A2(n_561),
.B(n_728),
.Y(n_1069)
);

OAI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_841),
.A2(n_580),
.B(n_513),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_846),
.B(n_339),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_886),
.B(n_512),
.Y(n_1072)
);

AND2x4_ASAP7_75t_L g1073 ( 
.A(n_747),
.B(n_495),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_876),
.B(n_209),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_886),
.Y(n_1075)
);

AND2x2_ASAP7_75t_L g1076 ( 
.A(n_874),
.B(n_331),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_905),
.B(n_331),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_902),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_847),
.B(n_459),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_796),
.B(n_231),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_902),
.B(n_512),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_860),
.A2(n_557),
.B(n_579),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_867),
.A2(n_557),
.B(n_579),
.Y(n_1083)
);

INVx3_ASAP7_75t_L g1084 ( 
.A(n_736),
.Y(n_1084)
);

BUFx4f_ASAP7_75t_L g1085 ( 
.A(n_736),
.Y(n_1085)
);

NAND2xp33_ASAP7_75t_L g1086 ( 
.A(n_796),
.B(n_346),
.Y(n_1086)
);

A2O1A1Ixp33_ASAP7_75t_L g1087 ( 
.A1(n_817),
.A2(n_350),
.B(n_212),
.C(n_216),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_893),
.B(n_210),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_740),
.B(n_743),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_870),
.A2(n_557),
.B(n_579),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_873),
.B(n_286),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_837),
.A2(n_354),
.B(n_356),
.Y(n_1092)
);

AOI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_837),
.A2(n_232),
.B1(n_393),
.B2(n_367),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_740),
.B(n_513),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_903),
.B(n_216),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_743),
.B(n_514),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_744),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_895),
.A2(n_557),
.B(n_579),
.Y(n_1098)
);

AOI21x1_ASAP7_75t_L g1099 ( 
.A1(n_924),
.A2(n_897),
.B(n_896),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_930),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_930),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_940),
.A2(n_875),
.B(n_890),
.Y(n_1102)
);

OAI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1034),
.A2(n_898),
.B(n_819),
.Y(n_1103)
);

AND2x4_ASAP7_75t_SL g1104 ( 
.A(n_987),
.B(n_744),
.Y(n_1104)
);

NOR2xp33_ASAP7_75t_L g1105 ( 
.A(n_941),
.B(n_777),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1025),
.Y(n_1106)
);

INVx5_ASAP7_75t_L g1107 ( 
.A(n_1002),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_907),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_940),
.A2(n_875),
.B(n_758),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_SL g1110 ( 
.A(n_912),
.B(n_758),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_1084),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1025),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_936),
.A2(n_891),
.B(n_884),
.C(n_881),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_945),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_940),
.A2(n_819),
.B(n_778),
.Y(n_1115)
);

INVxp67_ASAP7_75t_L g1116 ( 
.A(n_915),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_933),
.B(n_778),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1001),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_933),
.B(n_811),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_L g1120 ( 
.A1(n_908),
.A2(n_811),
.B1(n_231),
.B2(n_233),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_936),
.B(n_217),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_940),
.A2(n_1044),
.B(n_913),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_950),
.B(n_217),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_952),
.A2(n_891),
.B(n_884),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_915),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_964),
.A2(n_881),
.B(n_868),
.C(n_367),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1023),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_964),
.A2(n_868),
.B(n_232),
.C(n_238),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_935),
.A2(n_225),
.B(n_221),
.C(n_234),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_954),
.B(n_803),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_1004),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_987),
.B(n_495),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1041),
.Y(n_1133)
);

O2A1O1Ixp5_ASAP7_75t_SL g1134 ( 
.A1(n_916),
.A2(n_580),
.B(n_514),
.C(n_575),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_994),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_SL g1136 ( 
.A1(n_953),
.A2(n_354),
.B1(n_400),
.B2(n_395),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1004),
.A2(n_579),
.B(n_568),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_1004),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_960),
.B(n_331),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_994),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_962),
.B(n_293),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_R g1142 ( 
.A(n_991),
.B(n_375),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_1004),
.Y(n_1143)
);

NAND2xp33_ASAP7_75t_SL g1144 ( 
.A(n_1016),
.B(n_220),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_1016),
.A2(n_579),
.B(n_568),
.Y(n_1145)
);

AOI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_999),
.A2(n_948),
.B1(n_965),
.B2(n_1010),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1091),
.B(n_514),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1027),
.A2(n_937),
.B1(n_962),
.B2(n_1017),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_983),
.B(n_992),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1091),
.B(n_515),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1016),
.A2(n_568),
.B(n_221),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1077),
.B(n_375),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_1016),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1039),
.Y(n_1154)
);

AOI22xp33_ASAP7_75t_L g1155 ( 
.A1(n_1074),
.A2(n_291),
.B1(n_373),
.B2(n_376),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_910),
.B(n_220),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_919),
.A2(n_349),
.B1(n_350),
.B2(n_358),
.Y(n_1157)
);

NOR3xp33_ASAP7_75t_L g1158 ( 
.A(n_996),
.B(n_318),
.C(n_301),
.Y(n_1158)
);

AO22x1_ASAP7_75t_L g1159 ( 
.A1(n_1041),
.A2(n_379),
.B1(n_400),
.B2(n_369),
.Y(n_1159)
);

CKINVDCx8_ASAP7_75t_R g1160 ( 
.A(n_1060),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_995),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_910),
.B(n_234),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1085),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_983),
.B(n_310),
.Y(n_1164)
);

CKINVDCx6p67_ASAP7_75t_R g1165 ( 
.A(n_1009),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1038),
.A2(n_568),
.B(n_575),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_923),
.B(n_515),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_942),
.A2(n_349),
.B1(n_358),
.B2(n_364),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_992),
.B(n_311),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1009),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1085),
.Y(n_1171)
);

BUFx2_ASAP7_75t_L g1172 ( 
.A(n_1073),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_910),
.B(n_238),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_1037),
.A2(n_239),
.B(n_364),
.C(n_365),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_SL g1175 ( 
.A(n_910),
.B(n_951),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1080),
.B(n_315),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1084),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_966),
.A2(n_568),
.B(n_365),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_966),
.A2(n_568),
.B(n_575),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1029),
.B(n_1017),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1021),
.B(n_515),
.Y(n_1181)
);

NAND2x1p5_ASAP7_75t_L g1182 ( 
.A(n_922),
.B(n_929),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_978),
.A2(n_560),
.B(n_573),
.Y(n_1183)
);

OAI22x1_ASAP7_75t_L g1184 ( 
.A1(n_1020),
.A2(n_356),
.B1(n_395),
.B2(n_385),
.Y(n_1184)
);

INVx6_ASAP7_75t_L g1185 ( 
.A(n_1073),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1000),
.B(n_316),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1021),
.B(n_335),
.Y(n_1187)
);

NOR2xp67_ASAP7_75t_SL g1188 ( 
.A(n_922),
.B(n_233),
.Y(n_1188)
);

OR2x6_ASAP7_75t_L g1189 ( 
.A(n_1043),
.B(n_530),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1076),
.B(n_375),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_1043),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1088),
.A2(n_530),
.B(n_572),
.C(n_569),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_951),
.B(n_530),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_988),
.B(n_1022),
.Y(n_1194)
);

OR2x6_ASAP7_75t_L g1195 ( 
.A(n_961),
.B(n_534),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1031),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_972),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_978),
.A2(n_560),
.B(n_573),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_976),
.A2(n_338),
.B(n_337),
.C(n_379),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1049),
.A2(n_281),
.B1(n_291),
.B2(n_373),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_961),
.B(n_534),
.Y(n_1201)
);

BUFx3_ASAP7_75t_L g1202 ( 
.A(n_910),
.Y(n_1202)
);

AO32x1_ASAP7_75t_L g1203 ( 
.A1(n_939),
.A2(n_549),
.A3(n_572),
.B1(n_569),
.B2(n_534),
.Y(n_1203)
);

OAI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1074),
.A2(n_981),
.B1(n_918),
.B2(n_917),
.Y(n_1204)
);

INVx5_ASAP7_75t_L g1205 ( 
.A(n_973),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_984),
.A2(n_563),
.B(n_573),
.Y(n_1206)
);

HB1xp67_ASAP7_75t_L g1207 ( 
.A(n_973),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_944),
.A2(n_545),
.B(n_572),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_984),
.A2(n_560),
.B(n_569),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1005),
.A2(n_565),
.B(n_563),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_925),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1031),
.B(n_357),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1005),
.A2(n_565),
.B(n_563),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_986),
.B(n_539),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1046),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_989),
.B(n_539),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_1024),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_R g1218 ( 
.A(n_1086),
.B(n_357),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_943),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_985),
.A2(n_369),
.B1(n_381),
.B2(n_385),
.Y(n_1220)
);

INVx2_ASAP7_75t_SL g1221 ( 
.A(n_1088),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_976),
.A2(n_381),
.B(n_565),
.C(n_539),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1049),
.B(n_549),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1050),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_969),
.A2(n_1042),
.B(n_1079),
.C(n_1087),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_1095),
.A2(n_1092),
.B(n_997),
.C(n_970),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1079),
.B(n_549),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_910),
.B(n_376),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_929),
.A2(n_545),
.B1(n_576),
.B2(n_550),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1051),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1007),
.A2(n_545),
.B(n_576),
.Y(n_1231)
);

O2A1O1Ixp5_ASAP7_75t_L g1232 ( 
.A1(n_1071),
.A2(n_376),
.B(n_373),
.C(n_291),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1095),
.Y(n_1233)
);

INVx5_ASAP7_75t_SL g1234 ( 
.A(n_956),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_998),
.A2(n_576),
.B(n_550),
.C(n_24),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1071),
.A2(n_18),
.B(n_20),
.C(n_24),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1045),
.B(n_576),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1059),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1007),
.A2(n_576),
.B(n_550),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1061),
.B(n_576),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_SL g1241 ( 
.A1(n_1093),
.A2(n_18),
.B1(n_20),
.B2(n_26),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1063),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1066),
.B(n_576),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_974),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_928),
.A2(n_576),
.B1(n_550),
.B2(n_32),
.Y(n_1245)
);

NOR3xp33_ASAP7_75t_SL g1246 ( 
.A(n_1030),
.B(n_29),
.C(n_30),
.Y(n_1246)
);

O2A1O1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_947),
.A2(n_30),
.B(n_33),
.C(n_36),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1075),
.B(n_576),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1078),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_975),
.A2(n_1040),
.B1(n_1097),
.B2(n_1008),
.Y(n_1250)
);

NAND2x1_ASAP7_75t_L g1251 ( 
.A(n_1055),
.B(n_550),
.Y(n_1251)
);

NOR3xp33_ASAP7_75t_SL g1252 ( 
.A(n_938),
.B(n_36),
.C(n_37),
.Y(n_1252)
);

OAI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_949),
.A2(n_550),
.B1(n_39),
.B2(n_41),
.Y(n_1253)
);

NOR3xp33_ASAP7_75t_L g1254 ( 
.A(n_1014),
.B(n_37),
.C(n_39),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1011),
.B(n_41),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1089),
.Y(n_1256)
);

AND2x2_ASAP7_75t_SL g1257 ( 
.A(n_1018),
.B(n_42),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_957),
.A2(n_550),
.B(n_77),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_974),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1018),
.B(n_1015),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_920),
.A2(n_550),
.B(n_83),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1048),
.Y(n_1262)
);

AOI31xp67_ASAP7_75t_L g1263 ( 
.A1(n_1110),
.A2(n_1081),
.A3(n_1096),
.B(n_1094),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1204),
.A2(n_1225),
.A3(n_1253),
.B(n_1019),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1118),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1122),
.A2(n_1069),
.B(n_914),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1141),
.A2(n_1053),
.B1(n_1035),
.B2(n_927),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1166),
.A2(n_944),
.B(n_990),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1127),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1176),
.A2(n_1057),
.B(n_1070),
.C(n_931),
.Y(n_1270)
);

AOI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1105),
.A2(n_1035),
.B1(n_1072),
.B2(n_1062),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1204),
.A2(n_934),
.B(n_911),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1129),
.A2(n_931),
.B(n_1036),
.Y(n_1273)
);

NOR2xp67_ASAP7_75t_L g1274 ( 
.A(n_1116),
.B(n_993),
.Y(n_1274)
);

NOR4xp25_ASAP7_75t_L g1275 ( 
.A(n_1236),
.B(n_968),
.C(n_1065),
.D(n_1067),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1196),
.B(n_1012),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1260),
.A2(n_909),
.B(n_921),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1108),
.Y(n_1278)
);

AOI31xp67_ASAP7_75t_L g1279 ( 
.A1(n_1227),
.A2(n_1056),
.A3(n_1054),
.B(n_1058),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1256),
.B(n_1003),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1103),
.A2(n_977),
.B(n_979),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1163),
.Y(n_1282)
);

AOI221xp5_ASAP7_75t_SL g1283 ( 
.A1(n_1253),
.A2(n_1090),
.B1(n_1083),
.B2(n_1082),
.C(n_1098),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1212),
.A2(n_1057),
.B(n_1036),
.C(n_1047),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1148),
.A2(n_1047),
.B(n_1064),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1262),
.B(n_971),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1131),
.A2(n_932),
.B(n_921),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1148),
.A2(n_1006),
.A3(n_1068),
.B(n_1026),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1124),
.A2(n_946),
.B(n_955),
.Y(n_1289)
);

OR2x2_ASAP7_75t_L g1290 ( 
.A(n_1114),
.B(n_1125),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1099),
.A2(n_963),
.B(n_1013),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1102),
.A2(n_926),
.B(n_980),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1239),
.A2(n_1028),
.B(n_967),
.Y(n_1293)
);

AO21x2_ASAP7_75t_L g1294 ( 
.A1(n_1208),
.A2(n_959),
.B(n_958),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1194),
.B(n_1052),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1250),
.A2(n_982),
.B(n_1032),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1174),
.A2(n_1033),
.B(n_550),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1100),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1149),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1250),
.A2(n_191),
.B(n_189),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1186),
.A2(n_1199),
.B(n_1152),
.C(n_1158),
.Y(n_1301)
);

INVx1_ASAP7_75t_SL g1302 ( 
.A(n_1114),
.Y(n_1302)
);

AO21x1_ASAP7_75t_L g1303 ( 
.A1(n_1226),
.A2(n_44),
.B(n_45),
.Y(n_1303)
);

BUFx6f_ASAP7_75t_L g1304 ( 
.A(n_1163),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1180),
.B(n_45),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1146),
.A2(n_47),
.B(n_48),
.C(n_49),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1221),
.A2(n_49),
.B(n_50),
.C(n_52),
.Y(n_1307)
);

OAI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1258),
.A2(n_101),
.B(n_170),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1191),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1233),
.A2(n_50),
.B(n_55),
.C(n_56),
.Y(n_1310)
);

NOR2xp33_ASAP7_75t_L g1311 ( 
.A(n_1215),
.B(n_55),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1233),
.A2(n_57),
.B(n_59),
.C(n_61),
.Y(n_1312)
);

AO21x1_ASAP7_75t_L g1313 ( 
.A1(n_1223),
.A2(n_63),
.B(n_65),
.Y(n_1313)
);

O2A1O1Ixp33_ASAP7_75t_SL g1314 ( 
.A1(n_1222),
.A2(n_115),
.B(n_159),
.C(n_147),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1147),
.A2(n_107),
.B(n_140),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1107),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1200),
.A2(n_66),
.B(n_69),
.C(n_71),
.Y(n_1317)
);

INVxp67_ASAP7_75t_SL g1318 ( 
.A(n_1101),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1187),
.A2(n_66),
.B(n_69),
.C(n_73),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1217),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_SL g1321 ( 
.A1(n_1128),
.A2(n_116),
.B(n_136),
.C(n_131),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1231),
.A2(n_102),
.B(n_128),
.Y(n_1322)
);

BUFx2_ASAP7_75t_L g1323 ( 
.A(n_1170),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1120),
.A2(n_73),
.B(n_74),
.C(n_75),
.Y(n_1324)
);

OR2x2_ASAP7_75t_L g1325 ( 
.A(n_1106),
.B(n_86),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1107),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1257),
.A2(n_109),
.B1(n_126),
.B2(n_172),
.Y(n_1327)
);

NOR2xp67_ASAP7_75t_L g1328 ( 
.A(n_1133),
.B(n_1164),
.Y(n_1328)
);

INVxp67_ASAP7_75t_SL g1329 ( 
.A(n_1112),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1150),
.A2(n_1109),
.B(n_1115),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1161),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1134),
.A2(n_1235),
.B(n_1213),
.Y(n_1332)
);

BUFx2_ASAP7_75t_R g1333 ( 
.A(n_1160),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1139),
.B(n_1190),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_1165),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1155),
.A2(n_1241),
.B1(n_1130),
.B2(n_1123),
.Y(n_1336)
);

O2A1O1Ixp33_ASAP7_75t_SL g1337 ( 
.A1(n_1126),
.A2(n_1175),
.B(n_1173),
.C(n_1162),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1224),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1121),
.A2(n_1169),
.B1(n_1172),
.B2(n_1185),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1120),
.B(n_1167),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1242),
.Y(n_1341)
);

AO31x2_ASAP7_75t_L g1342 ( 
.A1(n_1261),
.A2(n_1255),
.A3(n_1203),
.B(n_1209),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1251),
.A2(n_1208),
.B(n_1179),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1183),
.A2(n_1210),
.B(n_1198),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1203),
.A2(n_1206),
.A3(n_1229),
.B(n_1178),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1228),
.A2(n_1156),
.B(n_1153),
.Y(n_1346)
);

A2O1A1Ixp33_ASAP7_75t_L g1347 ( 
.A1(n_1113),
.A2(n_1246),
.B(n_1232),
.C(n_1254),
.Y(n_1347)
);

NAND2x1_ASAP7_75t_L g1348 ( 
.A(n_1131),
.B(n_1153),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1249),
.Y(n_1349)
);

AO32x2_ASAP7_75t_L g1350 ( 
.A1(n_1220),
.A2(n_1203),
.A3(n_1229),
.B1(n_1136),
.B2(n_1142),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1245),
.A2(n_1252),
.B1(n_1189),
.B2(n_1195),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1238),
.B(n_1197),
.Y(n_1352)
);

AO31x2_ASAP7_75t_L g1353 ( 
.A1(n_1181),
.A2(n_1193),
.A3(n_1201),
.B(n_1243),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1182),
.A2(n_1202),
.B(n_1117),
.Y(n_1354)
);

AOI221xp5_ASAP7_75t_L g1355 ( 
.A1(n_1220),
.A2(n_1159),
.B1(n_1184),
.B2(n_1218),
.C(n_1247),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1192),
.A2(n_1248),
.B(n_1240),
.Y(n_1356)
);

BUFx8_ASAP7_75t_L g1357 ( 
.A(n_1163),
.Y(n_1357)
);

HB1xp67_ASAP7_75t_L g1358 ( 
.A(n_1189),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1237),
.A2(n_1216),
.B(n_1214),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1107),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1182),
.A2(n_1119),
.B(n_1244),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1137),
.A2(n_1145),
.B(n_1132),
.Y(n_1362)
);

AO31x2_ASAP7_75t_L g1363 ( 
.A1(n_1111),
.A2(n_1177),
.A3(n_1151),
.B(n_1195),
.Y(n_1363)
);

NOR2xp33_ASAP7_75t_SL g1364 ( 
.A(n_1171),
.B(n_1188),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1244),
.A2(n_1143),
.B(n_1138),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1189),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1138),
.A2(n_1143),
.B(n_1207),
.Y(n_1367)
);

INVx1_ASAP7_75t_SL g1368 ( 
.A(n_1132),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1144),
.A2(n_1259),
.B(n_1104),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1135),
.B(n_1140),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1157),
.A2(n_1168),
.B(n_1171),
.C(n_1205),
.Y(n_1371)
);

INVx1_ASAP7_75t_SL g1372 ( 
.A(n_1185),
.Y(n_1372)
);

NOR2xp33_ASAP7_75t_SL g1373 ( 
.A(n_1171),
.B(n_1154),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1135),
.B(n_1140),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1195),
.A2(n_1205),
.B1(n_1234),
.B2(n_1259),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_SL g1376 ( 
.A1(n_1234),
.A2(n_1205),
.B(n_1230),
.C(n_1259),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1211),
.Y(n_1377)
);

O2A1O1Ixp33_ASAP7_75t_L g1378 ( 
.A1(n_1234),
.A2(n_1211),
.B(n_1219),
.C(n_1135),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1140),
.Y(n_1379)
);

AOI21xp5_ASAP7_75t_L g1380 ( 
.A1(n_1219),
.A2(n_589),
.B(n_940),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1219),
.A2(n_935),
.B(n_1204),
.Y(n_1381)
);

OAI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1141),
.A2(n_615),
.B1(n_953),
.B2(n_570),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1099),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1141),
.B(n_783),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1204),
.A2(n_1225),
.A3(n_1253),
.B(n_935),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1099),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1141),
.A2(n_941),
.B(n_783),
.C(n_594),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1118),
.Y(n_1390)
);

BUFx2_ASAP7_75t_L g1391 ( 
.A(n_1108),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1110),
.A2(n_1122),
.B(n_1099),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1204),
.A2(n_1225),
.A3(n_1253),
.B(n_935),
.Y(n_1393)
);

AO31x2_ASAP7_75t_L g1394 ( 
.A1(n_1204),
.A2(n_1225),
.A3(n_1253),
.B(n_935),
.Y(n_1394)
);

OA21x2_ASAP7_75t_L g1395 ( 
.A1(n_1208),
.A2(n_935),
.B(n_1122),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1099),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1398)
);

BUFx2_ASAP7_75t_L g1399 ( 
.A(n_1108),
.Y(n_1399)
);

AOI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1110),
.A2(n_1122),
.B(n_1099),
.Y(n_1400)
);

BUFx3_ASAP7_75t_L g1401 ( 
.A(n_1108),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1141),
.A2(n_783),
.B(n_1194),
.C(n_746),
.Y(n_1402)
);

BUFx2_ASAP7_75t_SL g1403 ( 
.A(n_1108),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1204),
.A2(n_935),
.B(n_754),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_1152),
.B(n_832),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1118),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_L g1408 ( 
.A1(n_1204),
.A2(n_935),
.B(n_754),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1256),
.B(n_745),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1208),
.A2(n_935),
.B(n_1122),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1412)
);

OAI21xp5_ASAP7_75t_SL g1413 ( 
.A1(n_1141),
.A2(n_559),
.B(n_799),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1099),
.Y(n_1414)
);

AOI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1110),
.A2(n_1122),
.B(n_1099),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1122),
.A2(n_589),
.B(n_940),
.Y(n_1417)
);

NAND2xp33_ASAP7_75t_L g1418 ( 
.A(n_1163),
.B(n_1004),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_L g1419 ( 
.A(n_1116),
.B(n_793),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1256),
.B(n_745),
.Y(n_1420)
);

AO31x2_ASAP7_75t_L g1421 ( 
.A1(n_1204),
.A2(n_1225),
.A3(n_1253),
.B(n_935),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1099),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1204),
.A2(n_935),
.B(n_754),
.Y(n_1423)
);

O2A1O1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1141),
.A2(n_941),
.B(n_783),
.C(n_594),
.Y(n_1424)
);

O2A1O1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1141),
.A2(n_941),
.B(n_783),
.C(n_594),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1160),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1099),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1118),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1166),
.A2(n_1103),
.B(n_1099),
.Y(n_1429)
);

NAND2x1_ASAP7_75t_SL g1430 ( 
.A(n_1152),
.B(n_1009),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1108),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1384),
.A2(n_1382),
.B1(n_1336),
.B2(n_1355),
.Y(n_1432)
);

NAND2xp33_ASAP7_75t_SL g1433 ( 
.A(n_1430),
.B(n_1304),
.Y(n_1433)
);

INVx6_ASAP7_75t_L g1434 ( 
.A(n_1357),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1401),
.Y(n_1435)
);

AOI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1311),
.A2(n_1405),
.B1(n_1334),
.B2(n_1327),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1428),
.Y(n_1437)
);

OAI21xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1413),
.A2(n_1424),
.B(n_1389),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1320),
.Y(n_1439)
);

OAI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1340),
.A2(n_1299),
.B1(n_1351),
.B2(n_1423),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1402),
.A2(n_1425),
.B1(n_1276),
.B2(n_1339),
.Y(n_1441)
);

BUFx4f_ASAP7_75t_SL g1442 ( 
.A(n_1357),
.Y(n_1442)
);

INVx6_ASAP7_75t_L g1443 ( 
.A(n_1282),
.Y(n_1443)
);

AOI22xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1403),
.A2(n_1302),
.B1(n_1351),
.B2(n_1366),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1265),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1302),
.A2(n_1358),
.B1(n_1309),
.B2(n_1335),
.Y(n_1446)
);

BUFx6f_ASAP7_75t_SL g1447 ( 
.A(n_1431),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1404),
.A2(n_1408),
.B1(n_1423),
.B2(n_1303),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1269),
.Y(n_1449)
);

BUFx10_ASAP7_75t_L g1450 ( 
.A(n_1304),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1290),
.B(n_1278),
.Y(n_1451)
);

OAI21xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1301),
.A2(n_1324),
.B(n_1317),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1390),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1407),
.Y(n_1454)
);

OAI21xp33_ASAP7_75t_L g1455 ( 
.A1(n_1306),
.A2(n_1319),
.B(n_1347),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1404),
.A2(n_1408),
.B1(n_1313),
.B2(n_1381),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1426),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1391),
.Y(n_1458)
);

INVx6_ASAP7_75t_L g1459 ( 
.A(n_1282),
.Y(n_1459)
);

INVx6_ASAP7_75t_L g1460 ( 
.A(n_1360),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1373),
.A2(n_1364),
.B1(n_1305),
.B2(n_1368),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1331),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1338),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1399),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1335),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1341),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1323),
.B(n_1368),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1349),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_SL g1469 ( 
.A1(n_1318),
.A2(n_1329),
.B1(n_1372),
.B2(n_1375),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1352),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1352),
.Y(n_1471)
);

INVx8_ASAP7_75t_L g1472 ( 
.A(n_1418),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1373),
.A2(n_1364),
.B1(n_1305),
.B2(n_1420),
.Y(n_1473)
);

BUFx6f_ASAP7_75t_L g1474 ( 
.A(n_1379),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1286),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1381),
.A2(n_1395),
.B1(n_1411),
.B2(n_1409),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1395),
.A2(n_1411),
.B1(n_1409),
.B2(n_1420),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1298),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1271),
.A2(n_1328),
.B1(n_1325),
.B2(n_1295),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1286),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1385),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_SL g1482 ( 
.A1(n_1375),
.A2(n_1385),
.B1(n_1421),
.B2(n_1394),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1377),
.Y(n_1483)
);

OAI22x1_ASAP7_75t_L g1484 ( 
.A1(n_1267),
.A2(n_1372),
.B1(n_1295),
.B2(n_1400),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1274),
.A2(n_1362),
.B1(n_1315),
.B2(n_1419),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1280),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1310),
.B(n_1312),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1371),
.A2(n_1337),
.B1(n_1376),
.B2(n_1326),
.Y(n_1488)
);

INVx6_ASAP7_75t_L g1489 ( 
.A(n_1316),
.Y(n_1489)
);

BUFx8_ASAP7_75t_L g1490 ( 
.A(n_1333),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1367),
.Y(n_1491)
);

CKINVDCx11_ASAP7_75t_R g1492 ( 
.A(n_1370),
.Y(n_1492)
);

INVx1_ASAP7_75t_SL g1493 ( 
.A(n_1370),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1374),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1362),
.A2(n_1346),
.B1(n_1332),
.B2(n_1369),
.Y(n_1495)
);

INVx6_ASAP7_75t_L g1496 ( 
.A(n_1378),
.Y(n_1496)
);

INVx5_ASAP7_75t_L g1497 ( 
.A(n_1287),
.Y(n_1497)
);

BUFx12f_ASAP7_75t_L g1498 ( 
.A(n_1374),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1363),
.Y(n_1499)
);

BUFx12f_ASAP7_75t_L g1500 ( 
.A(n_1307),
.Y(n_1500)
);

BUFx4_ASAP7_75t_SL g1501 ( 
.A(n_1348),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1363),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1354),
.A2(n_1361),
.B1(n_1321),
.B2(n_1314),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1365),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1353),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1285),
.A2(n_1332),
.B1(n_1359),
.B2(n_1273),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1353),
.Y(n_1507)
);

BUFx4_ASAP7_75t_SL g1508 ( 
.A(n_1350),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1285),
.A2(n_1359),
.B1(n_1273),
.B2(n_1294),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1294),
.A2(n_1272),
.B1(n_1266),
.B2(n_1356),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1380),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1263),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1356),
.A2(n_1300),
.B1(n_1308),
.B2(n_1421),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1385),
.A2(n_1421),
.B1(n_1393),
.B2(n_1394),
.Y(n_1514)
);

BUFx8_ASAP7_75t_SL g1515 ( 
.A(n_1392),
.Y(n_1515)
);

BUFx3_ASAP7_75t_L g1516 ( 
.A(n_1322),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_SL g1517 ( 
.A1(n_1393),
.A2(n_1394),
.B1(n_1264),
.B2(n_1297),
.Y(n_1517)
);

CKINVDCx20_ASAP7_75t_R g1518 ( 
.A(n_1297),
.Y(n_1518)
);

OAI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1270),
.A2(n_1277),
.B1(n_1417),
.B2(n_1388),
.Y(n_1519)
);

INVx4_ASAP7_75t_L g1520 ( 
.A(n_1275),
.Y(n_1520)
);

OAI21xp33_ASAP7_75t_L g1521 ( 
.A1(n_1415),
.A2(n_1330),
.B(n_1386),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1396),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1398),
.A2(n_1406),
.B1(n_1416),
.B2(n_1412),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1283),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1350),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1410),
.A2(n_1344),
.B1(n_1343),
.B2(n_1296),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1284),
.A2(n_1292),
.B1(n_1289),
.B2(n_1264),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1264),
.A2(n_1350),
.B1(n_1279),
.B2(n_1283),
.Y(n_1528)
);

BUFx12f_ASAP7_75t_L g1529 ( 
.A(n_1288),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1293),
.A2(n_1291),
.B1(n_1268),
.B2(n_1281),
.Y(n_1530)
);

NAND2x1p5_ASAP7_75t_L g1531 ( 
.A(n_1383),
.B(n_1429),
.Y(n_1531)
);

BUFx4_ASAP7_75t_R g1532 ( 
.A(n_1342),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1387),
.A2(n_1427),
.B1(n_1397),
.B2(n_1414),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1422),
.A2(n_1342),
.B1(n_1345),
.B2(n_1288),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1342),
.A2(n_1384),
.B1(n_1402),
.B2(n_615),
.Y(n_1535)
);

BUFx6f_ASAP7_75t_L g1536 ( 
.A(n_1288),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1345),
.A2(n_1402),
.B(n_1016),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1384),
.A2(n_1141),
.B1(n_1241),
.B2(n_1257),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1384),
.B(n_783),
.Y(n_1539)
);

BUFx10_ASAP7_75t_L g1540 ( 
.A(n_1304),
.Y(n_1540)
);

AOI22xp33_ASAP7_75t_SL g1541 ( 
.A1(n_1384),
.A2(n_1257),
.B1(n_1141),
.B2(n_615),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1384),
.A2(n_1402),
.B1(n_615),
.B2(n_783),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1428),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1426),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1384),
.B(n_783),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1428),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1384),
.B(n_783),
.Y(n_1547)
);

BUFx6f_ASAP7_75t_SL g1548 ( 
.A(n_1401),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1428),
.Y(n_1549)
);

INVx6_ASAP7_75t_L g1550 ( 
.A(n_1357),
.Y(n_1550)
);

CKINVDCx20_ASAP7_75t_R g1551 ( 
.A(n_1426),
.Y(n_1551)
);

CKINVDCx11_ASAP7_75t_R g1552 ( 
.A(n_1426),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1428),
.Y(n_1553)
);

INVx1_ASAP7_75t_SL g1554 ( 
.A(n_1302),
.Y(n_1554)
);

OAI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1384),
.A2(n_1413),
.B1(n_1382),
.B2(n_1141),
.Y(n_1555)
);

OAI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1384),
.A2(n_1413),
.B1(n_1382),
.B2(n_1141),
.Y(n_1556)
);

CKINVDCx16_ASAP7_75t_R g1557 ( 
.A(n_1373),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1384),
.B(n_783),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1428),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1381),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1401),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_1426),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1428),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1304),
.Y(n_1564)
);

CKINVDCx11_ASAP7_75t_R g1565 ( 
.A(n_1426),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1384),
.B(n_783),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1384),
.A2(n_1257),
.B1(n_1141),
.B2(n_615),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1401),
.Y(n_1568)
);

BUFx12f_ASAP7_75t_L g1569 ( 
.A(n_1426),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1428),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1384),
.A2(n_1141),
.B1(n_1382),
.B2(n_1336),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1401),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1384),
.B(n_783),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1384),
.B(n_783),
.Y(n_1574)
);

CKINVDCx6p67_ASAP7_75t_R g1575 ( 
.A(n_1426),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_1426),
.Y(n_1576)
);

INVx6_ASAP7_75t_L g1577 ( 
.A(n_1357),
.Y(n_1577)
);

AOI22xp5_ASAP7_75t_L g1578 ( 
.A1(n_1384),
.A2(n_1413),
.B1(n_799),
.B2(n_746),
.Y(n_1578)
);

INVx5_ASAP7_75t_L g1579 ( 
.A(n_1304),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1405),
.B(n_1334),
.Y(n_1580)
);

CKINVDCx11_ASAP7_75t_R g1581 ( 
.A(n_1426),
.Y(n_1581)
);

OAI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1384),
.A2(n_1413),
.B1(n_1382),
.B2(n_1141),
.Y(n_1582)
);

CKINVDCx11_ASAP7_75t_R g1583 ( 
.A(n_1426),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1481),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1481),
.Y(n_1585)
);

AOI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1519),
.A2(n_1527),
.B(n_1441),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1554),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1534),
.A2(n_1506),
.B(n_1521),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1505),
.Y(n_1589)
);

INVx8_ASAP7_75t_L g1590 ( 
.A(n_1472),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1489),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1507),
.Y(n_1592)
);

BUFx4f_ASAP7_75t_SL g1593 ( 
.A(n_1569),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1578),
.A2(n_1571),
.B1(n_1556),
.B2(n_1555),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1499),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1502),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1449),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1560),
.B(n_1520),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1539),
.B(n_1545),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1453),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1520),
.B(n_1560),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1514),
.B(n_1524),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1445),
.Y(n_1603)
);

INVx2_ASAP7_75t_L g1604 ( 
.A(n_1462),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1489),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1463),
.Y(n_1606)
);

NAND2xp33_ASAP7_75t_L g1607 ( 
.A(n_1538),
.B(n_1432),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1468),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1454),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1514),
.B(n_1482),
.Y(n_1610)
);

AOI21x1_ASAP7_75t_L g1611 ( 
.A1(n_1535),
.A2(n_1484),
.B(n_1512),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1491),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1531),
.A2(n_1533),
.B(n_1530),
.Y(n_1613)
);

AO21x2_ASAP7_75t_L g1614 ( 
.A1(n_1537),
.A2(n_1528),
.B(n_1503),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1493),
.Y(n_1615)
);

AO31x2_ASAP7_75t_L g1616 ( 
.A1(n_1524),
.A2(n_1525),
.A3(n_1475),
.B(n_1480),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1448),
.A2(n_1510),
.B(n_1506),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1474),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_1474),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1494),
.B(n_1466),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1531),
.A2(n_1533),
.B(n_1530),
.Y(n_1621)
);

INVxp33_ASAP7_75t_L g1622 ( 
.A(n_1580),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1486),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1536),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1437),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1497),
.B(n_1546),
.Y(n_1626)
);

OR2x6_ASAP7_75t_L g1627 ( 
.A(n_1529),
.B(n_1472),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1559),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1517),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1517),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1563),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1547),
.B(n_1558),
.Y(n_1632)
);

OR2x2_ASAP7_75t_L g1633 ( 
.A(n_1509),
.B(n_1440),
.Y(n_1633)
);

BUFx6f_ASAP7_75t_L g1634 ( 
.A(n_1472),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1482),
.Y(n_1635)
);

OAI21x1_ASAP7_75t_L g1636 ( 
.A1(n_1526),
.A2(n_1523),
.B(n_1510),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1474),
.Y(n_1637)
);

OAI21x1_ASAP7_75t_L g1638 ( 
.A1(n_1526),
.A2(n_1523),
.B(n_1513),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1497),
.B(n_1570),
.Y(n_1639)
);

OAI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1513),
.A2(n_1534),
.B(n_1509),
.Y(n_1640)
);

INVx1_ASAP7_75t_SL g1641 ( 
.A(n_1451),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1448),
.B(n_1456),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1566),
.B(n_1573),
.Y(n_1643)
);

NAND2xp33_ASAP7_75t_SL g1644 ( 
.A(n_1538),
.B(n_1518),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1515),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1456),
.A2(n_1542),
.B(n_1555),
.Y(n_1646)
);

INVx11_ASAP7_75t_L g1647 ( 
.A(n_1490),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1470),
.Y(n_1648)
);

INVx2_ASAP7_75t_SL g1649 ( 
.A(n_1489),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1579),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1579),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1471),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1440),
.B(n_1476),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1532),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1477),
.B(n_1444),
.Y(n_1655)
);

NAND2x1_ASAP7_75t_L g1656 ( 
.A(n_1495),
.B(n_1485),
.Y(n_1656)
);

OA21x2_ASAP7_75t_L g1657 ( 
.A1(n_1438),
.A2(n_1452),
.B(n_1455),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1435),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1574),
.B(n_1432),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1508),
.Y(n_1660)
);

OR2x6_ASAP7_75t_L g1661 ( 
.A(n_1516),
.B(n_1496),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1543),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1549),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1553),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1488),
.A2(n_1483),
.B(n_1439),
.Y(n_1665)
);

CKINVDCx20_ASAP7_75t_R g1666 ( 
.A(n_1552),
.Y(n_1666)
);

NOR2x1_ASAP7_75t_SL g1667 ( 
.A(n_1497),
.B(n_1500),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1479),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1479),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1522),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1541),
.B(n_1567),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1469),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1496),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1541),
.B(n_1567),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1496),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1556),
.A2(n_1582),
.B(n_1473),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1504),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_SL g1678 ( 
.A(n_1562),
.B(n_1490),
.Y(n_1678)
);

HB1xp67_ASAP7_75t_L g1679 ( 
.A(n_1467),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1564),
.A2(n_1487),
.B(n_1436),
.Y(n_1680)
);

AOI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1473),
.A2(n_1458),
.B(n_1568),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1511),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1582),
.A2(n_1461),
.B1(n_1464),
.B2(n_1447),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1461),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1498),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1446),
.Y(n_1686)
);

HB1xp67_ASAP7_75t_L g1687 ( 
.A(n_1478),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1478),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1433),
.Y(n_1689)
);

BUFx2_ASAP7_75t_SL g1690 ( 
.A(n_1447),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1501),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1501),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1557),
.B(n_1564),
.Y(n_1693)
);

BUFx2_ASAP7_75t_L g1694 ( 
.A(n_1478),
.Y(n_1694)
);

INVx1_ASAP7_75t_SL g1695 ( 
.A(n_1492),
.Y(n_1695)
);

OAI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1561),
.A2(n_1572),
.B(n_1576),
.Y(n_1696)
);

CKINVDCx14_ASAP7_75t_R g1697 ( 
.A(n_1565),
.Y(n_1697)
);

OAI21x1_ASAP7_75t_SL g1698 ( 
.A1(n_1434),
.A2(n_1577),
.B(n_1550),
.Y(n_1698)
);

NAND2x1_ASAP7_75t_L g1699 ( 
.A(n_1443),
.B(n_1459),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_1443),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1450),
.B(n_1540),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1460),
.A2(n_1434),
.B(n_1577),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1459),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1434),
.B(n_1550),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1610),
.B(n_1629),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1702),
.B(n_1457),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1679),
.B(n_1465),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1601),
.B(n_1575),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1598),
.B(n_1550),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1598),
.B(n_1577),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1693),
.B(n_1460),
.Y(n_1711)
);

AO32x2_ASAP7_75t_L g1712 ( 
.A1(n_1616),
.A2(n_1548),
.A3(n_1460),
.B1(n_1442),
.B2(n_1581),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1607),
.A2(n_1548),
.B1(n_1544),
.B2(n_1551),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1693),
.B(n_1583),
.Y(n_1714)
);

AOI21xp5_ASAP7_75t_L g1715 ( 
.A1(n_1656),
.A2(n_1442),
.B(n_1646),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1641),
.B(n_1615),
.Y(n_1716)
);

OA21x2_ASAP7_75t_L g1717 ( 
.A1(n_1638),
.A2(n_1636),
.B(n_1640),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1587),
.B(n_1599),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1610),
.B(n_1629),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1609),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1657),
.B(n_1594),
.Y(n_1721)
);

AOI22xp5_ASAP7_75t_L g1722 ( 
.A1(n_1644),
.A2(n_1671),
.B1(n_1674),
.B2(n_1657),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1616),
.Y(n_1723)
);

OAI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1673),
.A2(n_1675),
.B1(n_1683),
.B2(n_1659),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1622),
.B(n_1670),
.Y(n_1725)
);

CKINVDCx20_ASAP7_75t_R g1726 ( 
.A(n_1666),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1657),
.B(n_1677),
.Y(n_1727)
);

AND2x4_ASAP7_75t_L g1728 ( 
.A(n_1702),
.B(n_1626),
.Y(n_1728)
);

CKINVDCx16_ASAP7_75t_R g1729 ( 
.A(n_1697),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1620),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_SL g1731 ( 
.A1(n_1645),
.A2(n_1657),
.B1(n_1676),
.B2(n_1682),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1626),
.B(n_1639),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1620),
.B(n_1655),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1671),
.A2(n_1674),
.B1(n_1617),
.B2(n_1642),
.C(n_1668),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1632),
.B(n_1643),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1655),
.B(n_1660),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_SL g1737 ( 
.A(n_1691),
.B(n_1692),
.C(n_1696),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1684),
.B(n_1625),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1677),
.A2(n_1682),
.B1(n_1656),
.B2(n_1684),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1586),
.A2(n_1669),
.B(n_1668),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1602),
.B(n_1654),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1642),
.A2(n_1633),
.B(n_1669),
.C(n_1653),
.Y(n_1742)
);

AOI22xp33_ASAP7_75t_L g1743 ( 
.A1(n_1633),
.A2(n_1653),
.B1(n_1686),
.B2(n_1645),
.Y(n_1743)
);

OR2x2_ASAP7_75t_L g1744 ( 
.A(n_1603),
.B(n_1630),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1677),
.B(n_1672),
.Y(n_1745)
);

OAI21xp5_ASAP7_75t_L g1746 ( 
.A1(n_1586),
.A2(n_1681),
.B(n_1680),
.Y(n_1746)
);

AOI22xp33_ASAP7_75t_L g1747 ( 
.A1(n_1635),
.A2(n_1630),
.B1(n_1680),
.B2(n_1690),
.Y(n_1747)
);

AOI21xp5_ASAP7_75t_L g1748 ( 
.A1(n_1614),
.A2(n_1667),
.B(n_1661),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1700),
.Y(n_1749)
);

NOR2x1_ASAP7_75t_SL g1750 ( 
.A(n_1661),
.B(n_1627),
.Y(n_1750)
);

OR2x6_ASAP7_75t_L g1751 ( 
.A(n_1661),
.B(n_1627),
.Y(n_1751)
);

NAND2x1_ASAP7_75t_L g1752 ( 
.A(n_1661),
.B(n_1627),
.Y(n_1752)
);

AO32x2_ASAP7_75t_L g1753 ( 
.A1(n_1616),
.A2(n_1651),
.A3(n_1650),
.B1(n_1649),
.B2(n_1605),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1625),
.B(n_1628),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1691),
.A2(n_1692),
.B1(n_1689),
.B2(n_1688),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1678),
.A2(n_1689),
.B1(n_1690),
.B2(n_1704),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1635),
.A2(n_1640),
.B(n_1636),
.C(n_1638),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1616),
.B(n_1631),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_L g1759 ( 
.A(n_1648),
.B(n_1652),
.Y(n_1759)
);

O2A1O1Ixp33_ASAP7_75t_SL g1760 ( 
.A1(n_1699),
.A2(n_1649),
.B(n_1605),
.C(n_1591),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1665),
.A2(n_1699),
.B(n_1590),
.C(n_1623),
.Y(n_1761)
);

OA21x2_ASAP7_75t_L g1762 ( 
.A1(n_1613),
.A2(n_1621),
.B(n_1611),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1687),
.B(n_1667),
.Y(n_1763)
);

AO32x2_ASAP7_75t_L g1764 ( 
.A1(n_1650),
.A2(n_1651),
.A3(n_1591),
.B1(n_1584),
.B2(n_1585),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1597),
.B(n_1608),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1662),
.A2(n_1664),
.B1(n_1663),
.B2(n_1614),
.C(n_1584),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1588),
.B(n_1604),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1767),
.B(n_1588),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1721),
.A2(n_1614),
.B1(n_1588),
.B2(n_1695),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1767),
.Y(n_1770)
);

NOR2x1_ASAP7_75t_SL g1771 ( 
.A(n_1751),
.B(n_1758),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1723),
.Y(n_1772)
);

AND2x6_ASAP7_75t_L g1773 ( 
.A(n_1732),
.B(n_1624),
.Y(n_1773)
);

NOR2xp67_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1606),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1705),
.B(n_1589),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1720),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1717),
.B(n_1589),
.Y(n_1777)
);

INVx3_ASAP7_75t_L g1778 ( 
.A(n_1728),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1705),
.B(n_1592),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1728),
.B(n_1621),
.Y(n_1780)
);

INVx4_ASAP7_75t_L g1781 ( 
.A(n_1751),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1757),
.B(n_1595),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1720),
.Y(n_1783)
);

AND2x2_ASAP7_75t_SL g1784 ( 
.A(n_1721),
.B(n_1585),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1757),
.B(n_1613),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1762),
.B(n_1764),
.Y(n_1786)
);

BUFx2_ASAP7_75t_L g1787 ( 
.A(n_1753),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1764),
.B(n_1596),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1731),
.A2(n_1704),
.B1(n_1685),
.B2(n_1593),
.Y(n_1789)
);

INVxp67_ASAP7_75t_L g1790 ( 
.A(n_1727),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_L g1791 ( 
.A(n_1751),
.B(n_1600),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1734),
.A2(n_1698),
.B1(n_1662),
.B2(n_1658),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1764),
.Y(n_1793)
);

INVx1_ASAP7_75t_SL g1794 ( 
.A(n_1745),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1764),
.B(n_1611),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1715),
.B(n_1694),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1765),
.Y(n_1797)
);

HB1xp67_ASAP7_75t_L g1798 ( 
.A(n_1759),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1754),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1722),
.A2(n_1698),
.B1(n_1658),
.B2(n_1606),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1727),
.B(n_1612),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1783),
.Y(n_1802)
);

INVx4_ASAP7_75t_L g1803 ( 
.A(n_1781),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1788),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1770),
.B(n_1719),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1783),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1768),
.B(n_1719),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1783),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1792),
.A2(n_1724),
.B1(n_1739),
.B2(n_1742),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1769),
.A2(n_1742),
.B1(n_1743),
.B2(n_1735),
.C(n_1718),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1790),
.B(n_1741),
.Y(n_1811)
);

HB1xp67_ASAP7_75t_L g1812 ( 
.A(n_1788),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1796),
.B(n_1708),
.Y(n_1813)
);

AOI21xp33_ASAP7_75t_SL g1814 ( 
.A1(n_1784),
.A2(n_1729),
.B(n_1713),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1798),
.B(n_1766),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1768),
.B(n_1733),
.Y(n_1816)
);

AOI31xp33_ASAP7_75t_L g1817 ( 
.A1(n_1769),
.A2(n_1743),
.A3(n_1706),
.B(n_1756),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1776),
.Y(n_1818)
);

INVx2_ASAP7_75t_L g1819 ( 
.A(n_1777),
.Y(n_1819)
);

OAI33xp33_ASAP7_75t_L g1820 ( 
.A1(n_1793),
.A2(n_1755),
.A3(n_1716),
.B1(n_1744),
.B2(n_1738),
.B3(n_1707),
.Y(n_1820)
);

INVx1_ASAP7_75t_SL g1821 ( 
.A(n_1798),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1789),
.A2(n_1737),
.B1(n_1747),
.B2(n_1746),
.C(n_1740),
.Y(n_1822)
);

OAI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1781),
.A2(n_1752),
.B1(n_1706),
.B2(n_1730),
.Y(n_1823)
);

OAI21xp33_ASAP7_75t_L g1824 ( 
.A1(n_1784),
.A2(n_1737),
.B(n_1747),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1768),
.B(n_1712),
.Y(n_1825)
);

OAI221xp5_ASAP7_75t_L g1826 ( 
.A1(n_1789),
.A2(n_1792),
.B1(n_1800),
.B2(n_1796),
.C(n_1761),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1787),
.B(n_1712),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1780),
.B(n_1750),
.Y(n_1828)
);

BUFx3_ASAP7_75t_L g1829 ( 
.A(n_1773),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1788),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1787),
.B(n_1712),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1787),
.B(n_1712),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1790),
.B(n_1799),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1780),
.B(n_1732),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1778),
.Y(n_1835)
);

INVx1_ASAP7_75t_SL g1836 ( 
.A(n_1794),
.Y(n_1836)
);

NAND2x1p5_ASAP7_75t_SL g1837 ( 
.A(n_1785),
.B(n_1791),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1786),
.B(n_1753),
.Y(n_1838)
);

OR2x2_ASAP7_75t_L g1839 ( 
.A(n_1797),
.B(n_1736),
.Y(n_1839)
);

NOR3xp33_ASAP7_75t_L g1840 ( 
.A(n_1785),
.B(n_1714),
.C(n_1703),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1786),
.B(n_1753),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1772),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1786),
.B(n_1753),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1802),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1815),
.B(n_1793),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1802),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1834),
.B(n_1778),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1821),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1834),
.B(n_1778),
.Y(n_1849)
);

OR2x2_ASAP7_75t_L g1850 ( 
.A(n_1815),
.B(n_1775),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1829),
.B(n_1771),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1833),
.B(n_1799),
.Y(n_1852)
);

OR2x2_ASAP7_75t_L g1853 ( 
.A(n_1821),
.B(n_1775),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1833),
.B(n_1801),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1806),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_SL g1856 ( 
.A(n_1814),
.B(n_1784),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1834),
.B(n_1807),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1806),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1810),
.B(n_1801),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1834),
.B(n_1807),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1810),
.B(n_1801),
.Y(n_1861)
);

AND2x2_ASAP7_75t_L g1862 ( 
.A(n_1834),
.B(n_1771),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1824),
.A2(n_1784),
.B1(n_1781),
.B2(n_1800),
.Y(n_1863)
);

NAND2xp67_ASAP7_75t_L g1864 ( 
.A(n_1827),
.B(n_1711),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1807),
.B(n_1771),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1811),
.B(n_1779),
.Y(n_1866)
);

NAND2x1_ASAP7_75t_L g1867 ( 
.A(n_1828),
.B(n_1791),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1819),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1808),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1811),
.B(n_1779),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1808),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1839),
.B(n_1797),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1842),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1813),
.B(n_1794),
.Y(n_1874)
);

NOR2xp33_ASAP7_75t_SL g1875 ( 
.A(n_1824),
.B(n_1781),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1842),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1818),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1819),
.Y(n_1878)
);

BUFx2_ASAP7_75t_L g1879 ( 
.A(n_1829),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1840),
.B(n_1797),
.Y(n_1880)
);

NAND3xp33_ASAP7_75t_L g1881 ( 
.A(n_1809),
.B(n_1795),
.C(n_1782),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1819),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1840),
.B(n_1782),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1803),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1818),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1844),
.Y(n_1886)
);

OAI211xp5_ASAP7_75t_L g1887 ( 
.A1(n_1881),
.A2(n_1814),
.B(n_1809),
.C(n_1822),
.Y(n_1887)
);

OAI21xp5_ASAP7_75t_L g1888 ( 
.A1(n_1881),
.A2(n_1817),
.B(n_1822),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1857),
.B(n_1816),
.Y(n_1889)
);

AND2x4_ASAP7_75t_L g1890 ( 
.A(n_1851),
.B(n_1829),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1850),
.B(n_1836),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1859),
.B(n_1820),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1844),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1846),
.Y(n_1894)
);

NAND3xp33_ASAP7_75t_SL g1895 ( 
.A(n_1875),
.B(n_1826),
.C(n_1726),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1857),
.B(n_1827),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1860),
.B(n_1827),
.Y(n_1897)
);

OAI21xp33_ASAP7_75t_L g1898 ( 
.A1(n_1875),
.A2(n_1861),
.B(n_1817),
.Y(n_1898)
);

AND2x4_ASAP7_75t_L g1899 ( 
.A(n_1851),
.B(n_1828),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1850),
.B(n_1805),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1868),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1846),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1860),
.B(n_1805),
.Y(n_1903)
);

O2A1O1Ixp5_ASAP7_75t_SL g1904 ( 
.A1(n_1856),
.A2(n_1835),
.B(n_1830),
.C(n_1804),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1866),
.B(n_1836),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1868),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1852),
.B(n_1805),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1855),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1855),
.Y(n_1909)
);

NOR2xp67_ASAP7_75t_L g1910 ( 
.A(n_1848),
.B(n_1803),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1858),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1858),
.Y(n_1912)
);

NAND2x1p5_ASAP7_75t_L g1913 ( 
.A(n_1867),
.B(n_1803),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1869),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1883),
.B(n_1825),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1870),
.B(n_1854),
.Y(n_1916)
);

HB1xp67_ASAP7_75t_L g1917 ( 
.A(n_1869),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1871),
.Y(n_1918)
);

OAI33xp33_ASAP7_75t_L g1919 ( 
.A1(n_1845),
.A2(n_1873),
.A3(n_1876),
.B1(n_1871),
.B2(n_1880),
.B3(n_1853),
.Y(n_1919)
);

OR2x2_ASAP7_75t_L g1920 ( 
.A(n_1872),
.B(n_1837),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1874),
.B(n_1825),
.Y(n_1921)
);

OAI211xp5_ASAP7_75t_L g1922 ( 
.A1(n_1863),
.A2(n_1826),
.B(n_1831),
.C(n_1832),
.Y(n_1922)
);

NOR2x1_ASAP7_75t_L g1923 ( 
.A(n_1867),
.B(n_1726),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1873),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1876),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1877),
.Y(n_1926)
);

AND2x4_ASAP7_75t_L g1927 ( 
.A(n_1851),
.B(n_1828),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1877),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1885),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1885),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_L g1931 ( 
.A(n_1884),
.B(n_1820),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1892),
.B(n_1845),
.Y(n_1932)
);

INVxp67_ASAP7_75t_L g1933 ( 
.A(n_1931),
.Y(n_1933)
);

AOI21xp33_ASAP7_75t_L g1934 ( 
.A1(n_1888),
.A2(n_1832),
.B(n_1831),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1892),
.B(n_1838),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1923),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1931),
.B(n_1838),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1887),
.B(n_1864),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1922),
.B(n_1838),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1898),
.B(n_1647),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1901),
.Y(n_1941)
);

NAND2xp33_ASAP7_75t_L g1942 ( 
.A(n_1913),
.B(n_1891),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1896),
.B(n_1862),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1896),
.B(n_1862),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1924),
.B(n_1841),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1897),
.B(n_1865),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1901),
.Y(n_1947)
);

OA21x2_ASAP7_75t_L g1948 ( 
.A1(n_1906),
.A2(n_1878),
.B(n_1868),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1917),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1900),
.B(n_1878),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1897),
.B(n_1865),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1913),
.B(n_1879),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1917),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1925),
.B(n_1841),
.Y(n_1954)
);

INVx4_ASAP7_75t_L g1955 ( 
.A(n_1890),
.Y(n_1955)
);

NAND3xp33_ASAP7_75t_L g1956 ( 
.A(n_1904),
.B(n_1832),
.C(n_1831),
.Y(n_1956)
);

AND2x2_ASAP7_75t_SL g1957 ( 
.A(n_1895),
.B(n_1706),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1910),
.B(n_1823),
.Y(n_1958)
);

INVx3_ASAP7_75t_L g1959 ( 
.A(n_1890),
.Y(n_1959)
);

AND3x2_ASAP7_75t_L g1960 ( 
.A(n_1895),
.B(n_1879),
.C(n_1647),
.Y(n_1960)
);

INVx2_ASAP7_75t_SL g1961 ( 
.A(n_1890),
.Y(n_1961)
);

NAND4xp75_ASAP7_75t_L g1962 ( 
.A(n_1919),
.B(n_1785),
.C(n_1841),
.D(n_1843),
.Y(n_1962)
);

INVx2_ASAP7_75t_L g1963 ( 
.A(n_1906),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1899),
.B(n_1851),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1899),
.B(n_1843),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1915),
.B(n_1878),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1899),
.B(n_1843),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1927),
.B(n_1847),
.Y(n_1968)
);

NAND3xp33_ASAP7_75t_L g1969 ( 
.A(n_1933),
.B(n_1920),
.C(n_1893),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1937),
.B(n_1916),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1957),
.B(n_1936),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1933),
.A2(n_1919),
.B1(n_1921),
.B2(n_1886),
.C(n_1909),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1938),
.A2(n_1905),
.B(n_1902),
.Y(n_1973)
);

AOI32xp33_ASAP7_75t_L g1974 ( 
.A1(n_1938),
.A2(n_1927),
.A3(n_1825),
.B1(n_1823),
.B2(n_1889),
.Y(n_1974)
);

AOI211x1_ASAP7_75t_SL g1975 ( 
.A1(n_1934),
.A2(n_1774),
.B(n_1907),
.C(n_1882),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1949),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1957),
.B(n_1927),
.Y(n_1977)
);

INVxp67_ASAP7_75t_L g1978 ( 
.A(n_1949),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1957),
.A2(n_1934),
.B1(n_1936),
.B2(n_1939),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1962),
.A2(n_1828),
.B1(n_1803),
.B2(n_1812),
.Y(n_1980)
);

NAND2xp5_ASAP7_75t_L g1981 ( 
.A(n_1932),
.B(n_1935),
.Y(n_1981)
);

AND2x2_ASAP7_75t_SL g1982 ( 
.A(n_1942),
.B(n_1781),
.Y(n_1982)
);

AOI31xp33_ASAP7_75t_L g1983 ( 
.A1(n_1940),
.A2(n_1709),
.A3(n_1710),
.B(n_1760),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1953),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1955),
.B(n_1959),
.Y(n_1985)
);

NAND4xp25_ASAP7_75t_L g1986 ( 
.A(n_1932),
.B(n_1763),
.C(n_1774),
.D(n_1911),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1962),
.A2(n_1828),
.B1(n_1912),
.B2(n_1918),
.Y(n_1987)
);

AOI221xp5_ASAP7_75t_L g1988 ( 
.A1(n_1937),
.A2(n_1894),
.B1(n_1908),
.B2(n_1914),
.C(n_1926),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1939),
.A2(n_1812),
.B1(n_1804),
.B2(n_1830),
.Y(n_1989)
);

HB1xp67_ASAP7_75t_L g1990 ( 
.A(n_1953),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1941),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1935),
.B(n_1961),
.Y(n_1992)
);

AOI21xp33_ASAP7_75t_L g1993 ( 
.A1(n_1961),
.A2(n_1928),
.B(n_1929),
.Y(n_1993)
);

NAND3xp33_ASAP7_75t_L g1994 ( 
.A(n_1956),
.B(n_1930),
.C(n_1763),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1961),
.B(n_1959),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1973),
.B(n_1959),
.Y(n_1996)
);

OAI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1979),
.A2(n_1956),
.B1(n_1958),
.B2(n_1955),
.Y(n_1997)
);

INVxp67_ASAP7_75t_L g1998 ( 
.A(n_1990),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1982),
.B(n_1955),
.Y(n_1999)
);

OAI21xp33_ASAP7_75t_L g2000 ( 
.A1(n_1971),
.A2(n_1952),
.B(n_1959),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1981),
.B(n_1955),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1987),
.A2(n_1955),
.B1(n_1959),
.B2(n_1952),
.Y(n_2002)
);

AOI22xp5_ASAP7_75t_L g2003 ( 
.A1(n_1977),
.A2(n_1960),
.B1(n_1952),
.B2(n_1964),
.Y(n_2003)
);

HB1xp67_ASAP7_75t_L g2004 ( 
.A(n_1990),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1991),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1976),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1982),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1985),
.B(n_1995),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1984),
.Y(n_2009)
);

AOI21xp33_ASAP7_75t_SL g2010 ( 
.A1(n_1969),
.A2(n_1960),
.B(n_1837),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1978),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1992),
.B(n_1968),
.Y(n_2012)
);

AOI22xp5_ASAP7_75t_L g2013 ( 
.A1(n_1980),
.A2(n_1964),
.B1(n_1968),
.B2(n_1967),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1978),
.B(n_1965),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1988),
.B(n_1965),
.Y(n_2015)
);

OAI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1994),
.A2(n_1945),
.B1(n_1954),
.B2(n_1966),
.Y(n_2016)
);

O2A1O1Ixp33_ASAP7_75t_L g2017 ( 
.A1(n_1998),
.A2(n_1993),
.B(n_1989),
.C(n_1972),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_L g2018 ( 
.A(n_2008),
.B(n_1970),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_2004),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2008),
.B(n_1974),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_2012),
.B(n_1975),
.Y(n_2021)
);

NAND3xp33_ASAP7_75t_L g2022 ( 
.A(n_1997),
.B(n_2010),
.C(n_1996),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_2004),
.Y(n_2023)
);

AOI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_2003),
.A2(n_1986),
.B1(n_1964),
.B2(n_1968),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1998),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_2014),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_2011),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_2005),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_2000),
.B(n_1983),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_1999),
.B(n_1943),
.Y(n_2030)
);

NOR3xp33_ASAP7_75t_SL g2031 ( 
.A(n_2022),
.B(n_2001),
.C(n_2002),
.Y(n_2031)
);

NOR2xp67_ASAP7_75t_L g2032 ( 
.A(n_2019),
.B(n_2006),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_2025),
.B(n_2015),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2023),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_2030),
.B(n_2009),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_2027),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_2029),
.B(n_2007),
.Y(n_2037)
);

NOR2x1_ASAP7_75t_L g2038 ( 
.A(n_2028),
.B(n_2016),
.Y(n_2038)
);

AOI211xp5_ASAP7_75t_L g2039 ( 
.A1(n_2017),
.A2(n_2016),
.B(n_2013),
.C(n_1966),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_SL g2040 ( 
.A(n_2017),
.B(n_2018),
.Y(n_2040)
);

NOR3xp33_ASAP7_75t_L g2041 ( 
.A(n_2026),
.B(n_1947),
.C(n_1941),
.Y(n_2041)
);

INVxp67_ASAP7_75t_L g2042 ( 
.A(n_2029),
.Y(n_2042)
);

O2A1O1Ixp5_ASAP7_75t_L g2043 ( 
.A1(n_2040),
.A2(n_2020),
.B(n_2021),
.C(n_1941),
.Y(n_2043)
);

CKINVDCx16_ASAP7_75t_R g2044 ( 
.A(n_2038),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2032),
.Y(n_2045)
);

OAI211xp5_ASAP7_75t_L g2046 ( 
.A1(n_2039),
.A2(n_2033),
.B(n_2031),
.C(n_2042),
.Y(n_2046)
);

AOI221xp5_ASAP7_75t_L g2047 ( 
.A1(n_2037),
.A2(n_2024),
.B1(n_1963),
.B2(n_1947),
.C(n_1954),
.Y(n_2047)
);

AOI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_2034),
.A2(n_1963),
.B1(n_1947),
.B2(n_1945),
.C(n_1943),
.Y(n_2048)
);

OAI211xp5_ASAP7_75t_SL g2049 ( 
.A1(n_2046),
.A2(n_2035),
.B(n_2036),
.C(n_2041),
.Y(n_2049)
);

NAND5xp2_ASAP7_75t_L g2050 ( 
.A(n_2047),
.B(n_1943),
.C(n_1944),
.D(n_1951),
.E(n_1946),
.Y(n_2050)
);

AOI22xp5_ASAP7_75t_L g2051 ( 
.A1(n_2044),
.A2(n_1963),
.B1(n_1967),
.B2(n_1965),
.Y(n_2051)
);

OAI21xp5_ASAP7_75t_SL g2052 ( 
.A1(n_2045),
.A2(n_1944),
.B(n_1951),
.Y(n_2052)
);

XNOR2xp5_ASAP7_75t_L g2053 ( 
.A(n_2043),
.B(n_1864),
.Y(n_2053)
);

AOI221xp5_ASAP7_75t_L g2054 ( 
.A1(n_2048),
.A2(n_1944),
.B1(n_1946),
.B2(n_1951),
.C(n_1967),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_2045),
.Y(n_2055)
);

XNOR2xp5_ASAP7_75t_L g2056 ( 
.A(n_2053),
.B(n_1694),
.Y(n_2056)
);

INVx2_ASAP7_75t_L g2057 ( 
.A(n_2055),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_2051),
.B(n_1966),
.Y(n_2058)
);

NAND4xp75_ASAP7_75t_L g2059 ( 
.A(n_2054),
.B(n_1948),
.C(n_1946),
.D(n_1701),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_2049),
.A2(n_1950),
.B1(n_1948),
.B2(n_1749),
.Y(n_2060)
);

NOR3xp33_ASAP7_75t_L g2061 ( 
.A(n_2050),
.B(n_1950),
.C(n_1725),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_SL g2062 ( 
.A(n_2060),
.B(n_1950),
.Y(n_2062)
);

OAI31xp33_ASAP7_75t_L g2063 ( 
.A1(n_2058),
.A2(n_2056),
.A3(n_2052),
.B(n_2057),
.Y(n_2063)
);

OAI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2059),
.A2(n_1853),
.B1(n_1948),
.B2(n_1882),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_2063),
.B(n_2058),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_SL g2066 ( 
.A1(n_2065),
.A2(n_2064),
.B1(n_2062),
.B2(n_2061),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2066),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2066),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_2067),
.B(n_1903),
.Y(n_2069)
);

XNOR2x1_ASAP7_75t_L g2070 ( 
.A(n_2068),
.B(n_1618),
.Y(n_2070)
);

OAI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_2069),
.A2(n_1948),
.B(n_1882),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_2070),
.Y(n_2072)
);

OAI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2072),
.A2(n_1948),
.B1(n_1618),
.B2(n_1619),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2073),
.B(n_2071),
.Y(n_2074)
);

XOR2xp5_ASAP7_75t_L g2075 ( 
.A(n_2074),
.B(n_1634),
.Y(n_2075)
);

OAI221xp5_ASAP7_75t_R g2076 ( 
.A1(n_2075),
.A2(n_1590),
.B1(n_1837),
.B2(n_1637),
.C(n_1619),
.Y(n_2076)
);

AOI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_2076),
.A2(n_1849),
.B1(n_1847),
.B2(n_1637),
.Y(n_2077)
);


endmodule