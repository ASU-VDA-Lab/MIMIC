module fake_netlist_6_3458_n_2447 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_507, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_396, n_495, n_350, n_78, n_84, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_468, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_466, n_506, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_493, n_397, n_155, n_109, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_472, n_270, n_239, n_126, n_414, n_97, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_154, n_456, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_455, n_83, n_363, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_406, n_483, n_102, n_204, n_482, n_474, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_33, n_477, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_436, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_487, n_128, n_241, n_30, n_275, n_43, n_276, n_441, n_221, n_444, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_514, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2447);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_507;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_468;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_493;
input n_397;
input n_155;
input n_109;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_154;
input n_456;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_455;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_33;
input n_477;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_441;
input n_221;
input n_444;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_514;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2447;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_539;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_2370;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_2073;
wire n_2273;
wire n_792;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_850;
wire n_690;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_2279;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_1139;
wire n_872;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_644;
wire n_682;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_1492;
wire n_987;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1966;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2025;
wire n_2357;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_2410;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_520;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_1617;
wire n_1470;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_736;
wire n_613;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_2016;
wire n_1905;
wire n_2343;
wire n_793;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_724;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_1037;
wire n_621;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2423;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_1974;
wire n_1720;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_533;
wire n_2390;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1949;
wire n_545;
wire n_1804;
wire n_1727;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_875;
wire n_680;
wire n_1678;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_2437;
wire n_839;
wire n_2444;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_1148;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_719;
wire n_1972;
wire n_1525;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1362;
wire n_1156;
wire n_984;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_583;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_1888;
wire n_1557;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2415;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_217),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_503),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_60),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_399),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_425),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_176),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_517),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_497),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_193),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_205),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_132),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_353),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_476),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_45),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_388),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_444),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_382),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_336),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_483),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_506),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_467),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_289),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_9),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_492),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_449),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_490),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_475),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_192),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_403),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_397),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_172),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_306),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_291),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_334),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_471),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_356),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_332),
.Y(n_556)
);

INVxp33_ASAP7_75t_L g557 ( 
.A(n_402),
.Y(n_557)
);

BUFx10_ASAP7_75t_L g558 ( 
.A(n_504),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_351),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_498),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_32),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_40),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_31),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_378),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_183),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_480),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_205),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_123),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_470),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_279),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_442),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_255),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_161),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_42),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_424),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_79),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_221),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_451),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_466),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_502),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_273),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_154),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_338),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_199),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_358),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_426),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_484),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_346),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_248),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_14),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_363),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_122),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_474),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_510),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_125),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_500),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_188),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_180),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_130),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_75),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_125),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_29),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_485),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_187),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_141),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_479),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_495),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_427),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_199),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_215),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_164),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_72),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_496),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_433),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_514),
.Y(n_615)
);

CKINVDCx16_ASAP7_75t_R g616 ( 
.A(n_187),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_478),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_499),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_168),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_450),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_355),
.Y(n_621)
);

BUFx8_ASAP7_75t_SL g622 ( 
.A(n_501),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_241),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_489),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_133),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_11),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_481),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_472),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_350),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_103),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_255),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_473),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_95),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_51),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_390),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_493),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_25),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_196),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_431),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_145),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_63),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_246),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_193),
.Y(n_643)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_491),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_184),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_422),
.Y(n_646)
);

BUFx5_ASAP7_75t_L g647 ( 
.A(n_505),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_12),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_171),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_488),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_90),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_153),
.Y(n_652)
);

HB1xp67_ASAP7_75t_L g653 ( 
.A(n_87),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_212),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_189),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_307),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_222),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_348),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_507),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_93),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_159),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_216),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_89),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_487),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_62),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_159),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_469),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_135),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_188),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_151),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_418),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_436),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_178),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_200),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_286),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_519),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_494),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_288),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_97),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_319),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_170),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_239),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_303),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_486),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_349),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_201),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_281),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_251),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_228),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_252),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_27),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_360),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_300),
.Y(n_693)
);

INVx1_ASAP7_75t_SL g694 ( 
.A(n_482),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_380),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_460),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_234),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_74),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_285),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_157),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_277),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_296),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_477),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_312),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_317),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_76),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_53),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_468),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_214),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_379),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_455),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_34),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_357),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_230),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_113),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_412),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_16),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_439),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_163),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_149),
.Y(n_720)
);

CKINVDCx16_ASAP7_75t_R g721 ( 
.A(n_129),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_44),
.Y(n_722)
);

BUFx2_ASAP7_75t_SL g723 ( 
.A(n_29),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_58),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_169),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_142),
.Y(n_726)
);

CKINVDCx20_ASAP7_75t_R g727 ( 
.A(n_48),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_92),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_392),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_345),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_374),
.Y(n_731)
);

BUFx10_ASAP7_75t_L g732 ( 
.A(n_268),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_1),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_56),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_96),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_18),
.Y(n_736)
);

INVx1_ASAP7_75t_SL g737 ( 
.A(n_163),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_204),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_157),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_90),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_103),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_420),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_377),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_458),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_97),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_333),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_342),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_166),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_198),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_707),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_707),
.Y(n_751)
);

INVxp33_ASAP7_75t_L g752 ( 
.A(n_525),
.Y(n_752)
);

INVxp33_ASAP7_75t_L g753 ( 
.A(n_653),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_749),
.Y(n_754)
);

INVxp33_ASAP7_75t_L g755 ( 
.A(n_577),
.Y(n_755)
);

INVxp33_ASAP7_75t_SL g756 ( 
.A(n_723),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_521),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_584),
.Y(n_758)
);

INVxp33_ASAP7_75t_L g759 ( 
.A(n_577),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_647),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_523),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_584),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_527),
.Y(n_763)
);

CKINVDCx16_ASAP7_75t_R g764 ( 
.A(n_616),
.Y(n_764)
);

INVxp67_ASAP7_75t_SL g765 ( 
.A(n_553),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_584),
.Y(n_766)
);

INVxp67_ASAP7_75t_L g767 ( 
.A(n_732),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_584),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_721),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_647),
.Y(n_771)
);

INVxp33_ASAP7_75t_L g772 ( 
.A(n_600),
.Y(n_772)
);

CKINVDCx20_ASAP7_75t_R g773 ( 
.A(n_520),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_602),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_538),
.Y(n_775)
);

BUFx10_ASAP7_75t_L g776 ( 
.A(n_624),
.Y(n_776)
);

INVxp67_ASAP7_75t_SL g777 ( 
.A(n_535),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_602),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_557),
.B(n_0),
.Y(n_779)
);

NOR2xp67_ASAP7_75t_L g780 ( 
.A(n_683),
.B(n_0),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_602),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_602),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_637),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_647),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_637),
.Y(n_785)
);

INVxp33_ASAP7_75t_L g786 ( 
.A(n_600),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_637),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_520),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_637),
.Y(n_789)
);

INVxp33_ASAP7_75t_SL g790 ( 
.A(n_529),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_663),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_663),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_663),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_530),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_663),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_522),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_528),
.Y(n_797)
);

INVxp67_ASAP7_75t_SL g798 ( 
.A(n_535),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_547),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_562),
.Y(n_800)
);

INVxp33_ASAP7_75t_SL g801 ( 
.A(n_533),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_565),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_567),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_541),
.Y(n_804)
);

INVxp67_ASAP7_75t_L g805 ( 
.A(n_732),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_572),
.Y(n_806)
);

INVxp67_ASAP7_75t_SL g807 ( 
.A(n_541),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_576),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_732),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_589),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_671),
.Y(n_811)
);

BUFx3_ASAP7_75t_L g812 ( 
.A(n_671),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_598),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_539),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_540),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_666),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_599),
.Y(n_817)
);

CKINVDCx20_ASAP7_75t_R g818 ( 
.A(n_666),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_543),
.Y(n_819)
);

INVxp67_ASAP7_75t_SL g820 ( 
.A(n_675),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_647),
.Y(n_821)
);

INVxp33_ASAP7_75t_SL g822 ( 
.A(n_542),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_545),
.Y(n_823)
);

INVxp33_ASAP7_75t_SL g824 ( 
.A(n_550),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_604),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_642),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_648),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_661),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_631),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_669),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_546),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_670),
.Y(n_832)
);

INVxp67_ASAP7_75t_SL g833 ( 
.A(n_675),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_679),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_548),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_647),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_559),
.Y(n_837)
);

INVxp33_ASAP7_75t_L g838 ( 
.A(n_631),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_647),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_702),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_638),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_681),
.Y(n_842)
);

INVxp33_ASAP7_75t_L g843 ( 
.A(n_638),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_686),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_560),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_564),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_697),
.Y(n_847)
);

INVxp33_ASAP7_75t_SL g848 ( 
.A(n_561),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_706),
.Y(n_849)
);

INVx3_ASAP7_75t_L g850 ( 
.A(n_841),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_757),
.B(n_552),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_841),
.Y(n_852)
);

INVx5_ASAP7_75t_L g853 ( 
.A(n_811),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_761),
.Y(n_854)
);

OA21x2_ASAP7_75t_L g855 ( 
.A1(n_760),
.A2(n_588),
.B(n_571),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_763),
.B(n_676),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_758),
.Y(n_857)
);

INVx5_ASAP7_75t_L g858 ( 
.A(n_811),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_762),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_811),
.Y(n_860)
);

BUFx6f_ASAP7_75t_L g861 ( 
.A(n_766),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_768),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_774),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_811),
.Y(n_864)
);

NOR2x1_ASAP7_75t_L g865 ( 
.A(n_780),
.B(n_683),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_778),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_781),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_782),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_783),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_785),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_760),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_770),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_787),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_777),
.B(n_557),
.Y(n_874)
);

INVxp67_ASAP7_75t_L g875 ( 
.A(n_794),
.Y(n_875)
);

CKINVDCx11_ASAP7_75t_R g876 ( 
.A(n_773),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_789),
.Y(n_877)
);

AND2x4_ASAP7_75t_L g878 ( 
.A(n_791),
.B(n_702),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_792),
.B(n_683),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_793),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_769),
.Y(n_881)
);

HB1xp67_ASAP7_75t_L g882 ( 
.A(n_764),
.Y(n_882)
);

OA21x2_ASAP7_75t_L g883 ( 
.A1(n_770),
.A2(n_784),
.B(n_771),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_795),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_771),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_784),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_775),
.B(n_678),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_821),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_798),
.B(n_840),
.Y(n_889)
);

INVx6_ASAP7_75t_L g890 ( 
.A(n_812),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_767),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_814),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_821),
.Y(n_893)
);

OAI21x1_ASAP7_75t_L g894 ( 
.A1(n_836),
.A2(n_839),
.B(n_588),
.Y(n_894)
);

BUFx6f_ASAP7_75t_L g895 ( 
.A(n_836),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_839),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_796),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_797),
.Y(n_898)
);

HB1xp67_ASAP7_75t_L g899 ( 
.A(n_815),
.Y(n_899)
);

INVxp67_ASAP7_75t_L g900 ( 
.A(n_809),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_812),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_779),
.A2(n_674),
.B1(n_714),
.B2(n_668),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_819),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_799),
.Y(n_904)
);

OA21x2_ASAP7_75t_L g905 ( 
.A1(n_800),
.A2(n_656),
.B(n_571),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_823),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_776),
.Y(n_907)
);

OAI22x1_ASAP7_75t_SL g908 ( 
.A1(n_773),
.A2(n_674),
.B1(n_714),
.B2(n_668),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_802),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_776),
.Y(n_910)
);

INVx3_ASAP7_75t_L g911 ( 
.A(n_803),
.Y(n_911)
);

INVx4_ASAP7_75t_L g912 ( 
.A(n_831),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_806),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_808),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_854),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_900),
.B(n_809),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_876),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_854),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_864),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_883),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_874),
.B(n_804),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_889),
.B(n_835),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_889),
.B(n_756),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_864),
.Y(n_924)
);

OA21x2_ASAP7_75t_L g925 ( 
.A1(n_894),
.A2(n_659),
.B(n_656),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_906),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_904),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_904),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_909),
.Y(n_929)
);

CKINVDCx20_ASAP7_75t_R g930 ( 
.A(n_881),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_874),
.B(n_807),
.Y(n_931)
);

NOR2xp67_ASAP7_75t_L g932 ( 
.A(n_912),
.B(n_837),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_883),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_906),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_892),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_889),
.B(n_659),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_889),
.B(n_845),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_883),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_881),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_909),
.Y(n_940)
);

INVxp67_ASAP7_75t_L g941 ( 
.A(n_891),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_883),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_898),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_898),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_898),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_875),
.B(n_820),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_882),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_898),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_891),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_899),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_885),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_898),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_914),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_914),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_890),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_914),
.Y(n_956)
);

AND2x4_ASAP7_75t_L g957 ( 
.A(n_878),
.B(n_833),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_914),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_903),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_912),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_912),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_871),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_886),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_886),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_914),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_912),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_907),
.B(n_846),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_911),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_890),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_901),
.B(n_684),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_890),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_902),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_R g973 ( 
.A(n_907),
.B(n_566),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_851),
.B(n_765),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_856),
.B(n_708),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_910),
.Y(n_976)
);

INVxp67_ASAP7_75t_L g977 ( 
.A(n_910),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_887),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_911),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_911),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_879),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_890),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_908),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_886),
.Y(n_984)
);

INVx3_ASAP7_75t_L g985 ( 
.A(n_871),
.Y(n_985)
);

AND2x6_ASAP7_75t_L g986 ( 
.A(n_865),
.B(n_684),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_902),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_908),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_878),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_879),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_897),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_879),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_879),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_878),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_897),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_901),
.B(n_790),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_913),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_878),
.Y(n_998)
);

AND2x4_ASAP7_75t_L g999 ( 
.A(n_901),
.B(n_810),
.Y(n_999)
);

HB1xp67_ASAP7_75t_L g1000 ( 
.A(n_867),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_901),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_901),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_901),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_941),
.B(n_805),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_962),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_SL g1006 ( 
.A(n_923),
.B(n_756),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_962),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_985),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_969),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_936),
.A2(n_905),
.B1(n_865),
.B2(n_855),
.Y(n_1010)
);

CKINVDCx16_ASAP7_75t_R g1011 ( 
.A(n_930),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_920),
.B(n_855),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_981),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_963),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_951),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_923),
.B(n_790),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_960),
.B(n_801),
.Y(n_1017)
);

NAND2xp33_ASAP7_75t_SL g1018 ( 
.A(n_973),
.B(n_976),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_990),
.Y(n_1019)
);

INVx2_ASAP7_75t_SL g1020 ( 
.A(n_916),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_992),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_917),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_920),
.B(n_855),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_993),
.Y(n_1024)
);

INVx5_ASAP7_75t_L g1025 ( 
.A(n_986),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_927),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_921),
.B(n_755),
.Y(n_1027)
);

AOI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_931),
.A2(n_569),
.B1(n_620),
.B2(n_551),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_957),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_951),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_961),
.B(n_801),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_933),
.B(n_855),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_936),
.A2(n_905),
.B1(n_888),
.B2(n_893),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_928),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_995),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_997),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_929),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_922),
.B(n_822),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_940),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_933),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_966),
.B(n_932),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_1000),
.Y(n_1042)
);

OAI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_937),
.A2(n_551),
.B1(n_620),
.B2(n_569),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_991),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_968),
.Y(n_1045)
);

AOI22xp33_ASAP7_75t_L g1046 ( 
.A1(n_957),
.A2(n_905),
.B1(n_888),
.B2(n_893),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_957),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_938),
.B(n_885),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_938),
.B(n_905),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_967),
.B(n_822),
.Y(n_1050)
);

BUFx3_ASAP7_75t_L g1051 ( 
.A(n_917),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_974),
.B(n_824),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_942),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_942),
.B(n_886),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_979),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_946),
.B(n_824),
.Y(n_1056)
);

AND3x2_ASAP7_75t_L g1057 ( 
.A(n_977),
.B(n_736),
.C(n_734),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_949),
.B(n_848),
.Y(n_1058)
);

INVx3_ASAP7_75t_L g1059 ( 
.A(n_963),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_980),
.A2(n_848),
.B1(n_526),
.B2(n_531),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_963),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_975),
.B(n_886),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_963),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_919),
.Y(n_1064)
);

INVx3_ASAP7_75t_L g1065 ( 
.A(n_964),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_986),
.B(n_895),
.Y(n_1066)
);

AND2x6_ASAP7_75t_L g1067 ( 
.A(n_924),
.B(n_524),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_978),
.B(n_998),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_964),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_964),
.Y(n_1070)
);

INVx8_ASAP7_75t_L g1071 ( 
.A(n_989),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_964),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_947),
.B(n_750),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_955),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_971),
.Y(n_1075)
);

CKINVDCx20_ASAP7_75t_R g1076 ( 
.A(n_930),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_984),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_982),
.Y(n_1078)
);

OAI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_994),
.A2(n_703),
.B1(n_746),
.B2(n_644),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_943),
.Y(n_1080)
);

INVx2_ASAP7_75t_SL g1081 ( 
.A(n_973),
.Y(n_1081)
);

NAND3xp33_ASAP7_75t_L g1082 ( 
.A(n_925),
.B(n_534),
.C(n_532),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_986),
.B(n_895),
.Y(n_1083)
);

INVxp67_ASAP7_75t_SL g1084 ( 
.A(n_984),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_935),
.B(n_829),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_SL g1086 ( 
.A1(n_972),
.A2(n_727),
.B1(n_816),
.B2(n_788),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_939),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_984),
.Y(n_1088)
);

NAND2xp33_ASAP7_75t_L g1089 ( 
.A(n_986),
.B(n_570),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_984),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_950),
.B(n_752),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_959),
.B(n_752),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_986),
.B(n_895),
.Y(n_1093)
);

OR2x6_ASAP7_75t_L g1094 ( 
.A(n_996),
.B(n_751),
.Y(n_1094)
);

BUFx3_ASAP7_75t_L g1095 ( 
.A(n_939),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_L g1096 ( 
.A(n_925),
.B(n_537),
.C(n_536),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_944),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_915),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_918),
.Y(n_1099)
);

INVxp67_ASAP7_75t_L g1100 ( 
.A(n_926),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_934),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_999),
.B(n_644),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_945),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_948),
.Y(n_1104)
);

INVxp33_ASAP7_75t_SL g1105 ( 
.A(n_983),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_999),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_952),
.Y(n_1107)
);

AOI22xp33_ASAP7_75t_L g1108 ( 
.A1(n_953),
.A2(n_549),
.B1(n_555),
.B2(n_544),
.Y(n_1108)
);

AND3x2_ASAP7_75t_L g1109 ( 
.A(n_972),
.B(n_745),
.C(n_739),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_987),
.A2(n_703),
.B1(n_746),
.B2(n_727),
.Y(n_1110)
);

INVx2_ASAP7_75t_SL g1111 ( 
.A(n_999),
.Y(n_1111)
);

AND2x6_ASAP7_75t_L g1112 ( 
.A(n_954),
.B(n_556),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_956),
.Y(n_1113)
);

INVx4_ASAP7_75t_L g1114 ( 
.A(n_1001),
.Y(n_1114)
);

AOI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_987),
.A2(n_694),
.B1(n_554),
.B2(n_583),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_988),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_958),
.Y(n_1117)
);

BUFx10_ASAP7_75t_L g1118 ( 
.A(n_965),
.Y(n_1118)
);

NOR2x1p5_ASAP7_75t_L g1119 ( 
.A(n_1002),
.B(n_754),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_970),
.B(n_753),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_925),
.B(n_759),
.Y(n_1121)
);

INVx3_ASAP7_75t_L g1122 ( 
.A(n_1002),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_970),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1003),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_981),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_981),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_915),
.Y(n_1127)
);

INVx2_ASAP7_75t_SL g1128 ( 
.A(n_916),
.Y(n_1128)
);

OAI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_922),
.A2(n_753),
.B1(n_759),
.B2(n_755),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_SL g1130 ( 
.A(n_927),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_922),
.B(n_776),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_969),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_947),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_962),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_962),
.Y(n_1135)
);

BUFx6f_ASAP7_75t_L g1136 ( 
.A(n_969),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_923),
.Y(n_1137)
);

AND2x6_ASAP7_75t_L g1138 ( 
.A(n_920),
.B(n_575),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_981),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_962),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1024),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1133),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_1076),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1053),
.Y(n_1144)
);

INVxp67_ASAP7_75t_L g1145 ( 
.A(n_1085),
.Y(n_1145)
);

BUFx2_ASAP7_75t_L g1146 ( 
.A(n_1087),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1053),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1099),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1137),
.B(n_1027),
.Y(n_1149)
);

BUFx10_ASAP7_75t_L g1150 ( 
.A(n_1091),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_1029),
.Y(n_1151)
);

AND2x6_ASAP7_75t_L g1152 ( 
.A(n_1029),
.B(n_585),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1024),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1137),
.B(n_586),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1139),
.Y(n_1155)
);

AOI22xp5_ASAP7_75t_L g1156 ( 
.A1(n_1029),
.A2(n_603),
.B1(n_613),
.B2(n_591),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_1052),
.B(n_788),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1139),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1019),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1013),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1040),
.B(n_614),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1021),
.Y(n_1162)
);

AND2x2_ASAP7_75t_SL g1163 ( 
.A(n_1011),
.B(n_816),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1073),
.Y(n_1164)
);

INVxp67_ASAP7_75t_L g1165 ( 
.A(n_1092),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1125),
.Y(n_1166)
);

BUFx3_ASAP7_75t_L g1167 ( 
.A(n_1132),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1020),
.B(n_772),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1126),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1026),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1019),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1034),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_1127),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1047),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1128),
.B(n_772),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1040),
.B(n_615),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1009),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1009),
.B(n_813),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1009),
.Y(n_1179)
);

AO22x2_ASAP7_75t_L g1180 ( 
.A1(n_1110),
.A2(n_605),
.B1(n_640),
.B2(n_573),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_1136),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_1019),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1015),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1039),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1121),
.B(n_1038),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1037),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_1095),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1058),
.B(n_786),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1045),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1079),
.B(n_818),
.Y(n_1190)
);

AND2x4_ASAP7_75t_L g1191 ( 
.A(n_1136),
.B(n_817),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1073),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1030),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1035),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1054),
.B(n_1046),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1136),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1036),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1106),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1055),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1005),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1117),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1016),
.A2(n_1006),
.B1(n_1094),
.B2(n_1131),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1028),
.B(n_786),
.Y(n_1203)
);

AND2x2_ASAP7_75t_SL g1204 ( 
.A(n_1028),
.B(n_1068),
.Y(n_1204)
);

BUFx4f_ASAP7_75t_L g1205 ( 
.A(n_1071),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1080),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1042),
.B(n_829),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1007),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1008),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1088),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1127),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1088),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1104),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1113),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1106),
.B(n_850),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1054),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1120),
.B(n_621),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1134),
.Y(n_1218)
);

OAI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1115),
.A2(n_688),
.B1(n_737),
.B2(n_728),
.C(n_682),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1048),
.Y(n_1220)
);

NAND2x1p5_ASAP7_75t_L g1221 ( 
.A(n_1081),
.B(n_850),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1044),
.B(n_838),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1074),
.B(n_825),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1135),
.Y(n_1224)
);

INVx4_ASAP7_75t_L g1225 ( 
.A(n_1088),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1140),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1056),
.B(n_838),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1048),
.Y(n_1228)
);

AND2x6_ASAP7_75t_L g1229 ( 
.A(n_1012),
.B(n_635),
.Y(n_1229)
);

BUFx6f_ASAP7_75t_L g1230 ( 
.A(n_1118),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1097),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1064),
.Y(n_1232)
);

AND2x4_ASAP7_75t_L g1233 ( 
.A(n_1075),
.B(n_826),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_1071),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_1118),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1103),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_SL g1237 ( 
.A1(n_1086),
.A2(n_738),
.B1(n_625),
.B2(n_634),
.Y(n_1237)
);

INVx1_ASAP7_75t_SL g1238 ( 
.A(n_1004),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1107),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1084),
.B(n_650),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_1070),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1084),
.B(n_664),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1012),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_SL g1244 ( 
.A(n_1018),
.B(n_578),
.Y(n_1244)
);

AOI222xp33_ASAP7_75t_L g1245 ( 
.A1(n_1043),
.A2(n_843),
.B1(n_748),
.B2(n_654),
.C1(n_828),
.C2(n_830),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1078),
.B(n_827),
.Y(n_1246)
);

INVxp67_ASAP7_75t_SL g1247 ( 
.A(n_1059),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1129),
.B(n_579),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1111),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1123),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1072),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1090),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1059),
.Y(n_1253)
);

BUFx6f_ASAP7_75t_L g1254 ( 
.A(n_1071),
.Y(n_1254)
);

INVx3_ASAP7_75t_L g1255 ( 
.A(n_1061),
.Y(n_1255)
);

BUFx2_ASAP7_75t_L g1256 ( 
.A(n_1073),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1061),
.Y(n_1257)
);

OR2x6_ASAP7_75t_L g1258 ( 
.A(n_1098),
.B(n_832),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1063),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1057),
.Y(n_1260)
);

AND2x6_ASAP7_75t_L g1261 ( 
.A(n_1023),
.B(n_692),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1063),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1014),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1065),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1050),
.B(n_843),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1014),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1065),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1069),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1069),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1032),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1062),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1041),
.B(n_580),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1138),
.Y(n_1273)
);

NAND2x1p5_ASAP7_75t_L g1274 ( 
.A(n_1025),
.B(n_1114),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1077),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1100),
.B(n_834),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1049),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1094),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1077),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1094),
.B(n_695),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1066),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1100),
.A2(n_730),
.B1(n_742),
.B2(n_718),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1066),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1119),
.B(n_842),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1083),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1124),
.B(n_1114),
.Y(n_1286)
);

NOR2xp33_ASAP7_75t_L g1287 ( 
.A(n_1017),
.B(n_622),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1010),
.B(n_743),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1101),
.Y(n_1289)
);

NAND3xp33_ASAP7_75t_L g1290 ( 
.A(n_1060),
.B(n_568),
.C(n_563),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1093),
.Y(n_1291)
);

BUFx6f_ASAP7_75t_L g1292 ( 
.A(n_1025),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1033),
.B(n_744),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1093),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_1025),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1022),
.Y(n_1296)
);

BUFx6f_ASAP7_75t_L g1297 ( 
.A(n_1067),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1122),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1067),
.B(n_871),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1122),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1082),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1051),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1082),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1109),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1096),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1102),
.B(n_844),
.Y(n_1306)
);

INVx8_ASAP7_75t_L g1307 ( 
.A(n_1130),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1031),
.B(n_847),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1067),
.B(n_872),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1096),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1112),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1112),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1130),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1109),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1089),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1108),
.A2(n_581),
.B1(n_593),
.B2(n_587),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1116),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1086),
.B(n_594),
.Y(n_1318)
);

AO22x2_ASAP7_75t_L g1319 ( 
.A1(n_1116),
.A2(n_849),
.B1(n_9),
.B2(n_17),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1105),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1053),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1052),
.B(n_622),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1053),
.B(n_872),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1053),
.B(n_872),
.Y(n_1324)
);

INVxp67_ASAP7_75t_L g1325 ( 
.A(n_1085),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1024),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1029),
.B(n_596),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1027),
.B(n_574),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1137),
.A2(n_895),
.B1(n_896),
.B2(n_558),
.Y(n_1329)
);

NAND3xp33_ASAP7_75t_SL g1330 ( 
.A(n_1157),
.B(n_590),
.C(n_582),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1144),
.B(n_867),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1165),
.B(n_592),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1177),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1160),
.Y(n_1334)
);

NAND2x1p5_ASAP7_75t_L g1335 ( 
.A(n_1151),
.B(n_894),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1144),
.A2(n_607),
.B1(n_608),
.B2(n_606),
.Y(n_1336)
);

OR2x2_ASAP7_75t_L g1337 ( 
.A(n_1149),
.B(n_868),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_SL g1338 ( 
.A(n_1202),
.B(n_1177),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_SL g1339 ( 
.A(n_1177),
.B(n_617),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1147),
.B(n_884),
.Y(n_1340)
);

AND2x4_ASAP7_75t_L g1341 ( 
.A(n_1286),
.B(n_868),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1147),
.B(n_884),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1188),
.B(n_595),
.Y(n_1343)
);

NAND2xp33_ASAP7_75t_L g1344 ( 
.A(n_1321),
.B(n_618),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1321),
.B(n_870),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1227),
.B(n_597),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1292),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1183),
.Y(n_1348)
);

AND2x2_ASAP7_75t_SL g1349 ( 
.A(n_1163),
.B(n_870),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1162),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1153),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1185),
.B(n_873),
.Y(n_1352)
);

AO22x1_ASAP7_75t_L g1353 ( 
.A1(n_1322),
.A2(n_601),
.B1(n_610),
.B2(n_609),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1216),
.B(n_1271),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1166),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1289),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1220),
.B(n_857),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1220),
.B(n_857),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_1238),
.B(n_1145),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_SL g1360 ( 
.A(n_1179),
.B(n_627),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1158),
.Y(n_1361)
);

INVx5_ASAP7_75t_L g1362 ( 
.A(n_1254),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1204),
.A2(n_558),
.B1(n_629),
.B2(n_628),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1169),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1228),
.B(n_859),
.Y(n_1365)
);

INVxp67_ASAP7_75t_L g1366 ( 
.A(n_1142),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1179),
.B(n_632),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_SL g1368 ( 
.A(n_1179),
.B(n_636),
.Y(n_1368)
);

NAND3xp33_ASAP7_75t_L g1369 ( 
.A(n_1217),
.B(n_863),
.C(n_859),
.Y(n_1369)
);

AND2x6_ASAP7_75t_SL g1370 ( 
.A(n_1190),
.B(n_558),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1326),
.Y(n_1371)
);

O2A1O1Ixp5_ASAP7_75t_L g1372 ( 
.A1(n_1315),
.A2(n_869),
.B(n_880),
.C(n_863),
.Y(n_1372)
);

AND2x6_ASAP7_75t_SL g1373 ( 
.A(n_1287),
.B(n_611),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1170),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1228),
.B(n_869),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1318),
.A2(n_646),
.B1(n_658),
.B2(n_639),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1195),
.A2(n_880),
.B(n_747),
.Y(n_1377)
);

INVx5_ASAP7_75t_L g1378 ( 
.A(n_1254),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1285),
.A2(n_672),
.B1(n_677),
.B2(n_667),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1277),
.B(n_850),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1325),
.B(n_612),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1203),
.A2(n_619),
.B1(n_626),
.B2(n_623),
.Y(n_1382)
);

NAND3xp33_ASAP7_75t_L g1383 ( 
.A(n_1245),
.B(n_685),
.C(n_680),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1181),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1281),
.A2(n_693),
.B1(n_696),
.B2(n_687),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1231),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1243),
.B(n_852),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1172),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1231),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1184),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1243),
.B(n_1270),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1283),
.A2(n_701),
.B1(n_704),
.B2(n_699),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1236),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1189),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1206),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1168),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_SL g1397 ( 
.A(n_1181),
.B(n_705),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1210),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_SL g1399 ( 
.A(n_1181),
.B(n_710),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1288),
.A2(n_713),
.B1(n_716),
.B2(n_711),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1196),
.B(n_1230),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_SL g1402 ( 
.A1(n_1273),
.A2(n_852),
.B(n_731),
.C(n_729),
.Y(n_1402)
);

XOR2xp5_ASAP7_75t_L g1403 ( 
.A(n_1296),
.B(n_1302),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1328),
.B(n_630),
.Y(n_1404)
);

NOR2x1p5_ASAP7_75t_L g1405 ( 
.A(n_1234),
.B(n_633),
.Y(n_1405)
);

INVx2_ASAP7_75t_SL g1406 ( 
.A(n_1196),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1250),
.B(n_641),
.Y(n_1407)
);

BUFx6f_ASAP7_75t_L g1408 ( 
.A(n_1210),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1236),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_SL g1410 ( 
.A1(n_1219),
.A2(n_645),
.B1(n_649),
.B2(n_643),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1239),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1154),
.B(n_651),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1291),
.B(n_652),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1294),
.A2(n_657),
.B1(n_660),
.B2(n_655),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1196),
.Y(n_1415)
);

INVx5_ASAP7_75t_L g1416 ( 
.A(n_1254),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1186),
.A2(n_862),
.B1(n_866),
.B2(n_861),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1175),
.B(n_662),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1213),
.Y(n_1419)
);

NAND2x1p5_ASAP7_75t_L g1420 ( 
.A(n_1151),
.B(n_853),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_SL g1421 ( 
.A(n_1230),
.B(n_853),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1306),
.A2(n_862),
.B1(n_866),
.B2(n_861),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1178),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1248),
.B(n_673),
.C(n_665),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_SL g1425 ( 
.A(n_1230),
.B(n_853),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1214),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1306),
.A2(n_862),
.B1(n_866),
.B2(n_861),
.Y(n_1427)
);

AND2x6_ASAP7_75t_SL g1428 ( 
.A(n_1320),
.B(n_1258),
.Y(n_1428)
);

NOR2xp33_ASAP7_75t_L g1429 ( 
.A(n_1150),
.B(n_689),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1222),
.B(n_690),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_SL g1431 ( 
.A(n_1235),
.B(n_853),
.Y(n_1431)
);

OR2x6_ASAP7_75t_L g1432 ( 
.A(n_1307),
.B(n_896),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1141),
.A2(n_698),
.B1(n_700),
.B2(n_691),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1232),
.A2(n_862),
.B1(n_866),
.B2(n_861),
.Y(n_1434)
);

OR2x6_ASAP7_75t_L g1435 ( 
.A(n_1307),
.B(n_896),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1265),
.B(n_709),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1193),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1148),
.Y(n_1438)
);

OR2x2_ASAP7_75t_SL g1439 ( 
.A(n_1320),
.B(n_1314),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_SL g1440 ( 
.A(n_1235),
.B(n_853),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1155),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1197),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1301),
.A2(n_858),
.B(n_853),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1182),
.B(n_712),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1199),
.Y(n_1445)
);

NOR2xp67_ASAP7_75t_L g1446 ( 
.A(n_1234),
.B(n_274),
.Y(n_1446)
);

OAI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1317),
.A2(n_717),
.B1(n_719),
.B2(n_715),
.Y(n_1447)
);

NAND2xp33_ASAP7_75t_L g1448 ( 
.A(n_1292),
.B(n_720),
.Y(n_1448)
);

NOR3xp33_ASAP7_75t_L g1449 ( 
.A(n_1237),
.B(n_724),
.C(n_722),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1194),
.A2(n_877),
.B1(n_726),
.B2(n_733),
.Y(n_1450)
);

AOI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1303),
.A2(n_735),
.B1(n_740),
.B2(n_725),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1207),
.B(n_741),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1182),
.B(n_896),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_SL g1454 ( 
.A(n_1235),
.B(n_858),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1150),
.B(n_1),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1167),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1201),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1198),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1286),
.B(n_275),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1143),
.B(n_2),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1292),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1210),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1198),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1241),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1276),
.B(n_2),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1251),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1159),
.B(n_877),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1171),
.B(n_877),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1323),
.B(n_1324),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1191),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1252),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1268),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1298),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1174),
.B(n_877),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1174),
.B(n_3),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1146),
.B(n_4),
.Y(n_1476)
);

AO22x1_ASAP7_75t_L g1477 ( 
.A1(n_1304),
.A2(n_6),
.B1(n_4),
.B2(n_5),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1187),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1278),
.A2(n_1229),
.B1(n_1261),
.B2(n_1308),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1249),
.B(n_5),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1308),
.B(n_6),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1295),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1191),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1200),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1305),
.B(n_7),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1310),
.B(n_7),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1240),
.B(n_8),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1242),
.B(n_10),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1295),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1280),
.B(n_11),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1208),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1209),
.B(n_12),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1173),
.B(n_276),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1293),
.A2(n_860),
.B1(n_278),
.B2(n_280),
.Y(n_1494)
);

OR2x2_ASAP7_75t_SL g1495 ( 
.A(n_1313),
.B(n_13),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1218),
.B(n_13),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1164),
.B(n_14),
.Y(n_1497)
);

NAND2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1297),
.B(n_15),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1192),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1224),
.B(n_15),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_SL g1501 ( 
.A(n_1205),
.B(n_282),
.Y(n_1501)
);

NOR2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1211),
.B(n_283),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1329),
.B(n_16),
.C(n_17),
.Y(n_1503)
);

BUFx4f_ASAP7_75t_L g1504 ( 
.A(n_1297),
.Y(n_1504)
);

INVx1_ASAP7_75t_SL g1505 ( 
.A(n_1256),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1226),
.B(n_18),
.Y(n_1506)
);

NAND2x1p5_ASAP7_75t_L g1507 ( 
.A(n_1263),
.B(n_284),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1255),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1275),
.B(n_19),
.Y(n_1509)
);

INVx3_ASAP7_75t_L g1510 ( 
.A(n_1295),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1275),
.B(n_19),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1300),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_SL g1513 ( 
.A(n_1205),
.B(n_287),
.Y(n_1513)
);

BUFx3_ASAP7_75t_L g1514 ( 
.A(n_1223),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1229),
.B(n_1261),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1261),
.B(n_20),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1255),
.Y(n_1517)
);

AOI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1261),
.A2(n_22),
.B1(n_20),
.B2(n_21),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1266),
.B(n_290),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1257),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1253),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1359),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1354),
.B(n_1396),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1391),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1386),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1334),
.Y(n_1526)
);

CKINVDCx8_ASAP7_75t_R g1527 ( 
.A(n_1428),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_SL g1528 ( 
.A(n_1349),
.B(n_1223),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1389),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1350),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1396),
.B(n_1233),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1457),
.Y(n_1532)
);

INVx2_ASAP7_75t_SL g1533 ( 
.A(n_1456),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1366),
.B(n_1258),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1355),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1364),
.Y(n_1536)
);

BUFx6f_ASAP7_75t_L g1537 ( 
.A(n_1362),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1393),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1438),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_SL g1540 ( 
.A(n_1356),
.B(n_1274),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1514),
.B(n_1233),
.Y(n_1541)
);

BUFx8_ASAP7_75t_L g1542 ( 
.A(n_1478),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1423),
.B(n_1246),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1505),
.Y(n_1544)
);

BUFx3_ASAP7_75t_L g1545 ( 
.A(n_1362),
.Y(n_1545)
);

CKINVDCx11_ASAP7_75t_R g1546 ( 
.A(n_1428),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1362),
.B(n_1378),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1409),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1374),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1388),
.Y(n_1550)
);

AO21x2_ASAP7_75t_L g1551 ( 
.A1(n_1443),
.A2(n_1176),
.B(n_1161),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1390),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1378),
.Y(n_1553)
);

BUFx3_ASAP7_75t_L g1554 ( 
.A(n_1378),
.Y(n_1554)
);

INVxp67_ASAP7_75t_L g1555 ( 
.A(n_1499),
.Y(n_1555)
);

NAND2xp33_ASAP7_75t_L g1556 ( 
.A(n_1416),
.B(n_1297),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_SL g1557 ( 
.A(n_1470),
.B(n_1246),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1416),
.Y(n_1558)
);

NOR2x1p5_ASAP7_75t_L g1559 ( 
.A(n_1330),
.B(n_1284),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1411),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1332),
.B(n_1290),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1394),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1395),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1419),
.Y(n_1564)
);

AO22x1_ASAP7_75t_L g1565 ( 
.A1(n_1449),
.A2(n_1152),
.B1(n_1284),
.B2(n_1260),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1426),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_SL g1567 ( 
.A(n_1410),
.B(n_1282),
.C(n_1244),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1333),
.Y(n_1568)
);

BUFx4f_ASAP7_75t_L g1569 ( 
.A(n_1459),
.Y(n_1569)
);

BUFx2_ASAP7_75t_L g1570 ( 
.A(n_1384),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_R g1571 ( 
.A(n_1416),
.B(n_1212),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1459),
.B(n_1279),
.Y(n_1572)
);

BUFx4f_ASAP7_75t_L g1573 ( 
.A(n_1493),
.Y(n_1573)
);

CKINVDCx8_ASAP7_75t_R g1574 ( 
.A(n_1373),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1505),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1520),
.Y(n_1576)
);

NOR3xp33_ASAP7_75t_SL g1577 ( 
.A(n_1410),
.B(n_1272),
.C(n_1327),
.Y(n_1577)
);

NOR3xp33_ASAP7_75t_SL g1578 ( 
.A(n_1455),
.B(n_1429),
.C(n_1465),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_L g1579 ( 
.A(n_1398),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1412),
.B(n_1337),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1442),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1445),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1483),
.Y(n_1583)
);

NOR3xp33_ASAP7_75t_SL g1584 ( 
.A(n_1447),
.B(n_1476),
.C(n_1497),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1352),
.B(n_1152),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_SL g1586 ( 
.A(n_1341),
.B(n_1212),
.Y(n_1586)
);

NOR3xp33_ASAP7_75t_SL g1587 ( 
.A(n_1383),
.B(n_1424),
.C(n_1481),
.Y(n_1587)
);

NOR3xp33_ASAP7_75t_SL g1588 ( 
.A(n_1424),
.B(n_1180),
.C(n_1319),
.Y(n_1588)
);

BUFx6f_ASAP7_75t_L g1589 ( 
.A(n_1398),
.Y(n_1589)
);

AND3x1_ASAP7_75t_SL g1590 ( 
.A(n_1502),
.B(n_1262),
.C(n_1259),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1436),
.B(n_1221),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1406),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1439),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_R g1594 ( 
.A(n_1504),
.B(n_1498),
.Y(n_1594)
);

BUFx2_ASAP7_75t_L g1595 ( 
.A(n_1341),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1437),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1382),
.B(n_1212),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1343),
.B(n_1152),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1387),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1338),
.A2(n_1346),
.B1(n_1381),
.B2(n_1452),
.Y(n_1600)
);

BUFx2_ASAP7_75t_L g1601 ( 
.A(n_1415),
.Y(n_1601)
);

BUFx6f_ASAP7_75t_L g1602 ( 
.A(n_1398),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1348),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1520),
.Y(n_1604)
);

BUFx4f_ASAP7_75t_L g1605 ( 
.A(n_1493),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1404),
.B(n_1316),
.Y(n_1606)
);

BUFx4f_ASAP7_75t_L g1607 ( 
.A(n_1493),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1484),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1491),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1403),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1430),
.B(n_1267),
.Y(n_1611)
);

AOI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1503),
.A2(n_1363),
.B1(n_1376),
.B2(n_1451),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1503),
.A2(n_1156),
.B1(n_1264),
.B2(n_1257),
.Y(n_1613)
);

INVx3_ASAP7_75t_SL g1614 ( 
.A(n_1460),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1413),
.B(n_1414),
.Y(n_1615)
);

AND2x6_ASAP7_75t_L g1616 ( 
.A(n_1347),
.B(n_1311),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1414),
.B(n_1247),
.Y(n_1617)
);

AND2x4_ASAP7_75t_L g1618 ( 
.A(n_1405),
.B(n_1257),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1466),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1418),
.B(n_1264),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1344),
.A2(n_1299),
.B1(n_1309),
.B2(n_1311),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1401),
.B(n_1264),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_R g1623 ( 
.A(n_1504),
.B(n_1312),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1407),
.B(n_1269),
.Y(n_1624)
);

INVx3_ASAP7_75t_L g1625 ( 
.A(n_1347),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1432),
.B(n_1225),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1490),
.B(n_1269),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1451),
.B(n_1215),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_R g1629 ( 
.A(n_1461),
.B(n_1312),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1485),
.B(n_1225),
.Y(n_1630)
);

NOR3xp33_ASAP7_75t_SL g1631 ( 
.A(n_1480),
.B(n_21),
.C(n_22),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1441),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1464),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_R g1634 ( 
.A(n_1461),
.B(n_292),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1471),
.Y(n_1635)
);

NOR2xp33_ASAP7_75t_R g1636 ( 
.A(n_1482),
.B(n_293),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1408),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1521),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1512),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1444),
.B(n_23),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1432),
.B(n_294),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1486),
.B(n_23),
.Y(n_1642)
);

INVx3_ASAP7_75t_L g1643 ( 
.A(n_1482),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1373),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1432),
.B(n_295),
.Y(n_1645)
);

BUFx6f_ASAP7_75t_L g1646 ( 
.A(n_1408),
.Y(n_1646)
);

NAND2xp33_ASAP7_75t_SL g1647 ( 
.A(n_1408),
.B(n_24),
.Y(n_1647)
);

INVx5_ASAP7_75t_L g1648 ( 
.A(n_1462),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1351),
.Y(n_1649)
);

CKINVDCx20_ASAP7_75t_R g1650 ( 
.A(n_1495),
.Y(n_1650)
);

AND3x1_ASAP7_75t_SL g1651 ( 
.A(n_1370),
.B(n_24),
.C(n_25),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1435),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_SL g1653 ( 
.A(n_1479),
.B(n_26),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1489),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1361),
.Y(n_1655)
);

AND2x6_ASAP7_75t_L g1656 ( 
.A(n_1510),
.B(n_297),
.Y(n_1656)
);

INVx3_ASAP7_75t_L g1657 ( 
.A(n_1510),
.Y(n_1657)
);

INVx3_ASAP7_75t_L g1658 ( 
.A(n_1462),
.Y(n_1658)
);

INVx1_ASAP7_75t_SL g1659 ( 
.A(n_1475),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1371),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1331),
.Y(n_1661)
);

BUFx4f_ASAP7_75t_L g1662 ( 
.A(n_1462),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1380),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1472),
.Y(n_1664)
);

INVx5_ASAP7_75t_L g1665 ( 
.A(n_1435),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1469),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1473),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1487),
.B(n_28),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1340),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1488),
.B(n_1342),
.Y(n_1670)
);

NOR2xp33_ASAP7_75t_L g1671 ( 
.A(n_1353),
.B(n_30),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1345),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1357),
.B(n_1358),
.Y(n_1673)
);

INVx2_ASAP7_75t_SL g1674 ( 
.A(n_1435),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1365),
.B(n_30),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1375),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1433),
.B(n_31),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1508),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1517),
.Y(n_1679)
);

INVx2_ASAP7_75t_L g1680 ( 
.A(n_1458),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1433),
.B(n_32),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_1370),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1463),
.B(n_33),
.Y(n_1683)
);

NOR3xp33_ASAP7_75t_SL g1684 ( 
.A(n_1339),
.B(n_33),
.C(n_34),
.Y(n_1684)
);

NOR3xp33_ASAP7_75t_L g1685 ( 
.A(n_1360),
.B(n_35),
.C(n_36),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1385),
.B(n_35),
.Y(n_1686)
);

BUFx6f_ASAP7_75t_L g1687 ( 
.A(n_1507),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1367),
.Y(n_1688)
);

BUFx3_ASAP7_75t_L g1689 ( 
.A(n_1507),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1492),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1496),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1420),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1392),
.B(n_36),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1379),
.B(n_37),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1368),
.B(n_518),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1500),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1506),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1509),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1511),
.B(n_1397),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1335),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1399),
.B(n_37),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1421),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1336),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1425),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1431),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1372),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_R g1707 ( 
.A(n_1448),
.B(n_298),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1450),
.B(n_38),
.Y(n_1708)
);

INVxp67_ASAP7_75t_SL g1709 ( 
.A(n_1453),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1706),
.A2(n_1377),
.B(n_1515),
.Y(n_1710)
);

OAI21x1_ASAP7_75t_L g1711 ( 
.A1(n_1706),
.A2(n_1474),
.B(n_1468),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1580),
.B(n_1477),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1575),
.Y(n_1713)
);

NOR2xp67_ASAP7_75t_L g1714 ( 
.A(n_1522),
.B(n_1369),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1700),
.A2(n_1467),
.B(n_1494),
.Y(n_1715)
);

AOI221x1_ASAP7_75t_L g1716 ( 
.A1(n_1666),
.A2(n_1516),
.B1(n_1369),
.B2(n_1400),
.C(n_1402),
.Y(n_1716)
);

INVx2_ASAP7_75t_SL g1717 ( 
.A(n_1542),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1561),
.B(n_1501),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1544),
.Y(n_1719)
);

A2O1A1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1606),
.A2(n_1513),
.B(n_1518),
.C(n_1519),
.Y(n_1720)
);

BUFx2_ASAP7_75t_L g1721 ( 
.A(n_1595),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1581),
.Y(n_1722)
);

AOI221xp5_ASAP7_75t_SL g1723 ( 
.A1(n_1612),
.A2(n_1454),
.B1(n_1440),
.B2(n_1427),
.C(n_1422),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1670),
.A2(n_1551),
.B(n_1524),
.Y(n_1724)
);

OAI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1621),
.A2(n_1420),
.B(n_1434),
.Y(n_1725)
);

OAI21x1_ASAP7_75t_L g1726 ( 
.A1(n_1673),
.A2(n_1417),
.B(n_1446),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1524),
.B(n_38),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1526),
.Y(n_1728)
);

AOI21xp5_ASAP7_75t_L g1729 ( 
.A1(n_1569),
.A2(n_516),
.B(n_301),
.Y(n_1729)
);

AOI221xp5_ASAP7_75t_L g1730 ( 
.A1(n_1578),
.A2(n_41),
.B1(n_39),
.B2(n_40),
.C(n_42),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1523),
.B(n_39),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1542),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1661),
.B(n_1669),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1672),
.B(n_41),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_SL g1735 ( 
.A1(n_1585),
.A2(n_43),
.B(n_44),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1532),
.Y(n_1736)
);

AOI21xp5_ASAP7_75t_L g1737 ( 
.A1(n_1569),
.A2(n_302),
.B(n_299),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1539),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1615),
.A2(n_305),
.B(n_304),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1630),
.A2(n_309),
.B(n_308),
.Y(n_1740)
);

AOI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1709),
.A2(n_311),
.B(n_310),
.Y(n_1741)
);

OAI21x1_ASAP7_75t_L g1742 ( 
.A1(n_1599),
.A2(n_314),
.B(n_313),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1677),
.B(n_43),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1699),
.A2(n_515),
.B(n_316),
.Y(n_1744)
);

OAI21x1_ASAP7_75t_L g1745 ( 
.A1(n_1599),
.A2(n_318),
.B(n_315),
.Y(n_1745)
);

OA21x2_ASAP7_75t_L g1746 ( 
.A1(n_1627),
.A2(n_321),
.B(n_320),
.Y(n_1746)
);

AOI21xp5_ASAP7_75t_L g1747 ( 
.A1(n_1624),
.A2(n_513),
.B(n_323),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1618),
.B(n_322),
.Y(n_1748)
);

AOI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1617),
.A2(n_325),
.B(n_324),
.Y(n_1749)
);

AOI21xp5_ASAP7_75t_L g1750 ( 
.A1(n_1591),
.A2(n_327),
.B(n_326),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1676),
.A2(n_329),
.B(n_328),
.Y(n_1751)
);

OAI21x1_ASAP7_75t_SL g1752 ( 
.A1(n_1675),
.A2(n_45),
.B(n_46),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1547),
.Y(n_1753)
);

OAI21x1_ASAP7_75t_L g1754 ( 
.A1(n_1663),
.A2(n_331),
.B(n_330),
.Y(n_1754)
);

AO31x2_ASAP7_75t_L g1755 ( 
.A1(n_1642),
.A2(n_48),
.A3(n_46),
.B(n_47),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1697),
.B(n_47),
.Y(n_1756)
);

HB1xp67_ASAP7_75t_L g1757 ( 
.A(n_1531),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1582),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_SL g1759 ( 
.A(n_1600),
.B(n_49),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1611),
.B(n_49),
.Y(n_1760)
);

AND2x4_ASAP7_75t_L g1761 ( 
.A(n_1618),
.B(n_1547),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1659),
.B(n_50),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1530),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1535),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1665),
.A2(n_512),
.B(n_337),
.Y(n_1765)
);

INVx4_ASAP7_75t_SL g1766 ( 
.A(n_1537),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1536),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1567),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_1768)
);

OAI21xp5_ASAP7_75t_L g1769 ( 
.A1(n_1584),
.A2(n_52),
.B(n_53),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1703),
.B(n_335),
.Y(n_1770)
);

INVx2_ASAP7_75t_SL g1771 ( 
.A(n_1533),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1549),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1690),
.B(n_54),
.Y(n_1773)
);

BUFx6f_ASAP7_75t_L g1774 ( 
.A(n_1537),
.Y(n_1774)
);

BUFx12f_ASAP7_75t_L g1775 ( 
.A(n_1546),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1681),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.C(n_57),
.Y(n_1776)
);

AO21x2_ASAP7_75t_L g1777 ( 
.A1(n_1587),
.A2(n_340),
.B(n_339),
.Y(n_1777)
);

OR2x6_ASAP7_75t_L g1778 ( 
.A(n_1641),
.B(n_341),
.Y(n_1778)
);

NAND2xp33_ASAP7_75t_L g1779 ( 
.A(n_1577),
.B(n_55),
.Y(n_1779)
);

INVx1_ASAP7_75t_SL g1780 ( 
.A(n_1614),
.Y(n_1780)
);

NOR2xp67_ASAP7_75t_L g1781 ( 
.A(n_1610),
.B(n_343),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1568),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1696),
.B(n_57),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1596),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1550),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1620),
.B(n_58),
.Y(n_1786)
);

AOI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1598),
.A2(n_59),
.B(n_60),
.Y(n_1787)
);

AO31x2_ASAP7_75t_L g1788 ( 
.A1(n_1668),
.A2(n_62),
.A3(n_59),
.B(n_61),
.Y(n_1788)
);

OAI21x1_ASAP7_75t_L g1789 ( 
.A1(n_1525),
.A2(n_347),
.B(n_344),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1665),
.A2(n_354),
.B(n_352),
.Y(n_1790)
);

NAND2x1p5_ASAP7_75t_L g1791 ( 
.A(n_1648),
.B(n_359),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1552),
.Y(n_1792)
);

BUFx8_ASAP7_75t_L g1793 ( 
.A(n_1570),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1556),
.A2(n_511),
.B(n_362),
.Y(n_1794)
);

BUFx5_ASAP7_75t_L g1795 ( 
.A(n_1616),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1698),
.B(n_63),
.Y(n_1796)
);

INVxp67_ASAP7_75t_SL g1797 ( 
.A(n_1555),
.Y(n_1797)
);

NOR2x1_ASAP7_75t_L g1798 ( 
.A(n_1689),
.B(n_361),
.Y(n_1798)
);

OAI21x1_ASAP7_75t_L g1799 ( 
.A1(n_1529),
.A2(n_365),
.B(n_364),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1573),
.A2(n_367),
.B(n_366),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1528),
.B(n_64),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1671),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.C(n_67),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1538),
.A2(n_369),
.B(n_368),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1537),
.Y(n_1804)
);

O2A1O1Ixp5_ASAP7_75t_L g1805 ( 
.A1(n_1693),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1558),
.Y(n_1806)
);

A2O1A1Ixp33_ASAP7_75t_L g1807 ( 
.A1(n_1686),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1807)
);

AOI221x1_ASAP7_75t_L g1808 ( 
.A1(n_1685),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.C(n_71),
.Y(n_1808)
);

AO31x2_ASAP7_75t_L g1809 ( 
.A1(n_1632),
.A2(n_1639),
.A3(n_1563),
.B(n_1564),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1583),
.B(n_71),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1597),
.B(n_1534),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1573),
.A2(n_371),
.B(n_370),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1572),
.B(n_72),
.Y(n_1813)
);

OAI21x1_ASAP7_75t_L g1814 ( 
.A1(n_1548),
.A2(n_373),
.B(n_372),
.Y(n_1814)
);

BUFx3_ASAP7_75t_L g1815 ( 
.A(n_1558),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1558),
.Y(n_1816)
);

OAI21x1_ASAP7_75t_SL g1817 ( 
.A1(n_1701),
.A2(n_73),
.B(n_74),
.Y(n_1817)
);

OAI21x1_ASAP7_75t_L g1818 ( 
.A1(n_1560),
.A2(n_376),
.B(n_375),
.Y(n_1818)
);

BUFx6f_ASAP7_75t_L g1819 ( 
.A(n_1662),
.Y(n_1819)
);

OAI22x1_ASAP7_75t_L g1820 ( 
.A1(n_1559),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_1820)
);

A2O1A1Ixp33_ASAP7_75t_L g1821 ( 
.A1(n_1694),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1572),
.B(n_77),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1541),
.B(n_1628),
.Y(n_1823)
);

AOI21xp5_ASAP7_75t_SL g1824 ( 
.A1(n_1641),
.A2(n_383),
.B(n_381),
.Y(n_1824)
);

A2O1A1Ixp33_ASAP7_75t_L g1825 ( 
.A1(n_1605),
.A2(n_1607),
.B(n_1588),
.C(n_1695),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1545),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1541),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_SL g1828 ( 
.A(n_1687),
.B(n_384),
.Y(n_1828)
);

INVx5_ASAP7_75t_L g1829 ( 
.A(n_1648),
.Y(n_1829)
);

INVx4_ASAP7_75t_L g1830 ( 
.A(n_1648),
.Y(n_1830)
);

AOI21x1_ASAP7_75t_L g1831 ( 
.A1(n_1565),
.A2(n_386),
.B(n_385),
.Y(n_1831)
);

NOR2xp67_ASAP7_75t_L g1832 ( 
.A(n_1679),
.B(n_387),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1562),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1566),
.Y(n_1834)
);

INVx2_ASAP7_75t_SL g1835 ( 
.A(n_1553),
.Y(n_1835)
);

O2A1O1Ixp5_ASAP7_75t_L g1836 ( 
.A1(n_1653),
.A2(n_1605),
.B(n_1607),
.C(n_1647),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1601),
.Y(n_1837)
);

AO31x2_ASAP7_75t_L g1838 ( 
.A1(n_1633),
.A2(n_81),
.A3(n_78),
.B(n_80),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1637),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1708),
.B(n_80),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_SL g1841 ( 
.A(n_1691),
.B(n_81),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1691),
.B(n_82),
.Y(n_1842)
);

BUFx6f_ASAP7_75t_L g1843 ( 
.A(n_1662),
.Y(n_1843)
);

BUFx4f_ASAP7_75t_SL g1844 ( 
.A(n_1554),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1684),
.B(n_82),
.C(n_83),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1691),
.B(n_83),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1638),
.Y(n_1847)
);

A2O1A1Ixp33_ASAP7_75t_L g1848 ( 
.A1(n_1695),
.A2(n_1640),
.B(n_1645),
.C(n_1631),
.Y(n_1848)
);

A2O1A1Ixp33_ASAP7_75t_L g1849 ( 
.A1(n_1645),
.A2(n_86),
.B(n_84),
.C(n_85),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_L g1850 ( 
.A(n_1576),
.B(n_389),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_SL g1851 ( 
.A1(n_1652),
.A2(n_84),
.B(n_85),
.Y(n_1851)
);

A2O1A1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1543),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_L g1853 ( 
.A1(n_1613),
.A2(n_509),
.B(n_393),
.Y(n_1853)
);

OAI21xp5_ASAP7_75t_L g1854 ( 
.A1(n_1557),
.A2(n_1702),
.B(n_1704),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1649),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1688),
.B(n_88),
.Y(n_1856)
);

A2O1A1Ixp33_ASAP7_75t_L g1857 ( 
.A1(n_1705),
.A2(n_1593),
.B(n_1586),
.C(n_1603),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1626),
.B(n_391),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1608),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1683),
.B(n_1609),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1687),
.A2(n_508),
.B(n_395),
.Y(n_1861)
);

OAI21x1_ASAP7_75t_L g1862 ( 
.A1(n_1576),
.A2(n_396),
.B(n_394),
.Y(n_1862)
);

OAI21x1_ASAP7_75t_L g1863 ( 
.A1(n_1604),
.A2(n_400),
.B(n_398),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1619),
.B(n_89),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1604),
.A2(n_404),
.B(n_401),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1635),
.Y(n_1866)
);

OAI22xp5_ASAP7_75t_L g1867 ( 
.A1(n_1718),
.A2(n_1527),
.B1(n_1650),
.B2(n_1574),
.Y(n_1867)
);

AOI221xp5_ASAP7_75t_L g1868 ( 
.A1(n_1730),
.A2(n_1682),
.B1(n_1644),
.B2(n_1707),
.C(n_1655),
.Y(n_1868)
);

AOI22xp33_ASAP7_75t_L g1869 ( 
.A1(n_1769),
.A2(n_1656),
.B1(n_1687),
.B2(n_1594),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1860),
.B(n_1678),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1757),
.B(n_1660),
.Y(n_1871)
);

AND2x4_ASAP7_75t_L g1872 ( 
.A(n_1761),
.B(n_1674),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1733),
.B(n_1664),
.Y(n_1873)
);

OAI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1848),
.A2(n_1592),
.B1(n_1626),
.B2(n_1622),
.Y(n_1874)
);

INVx3_ASAP7_75t_L g1875 ( 
.A(n_1793),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1722),
.Y(n_1876)
);

NAND2x1p5_ASAP7_75t_L g1877 ( 
.A(n_1829),
.B(n_1692),
.Y(n_1877)
);

INVx5_ASAP7_75t_L g1878 ( 
.A(n_1829),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1761),
.B(n_1622),
.Y(n_1879)
);

BUFx12f_ASAP7_75t_L g1880 ( 
.A(n_1793),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1827),
.B(n_1858),
.Y(n_1881)
);

INVx1_ASAP7_75t_SL g1882 ( 
.A(n_1719),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1724),
.A2(n_1540),
.B(n_1692),
.Y(n_1883)
);

NAND2x1p5_ASAP7_75t_L g1884 ( 
.A(n_1829),
.B(n_1625),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1809),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1858),
.B(n_1658),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_SL g1887 ( 
.A1(n_1779),
.A2(n_1656),
.B1(n_1651),
.B2(n_1634),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1809),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1809),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1736),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1844),
.Y(n_1891)
);

INVx3_ASAP7_75t_L g1892 ( 
.A(n_1819),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_L g1893 ( 
.A1(n_1759),
.A2(n_1656),
.B1(n_1667),
.B2(n_1636),
.Y(n_1893)
);

BUFx6f_ASAP7_75t_L g1894 ( 
.A(n_1819),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1823),
.B(n_1680),
.Y(n_1895)
);

NAND2x1_ASAP7_75t_L g1896 ( 
.A(n_1798),
.B(n_1656),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1712),
.B(n_1625),
.Y(n_1897)
);

BUFx6f_ASAP7_75t_L g1898 ( 
.A(n_1819),
.Y(n_1898)
);

OAI21xp33_ASAP7_75t_L g1899 ( 
.A1(n_1768),
.A2(n_1571),
.B(n_1623),
.Y(n_1899)
);

NOR2xp33_ASAP7_75t_R g1900 ( 
.A(n_1843),
.B(n_1658),
.Y(n_1900)
);

A2O1A1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1720),
.A2(n_1643),
.B(n_1657),
.C(n_1654),
.Y(n_1901)
);

INVxp67_ASAP7_75t_L g1902 ( 
.A(n_1713),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1839),
.B(n_1643),
.Y(n_1903)
);

OR2x6_ASAP7_75t_L g1904 ( 
.A(n_1778),
.B(n_1579),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1802),
.A2(n_1654),
.B1(n_1657),
.B2(n_1616),
.Y(n_1905)
);

AO21x1_ASAP7_75t_L g1906 ( 
.A1(n_1787),
.A2(n_1590),
.B(n_91),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1728),
.Y(n_1907)
);

INVx3_ASAP7_75t_L g1908 ( 
.A(n_1843),
.Y(n_1908)
);

INVx4_ASAP7_75t_L g1909 ( 
.A(n_1843),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1749),
.A2(n_1616),
.B(n_1629),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1763),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1753),
.B(n_1579),
.Y(n_1912)
);

BUFx6f_ASAP7_75t_L g1913 ( 
.A(n_1774),
.Y(n_1913)
);

NAND2xp33_ASAP7_75t_L g1914 ( 
.A(n_1825),
.B(n_1795),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1770),
.B(n_1589),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1738),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1758),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1778),
.B(n_1589),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1731),
.B(n_1602),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_SL g1920 ( 
.A(n_1836),
.B(n_1811),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_SL g1921 ( 
.A1(n_1845),
.A2(n_1646),
.B1(n_1602),
.B2(n_93),
.Y(n_1921)
);

NAND2x1_ASAP7_75t_L g1922 ( 
.A(n_1746),
.B(n_1602),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1727),
.B(n_1646),
.Y(n_1923)
);

AOI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1710),
.A2(n_406),
.B(n_405),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1764),
.Y(n_1925)
);

AND2x4_ASAP7_75t_L g1926 ( 
.A(n_1766),
.B(n_407),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1784),
.B(n_91),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1767),
.Y(n_1928)
);

OAI21x1_ASAP7_75t_SL g1929 ( 
.A1(n_1735),
.A2(n_92),
.B(n_94),
.Y(n_1929)
);

BUFx2_ASAP7_75t_SL g1930 ( 
.A(n_1771),
.Y(n_1930)
);

INVx4_ASAP7_75t_L g1931 ( 
.A(n_1766),
.Y(n_1931)
);

INVx3_ASAP7_75t_L g1932 ( 
.A(n_1815),
.Y(n_1932)
);

HB1xp67_ASAP7_75t_L g1933 ( 
.A(n_1772),
.Y(n_1933)
);

OAI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1857),
.A2(n_98),
.B1(n_94),
.B2(n_95),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1785),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1847),
.Y(n_1936)
);

INVx1_ASAP7_75t_SL g1937 ( 
.A(n_1782),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1786),
.B(n_98),
.Y(n_1938)
);

INVx3_ASAP7_75t_L g1939 ( 
.A(n_1774),
.Y(n_1939)
);

BUFx4f_ASAP7_75t_SL g1940 ( 
.A(n_1775),
.Y(n_1940)
);

BUFx2_ASAP7_75t_SL g1941 ( 
.A(n_1780),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1797),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1774),
.Y(n_1943)
);

OA21x2_ASAP7_75t_L g1944 ( 
.A1(n_1726),
.A2(n_1711),
.B(n_1716),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1792),
.Y(n_1945)
);

INVx2_ASAP7_75t_SL g1946 ( 
.A(n_1804),
.Y(n_1946)
);

AND2x2_ASAP7_75t_L g1947 ( 
.A(n_1760),
.B(n_408),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1859),
.B(n_99),
.Y(n_1948)
);

BUFx3_ASAP7_75t_L g1949 ( 
.A(n_1721),
.Y(n_1949)
);

BUFx2_ASAP7_75t_L g1950 ( 
.A(n_1833),
.Y(n_1950)
);

NOR2xp33_ASAP7_75t_L g1951 ( 
.A(n_1837),
.B(n_409),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1834),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1806),
.B(n_410),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_L g1954 ( 
.A(n_1804),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1866),
.B(n_100),
.Y(n_1955)
);

A2O1A1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1853),
.A2(n_104),
.B(n_101),
.C(n_102),
.Y(n_1956)
);

INVx6_ASAP7_75t_L g1957 ( 
.A(n_1804),
.Y(n_1957)
);

A2O1A1Ixp33_ASAP7_75t_L g1958 ( 
.A1(n_1805),
.A2(n_105),
.B(n_102),
.C(n_104),
.Y(n_1958)
);

BUFx3_ASAP7_75t_L g1959 ( 
.A(n_1826),
.Y(n_1959)
);

AOI21xp5_ASAP7_75t_L g1960 ( 
.A1(n_1741),
.A2(n_413),
.B(n_411),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1840),
.B(n_105),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1855),
.Y(n_1962)
);

NOR2xp33_ASAP7_75t_L g1963 ( 
.A(n_1856),
.B(n_414),
.Y(n_1963)
);

AND2x4_ASAP7_75t_L g1964 ( 
.A(n_1816),
.B(n_415),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1734),
.B(n_106),
.Y(n_1965)
);

OAI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1714),
.A2(n_108),
.B1(n_106),
.B2(n_107),
.Y(n_1966)
);

O2A1O1Ixp33_ASAP7_75t_SL g1967 ( 
.A1(n_1849),
.A2(n_109),
.B(n_107),
.C(n_108),
.Y(n_1967)
);

OAI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1801),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_1968)
);

AND2x4_ASAP7_75t_L g1969 ( 
.A(n_1854),
.B(n_1748),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_SL g1970 ( 
.A(n_1781),
.B(n_416),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1838),
.Y(n_1971)
);

HB1xp67_ASAP7_75t_L g1972 ( 
.A(n_1842),
.Y(n_1972)
);

OAI211xp5_ASAP7_75t_L g1973 ( 
.A1(n_1921),
.A2(n_1808),
.B(n_1807),
.C(n_1821),
.Y(n_1973)
);

BUFx2_ASAP7_75t_L g1974 ( 
.A(n_1890),
.Y(n_1974)
);

AOI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1920),
.A2(n_1831),
.B(n_1739),
.Y(n_1975)
);

OAI21x1_ASAP7_75t_L g1976 ( 
.A1(n_1924),
.A2(n_1715),
.B(n_1725),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1950),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1907),
.Y(n_1978)
);

OA21x2_ASAP7_75t_L g1979 ( 
.A1(n_1971),
.A2(n_1776),
.B(n_1745),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1911),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1950),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1913),
.Y(n_1982)
);

OAI21x1_ASAP7_75t_L g1983 ( 
.A1(n_1922),
.A2(n_1742),
.B(n_1754),
.Y(n_1983)
);

OR2x6_ASAP7_75t_L g1984 ( 
.A(n_1883),
.B(n_1824),
.Y(n_1984)
);

NAND3xp33_ASAP7_75t_L g1985 ( 
.A(n_1956),
.B(n_1852),
.C(n_1841),
.Y(n_1985)
);

AO21x2_ASAP7_75t_L g1986 ( 
.A1(n_1885),
.A2(n_1889),
.B(n_1888),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1925),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1887),
.A2(n_1743),
.B1(n_1783),
.B2(n_1773),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1903),
.Y(n_1989)
);

OAI21xp5_ASAP7_75t_L g1990 ( 
.A1(n_1960),
.A2(n_1958),
.B(n_1934),
.Y(n_1990)
);

OAI21x1_ASAP7_75t_L g1991 ( 
.A1(n_1944),
.A2(n_1863),
.B(n_1862),
.Y(n_1991)
);

OAI21x1_ASAP7_75t_SL g1992 ( 
.A1(n_1906),
.A2(n_1752),
.B(n_1817),
.Y(n_1992)
);

AOI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1901),
.A2(n_1794),
.B(n_1747),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1928),
.B(n_1717),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1933),
.B(n_1846),
.Y(n_1995)
);

AOI22xp33_ASAP7_75t_L g1996 ( 
.A1(n_1968),
.A2(n_1820),
.B1(n_1777),
.B2(n_1756),
.Y(n_1996)
);

OAI21x1_ASAP7_75t_L g1997 ( 
.A1(n_1944),
.A2(n_1865),
.B(n_1799),
.Y(n_1997)
);

AOI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1868),
.A2(n_1796),
.B1(n_1762),
.B2(n_1800),
.Y(n_1998)
);

NAND2x1p5_ASAP7_75t_L g1999 ( 
.A(n_1878),
.B(n_1746),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1880),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1935),
.B(n_1732),
.Y(n_2001)
);

BUFx2_ASAP7_75t_SL g2002 ( 
.A(n_1931),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1972),
.B(n_1864),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1945),
.Y(n_2004)
);

AND2x4_ASAP7_75t_L g2005 ( 
.A(n_1952),
.B(n_1835),
.Y(n_2005)
);

OAI21x1_ASAP7_75t_L g2006 ( 
.A1(n_1910),
.A2(n_1803),
.B(n_1789),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1959),
.Y(n_2007)
);

OAI21x1_ASAP7_75t_L g2008 ( 
.A1(n_1896),
.A2(n_1818),
.B(n_1814),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1962),
.Y(n_2009)
);

AND2x4_ASAP7_75t_L g2010 ( 
.A(n_1949),
.B(n_1838),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1870),
.B(n_1788),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1936),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1902),
.B(n_1838),
.Y(n_2013)
);

CKINVDCx20_ASAP7_75t_R g2014 ( 
.A(n_1940),
.Y(n_2014)
);

BUFx12f_ASAP7_75t_L g2015 ( 
.A(n_1891),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1876),
.Y(n_2016)
);

AO21x1_ASAP7_75t_L g2017 ( 
.A1(n_1966),
.A2(n_1744),
.B(n_1813),
.Y(n_2017)
);

OAI21x1_ASAP7_75t_SL g2018 ( 
.A1(n_1929),
.A2(n_1851),
.B(n_1828),
.Y(n_2018)
);

BUFx10_ASAP7_75t_L g2019 ( 
.A(n_1926),
.Y(n_2019)
);

AOI21xp5_ASAP7_75t_L g2020 ( 
.A1(n_1914),
.A2(n_1812),
.B(n_1737),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1871),
.B(n_1788),
.Y(n_2021)
);

OAI22xp5_ASAP7_75t_L g2022 ( 
.A1(n_1869),
.A2(n_1810),
.B1(n_1822),
.B2(n_1729),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1917),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1897),
.B(n_1788),
.Y(n_2024)
);

OAI21x1_ASAP7_75t_L g2025 ( 
.A1(n_1877),
.A2(n_1790),
.B(n_1765),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1873),
.Y(n_2026)
);

OAI21xp5_ASAP7_75t_L g2027 ( 
.A1(n_1893),
.A2(n_1750),
.B(n_1751),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1903),
.B(n_1755),
.Y(n_2028)
);

AND2x2_ASAP7_75t_L g2029 ( 
.A(n_1919),
.B(n_1755),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1948),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_R g2031 ( 
.A(n_2014),
.B(n_1875),
.Y(n_2031)
);

INVx4_ASAP7_75t_SL g2032 ( 
.A(n_1984),
.Y(n_2032)
);

AOI22xp5_ASAP7_75t_L g2033 ( 
.A1(n_1973),
.A2(n_1969),
.B1(n_1899),
.B2(n_1904),
.Y(n_2033)
);

AOI221xp5_ASAP7_75t_L g2034 ( 
.A1(n_1988),
.A2(n_1942),
.B1(n_1967),
.B2(n_1938),
.C(n_1965),
.Y(n_2034)
);

AOI22xp33_ASAP7_75t_SL g2035 ( 
.A1(n_1990),
.A2(n_1969),
.B1(n_1963),
.B2(n_1874),
.Y(n_2035)
);

OAI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_1985),
.A2(n_1904),
.B1(n_1923),
.B2(n_1878),
.Y(n_2036)
);

OAI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1985),
.A2(n_1878),
.B1(n_1937),
.B2(n_1882),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_2014),
.Y(n_2038)
);

OAI221xp5_ASAP7_75t_L g2039 ( 
.A1(n_1998),
.A2(n_1867),
.B1(n_1961),
.B2(n_1951),
.C(n_1970),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1978),
.Y(n_2040)
);

CKINVDCx5p33_ASAP7_75t_R g2041 ( 
.A(n_2000),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1978),
.Y(n_2042)
);

AND2x4_ASAP7_75t_L g2043 ( 
.A(n_2028),
.B(n_1916),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1974),
.B(n_1941),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1989),
.B(n_1930),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1980),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1980),
.Y(n_2047)
);

OAI21x1_ASAP7_75t_L g2048 ( 
.A1(n_1976),
.A2(n_1740),
.B(n_1850),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_SL g2049 ( 
.A(n_2020),
.B(n_1915),
.Y(n_2049)
);

AOI221xp5_ASAP7_75t_L g2050 ( 
.A1(n_1988),
.A2(n_1895),
.B1(n_1955),
.B2(n_1927),
.C(n_1947),
.Y(n_2050)
);

A2O1A1Ixp33_ASAP7_75t_L g2051 ( 
.A1(n_2020),
.A2(n_1861),
.B(n_1926),
.C(n_1918),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_2004),
.Y(n_2052)
);

AOI21xp5_ASAP7_75t_L g2053 ( 
.A1(n_1993),
.A2(n_1881),
.B(n_1884),
.Y(n_2053)
);

AND2x2_ASAP7_75t_SL g2054 ( 
.A(n_2010),
.B(n_1881),
.Y(n_2054)
);

INVx3_ASAP7_75t_L g2055 ( 
.A(n_1994),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_2013),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2026),
.B(n_1755),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1989),
.B(n_1932),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2009),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2026),
.B(n_1872),
.Y(n_2060)
);

BUFx2_ASAP7_75t_SL g2061 ( 
.A(n_2007),
.Y(n_2061)
);

OAI21x1_ASAP7_75t_L g2062 ( 
.A1(n_1991),
.A2(n_1791),
.B(n_1905),
.Y(n_2062)
);

AOI22xp5_ASAP7_75t_L g2063 ( 
.A1(n_1973),
.A2(n_1918),
.B1(n_1886),
.B2(n_1872),
.Y(n_2063)
);

AOI222xp33_ASAP7_75t_L g2064 ( 
.A1(n_1990),
.A2(n_1748),
.B1(n_1886),
.B2(n_1879),
.C1(n_1953),
.C2(n_1964),
.Y(n_2064)
);

OR2x6_ASAP7_75t_L g2065 ( 
.A(n_1984),
.B(n_1909),
.Y(n_2065)
);

OAI22xp5_ASAP7_75t_L g2066 ( 
.A1(n_1996),
.A2(n_1879),
.B1(n_1957),
.B2(n_1908),
.Y(n_2066)
);

INVx3_ASAP7_75t_L g2067 ( 
.A(n_1994),
.Y(n_2067)
);

NOR2xp33_ASAP7_75t_L g2068 ( 
.A(n_2030),
.B(n_1892),
.Y(n_2068)
);

INVx3_ASAP7_75t_L g2069 ( 
.A(n_2040),
.Y(n_2069)
);

INVxp67_ASAP7_75t_SL g2070 ( 
.A(n_2057),
.Y(n_2070)
);

HB1xp67_ASAP7_75t_L g2071 ( 
.A(n_2056),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2042),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2046),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2047),
.Y(n_2074)
);

BUFx3_ASAP7_75t_L g2075 ( 
.A(n_2065),
.Y(n_2075)
);

NOR2x1_ASAP7_75t_L g2076 ( 
.A(n_2065),
.B(n_2024),
.Y(n_2076)
);

NAND2x1p5_ASAP7_75t_L g2077 ( 
.A(n_2053),
.B(n_2010),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2043),
.B(n_2029),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_2052),
.Y(n_2079)
);

OAI21x1_ASAP7_75t_L g2080 ( 
.A1(n_2048),
.A2(n_1997),
.B(n_1999),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2059),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2060),
.Y(n_2082)
);

INVx3_ASAP7_75t_L g2083 ( 
.A(n_2065),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_2054),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2055),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_2032),
.Y(n_2086)
);

HB1xp67_ASAP7_75t_L g2087 ( 
.A(n_2043),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2044),
.B(n_2011),
.Y(n_2088)
);

INVxp67_ASAP7_75t_L g2089 ( 
.A(n_2049),
.Y(n_2089)
);

HB1xp67_ASAP7_75t_L g2090 ( 
.A(n_2055),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_2032),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_2084),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2084),
.B(n_2067),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_2089),
.A2(n_2035),
.B1(n_2017),
.B2(n_2049),
.Y(n_2094)
);

AOI22xp33_ASAP7_75t_L g2095 ( 
.A1(n_2089),
.A2(n_2066),
.B1(n_1984),
.B2(n_2027),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_2072),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2082),
.B(n_2024),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2082),
.B(n_2070),
.Y(n_2098)
);

HB1xp67_ASAP7_75t_L g2099 ( 
.A(n_2069),
.Y(n_2099)
);

AO21x2_ASAP7_75t_L g2100 ( 
.A1(n_2080),
.A2(n_2037),
.B(n_1986),
.Y(n_2100)
);

OAI22xp33_ASAP7_75t_L g2101 ( 
.A1(n_2077),
.A2(n_2066),
.B1(n_2033),
.B2(n_2039),
.Y(n_2101)
);

NAND3xp33_ASAP7_75t_L g2102 ( 
.A(n_2076),
.B(n_2050),
.C(n_2034),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2096),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_2098),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2102),
.B(n_2088),
.Y(n_2105)
);

BUFx6f_ASAP7_75t_L g2106 ( 
.A(n_2092),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2099),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_L g2108 ( 
.A(n_2101),
.B(n_2041),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2106),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2105),
.B(n_2094),
.Y(n_2110)
);

INVx2_ASAP7_75t_L g2111 ( 
.A(n_2106),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2103),
.Y(n_2112)
);

AO21x2_ASAP7_75t_L g2113 ( 
.A1(n_2107),
.A2(n_2101),
.B(n_2099),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2104),
.B(n_2093),
.Y(n_2114)
);

NAND3xp33_ASAP7_75t_L g2115 ( 
.A(n_2108),
.B(n_1998),
.C(n_1996),
.Y(n_2115)
);

OAI31xp33_ASAP7_75t_L g2116 ( 
.A1(n_2108),
.A2(n_2036),
.A3(n_2077),
.B(n_2075),
.Y(n_2116)
);

AOI221xp5_ASAP7_75t_L g2117 ( 
.A1(n_2105),
.A2(n_2095),
.B1(n_2068),
.B2(n_2100),
.C(n_1992),
.Y(n_2117)
);

NAND4xp75_ASAP7_75t_L g2118 ( 
.A(n_2117),
.B(n_2076),
.C(n_2027),
.D(n_1993),
.Y(n_2118)
);

NAND3xp33_ASAP7_75t_L g2119 ( 
.A(n_2115),
.B(n_2022),
.C(n_2013),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2109),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2111),
.Y(n_2121)
);

INVx3_ASAP7_75t_L g2122 ( 
.A(n_2113),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_2114),
.B(n_2113),
.Y(n_2123)
);

OA211x2_ASAP7_75t_L g2124 ( 
.A1(n_2116),
.A2(n_2031),
.B(n_2002),
.C(n_2000),
.Y(n_2124)
);

NAND4xp75_ASAP7_75t_L g2125 ( 
.A(n_2110),
.B(n_2091),
.C(n_2086),
.D(n_2063),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2115),
.B(n_2097),
.Y(n_2126)
);

NAND4xp75_ASAP7_75t_L g2127 ( 
.A(n_2112),
.B(n_2086),
.C(n_2091),
.D(n_2045),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_2110),
.B(n_2088),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2120),
.Y(n_2129)
);

BUFx2_ASAP7_75t_L g2130 ( 
.A(n_2123),
.Y(n_2130)
);

AOI222xp33_ASAP7_75t_L g2131 ( 
.A1(n_2122),
.A2(n_2022),
.B1(n_2075),
.B2(n_2083),
.C1(n_2003),
.C2(n_2032),
.Y(n_2131)
);

OAI222xp33_ASAP7_75t_L g2132 ( 
.A1(n_2126),
.A2(n_2077),
.B1(n_2083),
.B2(n_2091),
.C1(n_2086),
.C2(n_2075),
.Y(n_2132)
);

BUFx3_ASAP7_75t_L g2133 ( 
.A(n_2121),
.Y(n_2133)
);

NAND3xp33_ASAP7_75t_L g2134 ( 
.A(n_2119),
.B(n_1995),
.C(n_2051),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2128),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2127),
.B(n_2061),
.Y(n_2136)
);

AOI22xp5_ASAP7_75t_L g2137 ( 
.A1(n_2118),
.A2(n_2124),
.B1(n_2125),
.B2(n_2100),
.Y(n_2137)
);

NAND2x1_ASAP7_75t_L g2138 ( 
.A(n_2136),
.B(n_2083),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2130),
.Y(n_2139)
);

HB1xp67_ASAP7_75t_L g2140 ( 
.A(n_2133),
.Y(n_2140)
);

NOR2x1_ASAP7_75t_L g2141 ( 
.A(n_2133),
.B(n_2118),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2140),
.B(n_2129),
.Y(n_2142)
);

NOR4xp25_ASAP7_75t_SL g2143 ( 
.A(n_2139),
.B(n_2141),
.C(n_2135),
.D(n_2132),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2138),
.Y(n_2144)
);

NAND4xp25_ASAP7_75t_SL g2145 ( 
.A(n_2141),
.B(n_2137),
.C(n_2131),
.D(n_2134),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_2143),
.B(n_2038),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2144),
.B(n_2132),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2142),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2145),
.Y(n_2149)
);

INVx1_ASAP7_75t_SL g2150 ( 
.A(n_2142),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2142),
.Y(n_2151)
);

OAI211xp5_ASAP7_75t_L g2152 ( 
.A1(n_2146),
.A2(n_1900),
.B(n_2083),
.C(n_1830),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_2147),
.Y(n_2153)
);

OAI21xp5_ASAP7_75t_SL g2154 ( 
.A1(n_2149),
.A2(n_2064),
.B(n_2001),
.Y(n_2154)
);

OAI21xp33_ASAP7_75t_L g2155 ( 
.A1(n_2147),
.A2(n_2001),
.B(n_2005),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2148),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_2150),
.B(n_2071),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_2151),
.B(n_2015),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2147),
.Y(n_2159)
);

INVx1_ASAP7_75t_SL g2160 ( 
.A(n_2147),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2147),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_2153),
.B(n_2087),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2161),
.B(n_2078),
.Y(n_2163)
);

CKINVDCx16_ASAP7_75t_R g2164 ( 
.A(n_2160),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2159),
.B(n_2078),
.Y(n_2165)
);

XOR2x2_ASAP7_75t_L g2166 ( 
.A(n_2158),
.B(n_110),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2157),
.B(n_2090),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2156),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_2152),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2154),
.B(n_2079),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2155),
.Y(n_2171)
);

NAND2xp33_ASAP7_75t_SL g2172 ( 
.A(n_2153),
.B(n_1894),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2153),
.Y(n_2173)
);

O2A1O1Ixp33_ASAP7_75t_L g2174 ( 
.A1(n_2160),
.A2(n_113),
.B(n_111),
.C(n_112),
.Y(n_2174)
);

OAI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2164),
.A2(n_2085),
.B1(n_2067),
.B2(n_2069),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2173),
.Y(n_2176)
);

NOR4xp25_ASAP7_75t_SL g2177 ( 
.A(n_2172),
.B(n_2085),
.C(n_115),
.D(n_112),
.Y(n_2177)
);

INVx2_ASAP7_75t_SL g2178 ( 
.A(n_2162),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2165),
.Y(n_2179)
);

INVx3_ASAP7_75t_L g2180 ( 
.A(n_2163),
.Y(n_2180)
);

XNOR2xp5_ASAP7_75t_L g2181 ( 
.A(n_2166),
.B(n_114),
.Y(n_2181)
);

BUFx4f_ASAP7_75t_SL g2182 ( 
.A(n_2168),
.Y(n_2182)
);

CKINVDCx16_ASAP7_75t_R g2183 ( 
.A(n_2172),
.Y(n_2183)
);

AOI33xp33_ASAP7_75t_L g2184 ( 
.A1(n_2169),
.A2(n_2005),
.A3(n_1946),
.B1(n_1964),
.B2(n_1953),
.B3(n_1987),
.Y(n_2184)
);

OAI211xp5_ASAP7_75t_L g2185 ( 
.A1(n_2174),
.A2(n_1898),
.B(n_1894),
.C(n_2064),
.Y(n_2185)
);

INVx2_ASAP7_75t_SL g2186 ( 
.A(n_2167),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2171),
.B(n_2058),
.Y(n_2187)
);

AOI21xp33_ASAP7_75t_SL g2188 ( 
.A1(n_2174),
.A2(n_2170),
.B(n_114),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_2164),
.Y(n_2189)
);

NOR3xp33_ASAP7_75t_L g2190 ( 
.A(n_2189),
.B(n_1832),
.C(n_1975),
.Y(n_2190)
);

OAI222xp33_ASAP7_75t_L g2191 ( 
.A1(n_2182),
.A2(n_2069),
.B1(n_1999),
.B2(n_2074),
.C1(n_2073),
.C2(n_2072),
.Y(n_2191)
);

NOR3x1_ASAP7_75t_L g2192 ( 
.A(n_2186),
.B(n_115),
.C(n_116),
.Y(n_2192)
);

NOR2xp67_ASAP7_75t_L g2193 ( 
.A(n_2180),
.B(n_116),
.Y(n_2193)
);

NAND2xp5_ASAP7_75t_L g2194 ( 
.A(n_2180),
.B(n_2069),
.Y(n_2194)
);

NOR2xp33_ASAP7_75t_L g2195 ( 
.A(n_2188),
.B(n_2178),
.Y(n_2195)
);

NAND2xp33_ASAP7_75t_SL g2196 ( 
.A(n_2177),
.B(n_2181),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2183),
.B(n_2073),
.Y(n_2197)
);

OAI22xp5_ASAP7_75t_L g2198 ( 
.A1(n_2176),
.A2(n_1898),
.B1(n_1957),
.B2(n_2074),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2187),
.Y(n_2199)
);

NOR2xp67_ASAP7_75t_L g2200 ( 
.A(n_2179),
.B(n_117),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2184),
.Y(n_2201)
);

NOR2xp33_ASAP7_75t_L g2202 ( 
.A(n_2185),
.B(n_117),
.Y(n_2202)
);

AOI211xp5_ASAP7_75t_L g2203 ( 
.A1(n_2175),
.A2(n_120),
.B(n_118),
.C(n_119),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2193),
.Y(n_2204)
);

HB1xp67_ASAP7_75t_L g2205 ( 
.A(n_2200),
.Y(n_2205)
);

NOR2x1_ASAP7_75t_L g2206 ( 
.A(n_2195),
.B(n_118),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2199),
.B(n_119),
.Y(n_2207)
);

AOI22xp33_ASAP7_75t_L g2208 ( 
.A1(n_2196),
.A2(n_1982),
.B1(n_1943),
.B2(n_1954),
.Y(n_2208)
);

INVxp33_ASAP7_75t_SL g2209 ( 
.A(n_2192),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2202),
.B(n_120),
.Y(n_2210)
);

AOI21xp5_ASAP7_75t_L g2211 ( 
.A1(n_2197),
.A2(n_2018),
.B(n_121),
.Y(n_2211)
);

OAI211xp5_ASAP7_75t_L g2212 ( 
.A1(n_2203),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_2212)
);

NOR2x1_ASAP7_75t_L g2213 ( 
.A(n_2194),
.B(n_124),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2201),
.Y(n_2214)
);

AOI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2198),
.A2(n_1943),
.B1(n_1954),
.B2(n_1913),
.Y(n_2215)
);

NAND2xp5_ASAP7_75t_L g2216 ( 
.A(n_2190),
.B(n_124),
.Y(n_2216)
);

O2A1O1Ixp5_ASAP7_75t_L g2217 ( 
.A1(n_2191),
.A2(n_1939),
.B(n_128),
.C(n_126),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_2193),
.Y(n_2218)
);

NAND3xp33_ASAP7_75t_L g2219 ( 
.A(n_2203),
.B(n_126),
.C(n_127),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2193),
.B(n_127),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_2196),
.A2(n_128),
.B(n_129),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2193),
.B(n_130),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2193),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2193),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_2196),
.A2(n_1982),
.B1(n_2019),
.B2(n_2079),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2205),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2220),
.Y(n_2227)
);

NAND3xp33_ASAP7_75t_L g2228 ( 
.A(n_2221),
.B(n_131),
.C(n_132),
.Y(n_2228)
);

NOR3xp33_ASAP7_75t_L g2229 ( 
.A(n_2214),
.B(n_131),
.C(n_133),
.Y(n_2229)
);

HB1xp67_ASAP7_75t_L g2230 ( 
.A(n_2213),
.Y(n_2230)
);

AOI221xp5_ASAP7_75t_L g2231 ( 
.A1(n_2209),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.C(n_137),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2222),
.Y(n_2232)
);

AOI22xp5_ASAP7_75t_L g2233 ( 
.A1(n_2225),
.A2(n_1982),
.B1(n_2019),
.B2(n_2081),
.Y(n_2233)
);

AOI22xp5_ASAP7_75t_L g2234 ( 
.A1(n_2212),
.A2(n_1982),
.B1(n_2081),
.B2(n_1912),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2207),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_2204),
.B(n_2218),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2223),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_SL g2238 ( 
.A(n_2224),
.B(n_1912),
.Y(n_2238)
);

NOR2x1_ASAP7_75t_L g2239 ( 
.A(n_2206),
.B(n_134),
.Y(n_2239)
);

AO22x2_ASAP7_75t_L g2240 ( 
.A1(n_2219),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.Y(n_2240)
);

AOI221xp5_ASAP7_75t_L g2241 ( 
.A1(n_2217),
.A2(n_138),
.B1(n_139),
.B2(n_140),
.C(n_141),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_SL g2242 ( 
.A(n_2208),
.B(n_2080),
.Y(n_2242)
);

AOI22xp33_ASAP7_75t_L g2243 ( 
.A1(n_2210),
.A2(n_2080),
.B1(n_2021),
.B2(n_1977),
.Y(n_2243)
);

INVxp67_ASAP7_75t_L g2244 ( 
.A(n_2216),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2211),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2215),
.Y(n_2246)
);

AOI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2209),
.A2(n_1981),
.B1(n_2012),
.B2(n_2016),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2205),
.Y(n_2248)
);

OAI22xp5_ASAP7_75t_L g2249 ( 
.A1(n_2208),
.A2(n_2023),
.B1(n_1979),
.B2(n_142),
.Y(n_2249)
);

NOR4xp25_ASAP7_75t_L g2250 ( 
.A(n_2214),
.B(n_143),
.C(n_139),
.D(n_140),
.Y(n_2250)
);

AO22x2_ASAP7_75t_L g2251 ( 
.A1(n_2204),
.A2(n_145),
.B1(n_143),
.B2(n_144),
.Y(n_2251)
);

AO22x2_ASAP7_75t_L g2252 ( 
.A1(n_2204),
.A2(n_147),
.B1(n_144),
.B2(n_146),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2205),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2205),
.Y(n_2254)
);

OAI31xp33_ASAP7_75t_L g2255 ( 
.A1(n_2212),
.A2(n_148),
.A3(n_146),
.B(n_147),
.Y(n_2255)
);

AOI22xp5_ASAP7_75t_L g2256 ( 
.A1(n_2209),
.A2(n_2025),
.B1(n_1723),
.B2(n_2062),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2205),
.Y(n_2257)
);

OA22x2_ASAP7_75t_L g2258 ( 
.A1(n_2225),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2258)
);

AOI31xp33_ASAP7_75t_L g2259 ( 
.A1(n_2205),
.A2(n_152),
.A3(n_150),
.B(n_151),
.Y(n_2259)
);

NOR4xp25_ASAP7_75t_L g2260 ( 
.A(n_2214),
.B(n_154),
.C(n_152),
.D(n_153),
.Y(n_2260)
);

OAI22xp33_ASAP7_75t_SL g2261 ( 
.A1(n_2226),
.A2(n_158),
.B1(n_155),
.B2(n_156),
.Y(n_2261)
);

XNOR2xp5_ASAP7_75t_L g2262 ( 
.A(n_2240),
.B(n_155),
.Y(n_2262)
);

BUFx6f_ASAP7_75t_L g2263 ( 
.A(n_2248),
.Y(n_2263)
);

OAI21xp33_ASAP7_75t_SL g2264 ( 
.A1(n_2239),
.A2(n_156),
.B(n_158),
.Y(n_2264)
);

NOR3x1_ASAP7_75t_L g2265 ( 
.A(n_2228),
.B(n_160),
.C(n_161),
.Y(n_2265)
);

AOI22x1_ASAP7_75t_L g2266 ( 
.A1(n_2230),
.A2(n_164),
.B1(n_160),
.B2(n_162),
.Y(n_2266)
);

CKINVDCx12_ASAP7_75t_R g2267 ( 
.A(n_2259),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2251),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2260),
.B(n_162),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2252),
.Y(n_2270)
);

AND2x2_ASAP7_75t_L g2271 ( 
.A(n_2253),
.B(n_165),
.Y(n_2271)
);

AOI321xp33_ASAP7_75t_L g2272 ( 
.A1(n_2254),
.A2(n_165),
.A3(n_166),
.B1(n_167),
.B2(n_168),
.C(n_169),
.Y(n_2272)
);

NOR3xp33_ASAP7_75t_L g2273 ( 
.A(n_2236),
.B(n_167),
.C(n_170),
.Y(n_2273)
);

INVx1_ASAP7_75t_SL g2274 ( 
.A(n_2258),
.Y(n_2274)
);

A2O1A1Ixp33_ASAP7_75t_L g2275 ( 
.A1(n_2255),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_2257),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2237),
.Y(n_2277)
);

AOI21xp33_ASAP7_75t_SL g2278 ( 
.A1(n_2250),
.A2(n_173),
.B(n_174),
.Y(n_2278)
);

OA21x2_ASAP7_75t_L g2279 ( 
.A1(n_2227),
.A2(n_174),
.B(n_175),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2229),
.B(n_175),
.Y(n_2280)
);

CKINVDCx6p67_ASAP7_75t_R g2281 ( 
.A(n_2235),
.Y(n_2281)
);

NAND3xp33_ASAP7_75t_SL g2282 ( 
.A(n_2241),
.B(n_176),
.C(n_177),
.Y(n_2282)
);

OAI32xp33_ASAP7_75t_L g2283 ( 
.A1(n_2245),
.A2(n_177),
.A3(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2238),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_2232),
.Y(n_2285)
);

NAND4xp25_ASAP7_75t_SL g2286 ( 
.A(n_2233),
.B(n_182),
.C(n_179),
.D(n_181),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2234),
.A2(n_2246),
.B1(n_2244),
.B2(n_2247),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_R g2288 ( 
.A(n_2231),
.B(n_181),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2242),
.Y(n_2289)
);

NOR3xp33_ASAP7_75t_L g2290 ( 
.A(n_2276),
.B(n_2277),
.C(n_2287),
.Y(n_2290)
);

INVx3_ASAP7_75t_L g2291 ( 
.A(n_2279),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2279),
.Y(n_2292)
);

XNOR2xp5_ASAP7_75t_L g2293 ( 
.A(n_2262),
.B(n_2274),
.Y(n_2293)
);

INVxp67_ASAP7_75t_SL g2294 ( 
.A(n_2269),
.Y(n_2294)
);

XNOR2xp5_ASAP7_75t_L g2295 ( 
.A(n_2266),
.B(n_2249),
.Y(n_2295)
);

NAND2x1p5_ASAP7_75t_L g2296 ( 
.A(n_2263),
.B(n_2256),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2271),
.Y(n_2297)
);

NOR2x1p5_ASAP7_75t_L g2298 ( 
.A(n_2281),
.B(n_2243),
.Y(n_2298)
);

AND4x1_ASAP7_75t_L g2299 ( 
.A(n_2265),
.B(n_2273),
.C(n_2268),
.D(n_2270),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2267),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2263),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2278),
.B(n_182),
.Y(n_2302)
);

HB1xp67_ASAP7_75t_L g2303 ( 
.A(n_2264),
.Y(n_2303)
);

HB1xp67_ASAP7_75t_L g2304 ( 
.A(n_2261),
.Y(n_2304)
);

NOR2x1_ASAP7_75t_L g2305 ( 
.A(n_2280),
.B(n_183),
.Y(n_2305)
);

AND2x2_ASAP7_75t_L g2306 ( 
.A(n_2284),
.B(n_184),
.Y(n_2306)
);

AND2x2_ASAP7_75t_SL g2307 ( 
.A(n_2285),
.B(n_185),
.Y(n_2307)
);

OAI221xp5_ASAP7_75t_SL g2308 ( 
.A1(n_2275),
.A2(n_185),
.B1(n_186),
.B2(n_189),
.C(n_190),
.Y(n_2308)
);

INVx1_ASAP7_75t_SL g2309 ( 
.A(n_2288),
.Y(n_2309)
);

NOR2x1_ASAP7_75t_L g2310 ( 
.A(n_2282),
.B(n_2286),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2289),
.Y(n_2311)
);

NAND4xp75_ASAP7_75t_L g2312 ( 
.A(n_2283),
.B(n_186),
.C(n_190),
.D(n_191),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_2272),
.B(n_191),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_2271),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_2279),
.Y(n_2315)
);

NOR2x1_ASAP7_75t_L g2316 ( 
.A(n_2279),
.B(n_192),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_2271),
.Y(n_2317)
);

NOR2xp67_ASAP7_75t_L g2318 ( 
.A(n_2264),
.B(n_194),
.Y(n_2318)
);

NOR2xp33_ASAP7_75t_SL g2319 ( 
.A(n_2274),
.B(n_194),
.Y(n_2319)
);

NOR2x1_ASAP7_75t_L g2320 ( 
.A(n_2279),
.B(n_195),
.Y(n_2320)
);

NAND4xp75_ASAP7_75t_L g2321 ( 
.A(n_2265),
.B(n_195),
.C(n_196),
.D(n_197),
.Y(n_2321)
);

NOR3xp33_ASAP7_75t_L g2322 ( 
.A(n_2276),
.B(n_197),
.C(n_198),
.Y(n_2322)
);

NAND4xp75_ASAP7_75t_L g2323 ( 
.A(n_2265),
.B(n_200),
.C(n_201),
.D(n_202),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2271),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2264),
.B(n_202),
.Y(n_2325)
);

OAI211xp5_ASAP7_75t_L g2326 ( 
.A1(n_2264),
.A2(n_203),
.B(n_204),
.C(n_206),
.Y(n_2326)
);

NOR2xp67_ASAP7_75t_L g2327 ( 
.A(n_2291),
.B(n_203),
.Y(n_2327)
);

OAI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2326),
.A2(n_206),
.B(n_207),
.C(n_208),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_L g2329 ( 
.A(n_2307),
.B(n_207),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_2291),
.Y(n_2330)
);

OAI21xp33_ASAP7_75t_SL g2331 ( 
.A1(n_2316),
.A2(n_208),
.B(n_209),
.Y(n_2331)
);

AOI22xp33_ASAP7_75t_SL g2332 ( 
.A1(n_2319),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_2332)
);

OAI211xp5_ASAP7_75t_SL g2333 ( 
.A1(n_2300),
.A2(n_210),
.B(n_211),
.C(n_212),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2292),
.Y(n_2334)
);

XNOR2xp5_ASAP7_75t_L g2335 ( 
.A(n_2293),
.B(n_213),
.Y(n_2335)
);

XNOR2x1_ASAP7_75t_L g2336 ( 
.A(n_2321),
.B(n_2323),
.Y(n_2336)
);

AOI211xp5_ASAP7_75t_L g2337 ( 
.A1(n_2308),
.A2(n_213),
.B(n_214),
.C(n_215),
.Y(n_2337)
);

OAI322xp33_ASAP7_75t_L g2338 ( 
.A1(n_2301),
.A2(n_216),
.A3(n_217),
.B1(n_218),
.B2(n_219),
.C1(n_220),
.C2(n_221),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_2306),
.B(n_218),
.Y(n_2339)
);

AOI221xp5_ASAP7_75t_L g2340 ( 
.A1(n_2290),
.A2(n_219),
.B1(n_220),
.B2(n_222),
.C(n_223),
.Y(n_2340)
);

AOI221xp5_ASAP7_75t_L g2341 ( 
.A1(n_2313),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.C(n_226),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2303),
.B(n_224),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2315),
.Y(n_2343)
);

AND4x1_ASAP7_75t_L g2344 ( 
.A(n_2320),
.B(n_225),
.C(n_226),
.D(n_227),
.Y(n_2344)
);

OR3x2_ASAP7_75t_L g2345 ( 
.A(n_2297),
.B(n_227),
.C(n_228),
.Y(n_2345)
);

O2A1O1Ixp33_ASAP7_75t_L g2346 ( 
.A1(n_2302),
.A2(n_229),
.B(n_230),
.C(n_231),
.Y(n_2346)
);

NAND2x1_ASAP7_75t_L g2347 ( 
.A(n_2318),
.B(n_229),
.Y(n_2347)
);

AOI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2325),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_2348)
);

NOR3x2_ASAP7_75t_L g2349 ( 
.A(n_2312),
.B(n_232),
.C(n_233),
.Y(n_2349)
);

OAI221xp5_ASAP7_75t_L g2350 ( 
.A1(n_2299),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.C(n_237),
.Y(n_2350)
);

OAI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_2311),
.A2(n_2304),
.B1(n_2324),
.B2(n_2317),
.Y(n_2351)
);

AOI221xp5_ASAP7_75t_L g2352 ( 
.A1(n_2294),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.C(n_238),
.Y(n_2352)
);

HB1xp67_ASAP7_75t_L g2353 ( 
.A(n_2305),
.Y(n_2353)
);

AOI221xp5_ASAP7_75t_SL g2354 ( 
.A1(n_2309),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.C(n_241),
.Y(n_2354)
);

OR3x2_ASAP7_75t_L g2355 ( 
.A(n_2314),
.B(n_240),
.C(n_242),
.Y(n_2355)
);

AOI22xp5_ASAP7_75t_L g2356 ( 
.A1(n_2298),
.A2(n_2310),
.B1(n_2295),
.B2(n_2322),
.Y(n_2356)
);

OAI221xp5_ASAP7_75t_L g2357 ( 
.A1(n_2296),
.A2(n_242),
.B1(n_243),
.B2(n_244),
.C(n_245),
.Y(n_2357)
);

AOI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2290),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_2358)
);

AND2x4_ASAP7_75t_L g2359 ( 
.A(n_2327),
.B(n_246),
.Y(n_2359)
);

AOI22xp5_ASAP7_75t_L g2360 ( 
.A1(n_2351),
.A2(n_247),
.B1(n_248),
.B2(n_249),
.Y(n_2360)
);

XNOR2x1_ASAP7_75t_L g2361 ( 
.A(n_2335),
.B(n_247),
.Y(n_2361)
);

NOR3xp33_ASAP7_75t_L g2362 ( 
.A(n_2350),
.B(n_2347),
.C(n_2341),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2342),
.Y(n_2363)
);

HB1xp67_ASAP7_75t_L g2364 ( 
.A(n_2344),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2332),
.B(n_249),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2345),
.Y(n_2366)
);

AND2x2_ASAP7_75t_SL g2367 ( 
.A(n_2339),
.B(n_250),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2355),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2329),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2349),
.Y(n_2370)
);

OAI22xp5_ASAP7_75t_L g2371 ( 
.A1(n_2356),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_2371)
);

NAND4xp75_ASAP7_75t_L g2372 ( 
.A(n_2331),
.B(n_253),
.C(n_254),
.D(n_256),
.Y(n_2372)
);

INVx2_ASAP7_75t_L g2373 ( 
.A(n_2330),
.Y(n_2373)
);

OA22x2_ASAP7_75t_L g2374 ( 
.A1(n_2348),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_2374)
);

AND4x1_ASAP7_75t_L g2375 ( 
.A(n_2337),
.B(n_257),
.C(n_258),
.D(n_259),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2334),
.B(n_257),
.Y(n_2376)
);

XNOR2x1_ASAP7_75t_L g2377 ( 
.A(n_2336),
.B(n_258),
.Y(n_2377)
);

HB1xp67_ASAP7_75t_L g2378 ( 
.A(n_2353),
.Y(n_2378)
);

INVx1_ASAP7_75t_L g2379 ( 
.A(n_2343),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2328),
.B(n_2333),
.Y(n_2380)
);

XNOR2xp5_ASAP7_75t_L g2381 ( 
.A(n_2358),
.B(n_259),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_L g2382 ( 
.A(n_2354),
.B(n_260),
.Y(n_2382)
);

INVx2_ASAP7_75t_SL g2383 ( 
.A(n_2357),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2338),
.Y(n_2384)
);

AO21x2_ASAP7_75t_L g2385 ( 
.A1(n_2346),
.A2(n_260),
.B(n_261),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2340),
.Y(n_2386)
);

INVx2_ASAP7_75t_SL g2387 ( 
.A(n_2352),
.Y(n_2387)
);

XNOR2x1_ASAP7_75t_L g2388 ( 
.A(n_2335),
.B(n_261),
.Y(n_2388)
);

NOR3xp33_ASAP7_75t_L g2389 ( 
.A(n_2351),
.B(n_262),
.C(n_263),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2327),
.B(n_262),
.Y(n_2390)
);

OA22x2_ASAP7_75t_L g2391 ( 
.A1(n_2360),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_2363),
.Y(n_2392)
);

OAI221xp5_ASAP7_75t_L g2393 ( 
.A1(n_2389),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.C(n_267),
.Y(n_2393)
);

NAND3xp33_ASAP7_75t_SL g2394 ( 
.A(n_2390),
.B(n_267),
.C(n_268),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2359),
.Y(n_2395)
);

AND2x4_ASAP7_75t_L g2396 ( 
.A(n_2373),
.B(n_269),
.Y(n_2396)
);

NAND4xp25_ASAP7_75t_L g2397 ( 
.A(n_2380),
.B(n_269),
.C(n_270),
.D(n_271),
.Y(n_2397)
);

AOI22xp5_ASAP7_75t_L g2398 ( 
.A1(n_2379),
.A2(n_270),
.B1(n_271),
.B2(n_272),
.Y(n_2398)
);

CKINVDCx5p33_ASAP7_75t_R g2399 ( 
.A(n_2378),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2377),
.Y(n_2400)
);

HB1xp67_ASAP7_75t_L g2401 ( 
.A(n_2372),
.Y(n_2401)
);

CKINVDCx5p33_ASAP7_75t_R g2402 ( 
.A(n_2364),
.Y(n_2402)
);

CKINVDCx5p33_ASAP7_75t_R g2403 ( 
.A(n_2370),
.Y(n_2403)
);

OAI21xp33_ASAP7_75t_SL g2404 ( 
.A1(n_2382),
.A2(n_2365),
.B(n_2361),
.Y(n_2404)
);

HB1xp67_ASAP7_75t_L g2405 ( 
.A(n_2376),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2374),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2367),
.Y(n_2407)
);

AOI22xp33_ASAP7_75t_L g2408 ( 
.A1(n_2399),
.A2(n_2384),
.B1(n_2362),
.B2(n_2368),
.Y(n_2408)
);

INVxp67_ASAP7_75t_L g2409 ( 
.A(n_2393),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_2394),
.B(n_2385),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2391),
.Y(n_2411)
);

NOR2x1_ASAP7_75t_L g2412 ( 
.A(n_2407),
.B(n_2388),
.Y(n_2412)
);

OAI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2402),
.A2(n_2366),
.B1(n_2381),
.B2(n_2386),
.Y(n_2413)
);

OAI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2392),
.A2(n_2381),
.B1(n_2387),
.B2(n_2383),
.Y(n_2414)
);

AOI21xp5_ASAP7_75t_L g2415 ( 
.A1(n_2405),
.A2(n_2369),
.B(n_2371),
.Y(n_2415)
);

AOI22x1_ASAP7_75t_L g2416 ( 
.A1(n_2403),
.A2(n_2375),
.B1(n_272),
.B2(n_419),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2406),
.B(n_1979),
.Y(n_2417)
);

BUFx2_ASAP7_75t_L g2418 ( 
.A(n_2397),
.Y(n_2418)
);

INVx1_ASAP7_75t_SL g2419 ( 
.A(n_2396),
.Y(n_2419)
);

OA22x2_ASAP7_75t_L g2420 ( 
.A1(n_2395),
.A2(n_2008),
.B1(n_1983),
.B2(n_2006),
.Y(n_2420)
);

AND3x2_ASAP7_75t_L g2421 ( 
.A(n_2401),
.B(n_417),
.C(n_421),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2396),
.Y(n_2422)
);

OR2x2_ASAP7_75t_L g2423 ( 
.A(n_2410),
.B(n_2400),
.Y(n_2423)
);

AOI22xp33_ASAP7_75t_L g2424 ( 
.A1(n_2416),
.A2(n_2404),
.B1(n_2398),
.B2(n_1986),
.Y(n_2424)
);

NOR3xp33_ASAP7_75t_L g2425 ( 
.A(n_2413),
.B(n_423),
.C(n_428),
.Y(n_2425)
);

NAND3x1_ASAP7_75t_L g2426 ( 
.A(n_2412),
.B(n_429),
.C(n_430),
.Y(n_2426)
);

NAND3xp33_ASAP7_75t_SL g2427 ( 
.A(n_2419),
.B(n_432),
.C(n_434),
.Y(n_2427)
);

OR3x1_ASAP7_75t_L g2428 ( 
.A(n_2422),
.B(n_435),
.C(n_437),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2421),
.Y(n_2429)
);

OAI211xp5_ASAP7_75t_SL g2430 ( 
.A1(n_2408),
.A2(n_438),
.B(n_440),
.C(n_441),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2429),
.B(n_2411),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2428),
.B(n_2415),
.Y(n_2432)
);

INVxp33_ASAP7_75t_L g2433 ( 
.A(n_2425),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2432),
.Y(n_2434)
);

NAND2x1p5_ASAP7_75t_L g2435 ( 
.A(n_2431),
.B(n_2423),
.Y(n_2435)
);

CKINVDCx20_ASAP7_75t_R g2436 ( 
.A(n_2433),
.Y(n_2436)
);

AOI221xp5_ASAP7_75t_L g2437 ( 
.A1(n_2434),
.A2(n_2414),
.B1(n_2409),
.B2(n_2430),
.C(n_2424),
.Y(n_2437)
);

OAI221xp5_ASAP7_75t_L g2438 ( 
.A1(n_2435),
.A2(n_2418),
.B1(n_2427),
.B2(n_2417),
.C(n_2426),
.Y(n_2438)
);

OAI21xp5_ASAP7_75t_L g2439 ( 
.A1(n_2436),
.A2(n_2420),
.B(n_445),
.Y(n_2439)
);

XNOR2xp5_ASAP7_75t_L g2440 ( 
.A(n_2435),
.B(n_443),
.Y(n_2440)
);

INVxp67_ASAP7_75t_SL g2441 ( 
.A(n_2440),
.Y(n_2441)
);

AOI22xp33_ASAP7_75t_L g2442 ( 
.A1(n_2438),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.Y(n_2442)
);

OAI22xp5_ASAP7_75t_L g2443 ( 
.A1(n_2441),
.A2(n_2437),
.B1(n_2439),
.B2(n_454),
.Y(n_2443)
);

AOI22xp5_ASAP7_75t_SL g2444 ( 
.A1(n_2443),
.A2(n_2442),
.B1(n_453),
.B2(n_456),
.Y(n_2444)
);

OR2x2_ASAP7_75t_L g2445 ( 
.A(n_2444),
.B(n_452),
.Y(n_2445)
);

AOI221xp5_ASAP7_75t_L g2446 ( 
.A1(n_2445),
.A2(n_457),
.B1(n_459),
.B2(n_461),
.C(n_462),
.Y(n_2446)
);

AOI211xp5_ASAP7_75t_L g2447 ( 
.A1(n_2446),
.A2(n_463),
.B(n_464),
.C(n_465),
.Y(n_2447)
);


endmodule