module fake_jpeg_96_n_172 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_172);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_1),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_39),
.B(n_58),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_2),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_47),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_30),
.B(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_11),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_53),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_12),
.A2(n_3),
.B(n_4),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_52),
.Y(n_84)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_51),
.Y(n_87)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_4),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_12),
.B(n_10),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_57),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_31),
.B(n_10),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_56),
.B(n_17),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_63),
.A2(n_65),
.B1(n_67),
.B2(n_82),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_15),
.B1(n_18),
.B2(n_22),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_76),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_45),
.A2(n_19),
.B1(n_5),
.B2(n_6),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_66),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_6),
.B1(n_9),
.B2(n_38),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_74),
.A2(n_80),
.B1(n_69),
.B2(n_85),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_6),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_36),
.B(n_9),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_89),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_52),
.A2(n_39),
.B1(n_44),
.B2(n_37),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_79),
.A2(n_91),
.B(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_33),
.A2(n_35),
.B1(n_54),
.B2(n_58),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_34),
.A2(n_42),
.B1(n_43),
.B2(n_57),
.Y(n_88)
);

AO22x1_ASAP7_75t_L g93 ( 
.A1(n_88),
.A2(n_69),
.B1(n_68),
.B2(n_80),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_40),
.A2(n_48),
.B1(n_41),
.B2(n_50),
.Y(n_90)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_88),
.B(n_84),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_37),
.A2(n_38),
.B1(n_55),
.B2(n_39),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_61),
.C(n_60),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_100),
.C(n_102),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_99),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_97),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_79),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_77),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_83),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_101),
.A2(n_111),
.B(n_112),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_104),
.B(n_105),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_64),
.B(n_62),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_68),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_113),
.A2(n_80),
.B1(n_59),
.B2(n_86),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_93),
.B1(n_107),
.B2(n_111),
.Y(n_131)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

BUFx4f_ASAP7_75t_SL g138 ( 
.A(n_118),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_96),
.B(n_89),
.C(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_112),
.C(n_100),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_71),
.B(n_101),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_126),
.B(n_128),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_131),
.A2(n_132),
.B1(n_128),
.B2(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_126),
.A2(n_98),
.B1(n_113),
.B2(n_95),
.Y(n_132)
);

OAI32xp33_ASAP7_75t_L g133 ( 
.A1(n_117),
.A2(n_98),
.A3(n_99),
.B1(n_106),
.B2(n_108),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_133),
.A2(n_129),
.B(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_92),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_139),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_136),
.B(n_140),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_118),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_117),
.C(n_123),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_145),
.B(n_146),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_116),
.B(n_125),
.C(n_121),
.D(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_121),
.B(n_129),
.Y(n_148)
);

AO221x1_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_120),
.B1(n_128),
.B2(n_138),
.C(n_110),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_133),
.A2(n_103),
.B(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_132),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_146),
.B1(n_148),
.B2(n_145),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_143),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_144),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_140),
.C(n_136),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_100),
.C(n_102),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_124),
.B(n_102),
.Y(n_160)
);

AO221x1_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_118),
.B1(n_138),
.B2(n_119),
.C(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_156),
.B(n_138),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_158),
.B(n_161),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_159),
.B(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_154),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_164),
.A2(n_151),
.B(n_94),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_165),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_150),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_170),
.C(n_153),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_155),
.A3(n_153),
.B1(n_124),
.B2(n_94),
.C1(n_130),
.C2(n_127),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_130),
.Y(n_172)
);


endmodule