module fake_aes_11953_n_588 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_17, n_63, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_588);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_588;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_73;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_285;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_71;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g70 ( .A(n_37), .Y(n_70) );
CKINVDCx5p33_ASAP7_75t_R g71 ( .A(n_42), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_54), .Y(n_72) );
INVxp33_ASAP7_75t_L g73 ( .A(n_57), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_44), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_40), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_51), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_59), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_58), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_30), .Y(n_79) );
INVx2_ASAP7_75t_L g80 ( .A(n_25), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_47), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_36), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_66), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_69), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_6), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_34), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_49), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_63), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_43), .Y(n_89) );
INVxp67_ASAP7_75t_SL g90 ( .A(n_61), .Y(n_90) );
INVxp67_ASAP7_75t_SL g91 ( .A(n_3), .Y(n_91) );
INVx2_ASAP7_75t_L g92 ( .A(n_4), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_14), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_52), .Y(n_94) );
INVxp33_ASAP7_75t_SL g95 ( .A(n_22), .Y(n_95) );
INVxp33_ASAP7_75t_SL g96 ( .A(n_48), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
CKINVDCx14_ASAP7_75t_R g98 ( .A(n_60), .Y(n_98) );
INVxp67_ASAP7_75t_SL g99 ( .A(n_35), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_33), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_26), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_19), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_1), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_9), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_15), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_27), .Y(n_106) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_45), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_0), .Y(n_108) );
INVxp67_ASAP7_75t_SL g109 ( .A(n_2), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_9), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_23), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_80), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g114 ( .A(n_88), .B(n_0), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g115 ( .A(n_88), .B(n_1), .Y(n_115) );
INVx3_ASAP7_75t_L g116 ( .A(n_92), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_74), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_88), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_85), .B(n_104), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_105), .Y(n_124) );
OA21x2_ASAP7_75t_L g125 ( .A1(n_78), .A2(n_29), .B(n_67), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_88), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
BUFx6f_ASAP7_75t_L g128 ( .A(n_88), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_105), .Y(n_129) );
INVx3_ASAP7_75t_L g130 ( .A(n_92), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_104), .B(n_3), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_100), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_100), .Y(n_133) );
INVx4_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_70), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_103), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_72), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_75), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_76), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_77), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_86), .Y(n_141) );
OAI21x1_ASAP7_75t_L g142 ( .A1(n_87), .A2(n_24), .B(n_65), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_89), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_93), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_97), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_101), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_112), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_117), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_117), .Y(n_150) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_119), .B(n_71), .Y(n_151) );
NAND2xp5_ASAP7_75t_SL g152 ( .A(n_119), .B(n_71), .Y(n_152) );
NOR3xp33_ASAP7_75t_L g153 ( .A(n_121), .B(n_111), .C(n_109), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_122), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_120), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_118), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_122), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_118), .B(n_106), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_136), .B(n_110), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_132), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_133), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_133), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_113), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_113), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_120), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_137), .B(n_107), .Y(n_167) );
INVxp67_ASAP7_75t_L g168 ( .A(n_131), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_137), .B(n_73), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_139), .B(n_110), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_139), .B(n_79), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_123), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_141), .B(n_79), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_123), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_141), .B(n_83), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_144), .B(n_147), .Y(n_176) );
INVxp67_ASAP7_75t_SL g177 ( .A(n_127), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_144), .B(n_148), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_146), .B(n_83), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_146), .B(n_102), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_147), .B(n_102), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_124), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_124), .Y(n_183) );
HB1xp67_ASAP7_75t_L g184 ( .A(n_127), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_148), .B(n_98), .Y(n_185) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_135), .B(n_96), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_135), .B(n_96), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_127), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_138), .B(n_95), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_134), .B(n_95), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_145), .A2(n_91), .B1(n_108), .B2(n_143), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_134), .B(n_99), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_134), .B(n_90), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_120), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_134), .B(n_82), .Y(n_195) );
BUFx6f_ASAP7_75t_L g196 ( .A(n_120), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_129), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_156), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_197), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_164), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_156), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_197), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_188), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_184), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_168), .B(n_145), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_172), .Y(n_207) );
BUFx2_ASAP7_75t_L g208 ( .A(n_159), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_167), .A2(n_84), .B1(n_143), .B2(n_140), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_186), .B(n_140), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_187), .B(n_189), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_186), .B(n_169), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_182), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_183), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_149), .B(n_142), .Y(n_216) );
BUFx12f_ASAP7_75t_L g217 ( .A(n_191), .Y(n_217) );
BUFx2_ASAP7_75t_L g218 ( .A(n_195), .Y(n_218) );
BUFx8_ASAP7_75t_L g219 ( .A(n_150), .Y(n_219) );
AND3x1_ASAP7_75t_SL g220 ( .A(n_153), .B(n_4), .C(n_5), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_169), .B(n_138), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_177), .A2(n_125), .B(n_142), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_171), .B(n_130), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_178), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_187), .B(n_130), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_158), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_175), .B(n_130), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_170), .B(n_116), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_154), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_189), .B(n_116), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_155), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_179), .B(n_130), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_180), .Y(n_233) );
BUFx8_ASAP7_75t_L g234 ( .A(n_157), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g235 ( .A1(n_181), .A2(n_116), .B1(n_125), .B2(n_129), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_185), .B(n_116), .Y(n_236) );
CKINVDCx11_ASAP7_75t_R g237 ( .A(n_160), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_176), .B(n_115), .Y(n_238) );
AND2x4_ASAP7_75t_L g239 ( .A(n_173), .B(n_114), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_176), .B(n_125), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_173), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_151), .B(n_125), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_151), .Y(n_243) );
AND2x4_ASAP7_75t_L g244 ( .A(n_152), .B(n_5), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_161), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_162), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_163), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_192), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_226), .B(n_152), .Y(n_249) );
INVxp67_ASAP7_75t_L g250 ( .A(n_201), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_240), .A2(n_222), .B(n_216), .Y(n_251) );
CKINVDCx5p33_ASAP7_75t_R g252 ( .A(n_237), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_244), .A2(n_190), .B1(n_193), .B2(n_126), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_237), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_207), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_224), .B(n_6), .Y(n_256) );
BUFx12f_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_206), .B(n_7), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_229), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_213), .B(n_7), .Y(n_260) );
AND2x4_ASAP7_75t_L g261 ( .A(n_241), .B(n_8), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_246), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_207), .Y(n_263) );
INVxp67_ASAP7_75t_L g264 ( .A(n_208), .Y(n_264) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_229), .A2(n_128), .B(n_126), .C(n_120), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_247), .Y(n_266) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_216), .A2(n_194), .B(n_166), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_218), .B(n_8), .Y(n_268) );
AO21x2_ASAP7_75t_L g269 ( .A1(n_242), .A2(n_194), .B(n_166), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_233), .B(n_10), .Y(n_270) );
NOR2xp67_ASAP7_75t_L g271 ( .A(n_198), .B(n_10), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_246), .B(n_128), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_221), .A2(n_196), .B(n_155), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_212), .B(n_11), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_209), .A2(n_128), .B1(n_126), .B2(n_13), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_219), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_247), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_245), .Y(n_278) );
INVx3_ASAP7_75t_SL g279 ( .A(n_244), .Y(n_279) );
NOR2xp67_ASAP7_75t_SL g280 ( .A(n_205), .B(n_215), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_248), .B(n_11), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_200), .Y(n_282) );
BUFx12f_ASAP7_75t_L g283 ( .A(n_234), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_238), .A2(n_196), .B(n_155), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_207), .Y(n_285) );
BUFx10_ASAP7_75t_L g286 ( .A(n_244), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_228), .B(n_12), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_266), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_278), .B(n_204), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_251), .A2(n_236), .B(n_227), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_278), .B(n_214), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_266), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g293 ( .A1(n_270), .A2(n_217), .B1(n_243), .B2(n_239), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_277), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_277), .Y(n_295) );
NAND4xp25_ASAP7_75t_L g296 ( .A(n_249), .B(n_212), .C(n_225), .D(n_230), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_256), .B(n_210), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_282), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_282), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_259), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_255), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_264), .B(n_205), .Y(n_302) );
BUFx2_ASAP7_75t_L g303 ( .A(n_250), .Y(n_303) );
AND2x4_ASAP7_75t_L g304 ( .A(n_256), .B(n_230), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_260), .A2(n_235), .B(n_225), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_255), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_281), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_281), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_255), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_286), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_279), .B(n_217), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_255), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_292), .Y(n_314) );
AND2x2_ASAP7_75t_L g315 ( .A(n_289), .B(n_270), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_292), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_303), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
INVx2_ASAP7_75t_SL g319 ( .A(n_302), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_289), .B(n_268), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_297), .B(n_268), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_298), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_291), .B(n_287), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_288), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_298), .B(n_262), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_299), .B(n_287), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_299), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_288), .Y(n_329) );
AND2x4_ASAP7_75t_L g330 ( .A(n_294), .B(n_262), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_294), .B(n_279), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_302), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_300), .Y(n_334) );
BUFx2_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_296), .A2(n_261), .B1(n_286), .B2(n_239), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_318), .Y(n_338) );
OAI211xp5_ASAP7_75t_L g339 ( .A1(n_337), .A2(n_271), .B(n_293), .C(n_296), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_314), .A2(n_267), .B(n_290), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_314), .A2(n_267), .B(n_290), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_335), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_323), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_316), .B(n_308), .Y(n_344) );
AO21x2_ASAP7_75t_L g345 ( .A1(n_327), .A2(n_305), .B(n_269), .Y(n_345) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_324), .A2(n_220), .B1(n_275), .B2(n_308), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_314), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_336), .A2(n_261), .B1(n_304), .B2(n_286), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_327), .A2(n_313), .B(n_310), .Y(n_349) );
AO21x2_ASAP7_75t_L g350 ( .A1(n_323), .A2(n_269), .B(n_273), .Y(n_350) );
INVx2_ASAP7_75t_SL g351 ( .A(n_325), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_329), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_309), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_332), .B(n_309), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_328), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_328), .A2(n_284), .B(n_265), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_329), .B(n_297), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_329), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_320), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_320), .Y(n_360) );
NAND4xp25_ASAP7_75t_L g361 ( .A(n_322), .B(n_312), .C(n_261), .D(n_253), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_318), .A2(n_313), .B(n_301), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g363 ( .A1(n_324), .A2(n_274), .B(n_258), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_334), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_335), .Y(n_366) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
AOI221xp5_ASAP7_75t_L g368 ( .A1(n_332), .A2(n_211), .B1(n_230), .B2(n_304), .C(n_252), .Y(n_368) );
NAND3xp33_ASAP7_75t_SL g369 ( .A(n_346), .B(n_252), .C(n_254), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_338), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_366), .B(n_325), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_352), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_364), .Y(n_373) );
OAI33xp33_ASAP7_75t_L g374 ( .A1(n_361), .A2(n_317), .A3(n_254), .B1(n_331), .B2(n_220), .B3(n_232), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_352), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_352), .B(n_325), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_338), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_358), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_343), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_343), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_358), .B(n_321), .Y(n_381) );
AND2x4_ASAP7_75t_L g382 ( .A(n_360), .B(n_326), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_366), .B(n_319), .Y(n_383) );
CKINVDCx16_ASAP7_75t_R g384 ( .A(n_338), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_358), .B(n_321), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_355), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_364), .Y(n_388) );
NOR2xp33_ASAP7_75t_L g389 ( .A(n_367), .B(n_276), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_342), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_360), .B(n_315), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_347), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_360), .B(n_326), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_355), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_344), .B(n_315), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_357), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_347), .B(n_319), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_359), .B(n_336), .Y(n_398) );
INVx2_ASAP7_75t_SL g399 ( .A(n_351), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_365), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_359), .B(n_326), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_365), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_344), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_353), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_353), .B(n_326), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_357), .B(n_330), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_354), .B(n_330), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_354), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_346), .B(n_330), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_351), .B(n_331), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_361), .B(n_330), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_345), .B(n_307), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_368), .B(n_304), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_403), .B(n_345), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_403), .B(n_404), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_372), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_384), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_379), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_404), .B(n_345), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_376), .B(n_345), .Y(n_420) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_369), .A2(n_339), .B1(n_368), .B2(n_348), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_399), .B(n_234), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_379), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_372), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_396), .B(n_350), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_375), .Y(n_426) );
NAND3xp33_ASAP7_75t_SL g427 ( .A(n_389), .B(n_283), .C(n_257), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_391), .B(n_350), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_395), .B(n_350), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_377), .B(n_350), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_380), .Y(n_432) );
INVxp67_ASAP7_75t_L g433 ( .A(n_399), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_371), .B(n_341), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_371), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_386), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_391), .B(n_363), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_402), .B(n_340), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_370), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_381), .B(n_363), .Y(n_440) );
OR2x4_ASAP7_75t_L g441 ( .A(n_410), .B(n_126), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_381), .B(n_349), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_390), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_385), .B(n_408), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_376), .B(n_341), .Y(n_445) );
INVx2_ASAP7_75t_SL g446 ( .A(n_383), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_374), .B(n_12), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_375), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_411), .A2(n_283), .B1(n_257), .B2(n_311), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_385), .B(n_362), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_386), .B(n_340), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_383), .B(n_13), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_394), .B(n_356), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_394), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_378), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_402), .B(n_356), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_356), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_405), .B(n_356), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_373), .B(n_307), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_378), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_388), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_397), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_387), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_387), .Y(n_465) );
NOR4xp75_ASAP7_75t_L g466 ( .A(n_427), .B(n_409), .C(n_413), .D(n_406), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_458), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_462), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_418), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_446), .B(n_400), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_423), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_431), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_417), .B(n_382), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_439), .B(n_405), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_444), .B(n_398), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_433), .B(n_382), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_446), .B(n_392), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_432), .Y(n_478) );
INVxp67_ASAP7_75t_L g479 ( .A(n_430), .Y(n_479) );
AOI211x1_ASAP7_75t_SL g480 ( .A1(n_422), .A2(n_407), .B(n_392), .C(n_128), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_447), .B(n_412), .C(n_126), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_436), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_454), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_443), .Y(n_484) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_430), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_415), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_463), .B(n_401), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_435), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_437), .B(n_440), .Y(n_489) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_447), .B(n_128), .C(n_397), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_429), .B(n_398), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_450), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_442), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_428), .B(n_401), .Y(n_494) );
INVxp67_ASAP7_75t_SL g495 ( .A(n_425), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_420), .B(n_393), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_441), .Y(n_497) );
HB1xp67_ASAP7_75t_L g498 ( .A(n_434), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_441), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_452), .B(n_382), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_460), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_420), .B(n_393), .Y(n_502) );
OAI32xp33_ASAP7_75t_L g503 ( .A1(n_422), .A2(n_300), .A3(n_311), .B1(n_310), .B2(n_306), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_459), .B(n_393), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_459), .B(n_269), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_451), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_434), .B(n_306), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_414), .B(n_243), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_416), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_416), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_484), .B(n_449), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_474), .B(n_445), .Y(n_513) );
NAND4xp25_ASAP7_75t_L g514 ( .A(n_481), .B(n_421), .C(n_419), .D(n_457), .Y(n_514) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_490), .B(n_457), .C(n_453), .Y(n_515) );
AOI211x1_ASAP7_75t_SL g516 ( .A1(n_473), .A2(n_465), .B(n_464), .C(n_461), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_503), .A2(n_438), .B(n_464), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_468), .Y(n_518) );
NAND4xp25_ASAP7_75t_L g519 ( .A(n_500), .B(n_480), .C(n_473), .D(n_492), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_470), .Y(n_520) );
AOI31xp33_ASAP7_75t_L g521 ( .A1(n_476), .A2(n_445), .A3(n_453), .B(n_456), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_493), .B(n_456), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_500), .A2(n_438), .B(n_461), .C(n_455), .Y(n_523) );
NOR3xp33_ASAP7_75t_L g524 ( .A(n_497), .B(n_223), .C(n_239), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_467), .B(n_465), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_488), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_501), .B(n_438), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_489), .B(n_455), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_486), .B(n_448), .Y(n_529) );
OAI21xp5_ASAP7_75t_L g530 ( .A1(n_499), .A2(n_448), .B(n_426), .Y(n_530) );
NOR3xp33_ASAP7_75t_SL g531 ( .A(n_509), .B(n_476), .C(n_466), .Y(n_531) );
NAND4xp25_ASAP7_75t_L g532 ( .A(n_505), .B(n_426), .C(n_424), .D(n_272), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_498), .A2(n_424), .B1(n_301), .B2(n_262), .Y(n_533) );
NOR4xp25_ASAP7_75t_L g534 ( .A(n_479), .B(n_285), .C(n_202), .D(n_199), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_506), .B(n_16), .Y(n_535) );
AOI211xp5_ASAP7_75t_L g536 ( .A1(n_498), .A2(n_280), .B(n_203), .C(n_196), .Y(n_536) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_479), .A2(n_280), .B1(n_203), .B2(n_207), .C1(n_215), .C2(n_285), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_469), .Y(n_538) );
AOI211xp5_ASAP7_75t_SL g539 ( .A1(n_485), .A2(n_285), .B(n_18), .C(n_20), .Y(n_539) );
OAI21xp33_ASAP7_75t_L g540 ( .A1(n_485), .A2(n_155), .B(n_196), .Y(n_540) );
AOI211xp5_ASAP7_75t_L g541 ( .A1(n_470), .A2(n_203), .B(n_215), .C(n_255), .Y(n_541) );
AOI322xp5_ASAP7_75t_L g542 ( .A1(n_475), .A2(n_202), .A3(n_199), .B1(n_215), .B2(n_203), .C1(n_263), .C2(n_39), .Y(n_542) );
OAI22xp5_ASAP7_75t_SL g543 ( .A1(n_512), .A2(n_495), .B1(n_504), .B2(n_502), .Y(n_543) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_521), .A2(n_495), .B(n_496), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_513), .B(n_508), .Y(n_545) );
NOR2x1p5_ASAP7_75t_L g546 ( .A(n_519), .B(n_494), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_528), .B(n_487), .Y(n_547) );
AND4x2_ASAP7_75t_L g548 ( .A(n_517), .B(n_531), .C(n_516), .D(n_514), .Y(n_548) );
AOI211x1_ASAP7_75t_L g549 ( .A1(n_526), .A2(n_491), .B(n_471), .C(n_478), .Y(n_549) );
INVxp67_ASAP7_75t_L g550 ( .A(n_527), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_518), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_538), .Y(n_552) );
NOR3xp33_ASAP7_75t_L g553 ( .A(n_524), .B(n_483), .C(n_482), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_534), .B(n_477), .Y(n_554) );
OAI22xp5_ASAP7_75t_SL g555 ( .A1(n_515), .A2(n_472), .B1(n_510), .B2(n_511), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_520), .B(n_507), .Y(n_556) );
AOI22xp5_ASAP7_75t_L g557 ( .A1(n_531), .A2(n_263), .B1(n_231), .B2(n_31), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_522), .Y(n_558) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_525), .Y(n_559) );
OAI22xp33_ASAP7_75t_L g560 ( .A1(n_539), .A2(n_263), .B1(n_21), .B2(n_32), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_523), .A2(n_263), .B(n_38), .Y(n_561) );
NAND4xp75_ASAP7_75t_L g562 ( .A(n_557), .B(n_544), .C(n_549), .D(n_554), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_550), .B(n_530), .Y(n_563) );
NAND3xp33_ASAP7_75t_SL g564 ( .A(n_559), .B(n_541), .C(n_536), .Y(n_564) );
NAND4xp75_ASAP7_75t_L g565 ( .A(n_548), .B(n_535), .C(n_529), .D(n_524), .Y(n_565) );
NOR2x1_ASAP7_75t_L g566 ( .A(n_546), .B(n_540), .Y(n_566) );
NAND3x1_ASAP7_75t_L g567 ( .A(n_553), .B(n_542), .C(n_533), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_560), .B(n_532), .C(n_537), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_552), .Y(n_569) );
NOR4xp75_ASAP7_75t_SL g570 ( .A(n_547), .B(n_533), .C(n_41), .D(n_46), .Y(n_570) );
OAI21x1_ASAP7_75t_L g571 ( .A1(n_561), .A2(n_17), .B(n_50), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_551), .Y(n_572) );
AOI21xp5_ASAP7_75t_L g573 ( .A1(n_566), .A2(n_543), .B(n_555), .Y(n_573) );
XOR2xp5_ASAP7_75t_L g574 ( .A(n_565), .B(n_558), .Y(n_574) );
INVx3_ASAP7_75t_L g575 ( .A(n_562), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_569), .Y(n_576) );
OAI22xp33_ASAP7_75t_L g577 ( .A1(n_564), .A2(n_550), .B1(n_556), .B2(n_545), .Y(n_577) );
AOI211xp5_ASAP7_75t_L g578 ( .A1(n_568), .A2(n_263), .B(n_55), .C(n_56), .Y(n_578) );
XNOR2xp5_ASAP7_75t_SL g579 ( .A(n_574), .B(n_572), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_575), .A2(n_567), .B1(n_563), .B2(n_571), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_576), .Y(n_581) );
AOI221x1_ASAP7_75t_L g582 ( .A1(n_573), .A2(n_570), .B1(n_62), .B2(n_64), .C(n_68), .Y(n_582) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_580), .A2(n_577), .B1(n_578), .B2(n_570), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_581), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_584), .B(n_579), .Y(n_585) );
OAI21xp5_ASAP7_75t_L g586 ( .A1(n_583), .A2(n_582), .B(n_53), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_585), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g588 ( .A1(n_587), .A2(n_231), .B1(n_586), .B2(n_575), .C(n_585), .Y(n_588) );
endmodule