module fake_jpeg_18726_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_39),
.Y(n_65)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx2_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

FAx1_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_16),
.CI(n_23),
.CON(n_55),
.SN(n_55)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_16),
.B1(n_21),
.B2(n_28),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_49),
.A2(n_61),
.B1(n_39),
.B2(n_36),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_59),
.Y(n_67)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NAND2xp33_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_43),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_46),
.B(n_41),
.C(n_40),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_58),
.A2(n_43),
.B1(n_39),
.B2(n_36),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_35),
.B1(n_34),
.B2(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_64),
.Y(n_82)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_66),
.Y(n_70)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_42),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_71),
.A2(n_91),
.B(n_94),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_73),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_65),
.B(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_36),
.B1(n_45),
.B2(n_39),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

NAND3xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_44),
.C(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_77),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_52),
.C(n_55),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_84),
.C(n_87),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_29),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_78),
.A2(n_89),
.B1(n_103),
.B2(n_104),
.Y(n_126)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_79),
.B(n_93),
.Y(n_139)
);

AOI22x1_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_37),
.B1(n_43),
.B2(n_46),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_81),
.A2(n_91),
.B1(n_84),
.B2(n_85),
.Y(n_122)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_83),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_37),
.C(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_85),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_102),
.Y(n_132)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_47),
.B(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_90),
.Y(n_135)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_32),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_23),
.Y(n_94)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_56),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_107),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_29),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_96),
.Y(n_116)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_99),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_63),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_46),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_109),
.Y(n_118)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_60),
.A2(n_26),
.B1(n_19),
.B2(n_22),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_56),
.B(n_22),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_105),
.A2(n_108),
.B(n_0),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_56),
.A2(n_26),
.B1(n_19),
.B2(n_31),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_106),
.A2(n_17),
.B1(n_18),
.B2(n_25),
.Y(n_111)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_54),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_30),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_71),
.A2(n_41),
.B(n_40),
.C(n_38),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_110),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_111),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_94),
.A2(n_31),
.B1(n_33),
.B2(n_27),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_119),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_30),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_122),
.A2(n_131),
.B1(n_81),
.B2(n_101),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_128),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_86),
.A2(n_30),
.B(n_23),
.C(n_7),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_67),
.B(n_30),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_130),
.B(n_78),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_91),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_41),
.B1(n_40),
.B2(n_38),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_141),
.A2(n_95),
.B1(n_99),
.B2(n_102),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_134),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_142),
.B(n_148),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_165),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_108),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_144),
.Y(n_204)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_160),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_72),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_80),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_149),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_150),
.A2(n_152),
.B1(n_170),
.B2(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_67),
.C(n_94),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_157),
.C(n_164),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_80),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_155),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_87),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_87),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_163),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_104),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_122),
.B(n_82),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_166),
.Y(n_180)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_123),
.B(n_137),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_168),
.A2(n_138),
.B1(n_82),
.B2(n_114),
.Y(n_189)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_123),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_131),
.A2(n_126),
.B1(n_121),
.B2(n_137),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_SL g174 ( 
.A(n_171),
.B(n_120),
.C(n_117),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_132),
.B(n_125),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_191),
.B1(n_167),
.B2(n_166),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_174),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_132),
.C(n_130),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_202),
.C(n_30),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_147),
.A2(n_112),
.B(n_129),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_139),
.B(n_113),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_179),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_170),
.A2(n_126),
.B1(n_110),
.B2(n_140),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_185),
.A2(n_188),
.B1(n_200),
.B2(n_173),
.Y(n_232)
);

AND2x6_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_110),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_151),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_88),
.B1(n_90),
.B2(n_92),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_161),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_145),
.A2(n_138),
.B(n_114),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_201),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_169),
.A2(n_95),
.B1(n_124),
.B2(n_79),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_124),
.B1(n_70),
.B2(n_107),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_159),
.B1(n_146),
.B2(n_158),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_143),
.B(n_160),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_27),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_156),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_153),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_154),
.B(n_68),
.C(n_70),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_23),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_205),
.A2(n_232),
.B1(n_203),
.B2(n_199),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_206),
.A2(n_211),
.B1(n_179),
.B2(n_186),
.Y(n_237)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_220),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_218),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_151),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_172),
.B(n_229),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_157),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_225),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_222),
.C(n_224),
.Y(n_234)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_193),
.Y(n_215)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_193),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_219),
.B(n_231),
.Y(n_254)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_195),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_175),
.B(n_97),
.C(n_23),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_33),
.C(n_27),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_33),
.C(n_27),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_183),
.Y(n_244)
);

XOR2x2_ASAP7_75t_SL g228 ( 
.A(n_198),
.B(n_8),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_33),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g233 ( 
.A(n_221),
.Y(n_233)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_210),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_237),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_236),
.A2(n_247),
.B1(n_184),
.B2(n_195),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_207),
.A2(n_185),
.B1(n_226),
.B2(n_229),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_209),
.B1(n_227),
.B2(n_228),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_209),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_246),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_232),
.A2(n_194),
.B1(n_190),
.B2(n_182),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_245),
.A2(n_216),
.B1(n_211),
.B2(n_225),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_202),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_222),
.B(n_174),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_251),
.B(n_214),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_180),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_200),
.B(n_186),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_255),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_271),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_265),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_260),
.B(n_5),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_269),
.B1(n_275),
.B2(n_254),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_176),
.Y(n_263)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_263),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_264),
.A2(n_245),
.B1(n_243),
.B2(n_241),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_238),
.B(n_224),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_238),
.B(n_184),
.C(n_220),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_270),
.C(n_272),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_98),
.C(n_7),
.Y(n_270)
);

AND2x2_ASAP7_75t_SL g271 ( 
.A(n_240),
.B(n_0),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_234),
.B(n_7),
.C(n_14),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_9),
.Y(n_274)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_274),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_236),
.A2(n_9),
.B1(n_14),
.B2(n_13),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g277 ( 
.A(n_266),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_286),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_234),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_280),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_256),
.A2(n_247),
.B1(n_241),
.B2(n_249),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_281),
.A2(n_264),
.B1(n_263),
.B2(n_262),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_268),
.B(n_244),
.C(n_255),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_289),
.C(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_258),
.B(n_253),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_261),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_250),
.C(n_11),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_291),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_11),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_296),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_298),
.C(n_299),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_257),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_289),
.Y(n_299)
);

AOI211xp5_ASAP7_75t_SL g300 ( 
.A1(n_280),
.A2(n_259),
.B(n_271),
.C(n_273),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_302),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_271),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_288),
.C(n_13),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_284),
.B(n_4),
.C(n_13),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g304 ( 
.A(n_297),
.B(n_279),
.CI(n_300),
.CON(n_304),
.SN(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_283),
.C(n_279),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_307),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_283),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_311),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_14),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_311),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_15),
.Y(n_311)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_15),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_317),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_309),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_315),
.A2(n_306),
.B(n_303),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_319),
.A2(n_316),
.B(n_306),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_305),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_321),
.B(n_312),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_322),
.B(n_323),
.C(n_318),
.Y(n_324)
);

A2O1A1O1Ixp25_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_304),
.B(n_312),
.C(n_320),
.D(n_1),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_3),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_1),
.B(n_2),
.Y(n_328)
);


endmodule