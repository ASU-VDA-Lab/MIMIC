module fake_jpeg_31506_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_39),
.B(n_43),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_46),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx10_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_10),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_9),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_0),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_74),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_77),
.B(n_69),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_78),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_62),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_57),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_49),
.B1(n_63),
.B2(n_52),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_88),
.B1(n_21),
.B2(n_47),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_73),
.A2(n_65),
.B1(n_60),
.B2(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_91),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_90),
.B(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_63),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_70),
.A2(n_67),
.B(n_56),
.C(n_64),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_92),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_108)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx13_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_98),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_64),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_52),
.B1(n_66),
.B2(n_64),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_99),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_85),
.B(n_53),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_103),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_82),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_79),
.A2(n_78),
.B(n_66),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

AOI32xp33_ASAP7_75t_L g106 ( 
.A1(n_92),
.A2(n_59),
.A3(n_58),
.B1(n_54),
.B2(n_24),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_111),
.B1(n_13),
.B2(n_14),
.Y(n_130)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_88),
.B(n_93),
.C(n_3),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_112),
.B(n_93),
.C(n_2),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_117),
.B1(n_122),
.B2(n_44),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_111),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_116),
.A2(n_118),
.B(n_119),
.C(n_38),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_112),
.A2(n_104),
.B1(n_109),
.B2(n_98),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_96),
.A2(n_109),
.B1(n_108),
.B2(n_107),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_132),
.B1(n_116),
.B2(n_115),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_11),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_130),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_101),
.B(n_12),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_129),
.B(n_15),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_111),
.A2(n_13),
.B1(n_15),
.B2(n_18),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_131),
.B(n_32),
.C(n_22),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_135),
.C(n_136),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_138),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_26),
.C(n_28),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_29),
.C(n_30),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_128),
.A2(n_31),
.B(n_33),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_137),
.Y(n_150)
);

OA21x2_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_35),
.B(n_37),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_140),
.A2(n_141),
.B1(n_145),
.B2(n_146),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_45),
.C(n_48),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_120),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_127),
.B1(n_119),
.B2(n_118),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_147),
.B1(n_140),
.B2(n_139),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_155),
.B(n_156),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_133),
.C(n_135),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_138),
.Y(n_157)
);

OAI211xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_148),
.B(n_152),
.C(n_140),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_147),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_158),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_150),
.B(n_151),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_162),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_149),
.Y(n_164)
);


endmodule