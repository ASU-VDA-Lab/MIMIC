module fake_jpeg_30089_n_544 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_544);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_544;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_31),
.B(n_9),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_18),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_64),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_20),
.B(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_65),
.B(n_68),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_71),
.B(n_75),
.Y(n_133)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_74),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_31),
.B(n_18),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_91),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_83),
.Y(n_161)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_42),
.Y(n_85)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_97),
.Y(n_152)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_47),
.B(n_9),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_47),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_30),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_99),
.B(n_103),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_39),
.Y(n_100)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_101),
.Y(n_143)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_30),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_107),
.B(n_23),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_112),
.B(n_50),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_121),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g124 ( 
.A1(n_65),
.A2(n_58),
.B1(n_98),
.B2(n_102),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_85),
.B1(n_51),
.B2(n_19),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

BUFx24_ASAP7_75t_L g217 ( 
.A(n_125),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_65),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_145),
.Y(n_177)
);

INVx2_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_130),
.B(n_30),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_87),
.B(n_22),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_131),
.B(n_153),
.Y(n_174)
);

HAxp5_ASAP7_75t_SL g137 ( 
.A(n_84),
.B(n_29),
.CON(n_137),
.SN(n_137)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_137),
.A2(n_117),
.B(n_150),
.Y(n_184)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_52),
.Y(n_144)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_56),
.B(n_40),
.C(n_51),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_148),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_40),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_155),
.Y(n_187)
);

BUFx12_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_156),
.Y(n_171)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_59),
.Y(n_159)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_159),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_92),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_91),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_168),
.B(n_185),
.Y(n_253)
);

AND2x2_ASAP7_75t_SL g169 ( 
.A(n_106),
.B(n_0),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_169),
.B(n_156),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_130),
.A2(n_42),
.B1(n_91),
.B2(n_64),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_170),
.A2(n_193),
.B1(n_202),
.B2(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_172),
.Y(n_231)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_173),
.Y(n_236)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_131),
.A2(n_70),
.B1(n_100),
.B2(n_89),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_179),
.A2(n_208),
.B1(n_163),
.B2(n_157),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_137),
.A2(n_23),
.B1(n_19),
.B2(n_49),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_41),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_183),
.B(n_188),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_184),
.Y(n_259)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_133),
.B(n_41),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_108),
.B(n_49),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_189),
.B(n_209),
.Y(n_248)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_190),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_104),
.Y(n_191)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_108),
.B(n_26),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_192),
.B(n_198),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_122),
.A2(n_68),
.B1(n_64),
.B2(n_41),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_117),
.B(n_34),
.C(n_43),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_194),
.B(n_214),
.C(n_115),
.Y(n_246)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_195),
.Y(n_230)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_196),
.Y(n_270)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_150),
.B(n_41),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_127),
.Y(n_199)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_199),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_124),
.A2(n_73),
.B1(n_57),
.B2(n_82),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_200),
.A2(n_207),
.B1(n_202),
.B2(n_170),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_201),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_154),
.A2(n_68),
.B1(n_80),
.B2(n_74),
.Y(n_202)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_203),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_116),
.Y(n_204)
);

BUFx4f_ASAP7_75t_L g241 ( 
.A(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_205),
.Y(n_277)
);

O2A1O1Ixp33_ASAP7_75t_L g206 ( 
.A1(n_145),
.A2(n_124),
.B(n_120),
.C(n_147),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_206),
.A2(n_125),
.B(n_118),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_135),
.A2(n_53),
.B1(n_61),
.B2(n_101),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_152),
.A2(n_86),
.B1(n_43),
.B2(n_34),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_141),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_210),
.Y(n_235)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_211),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_213),
.B(n_220),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_30),
.C(n_11),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_215),
.Y(n_254)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_165),
.Y(n_216)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_216),
.Y(n_264)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_136),
.Y(n_218)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_218),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_132),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_219),
.A2(n_222),
.B1(n_226),
.B2(n_3),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_162),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_221),
.Y(n_280)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_138),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_138),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g224 ( 
.A(n_142),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_224),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_143),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_121),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_168),
.A2(n_123),
.B1(n_126),
.B2(n_111),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_229),
.A2(n_240),
.B1(n_242),
.B2(n_245),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_174),
.B(n_206),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_232),
.B(n_257),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_168),
.A2(n_157),
.B1(n_163),
.B2(n_139),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_200),
.A2(n_161),
.B1(n_114),
.B2(n_152),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_268),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_177),
.B(n_115),
.C(n_160),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_251),
.C(n_273),
.Y(n_288)
);

OR2x2_ASAP7_75t_SL g327 ( 
.A(n_249),
.B(n_267),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_149),
.C(n_155),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_169),
.A2(n_149),
.B1(n_13),
.B2(n_14),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_201),
.A2(n_2),
.B(n_3),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_180),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g269 ( 
.A1(n_219),
.A2(n_118),
.B(n_12),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_272),
.Y(n_289)
);

AOI32xp33_ASAP7_75t_L g272 ( 
.A1(n_199),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_8),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_204),
.A2(n_2),
.B(n_3),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_265),
.B1(n_171),
.B2(n_227),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_176),
.B(n_3),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_276),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_178),
.A2(n_15),
.B1(n_7),
.B2(n_8),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_279),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_193),
.A2(n_15),
.B1(n_7),
.B2(n_8),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_241),
.Y(n_281)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_281),
.B(n_293),
.Y(n_336)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

BUFx8_ASAP7_75t_L g330 ( 
.A(n_283),
.Y(n_330)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_286),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_182),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_290),
.B(n_316),
.Y(n_334)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_237),
.Y(n_291)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_291),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_224),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_292),
.B(n_294),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_255),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_224),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_295),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_296),
.A2(n_321),
.B1(n_234),
.B2(n_287),
.Y(n_370)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_297),
.Y(n_335)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_236),
.Y(n_299)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_299),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_231),
.B(n_212),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_300),
.B(n_301),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_230),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_230),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_302),
.B(n_303),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_270),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_167),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_305),
.B(n_306),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_244),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_307),
.Y(n_344)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_308),
.B(n_311),
.Y(n_331)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_175),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_312),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_270),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_313),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_239),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_318),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_239),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_315),
.Y(n_360)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_254),
.Y(n_316)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_254),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_322),
.Y(n_350)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_236),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_320),
.A2(n_324),
.B1(n_328),
.B2(n_187),
.Y(n_357)
);

OAI22x1_ASAP7_75t_SL g321 ( 
.A1(n_253),
.A2(n_226),
.B1(n_225),
.B2(n_217),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_253),
.B(n_225),
.Y(n_322)
);

AND2x6_ASAP7_75t_L g323 ( 
.A(n_259),
.B(n_217),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_323),
.A2(n_233),
.B(n_232),
.Y(n_337)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx13_ASAP7_75t_L g325 ( 
.A(n_260),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_325),
.Y(n_367)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_235),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_222),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_228),
.A2(n_187),
.B1(n_227),
.B2(n_203),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_256),
.B1(n_233),
.B2(n_265),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_332),
.A2(n_349),
.B1(n_354),
.B2(n_295),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_249),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_333),
.B(n_355),
.C(n_319),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_337),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_284),
.A2(n_242),
.B1(n_267),
.B2(n_247),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_340),
.A2(n_356),
.B1(n_362),
.B2(n_370),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_321),
.A2(n_279),
.B1(n_276),
.B2(n_263),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_289),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_276),
.B1(n_248),
.B2(n_250),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g351 ( 
.A1(n_322),
.A2(n_273),
.B(n_244),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_351),
.A2(n_353),
.B(n_363),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_298),
.A2(n_246),
.B(n_251),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_317),
.A2(n_250),
.B1(n_274),
.B2(n_261),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_258),
.C(n_252),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_309),
.A2(n_278),
.B1(n_257),
.B2(n_274),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_357),
.A2(n_307),
.B1(n_313),
.B2(n_303),
.Y(n_379)
);

AO22x1_ASAP7_75t_SL g361 ( 
.A1(n_290),
.A2(n_191),
.B1(n_223),
.B2(n_238),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_361),
.B(n_365),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_287),
.A2(n_195),
.B1(n_196),
.B2(n_218),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_298),
.A2(n_261),
.B(n_217),
.Y(n_363)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_364),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_285),
.B(n_7),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_285),
.B(n_7),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_281),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_293),
.B(n_187),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_369),
.B(n_314),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_371),
.A2(n_379),
.B(n_383),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_369),
.B(n_291),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_372),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_382),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_308),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_376),
.B(n_384),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_336),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_385),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_378),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_L g423 ( 
.A1(n_380),
.A2(n_341),
.B(n_367),
.Y(n_423)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_335),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

OA21x2_ASAP7_75t_L g382 ( 
.A1(n_351),
.A2(n_323),
.B(n_327),
.Y(n_382)
);

AND2x6_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_325),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_331),
.B(n_326),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_336),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_386),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_358),
.B(n_324),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_387),
.B(n_394),
.Y(n_416)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_346),
.Y(n_390)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_390),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_288),
.Y(n_391)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_364),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_393),
.B(n_395),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_352),
.B(n_320),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_350),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_347),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_396),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g397 ( 
.A1(n_332),
.A2(n_288),
.B1(n_302),
.B2(n_301),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_397),
.A2(n_349),
.B1(n_354),
.B2(n_359),
.Y(n_415)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_398),
.B(n_355),
.Y(n_413)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_399),
.Y(n_431)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_329),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_400),
.B(n_359),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_345),
.A2(n_297),
.B1(n_316),
.B2(n_307),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_401),
.A2(n_405),
.B1(n_356),
.B2(n_362),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g402 ( 
.A1(n_363),
.A2(n_312),
.B(n_310),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_402),
.A2(n_350),
.B(n_339),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_330),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_403),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_330),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_404),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_408),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_413),
.B(n_428),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_415),
.A2(n_401),
.B1(n_405),
.B2(n_371),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_396),
.B(n_366),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_418),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_419),
.A2(n_373),
.B1(n_375),
.B2(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

AO21x1_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_430),
.B(n_373),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_380),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_424),
.B(n_426),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_398),
.B(n_391),
.C(n_333),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_392),
.C(n_371),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_378),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_389),
.B(n_353),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_406),
.A2(n_377),
.B1(n_385),
.B2(n_392),
.Y(n_429)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

AND2x6_ASAP7_75t_L g430 ( 
.A(n_383),
.B(n_340),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_365),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_433),
.B(n_329),
.Y(n_457)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_438),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_440),
.C(n_441),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_413),
.B(n_406),
.C(n_393),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_374),
.C(n_395),
.Y(n_441)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g444 ( 
.A(n_412),
.B(n_404),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_454),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_445),
.A2(n_453),
.B1(n_456),
.B2(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_422),
.B(n_403),
.Y(n_448)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_448),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_390),
.Y(n_450)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_414),
.A2(n_381),
.B1(n_388),
.B2(n_386),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_421),
.A2(n_402),
.B(n_382),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_419),
.A2(n_382),
.B1(n_400),
.B2(n_343),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_457),
.B(n_430),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_433),
.A2(n_399),
.B1(n_344),
.B2(n_342),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_462),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_410),
.B(n_361),
.Y(n_459)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_459),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_428),
.B(n_361),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_460),
.B(n_417),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_409),
.B(n_338),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_461),
.B(n_408),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_435),
.A2(n_344),
.B1(n_342),
.B2(n_367),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_421),
.A2(n_368),
.B(n_360),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_463),
.B(n_436),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_439),
.B(n_435),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_464),
.B(n_484),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_467),
.A2(n_470),
.B1(n_458),
.B2(n_449),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_409),
.C(n_437),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_473),
.C(n_482),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_455),
.A2(n_416),
.B1(n_407),
.B2(n_434),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_437),
.C(n_436),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_476),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_477),
.B(n_442),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_478),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_452),
.B(n_411),
.C(n_427),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_441),
.B(n_434),
.C(n_427),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_443),
.C(n_450),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_457),
.B(n_407),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g485 ( 
.A(n_447),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_485),
.Y(n_487)
);

FAx1_ASAP7_75t_SL g489 ( 
.A(n_475),
.B(n_461),
.CI(n_460),
.CON(n_489),
.SN(n_489)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_489),
.B(n_496),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_491),
.B(n_496),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_492),
.B(n_495),
.Y(n_505)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_493),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_469),
.A2(n_463),
.B(n_454),
.Y(n_494)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_494),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_465),
.B(n_456),
.C(n_438),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_445),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_497),
.B(n_501),
.C(n_476),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g498 ( 
.A(n_471),
.B(n_446),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_498),
.B(n_499),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_465),
.B(n_462),
.C(n_459),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_479),
.B(n_482),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_431),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_451),
.C(n_432),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_486),
.A2(n_468),
.B(n_480),
.Y(n_504)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_504),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_500),
.A2(n_466),
.B1(n_481),
.B2(n_477),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_507),
.B(n_513),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_508),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_490),
.A2(n_474),
.B(n_484),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_509),
.A2(n_502),
.B(n_338),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_497),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_511),
.B(n_514),
.Y(n_523)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_499),
.B(n_432),
.CI(n_360),
.CON(n_514),
.SN(n_514)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_486),
.B(n_495),
.C(n_492),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_515),
.B(n_501),
.C(n_502),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_516),
.A2(n_368),
.B1(n_378),
.B2(n_299),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_518),
.B(n_511),
.C(n_505),
.Y(n_527)
);

AOI21x1_ASAP7_75t_L g521 ( 
.A1(n_510),
.A2(n_487),
.B(n_489),
.Y(n_521)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_521),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_488),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_522),
.B(n_525),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_506),
.A2(n_489),
.B1(n_488),
.B2(n_431),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_524),
.B(n_526),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_529),
.C(n_531),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_520),
.A2(n_516),
.B1(n_503),
.B2(n_508),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_514),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_532),
.A2(n_523),
.B1(n_519),
.B2(n_526),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_533),
.B(n_528),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_527),
.A2(n_519),
.B(n_509),
.Y(n_535)
);

AO21x1_ASAP7_75t_L g538 ( 
.A1(n_535),
.A2(n_536),
.B(n_522),
.Y(n_538)
);

MAJx2_ASAP7_75t_L g536 ( 
.A(n_530),
.B(n_528),
.C(n_517),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_537),
.B(n_538),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_539),
.B(n_534),
.C(n_536),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_540),
.B(n_512),
.C(n_304),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_315),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_542),
.A2(n_330),
.B1(n_318),
.B2(n_286),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_283),
.Y(n_544)
);


endmodule