module fake_netlist_6_514_n_1716 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1716);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1716;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_58),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_75),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_81),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_132),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_154),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_152),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_47),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_80),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_47),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_48),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_28),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_27),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_41),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_42),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_13),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_114),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_37),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_147),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_87),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_93),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_8),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_43),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_39),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_96),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_60),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_63),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_140),
.Y(n_189)
);

INVx4_ASAP7_75t_R g190 ( 
.A(n_66),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_146),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_62),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_88),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_30),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_13),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_134),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_3),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_49),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_119),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_121),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_44),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_153),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_4),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_92),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_99),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_20),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_55),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_111),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_4),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_11),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_24),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_36),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_118),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_73),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_128),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_90),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_106),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_83),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_8),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_34),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_43),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_58),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_5),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_55),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_112),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_102),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_40),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_137),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_1),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_20),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_34),
.Y(n_236)
);

BUFx10_ASAP7_75t_L g237 ( 
.A(n_70),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_104),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_74),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_2),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_7),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_79),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_68),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_57),
.Y(n_244)
);

INVxp67_ASAP7_75t_SL g245 ( 
.A(n_19),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_95),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_18),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_143),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_12),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_56),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_1),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_5),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_113),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_149),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_7),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_14),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_11),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_107),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_16),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_98),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_89),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_64),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_145),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_21),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_38),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_124),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_125),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_130),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_19),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_21),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_48),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_54),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_28),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_9),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_86),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_23),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_32),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_35),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_101),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_120),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_45),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_30),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_72),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_27),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_52),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_3),
.Y(n_290)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_69),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_12),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_57),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_110),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_133),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g296 ( 
.A(n_44),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_60),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_46),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_35),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_155),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_61),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_9),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_10),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_115),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_32),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_122),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_33),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_0),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_296),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_156),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_0),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_296),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_234),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_158),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_296),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_160),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_174),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_161),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_296),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_159),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_296),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_204),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_204),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_165),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_189),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_204),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_217),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_217),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_163),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_184),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_217),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_205),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_184),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_260),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_250),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_164),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_166),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_206),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_250),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_270),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_168),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_269),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_172),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_307),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_269),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_307),
.Y(n_353)
);

INVxp67_ASAP7_75t_SL g354 ( 
.A(n_263),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_290),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_176),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_178),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_290),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_173),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_305),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_179),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_172),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_172),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_266),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_180),
.Y(n_366)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_228),
.B(n_2),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_173),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_186),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_266),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_188),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_266),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_191),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_167),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_162),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_274),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_194),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_200),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_309),
.Y(n_379)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_350),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_312),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_312),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_314),
.B(n_316),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_314),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_231),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_317),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_317),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_322),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_L g391 ( 
.A(n_311),
.B(n_210),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_334),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

NAND2x1_ASAP7_75t_L g395 ( 
.A(n_311),
.B(n_190),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_325),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_325),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_326),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_326),
.B(n_231),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_375),
.B(n_162),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_327),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_203),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_331),
.B(n_295),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_319),
.B(n_203),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_332),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_335),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_338),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_338),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_342),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_347),
.B(n_264),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_347),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_349),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_349),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_351),
.B(n_264),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_353),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_363),
.B(n_295),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_319),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_337),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_360),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_364),
.B(n_295),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_344),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_339),
.A2(n_251),
.B1(n_171),
.B2(n_232),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_367),
.B(n_237),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_350),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_364),
.B(n_192),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_352),
.B(n_244),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_357),
.Y(n_443)
);

INVx6_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_401),
.B(n_315),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_318),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_435),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_410),
.B(n_320),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_430),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_392),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_392),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_388),
.B(n_333),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_403),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_388),
.B(n_340),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_435),
.B(n_339),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_391),
.A2(n_354),
.B1(n_313),
.B2(n_321),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_391),
.A2(n_274),
.B1(n_280),
.B2(n_359),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_382),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_382),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_392),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_410),
.B(n_341),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_393),
.B(n_346),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_392),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_412),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_383),
.Y(n_470)
);

INVxp33_ASAP7_75t_L g471 ( 
.A(n_442),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_388),
.B(n_356),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_388),
.B(n_366),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_383),
.Y(n_475)
);

OAI22xp33_ASAP7_75t_L g476 ( 
.A1(n_393),
.A2(n_157),
.B1(n_281),
.B2(n_367),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_443),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_403),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_403),
.A2(n_280),
.B1(n_274),
.B2(n_359),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_392),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_383),
.Y(n_482)
);

AND2x6_ASAP7_75t_L g483 ( 
.A(n_388),
.B(n_192),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_431),
.B(n_362),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_L g487 ( 
.A(n_387),
.B(n_210),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

INVxp67_ASAP7_75t_SL g489 ( 
.A(n_385),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_379),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_379),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_379),
.Y(n_494)
);

INVx11_ASAP7_75t_L g495 ( 
.A(n_381),
.Y(n_495)
);

NAND2xp33_ASAP7_75t_L g496 ( 
.A(n_387),
.B(n_210),
.Y(n_496)
);

NOR3xp33_ASAP7_75t_L g497 ( 
.A(n_437),
.B(n_245),
.C(n_292),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_431),
.B(n_369),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_379),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_389),
.Y(n_502)
);

BUFx4f_ASAP7_75t_L g503 ( 
.A(n_392),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_381),
.B(n_378),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_395),
.A2(n_377),
.B1(n_373),
.B2(n_371),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_438),
.B(n_374),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_398),
.B(n_380),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_438),
.B(n_376),
.Y(n_508)
);

NAND2xp33_ASAP7_75t_R g509 ( 
.A(n_384),
.B(n_376),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_398),
.B(n_365),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_392),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_429),
.B(n_365),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_398),
.Y(n_513)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_395),
.B(n_368),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_396),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_396),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_380),
.B(n_370),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_SL g518 ( 
.A(n_437),
.B(n_261),
.C(n_257),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_380),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_396),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_396),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_394),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_442),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_380),
.B(n_372),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_395),
.B(n_310),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_380),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_408),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_380),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_390),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_390),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_390),
.B(n_201),
.Y(n_531)
);

INVx4_ASAP7_75t_SL g532 ( 
.A(n_394),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_430),
.A2(n_215),
.B1(n_308),
.B2(n_302),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_397),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_394),
.Y(n_535)
);

BUFx10_ASAP7_75t_L g536 ( 
.A(n_443),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_390),
.B(n_211),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_397),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_381),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_385),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_429),
.B(n_368),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_390),
.B(n_218),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_408),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_390),
.B(n_219),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_429),
.B(n_434),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_385),
.B(n_220),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_397),
.B(n_222),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_394),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_SL g549 ( 
.A1(n_381),
.A2(n_328),
.B1(n_345),
.B2(n_343),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_397),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_394),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_429),
.B(n_434),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_404),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_381),
.B(n_237),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_434),
.B(n_223),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_440),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_404),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_434),
.Y(n_558)
);

OR2x6_ASAP7_75t_L g559 ( 
.A(n_384),
.B(n_280),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_440),
.B(n_237),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_408),
.B(n_233),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g562 ( 
.A(n_387),
.B(n_192),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_L g563 ( 
.A(n_413),
.B(n_238),
.Y(n_563)
);

CKINVDCx14_ASAP7_75t_R g564 ( 
.A(n_384),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_408),
.B(n_239),
.Y(n_565)
);

AND3x1_ASAP7_75t_L g566 ( 
.A(n_441),
.B(n_187),
.C(n_185),
.Y(n_566)
);

INVx5_ASAP7_75t_L g567 ( 
.A(n_394),
.Y(n_567)
);

BUFx8_ASAP7_75t_SL g568 ( 
.A(n_430),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_404),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_394),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_440),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_413),
.B(n_323),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_408),
.A2(n_202),
.B1(n_303),
.B2(n_299),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_404),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_408),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_405),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_394),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_394),
.B(n_243),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_405),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_440),
.B(n_237),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_405),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_441),
.B(n_221),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_394),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_441),
.A2(n_199),
.B1(n_303),
.B2(n_299),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_440),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_413),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_441),
.B(n_246),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_413),
.B(n_249),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_440),
.B(n_291),
.Y(n_589)
);

INVxp67_ASAP7_75t_L g590 ( 
.A(n_509),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_450),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_457),
.B(n_427),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_444),
.Y(n_593)
);

AND2x6_ASAP7_75t_SL g594 ( 
.A(n_485),
.B(n_185),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_457),
.B(n_427),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_527),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_489),
.B(n_440),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_527),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_459),
.Y(n_599)
);

AOI22xp5_ASAP7_75t_L g600 ( 
.A1(n_479),
.A2(n_336),
.B1(n_329),
.B2(n_265),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_450),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_543),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_446),
.B(n_442),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_543),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_540),
.B(n_413),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_545),
.A2(n_458),
.B(n_456),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_552),
.B(n_413),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_575),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_575),
.Y(n_609)
);

NOR3xp33_ASAP7_75t_L g610 ( 
.A(n_518),
.B(n_437),
.C(n_170),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_552),
.B(n_562),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_552),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_558),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_L g614 ( 
.A(n_582),
.B(n_210),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_444),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_562),
.B(n_546),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_562),
.A2(n_221),
.B1(n_287),
.B2(n_182),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_479),
.B(n_436),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_462),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_512),
.B(n_439),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_L g621 ( 
.A(n_448),
.B(n_400),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_462),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_508),
.B(n_436),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_463),
.B(n_436),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_512),
.B(n_439),
.Y(n_625)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_459),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_463),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_444),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_444),
.Y(n_629)
);

BUFx4f_ASAP7_75t_L g630 ( 
.A(n_514),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_470),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_470),
.B(n_436),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_586),
.B(n_210),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_586),
.B(n_210),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_586),
.B(n_287),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_475),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_506),
.B(n_221),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_475),
.B(n_436),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_482),
.B(n_436),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_466),
.B(n_255),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_473),
.B(n_268),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_482),
.B(n_402),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_486),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_467),
.B(n_169),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_474),
.B(n_279),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_512),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_568),
.Y(n_647)
);

INVx3_ASAP7_75t_L g648 ( 
.A(n_454),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_486),
.B(n_402),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_488),
.B(n_283),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_488),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_454),
.Y(n_652)
);

BUFx12f_ASAP7_75t_SL g653 ( 
.A(n_559),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_492),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_492),
.B(n_402),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_501),
.B(n_284),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_514),
.A2(n_306),
.B1(n_304),
.B2(n_301),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_501),
.B(n_402),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_502),
.B(n_402),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_502),
.B(n_402),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_513),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_445),
.B(n_175),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_447),
.B(n_400),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_541),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_513),
.B(n_417),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_561),
.B(n_300),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_587),
.B(n_417),
.Y(n_667)
);

AO22x2_ASAP7_75t_L g668 ( 
.A1(n_497),
.A2(n_254),
.B1(n_182),
.B2(n_193),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_469),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_565),
.B(n_181),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_510),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_517),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_469),
.B(n_181),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_572),
.B(n_177),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_472),
.B(n_193),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_533),
.B(n_183),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_524),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_519),
.B(n_417),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_L g679 ( 
.A1(n_480),
.A2(n_199),
.B(n_187),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_519),
.B(n_417),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_498),
.Y(n_681)
);

AOI22xp5_ASAP7_75t_L g682 ( 
.A1(n_514),
.A2(n_242),
.B1(n_259),
.B2(n_294),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_526),
.B(n_417),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_526),
.B(n_528),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_528),
.B(n_417),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_472),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_477),
.B(n_197),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_582),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_477),
.B(n_197),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_529),
.B(n_399),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_490),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_490),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_529),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_553),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_582),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_530),
.B(n_399),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_530),
.B(n_208),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_507),
.Y(n_698)
);

INVxp67_ASAP7_75t_L g699 ( 
.A(n_559),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_541),
.B(n_427),
.Y(n_700)
);

NAND3xp33_ASAP7_75t_L g701 ( 
.A(n_460),
.B(n_216),
.C(n_196),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_531),
.B(n_208),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_555),
.B(n_399),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_557),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_557),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_547),
.B(n_407),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_541),
.B(n_439),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_559),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_478),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_541),
.B(n_207),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_514),
.A2(n_230),
.B1(n_294),
.B2(n_262),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_559),
.B(n_195),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_525),
.B(n_198),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_537),
.B(n_213),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_523),
.B(n_229),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_582),
.B(n_407),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_569),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_582),
.B(n_407),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_582),
.B(n_411),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_582),
.B(n_411),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_588),
.B(n_411),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_542),
.B(n_414),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_574),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_574),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_483),
.A2(n_213),
.B1(n_230),
.B2(n_262),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_544),
.B(n_242),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_487),
.A2(n_418),
.B(n_422),
.C(n_289),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_576),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_563),
.B(n_414),
.Y(n_729)
);

BUFx8_ASAP7_75t_L g730 ( 
.A(n_449),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_576),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_481),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_483),
.A2(n_259),
.B1(n_254),
.B2(n_409),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_505),
.B(n_209),
.Y(n_734)
);

AOI221xp5_ASAP7_75t_L g735 ( 
.A1(n_476),
.A2(n_236),
.B1(n_241),
.B2(n_256),
.C(n_267),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_487),
.A2(n_496),
.B(n_589),
.C(n_580),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_564),
.B(n_212),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_566),
.B(n_285),
.C(n_225),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_579),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_579),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_563),
.B(n_414),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_581),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_453),
.B(n_419),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_453),
.B(n_419),
.Y(n_744)
);

INVx2_ASAP7_75t_SL g745 ( 
.A(n_483),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_464),
.B(n_236),
.Y(n_746)
);

INVx3_ASAP7_75t_L g747 ( 
.A(n_481),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_483),
.A2(n_409),
.B1(n_256),
.B2(n_288),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_453),
.B(n_465),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_461),
.B(n_428),
.Y(n_750)
);

OR2x2_ASAP7_75t_L g751 ( 
.A(n_471),
.B(n_241),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_584),
.B(n_428),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_478),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_L g754 ( 
.A(n_483),
.B(n_418),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_581),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_465),
.B(n_419),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_621),
.A2(n_504),
.B1(n_554),
.B2(n_560),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_648),
.Y(n_758)
);

O2A1O1Ixp5_ASAP7_75t_L g759 ( 
.A1(n_637),
.A2(n_578),
.B(n_503),
.C(n_484),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_754),
.A2(n_503),
.B(n_455),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_671),
.B(n_465),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_612),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_648),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_592),
.B(n_468),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_754),
.A2(n_503),
.B(n_455),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_616),
.B(n_571),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_592),
.B(n_468),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_614),
.A2(n_455),
.B(n_452),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_648),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_614),
.A2(n_522),
.B(n_452),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_595),
.B(n_468),
.Y(n_771)
);

AOI21x1_ASAP7_75t_L g772 ( 
.A1(n_635),
.A2(n_570),
.B(n_551),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_607),
.A2(n_522),
.B(n_452),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_667),
.A2(n_522),
.B(n_496),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_595),
.B(n_674),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_644),
.B(n_484),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_605),
.A2(n_570),
.B(n_551),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_652),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_681),
.B(n_549),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_606),
.A2(n_550),
.B(n_577),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_698),
.B(n_484),
.Y(n_781)
);

OAI21xp5_ASAP7_75t_L g782 ( 
.A1(n_611),
.A2(n_550),
.B(n_577),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_703),
.B(n_535),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_620),
.B(n_535),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_590),
.B(n_451),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_593),
.A2(n_535),
.B(n_548),
.Y(n_786)
);

AOI21x1_ASAP7_75t_L g787 ( 
.A1(n_635),
.A2(n_534),
.B(n_494),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_620),
.B(n_548),
.Y(n_788)
);

AOI21x1_ASAP7_75t_L g789 ( 
.A1(n_633),
.A2(n_634),
.B(n_729),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_625),
.B(n_548),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_617),
.A2(n_556),
.B1(n_571),
.B2(n_585),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_625),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_593),
.A2(n_500),
.B(n_583),
.Y(n_793)
);

A2O1A1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_662),
.A2(n_556),
.B(n_573),
.C(n_539),
.Y(n_794)
);

O2A1O1Ixp33_ASAP7_75t_SL g795 ( 
.A1(n_637),
.A2(n_267),
.B(n_288),
.C(n_289),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_646),
.A2(n_483),
.B1(n_451),
.B2(n_539),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_626),
.B(n_536),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_593),
.A2(n_500),
.B(n_583),
.Y(n_798)
);

AOI21x1_ASAP7_75t_L g799 ( 
.A1(n_633),
.A2(n_499),
.B(n_494),
.Y(n_799)
);

BUFx6f_ASAP7_75t_L g800 ( 
.A(n_602),
.Y(n_800)
);

CKINVDCx10_ASAP7_75t_R g801 ( 
.A(n_647),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_630),
.A2(n_585),
.B1(n_495),
.B2(n_538),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_602),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_652),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_599),
.B(n_536),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_700),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_672),
.B(n_491),
.Y(n_807)
);

INVx4_ASAP7_75t_L g808 ( 
.A(n_602),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_630),
.B(n_481),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_603),
.B(n_227),
.C(n_273),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_602),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_700),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_677),
.B(n_491),
.Y(n_813)
);

AO21x1_ASAP7_75t_L g814 ( 
.A1(n_736),
.A2(n_422),
.B(n_293),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_750),
.B(n_493),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_652),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_750),
.B(n_493),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_706),
.A2(n_500),
.B(n_481),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_646),
.B(n_499),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_722),
.A2(n_583),
.B(n_481),
.Y(n_820)
);

CKINVDCx6p67_ASAP7_75t_R g821 ( 
.A(n_751),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_630),
.B(n_500),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_SL g823 ( 
.A1(n_711),
.A2(n_293),
.B(n_297),
.C(n_534),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_591),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_643),
.B(n_515),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_709),
.B(n_536),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_713),
.A2(n_516),
.B(n_515),
.C(n_538),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_654),
.B(n_516),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_664),
.B(n_428),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_661),
.B(n_520),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_721),
.A2(n_684),
.B(n_618),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_615),
.B(n_500),
.Y(n_832)
);

AOI21x1_ASAP7_75t_L g833 ( 
.A1(n_634),
.A2(n_521),
.B(n_520),
.Y(n_833)
);

NOR3xp33_ASAP7_75t_L g834 ( 
.A(n_734),
.B(n_276),
.C(n_275),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_615),
.B(n_597),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_752),
.B(n_521),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_663),
.B(n_224),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_615),
.B(n_583),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_615),
.B(n_583),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_752),
.B(n_483),
.Y(n_840)
);

OAI21xp5_ASAP7_75t_L g841 ( 
.A1(n_716),
.A2(n_567),
.B(n_511),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_623),
.B(n_532),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_746),
.B(n_532),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_601),
.B(n_532),
.Y(n_844)
);

INVx4_ASAP7_75t_L g845 ( 
.A(n_688),
.Y(n_845)
);

O2A1O1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_640),
.A2(n_432),
.B(n_423),
.C(n_425),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_601),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_619),
.B(n_532),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_619),
.Y(n_849)
);

BUFx3_ASAP7_75t_L g850 ( 
.A(n_709),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_741),
.A2(n_567),
.B(n_511),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_688),
.A2(n_298),
.B1(n_235),
.B2(n_240),
.Y(n_852)
);

OAI321xp33_ASAP7_75t_L g853 ( 
.A1(n_676),
.A2(n_735),
.A3(n_701),
.B1(n_679),
.B2(n_738),
.C(n_682),
.Y(n_853)
);

NAND2x1p5_ASAP7_75t_L g854 ( 
.A(n_695),
.B(n_511),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_622),
.B(n_423),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_715),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_749),
.A2(n_567),
.B(n_511),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_718),
.A2(n_567),
.B(n_511),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_707),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_719),
.A2(n_567),
.B(n_406),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_746),
.B(n_409),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_695),
.B(n_409),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_720),
.A2(n_424),
.B(n_425),
.Y(n_863)
);

INVx11_ASAP7_75t_L g864 ( 
.A(n_730),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_628),
.A2(n_406),
.B(n_405),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_664),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_629),
.A2(n_406),
.B(n_415),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_622),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_745),
.A2(n_406),
.B(n_415),
.Y(n_869)
);

OAI21xp5_ASAP7_75t_L g870 ( 
.A1(n_642),
.A2(n_424),
.B(n_425),
.Y(n_870)
);

NOR2x1_ASAP7_75t_L g871 ( 
.A(n_613),
.B(n_432),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_745),
.A2(n_420),
.B(n_415),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_649),
.A2(n_424),
.B(n_421),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_627),
.B(n_433),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_743),
.A2(n_420),
.B(n_415),
.Y(n_875)
);

O2A1O1Ixp33_ASAP7_75t_L g876 ( 
.A1(n_670),
.A2(n_697),
.B(n_687),
.C(n_689),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_647),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_744),
.A2(n_420),
.B(n_421),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_756),
.A2(n_420),
.B(n_421),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_627),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_596),
.A2(n_277),
.B1(n_214),
.B2(n_226),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_631),
.B(n_426),
.Y(n_882)
);

AOI33xp33_ASAP7_75t_L g883 ( 
.A1(n_600),
.A2(n_361),
.A3(n_224),
.B1(n_433),
.B2(n_426),
.B3(n_271),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_669),
.A2(n_421),
.B(n_416),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_631),
.B(n_426),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_669),
.A2(n_421),
.B(n_416),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_691),
.A2(n_747),
.B(n_732),
.Y(n_887)
);

OAI21xp33_ASAP7_75t_L g888 ( 
.A1(n_610),
.A2(n_272),
.B(n_247),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_707),
.A2(n_433),
.B(n_426),
.C(n_278),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_636),
.B(n_433),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_636),
.B(n_416),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_651),
.B(n_598),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_651),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_691),
.A2(n_416),
.B(n_190),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_715),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_732),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_604),
.B(n_409),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_737),
.B(n_224),
.Y(n_898)
);

NOR2xp67_ASAP7_75t_SL g899 ( 
.A(n_732),
.B(n_258),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_608),
.B(n_416),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_710),
.B(n_248),
.Y(n_901)
);

OAI22xp5_ASAP7_75t_L g902 ( 
.A1(n_609),
.A2(n_286),
.B1(n_282),
.B2(n_253),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_710),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_693),
.A2(n_252),
.B1(n_409),
.B2(n_291),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_650),
.B(n_409),
.Y(n_905)
);

AO21x1_ASAP7_75t_L g906 ( 
.A1(n_702),
.A2(n_291),
.B(n_10),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_697),
.A2(n_291),
.B(n_224),
.C(n_16),
.Y(n_907)
);

AND2x2_ASAP7_75t_SL g908 ( 
.A(n_725),
.B(n_409),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_653),
.Y(n_909)
);

INVx11_ASAP7_75t_L g910 ( 
.A(n_730),
.Y(n_910)
);

AO21x1_ASAP7_75t_L g911 ( 
.A1(n_702),
.A2(n_6),
.B(n_15),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_712),
.A2(n_409),
.B(n_15),
.C(n_17),
.Y(n_912)
);

OAI22xp5_ASAP7_75t_L g913 ( 
.A1(n_657),
.A2(n_409),
.B1(n_150),
.B2(n_141),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_650),
.B(n_656),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_666),
.A2(n_139),
.B1(n_135),
.B2(n_131),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_747),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_747),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_656),
.B(n_6),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_655),
.A2(n_129),
.B(n_127),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_666),
.A2(n_126),
.B1(n_123),
.B2(n_116),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_694),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_641),
.B(n_17),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_686),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_699),
.B(n_18),
.C(n_22),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_704),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_668),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_708),
.A2(n_109),
.B1(n_108),
.B2(n_105),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_733),
.A2(n_103),
.B1(n_94),
.B2(n_84),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_641),
.B(n_22),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_645),
.B(n_692),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_624),
.A2(n_82),
.B(n_78),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_653),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_645),
.B(n_23),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_753),
.B(n_24),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_632),
.A2(n_77),
.B(n_76),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_638),
.A2(n_71),
.B(n_67),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_704),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_705),
.B(n_25),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_748),
.A2(n_65),
.B1(n_26),
.B2(n_29),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_639),
.A2(n_25),
.B(n_26),
.Y(n_940)
);

OAI22x1_ASAP7_75t_L g941 ( 
.A1(n_779),
.A2(n_594),
.B1(n_668),
.B2(n_730),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_775),
.B(n_668),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_757),
.A2(n_714),
.B1(n_726),
.B2(n_696),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_929),
.A2(n_726),
.B(n_714),
.C(n_727),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_800),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_856),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_760),
.A2(n_658),
.B(n_659),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_800),
.Y(n_948)
);

OAI22xp5_ASAP7_75t_L g949 ( 
.A1(n_908),
.A2(n_690),
.B1(n_660),
.B2(n_665),
.Y(n_949)
);

INVx1_ASAP7_75t_SL g950 ( 
.A(n_895),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_800),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_821),
.Y(n_952)
);

INVxp67_ASAP7_75t_L g953 ( 
.A(n_934),
.Y(n_953)
);

O2A1O1Ixp33_ASAP7_75t_L g954 ( 
.A1(n_929),
.A2(n_673),
.B(n_689),
.C(n_687),
.Y(n_954)
);

NAND2x1_ASAP7_75t_L g955 ( 
.A(n_808),
.B(n_717),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_792),
.B(n_717),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_834),
.A2(n_673),
.B(n_675),
.C(n_683),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_831),
.B(n_705),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_800),
.Y(n_959)
);

AOI22xp33_ASAP7_75t_L g960 ( 
.A1(n_834),
.A2(n_675),
.B1(n_742),
.B2(n_740),
.Y(n_960)
);

INVx4_ASAP7_75t_L g961 ( 
.A(n_811),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_806),
.B(n_728),
.Y(n_962)
);

INVx4_ASAP7_75t_SL g963 ( 
.A(n_811),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_765),
.A2(n_678),
.B(n_680),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_903),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_837),
.B(n_731),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_768),
.A2(n_770),
.B(n_776),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_762),
.B(n_755),
.Y(n_968)
);

OR2x2_ASAP7_75t_L g969 ( 
.A(n_903),
.B(n_739),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_783),
.A2(n_685),
.B(n_723),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_779),
.B(n_724),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_914),
.B(n_29),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_840),
.A2(n_31),
.B(n_36),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_810),
.A2(n_59),
.B1(n_37),
.B2(n_38),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_806),
.B(n_31),
.Y(n_975)
);

CKINVDCx10_ASAP7_75t_R g976 ( 
.A(n_801),
.Y(n_976)
);

NOR2xp67_ASAP7_75t_SL g977 ( 
.A(n_811),
.B(n_850),
.Y(n_977)
);

OAI21xp33_ASAP7_75t_L g978 ( 
.A1(n_898),
.A2(n_39),
.B(n_40),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_759),
.A2(n_41),
.B(n_42),
.Y(n_979)
);

INVx5_ASAP7_75t_L g980 ( 
.A(n_811),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_812),
.B(n_45),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_812),
.B(n_46),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_787),
.A2(n_50),
.B(n_51),
.Y(n_983)
);

CKINVDCx6p67_ASAP7_75t_R g984 ( 
.A(n_877),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_785),
.B(n_50),
.C(n_51),
.Y(n_985)
);

CKINVDCx6p67_ASAP7_75t_R g986 ( 
.A(n_932),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_868),
.Y(n_987)
);

HB1xp67_ASAP7_75t_L g988 ( 
.A(n_859),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_R g989 ( 
.A(n_826),
.B(n_785),
.Y(n_989)
);

O2A1O1Ixp5_ASAP7_75t_SL g990 ( 
.A1(n_835),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_859),
.B(n_797),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_815),
.A2(n_817),
.B(n_798),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_793),
.A2(n_774),
.B(n_773),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_866),
.B(n_871),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_853),
.B(n_810),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_836),
.B(n_829),
.Y(n_996)
);

OAI22x1_ASAP7_75t_L g997 ( 
.A1(n_926),
.A2(n_934),
.B1(n_805),
.B2(n_797),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_764),
.A2(n_771),
.B(n_767),
.Y(n_998)
);

NOR3xp33_ASAP7_75t_SL g999 ( 
.A(n_909),
.B(n_805),
.C(n_888),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_866),
.B(n_826),
.Y(n_1000)
);

OR2x6_ASAP7_75t_L g1001 ( 
.A(n_808),
.B(n_866),
.Y(n_1001)
);

AO22x1_ASAP7_75t_L g1002 ( 
.A1(n_924),
.A2(n_922),
.B1(n_933),
.B2(n_918),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_863),
.A2(n_820),
.B(n_818),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_835),
.A2(n_782),
.B(n_858),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_893),
.Y(n_1005)
);

OAI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_908),
.A2(n_794),
.B1(n_843),
.B2(n_845),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_843),
.A2(n_845),
.B1(n_796),
.B2(n_880),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_824),
.B(n_847),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_912),
.A2(n_907),
.B(n_924),
.C(n_795),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_901),
.B(n_829),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_SL g1011 ( 
.A1(n_899),
.A2(n_919),
.B(n_780),
.C(n_841),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_809),
.A2(n_822),
.B(n_781),
.Y(n_1012)
);

NAND2x1_ASAP7_75t_L g1013 ( 
.A(n_896),
.B(n_803),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_852),
.B(n_881),
.Y(n_1014)
);

AO32x2_ASAP7_75t_L g1015 ( 
.A1(n_913),
.A2(n_791),
.A3(n_939),
.B1(n_802),
.B2(n_904),
.Y(n_1015)
);

AO21x1_ASAP7_75t_L g1016 ( 
.A1(n_766),
.A2(n_822),
.B(n_809),
.Y(n_1016)
);

AOI221xp5_ASAP7_75t_L g1017 ( 
.A1(n_902),
.A2(n_823),
.B1(n_795),
.B2(n_906),
.C(n_940),
.Y(n_1017)
);

O2A1O1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_766),
.A2(n_823),
.B(n_889),
.C(n_938),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_864),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_799),
.A2(n_833),
.B(n_772),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_849),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_866),
.B(n_883),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_784),
.A2(n_790),
.B(n_788),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_876),
.A2(n_930),
.B(n_892),
.C(n_761),
.Y(n_1024)
);

O2A1O1Ixp5_ASAP7_75t_L g1025 ( 
.A1(n_814),
.A2(n_861),
.B(n_842),
.C(n_789),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_915),
.A2(n_920),
.B(n_846),
.C(n_905),
.Y(n_1026)
);

A2O1A1Ixp33_ASAP7_75t_SL g1027 ( 
.A1(n_894),
.A2(n_870),
.B(n_873),
.C(n_803),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_807),
.A2(n_813),
.B(n_862),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_916),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_911),
.Y(n_1030)
);

INVx4_ASAP7_75t_L g1031 ( 
.A(n_916),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_937),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_910),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_923),
.B(n_925),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_923),
.B(n_855),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_921),
.B(n_830),
.Y(n_1036)
);

HB1xp67_ASAP7_75t_L g1037 ( 
.A(n_921),
.Y(n_1037)
);

AO22x1_ASAP7_75t_L g1038 ( 
.A1(n_927),
.A2(n_928),
.B1(n_896),
.B2(n_916),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_819),
.B(n_828),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_825),
.B(n_758),
.Y(n_1040)
);

BUFx12f_ASAP7_75t_L g1041 ( 
.A(n_916),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_917),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_763),
.Y(n_1043)
);

O2A1O1Ixp5_ASAP7_75t_L g1044 ( 
.A1(n_861),
.A2(n_838),
.B(n_832),
.C(n_839),
.Y(n_1044)
);

A2O1A1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_777),
.A2(n_869),
.B(n_872),
.C(n_887),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_862),
.A2(n_786),
.B(n_832),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_900),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_838),
.A2(n_839),
.B(n_848),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_921),
.B(n_769),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_874),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_778),
.B(n_804),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_921),
.B(n_816),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_897),
.A2(n_917),
.B1(n_844),
.B2(n_890),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_917),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_917),
.B(n_897),
.Y(n_1055)
);

AND2x4_ASAP7_75t_L g1056 ( 
.A(n_827),
.B(n_882),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_885),
.B(n_891),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_865),
.A2(n_867),
.B1(n_875),
.B2(n_879),
.Y(n_1058)
);

NAND2x1_ASAP7_75t_L g1059 ( 
.A(n_884),
.B(n_886),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_878),
.B(n_854),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_860),
.A2(n_931),
.B(n_935),
.C(n_936),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_854),
.B(n_857),
.Y(n_1062)
);

XOR2xp5_ASAP7_75t_L g1063 ( 
.A(n_851),
.B(n_451),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_SL g1064 ( 
.A1(n_899),
.A2(n_674),
.B(n_713),
.C(n_644),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_929),
.A2(n_834),
.B1(n_810),
.B2(n_644),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_792),
.B(n_806),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_868),
.Y(n_1067)
);

INVxp33_ASAP7_75t_SL g1068 ( 
.A(n_826),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_760),
.A2(n_593),
.B(n_765),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_856),
.Y(n_1070)
);

BUFx12f_ASAP7_75t_L g1071 ( 
.A(n_909),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_850),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_760),
.A2(n_593),
.B(n_765),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_775),
.B(n_489),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_929),
.A2(n_834),
.B(n_637),
.C(n_644),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_800),
.Y(n_1076)
);

BUFx3_ASAP7_75t_L g1077 ( 
.A(n_850),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_909),
.B(n_478),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_775),
.B(n_489),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_856),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_800),
.Y(n_1081)
);

HB1xp67_ASAP7_75t_L g1082 ( 
.A(n_946),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_1016),
.A2(n_1006),
.A3(n_1004),
.B(n_943),
.Y(n_1083)
);

NOR2xp67_ASAP7_75t_L g1084 ( 
.A(n_1080),
.B(n_1070),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1032),
.Y(n_1085)
);

OAI21x1_ASAP7_75t_L g1086 ( 
.A1(n_1020),
.A2(n_1073),
.B(n_1069),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_995),
.A2(n_1025),
.B(n_1075),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1088)
);

INVx2_ASAP7_75t_SL g1089 ( 
.A(n_1072),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_993),
.A2(n_1046),
.B(n_1048),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_1077),
.Y(n_1091)
);

OAI21x1_ASAP7_75t_L g1092 ( 
.A1(n_964),
.A2(n_947),
.B(n_967),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_992),
.A2(n_998),
.B(n_1023),
.Y(n_1093)
);

INVxp67_ASAP7_75t_L g1094 ( 
.A(n_946),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1065),
.A2(n_1010),
.B1(n_1014),
.B2(n_971),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_984),
.Y(n_1096)
);

NAND3xp33_ASAP7_75t_L g1097 ( 
.A(n_974),
.B(n_978),
.C(n_944),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_1066),
.B(n_994),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1026),
.A2(n_1024),
.B(n_1006),
.Y(n_1099)
);

AOI221xp5_ASAP7_75t_L g1100 ( 
.A1(n_941),
.A2(n_953),
.B1(n_1009),
.B2(n_997),
.C(n_1002),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1021),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1041),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_954),
.A2(n_1018),
.B(n_957),
.C(n_1064),
.Y(n_1103)
);

O2A1O1Ixp33_ASAP7_75t_SL g1104 ( 
.A1(n_1011),
.A2(n_1022),
.B(n_942),
.C(n_979),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1003),
.A2(n_1079),
.B(n_1074),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1066),
.B(n_994),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_972),
.A2(n_943),
.B(n_979),
.C(n_1017),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_SL g1108 ( 
.A(n_1068),
.B(n_977),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1027),
.A2(n_1028),
.B(n_1039),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1012),
.A2(n_991),
.B(n_999),
.C(n_1030),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_996),
.B(n_966),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_958),
.A2(n_1061),
.B(n_1045),
.Y(n_1112)
);

AOI21x1_ASAP7_75t_L g1113 ( 
.A1(n_1062),
.A2(n_1060),
.B(n_1038),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1008),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_1078),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_969),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_962),
.B(n_1050),
.Y(n_1117)
);

NAND3xp33_ASAP7_75t_L g1118 ( 
.A(n_985),
.B(n_973),
.C(n_989),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1035),
.A2(n_1060),
.B(n_970),
.Y(n_1119)
);

OAI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_949),
.A2(n_1044),
.B(n_1056),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1059),
.A2(n_983),
.B(n_1058),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1036),
.A2(n_1057),
.B(n_1053),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1063),
.A2(n_981),
.B1(n_962),
.B2(n_988),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1047),
.B(n_950),
.Y(n_1124)
);

INVxp67_ASAP7_75t_L g1125 ( 
.A(n_950),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1035),
.B(n_975),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_1019),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_949),
.A2(n_1056),
.B(n_1007),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_982),
.A2(n_1000),
.B(n_965),
.C(n_981),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_945),
.Y(n_1130)
);

AO32x2_ASAP7_75t_L g1131 ( 
.A1(n_990),
.A2(n_1081),
.A3(n_961),
.B1(n_1015),
.B2(n_1031),
.Y(n_1131)
);

OAI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1040),
.A2(n_960),
.B(n_1034),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_980),
.A2(n_1052),
.B(n_1049),
.Y(n_1133)
);

BUFx10_ASAP7_75t_L g1134 ( 
.A(n_1033),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_987),
.Y(n_1135)
);

AOI221x1_ASAP7_75t_L g1136 ( 
.A1(n_1015),
.A2(n_1055),
.B1(n_968),
.B2(n_956),
.C(n_1076),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_952),
.Y(n_1137)
);

INVx2_ASAP7_75t_SL g1138 ( 
.A(n_986),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1054),
.B(n_980),
.Y(n_1139)
);

O2A1O1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1005),
.A2(n_1067),
.B(n_1037),
.C(n_1043),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_980),
.A2(n_1001),
.B(n_955),
.Y(n_1141)
);

AOI221x1_ASAP7_75t_L g1142 ( 
.A1(n_1015),
.A2(n_1076),
.B1(n_951),
.B2(n_961),
.C(n_1081),
.Y(n_1142)
);

NAND2x1p5_ASAP7_75t_L g1143 ( 
.A(n_980),
.B(n_1031),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_1029),
.B(n_945),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_1051),
.B(n_1001),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_951),
.B(n_1001),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1013),
.A2(n_1042),
.B(n_948),
.Y(n_1147)
);

O2A1O1Ixp33_ASAP7_75t_L g1148 ( 
.A1(n_1071),
.A2(n_963),
.B(n_1042),
.C(n_1029),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_1029),
.B(n_945),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_963),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_948),
.A2(n_959),
.B(n_963),
.Y(n_1151)
);

OR2x6_ASAP7_75t_L g1152 ( 
.A(n_948),
.B(n_959),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_959),
.A2(n_1075),
.B(n_1065),
.C(n_1014),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_976),
.B(n_1074),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1016),
.A2(n_814),
.A3(n_1006),
.B(n_1004),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_995),
.A2(n_603),
.B1(n_834),
.B2(n_1065),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_995),
.A2(n_1025),
.B(n_1004),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_995),
.A2(n_1025),
.B(n_1004),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_1001),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_984),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1070),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1162)
);

AO21x2_ASAP7_75t_L g1163 ( 
.A1(n_1011),
.A2(n_1004),
.B(n_1003),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_1065),
.A2(n_1079),
.B1(n_1074),
.B2(n_995),
.Y(n_1164)
);

OAI22x1_ASAP7_75t_L g1165 ( 
.A1(n_995),
.A2(n_779),
.B1(n_974),
.B2(n_603),
.Y(n_1165)
);

BUFx4f_ASAP7_75t_L g1166 ( 
.A(n_984),
.Y(n_1166)
);

AOI21x1_ASAP7_75t_SL g1167 ( 
.A1(n_942),
.A2(n_597),
.B(n_972),
.Y(n_1167)
);

OAI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_995),
.A2(n_1025),
.B(n_1004),
.Y(n_1168)
);

AOI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1002),
.A2(n_835),
.B(n_1004),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_962),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1020),
.A2(n_1073),
.B(n_1069),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1065),
.A2(n_603),
.B1(n_323),
.B2(n_328),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_995),
.A2(n_1025),
.B(n_1004),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_946),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1177)
);

NOR3xp33_ASAP7_75t_L g1178 ( 
.A(n_995),
.B(n_603),
.C(n_466),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_1019),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_1065),
.B(n_590),
.Y(n_1181)
);

NAND3xp33_ASAP7_75t_L g1182 ( 
.A(n_1065),
.B(n_674),
.C(n_644),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1183)
);

BUFx3_ASAP7_75t_L g1184 ( 
.A(n_1072),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1032),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_1080),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1188)
);

AOI221x1_ASAP7_75t_L g1189 ( 
.A1(n_997),
.A2(n_834),
.B1(n_1006),
.B2(n_1026),
.C(n_979),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1032),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1020),
.A2(n_1073),
.B(n_1069),
.Y(n_1191)
);

AO31x2_ASAP7_75t_L g1192 ( 
.A1(n_1016),
.A2(n_814),
.A3(n_1006),
.B(n_1004),
.Y(n_1192)
);

INVx3_ASAP7_75t_L g1193 ( 
.A(n_1031),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1025),
.A2(n_1004),
.B(n_979),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1196)
);

AOI221x1_ASAP7_75t_L g1197 ( 
.A1(n_997),
.A2(n_834),
.B1(n_1006),
.B2(n_1026),
.C(n_979),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1065),
.B(n_590),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1016),
.A2(n_814),
.A3(n_1006),
.B(n_1004),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1032),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_946),
.B(n_856),
.Y(n_1201)
);

NOR2x1_ASAP7_75t_SL g1202 ( 
.A(n_980),
.B(n_1001),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1016),
.A2(n_814),
.A3(n_1006),
.B(n_1004),
.Y(n_1203)
);

NAND2x1p5_ASAP7_75t_L g1204 ( 
.A(n_980),
.B(n_808),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_981),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1065),
.B(n_590),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_995),
.A2(n_603),
.B(n_681),
.C(n_644),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1210)
);

AOI221xp5_ASAP7_75t_SL g1211 ( 
.A1(n_995),
.A2(n_1065),
.B1(n_978),
.B2(n_929),
.C(n_1075),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_962),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_953),
.B(n_603),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1020),
.A2(n_1073),
.B(n_1069),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1074),
.B(n_1079),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_952),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_976),
.Y(n_1218)
);

NOR2xp67_ASAP7_75t_L g1219 ( 
.A(n_1080),
.B(n_753),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_962),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_967),
.A2(n_1073),
.B(n_1069),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1178),
.A2(n_1156),
.B1(n_1182),
.B2(n_1165),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1082),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_1175),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1101),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1182),
.A2(n_1097),
.B1(n_1099),
.B2(n_1164),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1102),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_1218),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1185),
.Y(n_1229)
);

CKINVDCx20_ASAP7_75t_R g1230 ( 
.A(n_1115),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_SL g1231 ( 
.A1(n_1172),
.A2(n_1154),
.B1(n_1213),
.B2(n_1123),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_1152),
.Y(n_1232)
);

BUFx2_ASAP7_75t_SL g1233 ( 
.A(n_1084),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_L g1234 ( 
.A1(n_1097),
.A2(n_1095),
.B1(n_1181),
.B2(n_1206),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1184),
.Y(n_1235)
);

OAI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1153),
.A2(n_1209),
.B1(n_1177),
.B2(n_1174),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1190),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1200),
.Y(n_1238)
);

INVx5_ASAP7_75t_L g1239 ( 
.A(n_1152),
.Y(n_1239)
);

INVx1_ASAP7_75t_SL g1240 ( 
.A(n_1201),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1159),
.B(n_1139),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_1127),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1111),
.B(n_1126),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_1102),
.Y(n_1244)
);

OAI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1189),
.A2(n_1197),
.B1(n_1164),
.B2(n_1177),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_1116),
.Y(n_1246)
);

OAI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1099),
.A2(n_1187),
.B1(n_1194),
.B2(n_1210),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_1179),
.Y(n_1248)
);

OAI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1088),
.A2(n_1208),
.B1(n_1196),
.B2(n_1216),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1124),
.A2(n_1111),
.B1(n_1108),
.B2(n_1142),
.Y(n_1250)
);

BUFx12f_ASAP7_75t_L g1251 ( 
.A(n_1134),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1135),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1117),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1170),
.Y(n_1254)
);

BUFx8_ASAP7_75t_L g1255 ( 
.A(n_1102),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1114),
.Y(n_1256)
);

OAI22xp5_ASAP7_75t_L g1257 ( 
.A1(n_1107),
.A2(n_1110),
.B1(n_1198),
.B2(n_1186),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1118),
.A2(n_1100),
.B1(n_1129),
.B2(n_1125),
.Y(n_1258)
);

INVx3_ASAP7_75t_SL g1259 ( 
.A(n_1160),
.Y(n_1259)
);

INVx4_ASAP7_75t_SL g1260 ( 
.A(n_1152),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1212),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1118),
.A2(n_1094),
.B1(n_1159),
.B2(n_1219),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_SL g1263 ( 
.A(n_1134),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1220),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1217),
.Y(n_1265)
);

INVx4_ASAP7_75t_L g1266 ( 
.A(n_1159),
.Y(n_1266)
);

INVx3_ASAP7_75t_SL g1267 ( 
.A(n_1089),
.Y(n_1267)
);

AND2x4_ASAP7_75t_SL g1268 ( 
.A(n_1205),
.B(n_1098),
.Y(n_1268)
);

BUFx4_ASAP7_75t_R g1269 ( 
.A(n_1205),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1096),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1091),
.Y(n_1271)
);

INVxp67_ASAP7_75t_SL g1272 ( 
.A(n_1105),
.Y(n_1272)
);

OAI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1108),
.A2(n_1087),
.B1(n_1128),
.B2(n_1159),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1211),
.B(n_1098),
.Y(n_1274)
);

INVx6_ASAP7_75t_L g1275 ( 
.A(n_1217),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1161),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_L g1277 ( 
.A1(n_1087),
.A2(n_1106),
.B1(n_1145),
.B2(n_1120),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1144),
.Y(n_1278)
);

OAI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1136),
.A2(n_1132),
.B1(n_1157),
.B2(n_1173),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1140),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_SL g1281 ( 
.A1(n_1106),
.A2(n_1137),
.B1(n_1138),
.B2(n_1146),
.Y(n_1281)
);

NAND2x1p5_ASAP7_75t_L g1282 ( 
.A(n_1193),
.B(n_1166),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1120),
.A2(n_1132),
.B1(n_1168),
.B2(n_1158),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1211),
.B(n_1158),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_SL g1285 ( 
.A1(n_1157),
.A2(n_1173),
.B1(n_1168),
.B2(n_1195),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1163),
.A2(n_1195),
.B1(n_1112),
.B2(n_1093),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1163),
.A2(n_1093),
.B1(n_1109),
.B2(n_1119),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1103),
.A2(n_1166),
.B1(n_1133),
.B2(n_1113),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1169),
.A2(n_1193),
.B1(n_1204),
.B2(n_1150),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1149),
.Y(n_1290)
);

OAI22xp5_ASAP7_75t_L g1291 ( 
.A1(n_1204),
.A2(n_1143),
.B1(n_1148),
.B2(n_1141),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1122),
.A2(n_1221),
.B1(n_1176),
.B2(n_1183),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_1130),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1202),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1083),
.B(n_1104),
.Y(n_1295)
);

INVx6_ASAP7_75t_L g1296 ( 
.A(n_1151),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1147),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1131),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1162),
.A2(n_1215),
.B1(n_1207),
.B2(n_1188),
.Y(n_1299)
);

BUFx2_ASAP7_75t_SL g1300 ( 
.A(n_1180),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1083),
.A2(n_1090),
.B1(n_1092),
.B2(n_1192),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1121),
.A2(n_1171),
.B1(n_1086),
.B2(n_1191),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1131),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1131),
.Y(n_1304)
);

INVx5_ASAP7_75t_L g1305 ( 
.A(n_1167),
.Y(n_1305)
);

CKINVDCx6p67_ASAP7_75t_R g1306 ( 
.A(n_1155),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1083),
.Y(n_1307)
);

INVxp67_ASAP7_75t_SL g1308 ( 
.A(n_1214),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1192),
.A2(n_1156),
.B1(n_603),
.B2(n_1065),
.Y(n_1309)
);

BUFx8_ASAP7_75t_L g1310 ( 
.A(n_1199),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1199),
.A2(n_603),
.B1(n_437),
.B2(n_1182),
.Y(n_1311)
);

BUFx12f_ASAP7_75t_L g1312 ( 
.A(n_1199),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1203),
.B(n_1213),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1203),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1156),
.A2(n_603),
.B1(n_1065),
.B2(n_1095),
.Y(n_1315)
);

BUFx12f_ASAP7_75t_L g1316 ( 
.A(n_1134),
.Y(n_1316)
);

BUFx2_ASAP7_75t_L g1317 ( 
.A(n_1082),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1178),
.A2(n_603),
.B1(n_1156),
.B2(n_1182),
.Y(n_1318)
);

OAI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1095),
.A2(n_974),
.B1(n_1097),
.B2(n_1165),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1178),
.A2(n_1165),
.B1(n_1156),
.B2(n_995),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_SL g1321 ( 
.A1(n_1182),
.A2(n_603),
.B1(n_437),
.B2(n_1097),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1156),
.A2(n_603),
.B1(n_1065),
.B2(n_1095),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1159),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1178),
.A2(n_603),
.B1(n_1156),
.B2(n_1182),
.Y(n_1324)
);

BUFx8_ASAP7_75t_SL g1325 ( 
.A(n_1218),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1218),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1218),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1082),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1085),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1178),
.A2(n_603),
.B1(n_1156),
.B2(n_1182),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1213),
.B(n_1178),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1201),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1156),
.A2(n_603),
.B1(n_1065),
.B2(n_1095),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1178),
.A2(n_603),
.B1(n_1156),
.B2(n_1182),
.Y(n_1334)
);

OAI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1095),
.A2(n_974),
.B1(n_1097),
.B2(n_1165),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1178),
.A2(n_1165),
.B1(n_1156),
.B2(n_995),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1159),
.Y(n_1337)
);

BUFx12f_ASAP7_75t_L g1338 ( 
.A(n_1134),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1156),
.A2(n_603),
.B1(n_1065),
.B2(n_1095),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1213),
.B(n_903),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1178),
.A2(n_1165),
.B1(n_1156),
.B2(n_995),
.Y(n_1341)
);

AND2x4_ASAP7_75t_L g1342 ( 
.A(n_1294),
.B(n_1337),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1223),
.Y(n_1343)
);

NOR2xp33_ASAP7_75t_L g1344 ( 
.A(n_1331),
.B(n_1240),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1307),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1315),
.A2(n_1322),
.B1(n_1339),
.B2(n_1333),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1314),
.A2(n_1295),
.A3(n_1309),
.B(n_1298),
.Y(n_1347)
);

OAI222xp33_ASAP7_75t_L g1348 ( 
.A1(n_1321),
.A2(n_1226),
.B1(n_1311),
.B2(n_1318),
.C1(n_1324),
.C2(n_1330),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1325),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1302),
.A2(n_1292),
.B(n_1299),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1306),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_SL g1352 ( 
.A1(n_1249),
.A2(n_1236),
.B(n_1273),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1247),
.B(n_1243),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1323),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1224),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1313),
.B(n_1226),
.Y(n_1356)
);

NAND2xp5_ASAP7_75t_L g1357 ( 
.A(n_1247),
.B(n_1284),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1310),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1310),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1312),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1317),
.Y(n_1361)
);

HB1xp67_ASAP7_75t_L g1362 ( 
.A(n_1328),
.Y(n_1362)
);

OR2x2_ASAP7_75t_L g1363 ( 
.A(n_1283),
.B(n_1274),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1246),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1321),
.A2(n_1334),
.B1(n_1319),
.B2(n_1335),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1303),
.Y(n_1366)
);

BUFx3_ASAP7_75t_L g1367 ( 
.A(n_1241),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1272),
.Y(n_1368)
);

AND2x4_ASAP7_75t_L g1369 ( 
.A(n_1260),
.B(n_1266),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1304),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1256),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1272),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1279),
.Y(n_1373)
);

AND2x4_ASAP7_75t_L g1374 ( 
.A(n_1260),
.B(n_1266),
.Y(n_1374)
);

OR2x6_ASAP7_75t_L g1375 ( 
.A(n_1300),
.B(n_1288),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1225),
.Y(n_1376)
);

NAND2x1_ASAP7_75t_L g1377 ( 
.A(n_1296),
.B(n_1292),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1287),
.A2(n_1286),
.B(n_1299),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1290),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1237),
.Y(n_1380)
);

HB1xp67_ASAP7_75t_L g1381 ( 
.A(n_1332),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1238),
.Y(n_1382)
);

NOR2xp33_ASAP7_75t_L g1383 ( 
.A(n_1231),
.B(n_1340),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1311),
.B(n_1285),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1329),
.Y(n_1385)
);

AOI21xp5_ASAP7_75t_SL g1386 ( 
.A1(n_1273),
.A2(n_1257),
.B(n_1291),
.Y(n_1386)
);

INVx2_ASAP7_75t_L g1387 ( 
.A(n_1229),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1245),
.A2(n_1289),
.B(n_1308),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1302),
.A2(n_1287),
.B(n_1286),
.Y(n_1389)
);

OR2x2_ASAP7_75t_L g1390 ( 
.A(n_1250),
.B(n_1258),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1252),
.Y(n_1391)
);

AOI21xp33_ASAP7_75t_L g1392 ( 
.A1(n_1319),
.A2(n_1335),
.B(n_1336),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1245),
.Y(n_1393)
);

AO21x1_ASAP7_75t_L g1394 ( 
.A1(n_1250),
.A2(n_1280),
.B(n_1289),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1305),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1305),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1222),
.A2(n_1341),
.B(n_1336),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1305),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1277),
.A2(n_1241),
.B(n_1320),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1234),
.B(n_1341),
.Y(n_1400)
);

BUFx6f_ASAP7_75t_L g1401 ( 
.A(n_1232),
.Y(n_1401)
);

BUFx2_ASAP7_75t_SL g1402 ( 
.A(n_1297),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1320),
.B(n_1253),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1262),
.A2(n_1276),
.B1(n_1263),
.B2(n_1338),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1301),
.B(n_1264),
.Y(n_1405)
);

AO21x1_ASAP7_75t_L g1406 ( 
.A1(n_1278),
.A2(n_1261),
.B(n_1254),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1296),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1281),
.A2(n_1268),
.B(n_1232),
.C(n_1239),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1296),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1282),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1282),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1269),
.A2(n_1263),
.B(n_1293),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1233),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1227),
.Y(n_1414)
);

INVx4_ASAP7_75t_L g1415 ( 
.A(n_1244),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1244),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1365),
.A2(n_1275),
.B1(n_1267),
.B2(n_1271),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1384),
.B(n_1259),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1384),
.B(n_1356),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1346),
.A2(n_1275),
.B1(n_1316),
.B2(n_1251),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_SL g1421 ( 
.A1(n_1348),
.A2(n_1265),
.B(n_1275),
.C(n_1255),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1392),
.A2(n_1267),
.B(n_1259),
.C(n_1235),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1353),
.B(n_1255),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1363),
.B(n_1242),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_SL g1425 ( 
.A(n_1375),
.B(n_1270),
.Y(n_1425)
);

INVx3_ASAP7_75t_L g1426 ( 
.A(n_1342),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1344),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1356),
.B(n_1248),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1360),
.B(n_1230),
.Y(n_1429)
);

NAND4xp25_ASAP7_75t_L g1430 ( 
.A(n_1392),
.B(n_1228),
.C(n_1326),
.D(n_1327),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1360),
.B(n_1228),
.Y(n_1431)
);

OAI22xp5_ASAP7_75t_L g1432 ( 
.A1(n_1390),
.A2(n_1383),
.B1(n_1404),
.B2(n_1400),
.Y(n_1432)
);

AND2x2_ASAP7_75t_SL g1433 ( 
.A(n_1390),
.B(n_1397),
.Y(n_1433)
);

NOR2x1_ASAP7_75t_L g1434 ( 
.A(n_1402),
.B(n_1352),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1363),
.B(n_1381),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1373),
.B(n_1376),
.Y(n_1436)
);

AOI221xp5_ASAP7_75t_L g1437 ( 
.A1(n_1348),
.A2(n_1352),
.B1(n_1400),
.B2(n_1386),
.C(n_1393),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1376),
.B(n_1382),
.Y(n_1438)
);

A2O1A1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1399),
.A2(n_1353),
.B(n_1377),
.C(n_1357),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1403),
.B(n_1397),
.Y(n_1440)
);

AO21x2_ASAP7_75t_L g1441 ( 
.A1(n_1394),
.A2(n_1389),
.B(n_1350),
.Y(n_1441)
);

AOI221xp5_ASAP7_75t_L g1442 ( 
.A1(n_1386),
.A2(n_1394),
.B1(n_1403),
.B2(n_1361),
.C(n_1364),
.Y(n_1442)
);

NAND4xp25_ASAP7_75t_L g1443 ( 
.A(n_1361),
.B(n_1413),
.C(n_1391),
.D(n_1380),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1382),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1343),
.B(n_1355),
.Y(n_1445)
);

A2O1A1Ixp33_ASAP7_75t_L g1446 ( 
.A1(n_1399),
.A2(n_1402),
.B(n_1408),
.C(n_1368),
.Y(n_1446)
);

AOI211xp5_ASAP7_75t_L g1447 ( 
.A1(n_1358),
.A2(n_1359),
.B(n_1351),
.C(n_1411),
.Y(n_1447)
);

NAND3xp33_ASAP7_75t_L g1448 ( 
.A(n_1397),
.B(n_1407),
.C(n_1409),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1368),
.A2(n_1372),
.B(n_1350),
.C(n_1389),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1362),
.B(n_1379),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1397),
.A2(n_1359),
.B1(n_1358),
.B2(n_1375),
.Y(n_1451)
);

NAND2x1_ASAP7_75t_L g1452 ( 
.A(n_1375),
.B(n_1369),
.Y(n_1452)
);

AND2x6_ASAP7_75t_L g1453 ( 
.A(n_1369),
.B(n_1374),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_R g1454 ( 
.A(n_1349),
.B(n_1415),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1385),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1354),
.Y(n_1456)
);

OAI21xp5_ASAP7_75t_L g1457 ( 
.A1(n_1412),
.A2(n_1395),
.B(n_1396),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1347),
.B(n_1366),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1433),
.A2(n_1388),
.B1(n_1378),
.B2(n_1401),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1452),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1458),
.B(n_1378),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1437),
.A2(n_1378),
.B1(n_1388),
.B2(n_1406),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1458),
.B(n_1378),
.Y(n_1463)
);

INVx4_ASAP7_75t_R g1464 ( 
.A(n_1456),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1423),
.B(n_1410),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1429),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1444),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1457),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1432),
.A2(n_1378),
.B1(n_1388),
.B2(n_1406),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1441),
.B(n_1388),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1444),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1441),
.B(n_1449),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1449),
.B(n_1345),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1440),
.B(n_1347),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1455),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1438),
.B(n_1347),
.Y(n_1476)
);

BUFx3_ASAP7_75t_L g1477 ( 
.A(n_1453),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1435),
.B(n_1347),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1438),
.B(n_1347),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1442),
.A2(n_1367),
.B1(n_1405),
.B2(n_1396),
.C(n_1398),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1445),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1434),
.A2(n_1391),
.B1(n_1371),
.B2(n_1387),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1440),
.B(n_1371),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1448),
.B(n_1370),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1433),
.A2(n_1419),
.B1(n_1417),
.B2(n_1425),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1453),
.Y(n_1486)
);

AND2x4_ASAP7_75t_SL g1487 ( 
.A(n_1460),
.B(n_1401),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1461),
.B(n_1463),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1471),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1467),
.Y(n_1490)
);

OAI21xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1462),
.A2(n_1443),
.B(n_1418),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1471),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1477),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1467),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1467),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1461),
.B(n_1426),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1461),
.B(n_1426),
.Y(n_1497)
);

NAND2x1_ASAP7_75t_L g1498 ( 
.A(n_1464),
.B(n_1453),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1459),
.A2(n_1421),
.B(n_1446),
.Y(n_1499)
);

INVx5_ASAP7_75t_L g1500 ( 
.A(n_1472),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1477),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_SL g1502 ( 
.A(n_1477),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1483),
.B(n_1439),
.Y(n_1503)
);

AND2x2_ASAP7_75t_SL g1504 ( 
.A(n_1468),
.B(n_1469),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1486),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1483),
.B(n_1424),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1474),
.B(n_1450),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1475),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1462),
.A2(n_1430),
.B1(n_1427),
.B2(n_1420),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1480),
.A2(n_1428),
.B1(n_1451),
.B2(n_1429),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1474),
.B(n_1439),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1476),
.B(n_1436),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1488),
.B(n_1472),
.Y(n_1513)
);

AOI22xp33_ASAP7_75t_L g1514 ( 
.A1(n_1504),
.A2(n_1509),
.B1(n_1510),
.B2(n_1491),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1508),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1488),
.B(n_1472),
.Y(n_1516)
);

HB1xp67_ASAP7_75t_L g1517 ( 
.A(n_1490),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1500),
.B(n_1468),
.Y(n_1518)
);

NAND2x1p5_ASAP7_75t_L g1519 ( 
.A(n_1500),
.B(n_1470),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1511),
.B(n_1476),
.Y(n_1520)
);

INVx4_ASAP7_75t_L g1521 ( 
.A(n_1500),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1511),
.B(n_1476),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1500),
.B(n_1496),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1490),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1500),
.B(n_1468),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1500),
.B(n_1496),
.Y(n_1526)
);

INVx3_ASAP7_75t_L g1527 ( 
.A(n_1500),
.Y(n_1527)
);

AND2x4_ASAP7_75t_L g1528 ( 
.A(n_1500),
.B(n_1486),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1489),
.B(n_1484),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1503),
.B(n_1479),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1503),
.B(n_1479),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1508),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1500),
.B(n_1496),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1494),
.Y(n_1534)
);

AND2x4_ASAP7_75t_SL g1535 ( 
.A(n_1501),
.B(n_1460),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1501),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1495),
.Y(n_1537)
);

OR2x2_ASAP7_75t_L g1538 ( 
.A(n_1489),
.B(n_1484),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1489),
.B(n_1484),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1497),
.B(n_1473),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1487),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1492),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1536),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1514),
.B(n_1504),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1530),
.B(n_1431),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1528),
.B(n_1505),
.Y(n_1546)
);

AND2x4_ASAP7_75t_L g1547 ( 
.A(n_1521),
.B(n_1493),
.Y(n_1547)
);

NOR2x1p5_ASAP7_75t_SL g1548 ( 
.A(n_1515),
.B(n_1489),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1517),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1514),
.B(n_1506),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1517),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1521),
.B(n_1504),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1530),
.B(n_1507),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1528),
.B(n_1505),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1530),
.B(n_1506),
.Y(n_1555)
);

OAI21xp33_ASAP7_75t_L g1556 ( 
.A1(n_1531),
.A2(n_1504),
.B(n_1491),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1537),
.Y(n_1558)
);

AOI21xp33_ASAP7_75t_SL g1559 ( 
.A1(n_1519),
.A2(n_1466),
.B(n_1541),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1531),
.B(n_1507),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1515),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1536),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1520),
.B(n_1512),
.Y(n_1563)
);

OR2x2_ASAP7_75t_L g1564 ( 
.A(n_1520),
.B(n_1512),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1537),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1524),
.Y(n_1566)
);

INVx1_ASAP7_75t_SL g1567 ( 
.A(n_1536),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1520),
.B(n_1522),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1524),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1522),
.B(n_1481),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1515),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1522),
.B(n_1478),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1528),
.B(n_1505),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1529),
.B(n_1478),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1540),
.B(n_1481),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1540),
.B(n_1509),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1518),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1524),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1534),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1521),
.B(n_1493),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1529),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1515),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_SL g1583 ( 
.A1(n_1521),
.A2(n_1510),
.B(n_1499),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1540),
.B(n_1465),
.Y(n_1584)
);

NAND4xp25_ASAP7_75t_L g1585 ( 
.A(n_1544),
.B(n_1499),
.C(n_1422),
.D(n_1421),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1550),
.B(n_1513),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1555),
.B(n_1513),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1543),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1546),
.B(n_1541),
.Y(n_1589)
);

INVx1_ASAP7_75t_SL g1590 ( 
.A(n_1562),
.Y(n_1590)
);

OAI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1544),
.A2(n_1485),
.B(n_1480),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1546),
.B(n_1541),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1553),
.B(n_1529),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1566),
.Y(n_1594)
);

AND2x4_ASAP7_75t_L g1595 ( 
.A(n_1547),
.B(n_1521),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1554),
.B(n_1541),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1576),
.B(n_1549),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1562),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1554),
.B(n_1535),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1553),
.B(n_1529),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1573),
.B(n_1535),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1569),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1560),
.B(n_1538),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1573),
.B(n_1535),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1578),
.Y(n_1605)
);

AND2x4_ASAP7_75t_L g1606 ( 
.A(n_1547),
.B(n_1521),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1579),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1547),
.B(n_1535),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1561),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1567),
.Y(n_1610)
);

OAI31xp33_ASAP7_75t_L g1611 ( 
.A1(n_1556),
.A2(n_1552),
.A3(n_1446),
.B(n_1525),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1551),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1581),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1560),
.B(n_1538),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1558),
.B(n_1513),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1565),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1580),
.B(n_1528),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1561),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1528),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1608),
.B(n_1545),
.Y(n_1620)
);

OAI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1591),
.A2(n_1583),
.B(n_1552),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1591),
.A2(n_1485),
.B1(n_1459),
.B2(n_1469),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1608),
.B(n_1580),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1585),
.A2(n_1559),
.B(n_1525),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1617),
.B(n_1619),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1590),
.B(n_1584),
.Y(n_1626)
);

NOR2xp33_ASAP7_75t_L g1627 ( 
.A(n_1597),
.B(n_1431),
.Y(n_1627)
);

INVxp67_ASAP7_75t_SL g1628 ( 
.A(n_1613),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1613),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1594),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1594),
.Y(n_1631)
);

OAI211xp5_ASAP7_75t_L g1632 ( 
.A1(n_1611),
.A2(n_1577),
.B(n_1518),
.C(n_1525),
.Y(n_1632)
);

NAND2x1p5_ASAP7_75t_L g1633 ( 
.A(n_1590),
.B(n_1498),
.Y(n_1633)
);

AOI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1585),
.A2(n_1528),
.B1(n_1518),
.B2(n_1525),
.Y(n_1634)
);

NAND2x1_ASAP7_75t_L g1635 ( 
.A(n_1595),
.B(n_1527),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1611),
.A2(n_1518),
.B1(n_1568),
.B2(n_1557),
.Y(n_1636)
);

OAI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1597),
.A2(n_1519),
.B(n_1527),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1602),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1602),
.Y(n_1639)
);

AOI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1586),
.A2(n_1528),
.B(n_1527),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1586),
.A2(n_1568),
.B1(n_1527),
.B2(n_1519),
.C(n_1575),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1587),
.B(n_1563),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1598),
.B(n_1527),
.Y(n_1643)
);

AOI32xp33_ASAP7_75t_L g1644 ( 
.A1(n_1610),
.A2(n_1533),
.A3(n_1526),
.B1(n_1523),
.B2(n_1527),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1621),
.A2(n_1610),
.B(n_1617),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1629),
.B(n_1598),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1635),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1628),
.Y(n_1648)
);

OAI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1634),
.A2(n_1519),
.B1(n_1587),
.B2(n_1615),
.Y(n_1649)
);

OAI21xp33_ASAP7_75t_L g1650 ( 
.A1(n_1636),
.A2(n_1598),
.B(n_1615),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1628),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1627),
.B(n_1588),
.Y(n_1652)
);

AOI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1636),
.A2(n_1588),
.B(n_1612),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_L g1654 ( 
.A(n_1632),
.B(n_1616),
.C(n_1612),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1627),
.B(n_1616),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1624),
.A2(n_1519),
.B1(n_1498),
.B2(n_1501),
.Y(n_1656)
);

INVxp67_ASAP7_75t_SL g1657 ( 
.A(n_1643),
.Y(n_1657)
);

OAI22xp33_ASAP7_75t_L g1658 ( 
.A1(n_1633),
.A2(n_1498),
.B1(n_1501),
.B2(n_1563),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1622),
.A2(n_1564),
.B1(n_1599),
.B2(n_1601),
.Y(n_1659)
);

NOR2xp33_ASAP7_75t_L g1660 ( 
.A(n_1626),
.B(n_1595),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_L g1661 ( 
.A1(n_1622),
.A2(n_1564),
.B1(n_1599),
.B2(n_1601),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1625),
.B(n_1589),
.Y(n_1662)
);

AOI222xp33_ASAP7_75t_L g1663 ( 
.A1(n_1641),
.A2(n_1548),
.B1(n_1619),
.B2(n_1606),
.C1(n_1595),
.C2(n_1589),
.Y(n_1663)
);

AOI22xp33_ASAP7_75t_L g1664 ( 
.A1(n_1653),
.A2(n_1623),
.B1(n_1631),
.B2(n_1630),
.Y(n_1664)
);

AOI21xp33_ASAP7_75t_L g1665 ( 
.A1(n_1650),
.A2(n_1643),
.B(n_1633),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1657),
.Y(n_1666)
);

NAND2xp33_ASAP7_75t_L g1667 ( 
.A(n_1652),
.B(n_1644),
.Y(n_1667)
);

AOI222xp33_ASAP7_75t_L g1668 ( 
.A1(n_1645),
.A2(n_1638),
.B1(n_1639),
.B2(n_1637),
.C1(n_1548),
.C2(n_1606),
.Y(n_1668)
);

OAI21xp33_ASAP7_75t_SL g1669 ( 
.A1(n_1663),
.A2(n_1620),
.B(n_1604),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1648),
.B(n_1643),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1657),
.Y(n_1671)
);

OAI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1654),
.A2(n_1660),
.B(n_1659),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1651),
.B(n_1646),
.Y(n_1673)
);

O2A1O1Ixp5_ASAP7_75t_L g1674 ( 
.A1(n_1658),
.A2(n_1595),
.B(n_1606),
.C(n_1640),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1661),
.A2(n_1606),
.B(n_1642),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1672),
.A2(n_1655),
.B(n_1647),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1664),
.B(n_1662),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1666),
.Y(n_1678)
);

O2A1O1Ixp33_ASAP7_75t_L g1679 ( 
.A1(n_1667),
.A2(n_1649),
.B(n_1656),
.C(n_1605),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1664),
.B(n_1607),
.C(n_1605),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1671),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1670),
.B(n_1592),
.Y(n_1682)
);

NOR3xp33_ASAP7_75t_L g1683 ( 
.A(n_1673),
.B(n_1675),
.C(n_1669),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1665),
.B(n_1592),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_SL g1685 ( 
.A1(n_1678),
.A2(n_1607),
.B(n_1674),
.C(n_1668),
.Y(n_1685)
);

AOI211xp5_ASAP7_75t_L g1686 ( 
.A1(n_1683),
.A2(n_1604),
.B(n_1596),
.C(n_1454),
.Y(n_1686)
);

OAI211xp5_ASAP7_75t_SL g1687 ( 
.A1(n_1677),
.A2(n_1593),
.B(n_1614),
.C(n_1600),
.Y(n_1687)
);

XOR2x2_ASAP7_75t_L g1688 ( 
.A(n_1676),
.B(n_1431),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1681),
.B(n_1596),
.Y(n_1689)
);

AOI221xp5_ASAP7_75t_SL g1690 ( 
.A1(n_1686),
.A2(n_1679),
.B1(n_1684),
.B2(n_1682),
.C(n_1680),
.Y(n_1690)
);

NAND4xp75_ASAP7_75t_L g1691 ( 
.A(n_1689),
.B(n_1618),
.C(n_1609),
.D(n_1533),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1687),
.A2(n_1618),
.B1(n_1609),
.B2(n_1523),
.Y(n_1692)
);

AOI31xp33_ASAP7_75t_L g1693 ( 
.A1(n_1685),
.A2(n_1466),
.A3(n_1603),
.B(n_1600),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_SL g1694 ( 
.A1(n_1688),
.A2(n_1502),
.B1(n_1614),
.B2(n_1603),
.Y(n_1694)
);

OAI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1686),
.A2(n_1593),
.B1(n_1609),
.B2(n_1447),
.C(n_1493),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1691),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1692),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1693),
.Y(n_1698)
);

NAND4xp75_ASAP7_75t_L g1699 ( 
.A(n_1690),
.B(n_1533),
.C(n_1526),
.D(n_1523),
.Y(n_1699)
);

NAND3xp33_ASAP7_75t_L g1700 ( 
.A(n_1694),
.B(n_1582),
.C(n_1571),
.Y(n_1700)
);

NOR4xp25_ASAP7_75t_L g1701 ( 
.A(n_1696),
.B(n_1695),
.C(n_1582),
.D(n_1571),
.Y(n_1701)
);

NOR3xp33_ASAP7_75t_L g1702 ( 
.A(n_1698),
.B(n_1429),
.C(n_1501),
.Y(n_1702)
);

AOI322xp5_ASAP7_75t_L g1703 ( 
.A1(n_1697),
.A2(n_1513),
.A3(n_1516),
.B1(n_1523),
.B2(n_1533),
.C1(n_1526),
.C2(n_1542),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1702),
.A2(n_1699),
.B1(n_1700),
.B2(n_1526),
.Y(n_1704)
);

AOI211xp5_ASAP7_75t_SL g1705 ( 
.A1(n_1704),
.A2(n_1701),
.B(n_1703),
.C(n_1465),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1705),
.Y(n_1706)
);

AOI22xp5_ASAP7_75t_L g1707 ( 
.A1(n_1706),
.A2(n_1574),
.B1(n_1542),
.B2(n_1516),
.Y(n_1707)
);

OAI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1707),
.A2(n_1570),
.B(n_1572),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1708),
.A2(n_1574),
.B1(n_1572),
.B2(n_1538),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1708),
.A2(n_1516),
.B(n_1532),
.Y(n_1710)
);

OR2x6_ASAP7_75t_L g1711 ( 
.A(n_1710),
.B(n_1415),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1709),
.A2(n_1516),
.B(n_1532),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_1711),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1712),
.Y(n_1714)
);

OAI221xp5_ASAP7_75t_R g1715 ( 
.A1(n_1713),
.A2(n_1482),
.B1(n_1539),
.B2(n_1538),
.C(n_1502),
.Y(n_1715)
);

AOI211xp5_ASAP7_75t_L g1716 ( 
.A1(n_1715),
.A2(n_1714),
.B(n_1414),
.C(n_1416),
.Y(n_1716)
);


endmodule