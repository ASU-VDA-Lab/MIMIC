module fake_jpeg_31956_n_502 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_502);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_502;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_8),
.B(n_13),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_52),
.B(n_26),
.C(n_48),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx3_ASAP7_75t_SL g54 ( 
.A(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_56),
.B(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_17),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_57),
.B(n_98),
.Y(n_155)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_64),
.Y(n_127)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_17),
.B(n_7),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_69),
.B(n_71),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_25),
.Y(n_70)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_21),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_72),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx2_ASAP7_75t_SL g141 ( 
.A(n_73),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_74),
.B(n_77),
.Y(n_148)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_76),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_27),
.B(n_9),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_9),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_9),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_81),
.B(n_88),
.Y(n_152)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_39),
.A2(n_9),
.B1(n_13),
.B2(n_12),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_99),
.B1(n_80),
.B2(n_43),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_31),
.Y(n_88)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx6_ASAP7_75t_SL g144 ( 
.A(n_93),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx4_ASAP7_75t_SL g95 ( 
.A(n_40),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_22),
.B(n_6),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_33),
.Y(n_108)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_34),
.B(n_6),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_95),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_106),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_107),
.A2(n_125),
.B1(n_137),
.B2(n_140),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_108),
.B(n_142),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_65),
.A2(n_22),
.B1(n_30),
.B2(n_33),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_54),
.A2(n_40),
.B1(n_49),
.B2(n_98),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_49),
.B1(n_45),
.B2(n_38),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_51),
.A2(n_49),
.B1(n_45),
.B2(n_38),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_138),
.B1(n_96),
.B2(n_73),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_52),
.A2(n_30),
.B1(n_43),
.B2(n_44),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_129),
.A2(n_16),
.B(n_13),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_53),
.A2(n_44),
.B1(n_48),
.B2(n_47),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_130),
.B(n_83),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_55),
.B(n_21),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_74),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_87),
.A2(n_49),
.B1(n_23),
.B2(n_46),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_63),
.A2(n_38),
.B1(n_45),
.B2(n_35),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_58),
.A2(n_23),
.B1(n_46),
.B2(n_47),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_64),
.B(n_37),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_72),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_71),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_157),
.A2(n_175),
.B1(n_191),
.B2(n_109),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_126),
.B(n_62),
.C(n_56),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_158),
.B(n_190),
.C(n_200),
.Y(n_218)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx4_ASAP7_75t_SL g251 ( 
.A(n_159),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_160),
.A2(n_205),
.B1(n_144),
.B2(n_123),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_100),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_161),
.B(n_162),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_141),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_163),
.B(n_167),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_126),
.A2(n_37),
.B(n_35),
.C(n_29),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_164),
.B(n_198),
.Y(n_244)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_103),
.Y(n_165)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_172),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_113),
.A2(n_29),
.B1(n_26),
.B2(n_93),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_129),
.B(n_21),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_180),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_113),
.A2(n_78),
.B1(n_82),
.B2(n_89),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_60),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_183),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_107),
.B(n_21),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

BUFx24_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_132),
.Y(n_182)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_152),
.B(n_96),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_155),
.B(n_59),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_192),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_61),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_187),
.Y(n_224)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_94),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_147),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_189),
.B(n_203),
.Y(n_252)
);

AND2x2_ASAP7_75t_SL g190 ( 
.A(n_134),
.B(n_66),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_102),
.A2(n_75),
.B1(n_67),
.B2(n_90),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_102),
.Y(n_192)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_194),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_117),
.B(n_92),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_128),
.Y(n_237)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_101),
.Y(n_196)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_196),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_101),
.Y(n_197)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_197),
.Y(n_236)
);

A2O1A1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_137),
.A2(n_86),
.B(n_73),
.C(n_31),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_110),
.Y(n_199)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_104),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_104),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_116),
.B(n_86),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_207),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_124),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_105),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_206),
.Y(n_233)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_105),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_162),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_219),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_168),
.A2(n_150),
.B1(n_149),
.B2(n_76),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_222),
.A2(n_226),
.B1(n_238),
.B2(n_248),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_168),
.A2(n_150),
.B1(n_149),
.B2(n_91),
.Y(n_226)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_144),
.C(n_145),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_118),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_156),
.A2(n_123),
.B(n_118),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_231),
.A2(n_195),
.B(n_198),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_161),
.B(n_114),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_247),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_240),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_171),
.A2(n_180),
.B1(n_167),
.B2(n_158),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_177),
.B1(n_163),
.B2(n_205),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_185),
.B(n_151),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_84),
.B1(n_151),
.B2(n_124),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_253),
.B1(n_205),
.B2(n_187),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_245),
.A2(n_179),
.B1(n_190),
.B2(n_199),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_166),
.B(n_114),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_157),
.A2(n_139),
.B1(n_143),
.B2(n_85),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_178),
.A2(n_143),
.B1(n_139),
.B2(n_109),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_255),
.A2(n_259),
.B(n_31),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_252),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_272),
.Y(n_307)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_260),
.A2(n_286),
.B1(n_255),
.B2(n_273),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_261),
.B(n_274),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_210),
.A2(n_183),
.B(n_164),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_262),
.A2(n_270),
.B(n_177),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_238),
.B(n_190),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_263),
.B(n_268),
.Y(n_315)
);

INVx13_ASAP7_75t_L g264 ( 
.A(n_212),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_264),
.Y(n_326)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_213),
.Y(n_266)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_266),
.Y(n_305)
);

AOI221xp5_ASAP7_75t_L g267 ( 
.A1(n_216),
.A2(n_220),
.B1(n_224),
.B2(n_229),
.C(n_240),
.Y(n_267)
);

XOR2x2_ASAP7_75t_SL g304 ( 
.A(n_267),
.B(n_279),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_217),
.B(n_203),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_210),
.A2(n_181),
.B(n_206),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_224),
.B(n_220),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_271),
.B(n_273),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_252),
.Y(n_272)
);

NAND2x1_ASAP7_75t_SL g274 ( 
.A(n_244),
.B(n_207),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_169),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_275),
.B(n_280),
.Y(n_313)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_276),
.Y(n_308)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_227),
.A2(n_170),
.B(n_186),
.C(n_188),
.D(n_165),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_252),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_230),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_287),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_242),
.A2(n_201),
.B(n_202),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_282),
.A2(n_45),
.B(n_38),
.Y(n_327)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_283),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_222),
.A2(n_182),
.B1(n_145),
.B2(n_196),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_284),
.A2(n_293),
.B1(n_294),
.B2(n_193),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_218),
.B(n_119),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_285),
.B(n_235),
.C(n_215),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_218),
.A2(n_226),
.B1(n_231),
.B2(n_237),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_225),
.B(n_189),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_242),
.B(n_159),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_290),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_242),
.A2(n_194),
.B(n_177),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_289),
.A2(n_0),
.B(n_1),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_249),
.B(n_31),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_249),
.Y(n_291)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_291),
.Y(n_333)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_212),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_295),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_146),
.B1(n_136),
.B2(n_135),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_146),
.B1(n_136),
.B2(n_119),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_281),
.A2(n_250),
.B1(n_236),
.B2(n_232),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_258),
.A2(n_233),
.B1(n_236),
.B2(n_251),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_297),
.A2(n_310),
.B1(n_318),
.B2(n_321),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_298),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_250),
.B1(n_235),
.B2(n_241),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_302),
.A2(n_322),
.B1(n_290),
.B2(n_274),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_332),
.C(n_289),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_262),
.A2(n_215),
.B(n_221),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_306),
.A2(n_316),
.B(n_323),
.Y(n_339)
);

OAI32xp33_ASAP7_75t_L g309 ( 
.A1(n_271),
.A2(n_246),
.A3(n_223),
.B1(n_214),
.B2(n_128),
.Y(n_309)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_309),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_258),
.A2(n_251),
.B1(n_208),
.B2(n_223),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_221),
.B(n_241),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_261),
.A2(n_208),
.B1(n_246),
.B2(n_228),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_221),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_324),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_260),
.A2(n_228),
.B1(n_79),
.B2(n_2),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_269),
.A2(n_45),
.B1(n_38),
.B2(n_31),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_327),
.A2(n_329),
.B(n_330),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_282),
.A2(n_5),
.B(n_11),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_268),
.B(n_6),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_292),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_275),
.C(n_269),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_312),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_334),
.B(n_335),
.C(n_337),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_312),
.B(n_279),
.Y(n_335)
);

OAI22x1_ASAP7_75t_L g338 ( 
.A1(n_323),
.A2(n_274),
.B1(n_270),
.B2(n_265),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_338),
.A2(n_340),
.B1(n_345),
.B2(n_363),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_265),
.B1(n_287),
.B2(n_294),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_308),
.Y(n_341)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_341),
.Y(n_368)
);

INVxp33_ASAP7_75t_SL g342 ( 
.A(n_326),
.Y(n_342)
);

CKINVDCx14_ASAP7_75t_R g371 ( 
.A(n_342),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_328),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_344),
.B(n_350),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_284),
.B1(n_293),
.B2(n_280),
.Y(n_345)
);

BUFx5_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_256),
.C(n_288),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_349),
.B(n_362),
.C(n_316),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_315),
.B(n_254),
.Y(n_350)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_300),
.Y(n_352)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_328),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_355),
.B(n_360),
.Y(n_384)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_356),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_309),
.Y(n_357)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_359),
.A2(n_364),
.B1(n_318),
.B2(n_310),
.Y(n_385)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_361),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_291),
.C(n_283),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_322),
.A2(n_278),
.B1(n_277),
.B2(n_276),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_301),
.A2(n_295),
.B1(n_266),
.B2(n_257),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_299),
.A2(n_264),
.B(n_10),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_365),
.A2(n_330),
.B(n_329),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_315),
.B(n_264),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_366),
.B(n_344),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_339),
.A2(n_299),
.B(n_298),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_367),
.A2(n_327),
.B(n_360),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_334),
.B(n_299),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_372),
.B(n_395),
.Y(n_418)
);

XNOR2x1_ASAP7_75t_L g373 ( 
.A(n_335),
.B(n_338),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_393),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_379),
.C(n_347),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_337),
.B(n_311),
.C(n_304),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_339),
.A2(n_353),
.B(n_347),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_380),
.A2(n_367),
.B(n_346),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_336),
.A2(n_304),
.B1(n_313),
.B2(n_306),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_381),
.A2(n_354),
.B1(n_357),
.B2(n_353),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_336),
.A2(n_331),
.B1(n_296),
.B2(n_313),
.Y(n_383)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_383),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_385),
.A2(n_389),
.B1(n_351),
.B2(n_354),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_351),
.A2(n_333),
.B1(n_325),
.B2(n_317),
.Y(n_386)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_386),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_346),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_357),
.A2(n_297),
.B1(n_321),
.B2(n_311),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_390),
.B(n_355),
.Y(n_405)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_348),
.Y(n_391)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_391),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_349),
.B(n_307),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_362),
.B(n_307),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_394),
.B(n_365),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_359),
.B(n_327),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_400),
.Y(n_435)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_397),
.Y(n_422)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_384),
.Y(n_398)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_398),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_401),
.A2(n_385),
.B1(n_389),
.B2(n_378),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_402),
.A2(n_395),
.B1(n_393),
.B2(n_371),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_403),
.Y(n_430)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_404),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_405),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_343),
.C(n_319),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_407),
.B(n_409),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_408),
.A2(n_412),
.B(n_414),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_343),
.C(n_319),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_387),
.B(n_381),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_417),
.Y(n_423)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_368),
.Y(n_415)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_415),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_378),
.A2(n_341),
.B1(n_361),
.B2(n_358),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_392),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_379),
.B(n_364),
.C(n_356),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g419 ( 
.A(n_377),
.B(n_333),
.C(n_325),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_394),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g420 ( 
.A(n_390),
.B(n_254),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_420),
.B(n_376),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_421),
.A2(n_402),
.B1(n_413),
.B2(n_398),
.Y(n_441)
);

AOI322xp5_ASAP7_75t_SL g424 ( 
.A1(n_414),
.A2(n_373),
.A3(n_382),
.B1(n_380),
.B2(n_388),
.C1(n_372),
.C2(n_324),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_440),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_418),
.Y(n_443)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_429),
.A2(n_417),
.B1(n_401),
.B2(n_409),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_405),
.B(n_374),
.Y(n_434)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_434),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_SL g436 ( 
.A(n_418),
.B(n_330),
.C(n_370),
.Y(n_436)
);

OAI21xp33_ASAP7_75t_SL g445 ( 
.A1(n_436),
.A2(n_412),
.B(n_406),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_411),
.A2(n_392),
.B1(n_375),
.B2(n_374),
.Y(n_437)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_437),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_397),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_441),
.A2(n_452),
.B1(n_428),
.B2(n_431),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_443),
.B(n_446),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_429),
.Y(n_459)
);

XOR2x2_ASAP7_75t_L g463 ( 
.A(n_445),
.B(n_427),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_436),
.A2(n_407),
.B1(n_399),
.B2(n_419),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_396),
.C(n_399),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_448),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_435),
.B(n_400),
.C(n_404),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_415),
.Y(n_449)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_449),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_421),
.A2(n_422),
.B1(n_431),
.B2(n_430),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_432),
.Y(n_455)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_455),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_430),
.B(n_375),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_456),
.B(n_406),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_459),
.B(n_460),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_11),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_453),
.A2(n_434),
.B(n_422),
.Y(n_462)
);

AND2x2_ASAP7_75t_SL g471 ( 
.A(n_462),
.B(n_463),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_454),
.A2(n_423),
.B1(n_439),
.B2(n_432),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_464),
.A2(n_469),
.B1(n_300),
.B2(n_10),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_439),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_466),
.B(n_305),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_435),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_468),
.B(n_448),
.C(n_447),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_451),
.A2(n_450),
.B1(n_352),
.B2(n_449),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_441),
.A2(n_427),
.B1(n_317),
.B2(n_425),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_470),
.B(n_446),
.C(n_305),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_457),
.A2(n_463),
.B(n_456),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_472),
.B(n_474),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_458),
.B(n_452),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_473),
.B(n_475),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_477),
.B(n_478),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_467),
.B(n_10),
.C(n_11),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_479),
.B(n_480),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_462),
.A2(n_16),
.B(n_1),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_482),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_467),
.A2(n_458),
.B(n_459),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_464),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_484),
.Y(n_494)
);

NOR3xp33_ASAP7_75t_SL g487 ( 
.A(n_471),
.B(n_468),
.C(n_465),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_487),
.B(n_473),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_474),
.B(n_476),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_490),
.B(n_16),
.Y(n_493)
);

AOI21x1_ASAP7_75t_L g498 ( 
.A1(n_491),
.A2(n_484),
.B(n_486),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_485),
.A2(n_480),
.B1(n_465),
.B2(n_16),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_492),
.A2(n_495),
.B1(n_483),
.B2(n_488),
.Y(n_497)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_493),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_489),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_497),
.A2(n_498),
.B(n_494),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_494),
.C(n_496),
.Y(n_500)
);

AOI221xp5_ASAP7_75t_L g501 ( 
.A1(n_500),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.C(n_494),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_501),
.A2(n_3),
.B(n_499),
.Y(n_502)
);


endmodule