module fake_jpeg_5906_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_36),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_17),
.B(n_1),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_21),
.B1(n_26),
.B2(n_19),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

OR2x4_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_1),
.Y(n_42)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_26),
.B1(n_21),
.B2(n_19),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_43),
.A2(n_27),
.B(n_29),
.C(n_28),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_51),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_46),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_16),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_29),
.Y(n_83)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_39),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_21),
.B1(n_20),
.B2(n_17),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_57),
.B1(n_52),
.B2(n_31),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_27),
.B1(n_20),
.B2(n_25),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_37),
.B1(n_41),
.B2(n_36),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_62),
.B1(n_74),
.B2(n_82),
.Y(n_94)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_41),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_75),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_39),
.B1(n_25),
.B2(n_33),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_18),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_66),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_68),
.Y(n_95)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_69),
.A2(n_53),
.B(n_48),
.C(n_29),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_73),
.Y(n_102)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_33),
.B(n_35),
.C(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_35),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_77),
.B1(n_28),
.B2(n_2),
.Y(n_99)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_78),
.B(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_35),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_30),
.B1(n_18),
.B2(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_98),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_78),
.A2(n_53),
.B1(n_36),
.B2(n_48),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_54),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_33),
.B1(n_55),
.B2(n_47),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_96),
.B1(n_104),
.B2(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_55),
.B1(n_47),
.B2(n_35),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_101),
.B(n_103),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_59),
.A2(n_55),
.B1(n_40),
.B2(n_22),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_40),
.B1(n_22),
.B2(n_54),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_72),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_70),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_100),
.A2(n_65),
.B1(n_68),
.B2(n_73),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_108),
.A2(n_117),
.B(n_127),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_75),
.C(n_61),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_122),
.C(n_4),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_74),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_111),
.A2(n_88),
.B(n_98),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_60),
.B(n_83),
.C(n_74),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_112),
.B(n_92),
.Y(n_140)
);

O2A1O1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_97),
.A2(n_58),
.B(n_83),
.C(n_60),
.Y(n_113)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_40),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_120),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_101),
.A2(n_40),
.B(n_54),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_22),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_22),
.C(n_28),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_88),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_120),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_1),
.B(n_2),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_85),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_88),
.A2(n_3),
.B(n_4),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_127),
.B(n_117),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_96),
.B(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_133),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_131),
.B(n_6),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_134),
.B(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

XNOR2x1_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_95),
.Y(n_138)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_114),
.C(n_119),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_109),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_142),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_113),
.B1(n_111),
.B2(n_124),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_92),
.B1(n_89),
.B2(n_91),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_141),
.A2(n_114),
.B1(n_110),
.B2(n_115),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_126),
.B(n_89),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_102),
.B(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_123),
.B(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_147),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_129),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_122),
.C(n_118),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_134),
.B(n_147),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_158),
.C(n_160),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_159),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_156),
.A2(n_130),
.B1(n_135),
.B2(n_146),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_136),
.A2(n_110),
.B1(n_86),
.B2(n_128),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_157),
.B(n_143),
.Y(n_169)
);

AOI322xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_86),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C1(n_8),
.C2(n_9),
.Y(n_158)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_4),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_5),
.C(n_6),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_148),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_165),
.B(n_176),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_166),
.A2(n_132),
.B1(n_133),
.B2(n_144),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_140),
.B1(n_130),
.B2(n_134),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_167),
.A2(n_173),
.B1(n_163),
.B2(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_164),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_175),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_130),
.B1(n_141),
.B2(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_149),
.Y(n_176)
);

AOI211xp5_ASAP7_75t_SL g189 ( 
.A1(n_177),
.A2(n_178),
.B(n_180),
.C(n_182),
.Y(n_189)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_174),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_185),
.Y(n_187)
);

AOI31xp67_ASAP7_75t_L g182 ( 
.A1(n_166),
.A2(n_159),
.A3(n_135),
.B(n_139),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_171),
.B(n_161),
.C(n_152),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_183),
.B(n_170),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_188),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_167),
.B(n_132),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_181),
.B(n_144),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_190),
.B(n_172),
.C(n_165),
.Y(n_197)
);

OAI21x1_ASAP7_75t_L g191 ( 
.A1(n_182),
.A2(n_168),
.B(n_146),
.Y(n_191)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_191),
.B(n_185),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_149),
.B1(n_151),
.B2(n_168),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_192),
.A2(n_160),
.B1(n_142),
.B2(n_172),
.Y(n_195)
);

AO21x1_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_186),
.B(n_15),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_195),
.B(n_197),
.C(n_187),
.Y(n_198)
);

NAND3xp33_ASAP7_75t_SL g196 ( 
.A(n_189),
.B(n_165),
.C(n_9),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_14),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_201),
.C(n_194),
.Y(n_202)
);

AOI31xp33_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_200),
.A3(n_196),
.B(n_11),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_7),
.C(n_10),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.C(n_10),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_12),
.Y(n_205)
);


endmodule