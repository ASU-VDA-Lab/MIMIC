module fake_jpeg_20583_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_50),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_22),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_28),
.Y(n_79)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_55),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_19),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_63),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_0),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_61),
.B(n_64),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_18),
.B(n_15),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_65),
.A2(n_32),
.B1(n_30),
.B2(n_38),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_18),
.B(n_15),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_66),
.B(n_67),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_28),
.B(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx3_ASAP7_75t_SL g71 ( 
.A(n_24),
.Y(n_71)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

BUFx16f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_72),
.B(n_75),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_73),
.Y(n_115)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_33),
.Y(n_74)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_26),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_32),
.B1(n_38),
.B2(n_30),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_76),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_79),
.B(n_84),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_67),
.B1(n_65),
.B2(n_71),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_83),
.A2(n_87),
.B1(n_96),
.B2(n_110),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_32),
.B1(n_38),
.B2(n_30),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_91),
.A2(n_74),
.B1(n_75),
.B2(n_68),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_39),
.B1(n_37),
.B2(n_17),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_41),
.A2(n_39),
.B1(n_37),
.B2(n_17),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_67),
.A2(n_36),
.B1(n_27),
.B2(n_29),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_43),
.A2(n_25),
.B1(n_29),
.B2(n_27),
.Y(n_97)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_54),
.B(n_25),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_31),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_71),
.A2(n_36),
.B1(n_27),
.B2(n_31),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_74),
.A2(n_36),
.B1(n_31),
.B2(n_14),
.Y(n_111)
);

AO22x1_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_23),
.B1(n_69),
.B2(n_62),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_117),
.A2(n_136),
.B1(n_137),
.B2(n_141),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_56),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_121),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_81),
.C(n_86),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_122),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_55),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_63),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_83),
.A2(n_50),
.B(n_46),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_140),
.B(n_143),
.Y(n_157)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_80),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_146),
.B1(n_78),
.B2(n_85),
.Y(n_161)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_127),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_90),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_129),
.Y(n_172)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_105),
.A2(n_40),
.B1(n_53),
.B2(n_31),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_131),
.A2(n_90),
.B(n_28),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_134),
.B(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_135),
.B(n_138),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_100),
.A2(n_60),
.B1(n_16),
.B2(n_20),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_100),
.A2(n_20),
.B1(n_16),
.B2(n_50),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_76),
.B(n_58),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_103),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_87),
.B(n_42),
.Y(n_140)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_101),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_109),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_88),
.B(n_45),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_28),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_77),
.A2(n_20),
.B1(n_16),
.B2(n_50),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_147),
.B(n_154),
.Y(n_171)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_148),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_110),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_149),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_72),
.C(n_70),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_151),
.C(n_99),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g151 ( 
.A(n_101),
.B(n_47),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_58),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_73),
.B1(n_57),
.B2(n_59),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_156),
.A2(n_85),
.B1(n_114),
.B2(n_113),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_89),
.B(n_94),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_179),
.B(n_180),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_169),
.B1(n_173),
.B2(n_182),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_77),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_168),
.B(n_90),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_138),
.A2(n_114),
.B1(n_116),
.B2(n_104),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_122),
.B(n_116),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_177),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_45),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_0),
.B(n_1),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_150),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_123),
.B1(n_128),
.B2(n_152),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_128),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_126),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_151),
.B1(n_117),
.B2(n_148),
.Y(n_210)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_131),
.B(n_99),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_186),
.A2(n_192),
.B(n_129),
.Y(n_221)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_189),
.Y(n_199)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_151),
.A2(n_51),
.B(n_28),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_139),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_195),
.B(n_196),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_159),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_147),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_124),
.Y(n_201)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_201),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_202),
.B(n_225),
.C(n_181),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_124),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_204),
.Y(n_233)
);

MAJx2_ASAP7_75t_L g205 ( 
.A(n_157),
.B(n_168),
.C(n_158),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_205),
.B(n_225),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_159),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_207),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_165),
.B(n_174),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_193),
.Y(n_209)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_210),
.B(n_221),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_160),
.B(n_155),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_213),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_171),
.B(n_142),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_185),
.Y(n_216)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_174),
.B(n_130),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_218),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_176),
.B(n_189),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_182),
.B(n_126),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_223),
.Y(n_249)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_220),
.Y(n_260)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_164),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_183),
.B(n_143),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_175),
.B(n_52),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_172),
.B(n_132),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_162),
.A2(n_141),
.B1(n_112),
.B2(n_104),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_228),
.A2(n_188),
.B1(n_178),
.B2(n_170),
.Y(n_245)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_209),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_230),
.B(n_250),
.C(n_199),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_219),
.A2(n_177),
.B1(n_208),
.B2(n_197),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_232),
.A2(n_248),
.B1(n_254),
.B2(n_261),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_161),
.B1(n_175),
.B2(n_186),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_238),
.A2(n_203),
.B1(n_166),
.B2(n_193),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_157),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_239),
.B(n_243),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_221),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_245),
.A2(n_229),
.B1(n_203),
.B2(n_220),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_214),
.A2(n_184),
.B1(n_179),
.B2(n_173),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_163),
.C(n_192),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_218),
.B(n_180),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_211),
.Y(n_275)
);

OA21x2_ASAP7_75t_SL g253 ( 
.A1(n_217),
.A2(n_163),
.B(n_180),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_213),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_208),
.A2(n_125),
.B1(n_172),
.B2(n_190),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_259),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_194),
.A2(n_190),
.B1(n_188),
.B2(n_170),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_194),
.A2(n_170),
.B1(n_166),
.B2(n_178),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_209),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_205),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_275),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_257),
.A2(n_202),
.B(n_226),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_264),
.A2(n_272),
.B(n_282),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_265),
.A2(n_283),
.B1(n_254),
.B2(n_256),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_268),
.Y(n_294)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_231),
.B(n_198),
.Y(n_269)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_269),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_271),
.B(n_257),
.CI(n_238),
.CON(n_302),
.SN(n_302)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_278),
.C(n_286),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_275),
.B(n_267),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_199),
.A3(n_205),
.B1(n_224),
.B2(n_222),
.C1(n_196),
.C2(n_206),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_246),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_230),
.B(n_216),
.C(n_215),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_240),
.Y(n_280)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_233),
.B(n_200),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_281),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_240),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_284),
.A2(n_287),
.B(n_288),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_187),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_285),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_251),
.B(n_132),
.C(n_119),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_236),
.B(n_33),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_119),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_293),
.A2(n_310),
.B1(n_280),
.B2(n_291),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_243),
.C(n_250),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_296),
.B(n_297),
.C(n_301),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_239),
.C(n_252),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_257),
.C(n_237),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_302),
.B(n_304),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_242),
.C(n_236),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_307),
.B(n_234),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_264),
.A2(n_249),
.B(n_246),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_269),
.B(n_289),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_266),
.A2(n_249),
.B1(n_242),
.B2(n_235),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_288),
.A2(n_232),
.B1(n_235),
.B2(n_241),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_277),
.B1(n_287),
.B2(n_270),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_241),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_315),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_72),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_317),
.A2(n_326),
.B(n_331),
.Y(n_348)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_306),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_327),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_306),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_325),
.B(n_328),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_SL g326 ( 
.A(n_302),
.B(n_272),
.C(n_282),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_283),
.B1(n_270),
.B2(n_273),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_303),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g329 ( 
.A(n_314),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_329),
.B(n_330),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_303),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_299),
.B(n_284),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_331),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_332),
.A2(n_333),
.B1(n_293),
.B2(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_334),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_336),
.B(n_307),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_309),
.Y(n_337)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_337),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_234),
.Y(n_338)
);

AOI32xp33_ASAP7_75t_L g341 ( 
.A1(n_338),
.A2(n_308),
.A3(n_302),
.B1(n_312),
.B2(n_315),
.Y(n_341)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_341),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_SL g342 ( 
.A(n_326),
.B(n_301),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_342),
.B(n_324),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_295),
.C(n_296),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_346),
.C(n_322),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_344),
.A2(n_327),
.B1(n_324),
.B2(n_329),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_345),
.B(n_320),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_295),
.C(n_297),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_349),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_330),
.A2(n_304),
.B(n_298),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_319),
.A2(n_305),
.B(n_13),
.C(n_2),
.Y(n_354)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_354),
.B(n_317),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_347),
.A2(n_332),
.B1(n_321),
.B2(n_340),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_356),
.A2(n_366),
.B1(n_344),
.B2(n_342),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_360),
.Y(n_372)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_359),
.Y(n_370)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_348),
.A2(n_318),
.B1(n_323),
.B2(n_334),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_349),
.B(n_354),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_362),
.B(n_363),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_353),
.B(n_322),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_364),
.B(n_367),
.C(n_369),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_347),
.A2(n_340),
.B1(n_352),
.B2(n_351),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_132),
.C(n_119),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_13),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_368),
.B(n_0),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_70),
.C(n_33),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_371),
.B(n_378),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_359),
.A2(n_350),
.B1(n_355),
.B2(n_339),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_375),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_366),
.B(n_350),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_380),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g379 ( 
.A(n_358),
.B(n_345),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_379),
.B(n_13),
.C(n_2),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_356),
.A2(n_365),
.B1(n_358),
.B2(n_361),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_367),
.A2(n_364),
.B(n_369),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_381),
.A2(n_370),
.B1(n_374),
.B2(n_377),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_382),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_384),
.B(n_385),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_1),
.C(n_2),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_1),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_387),
.B(n_388),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_380),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_381),
.B(n_2),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_389),
.B(n_4),
.Y(n_393)
);

OAI221xp5_ASAP7_75t_L g391 ( 
.A1(n_379),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_382),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_392),
.B(n_9),
.C(n_10),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_393),
.B(n_395),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_383),
.A2(n_5),
.B(n_8),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_396),
.A2(n_397),
.B(n_9),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_386),
.A2(n_5),
.B(n_9),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_384),
.A2(n_390),
.B1(n_385),
.B2(n_11),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_11),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_399),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_400),
.B(n_401),
.Y(n_407)
);

AO21x1_ASAP7_75t_L g406 ( 
.A1(n_403),
.A2(n_404),
.B(n_11),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_L g405 ( 
.A1(n_402),
.A2(n_394),
.B(n_393),
.Y(n_405)
);

INVxp33_ASAP7_75t_L g408 ( 
.A(n_405),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_407),
.B(n_406),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_12),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_12),
.Y(n_411)
);


endmodule