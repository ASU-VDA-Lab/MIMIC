module fake_jpeg_2311_n_210 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_210);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_210;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx2_ASAP7_75t_L g51 ( 
.A(n_5),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_42),
.Y(n_60)
);

INVx8_ASAP7_75t_SL g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_8),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_28),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_31),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_61),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_73),
.B(n_77),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_67),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_67),
.B1(n_58),
.B2(n_52),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_83),
.A2(n_71),
.B1(n_56),
.B2(n_66),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_53),
.B(n_54),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_87),
.A2(n_94),
.B(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_53),
.B1(n_62),
.B2(n_69),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_59),
.B1(n_65),
.B2(n_60),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_62),
.B1(n_69),
.B2(n_59),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_71),
.B1(n_66),
.B2(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_73),
.A2(n_76),
.B(n_54),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_72),
.B(n_49),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_57),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_98),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_68),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_84),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_68),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_102),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_64),
.B1(n_55),
.B2(n_70),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_63),
.Y(n_105)
);

OAI32xp33_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_109),
.A3(n_72),
.B1(n_89),
.B2(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_106),
.Y(n_132)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_108),
.A2(n_97),
.B1(n_109),
.B2(n_110),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_63),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_65),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_111),
.Y(n_114)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_89),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_88),
.Y(n_116)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_90),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_46),
.C(n_45),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_5),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_124),
.Y(n_148)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_95),
.A2(n_111),
.B1(n_106),
.B2(n_100),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_41),
.B1(n_40),
.B2(n_39),
.Y(n_139)
);

HAxp5_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_88),
.CON(n_123),
.SN(n_123)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_123),
.A2(n_116),
.B(n_126),
.Y(n_134)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_133),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_35),
.B(n_33),
.Y(n_142)
);

AOI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_107),
.A2(n_112),
.B(n_48),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_0),
.Y(n_137)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_134),
.A2(n_141),
.B(n_142),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_125),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_138),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_140),
.C(n_146),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_151),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_0),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_139),
.A2(n_147),
.B1(n_154),
.B2(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_38),
.C(n_37),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_122),
.A2(n_1),
.B(n_2),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_114),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_19),
.Y(n_172)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_32),
.C(n_29),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_24),
.B1(n_6),
.B2(n_7),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_149),
.A2(n_16),
.B(n_17),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_6),
.C(n_7),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_15),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_124),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_148),
.A2(n_128),
.B1(n_120),
.B2(n_133),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_157),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_123),
.B1(n_127),
.B2(n_131),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_158),
.A2(n_161),
.B(n_163),
.Y(n_177)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_171),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_149),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.C(n_172),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_16),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_174),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_169),
.B(n_173),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_143),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_145),
.B(n_147),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_144),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_150),
.B(n_20),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_136),
.B(n_21),
.Y(n_174)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_162),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_179),
.B(n_160),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_140),
.C(n_164),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_180),
.B(n_186),
.C(n_156),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_181),
.A2(n_161),
.B1(n_168),
.B2(n_142),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_182),
.B(n_184),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_156),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_187),
.B(n_191),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_188),
.B(n_186),
.Y(n_199)
);

CKINVDCx11_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_190),
.B(n_192),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_180),
.B(n_160),
.C(n_146),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_176),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_193),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_195),
.B(n_175),
.Y(n_198)
);

AOI21x1_ASAP7_75t_L g201 ( 
.A1(n_198),
.A2(n_192),
.B(n_177),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_194),
.C(n_185),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_201),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_200),
.B(n_189),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_202),
.B(n_203),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_197),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_206),
.A2(n_196),
.B1(n_199),
.B2(n_204),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_163),
.A3(n_137),
.B1(n_170),
.B2(n_22),
.C1(n_21),
.C2(n_23),
.Y(n_208)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_208),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_209),
.B(n_22),
.Y(n_210)
);


endmodule