module real_jpeg_18706_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_513),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_0),
.B(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_1),
.B(n_76),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_1),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_1),
.B(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g323 ( 
.A(n_1),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g416 ( 
.A(n_1),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_1),
.B(n_273),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_2),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_2),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_3),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_3),
.B(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_3),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_3),
.B(n_115),
.Y(n_114)
);

NAND2xp67_ASAP7_75t_L g197 ( 
.A(n_3),
.B(n_101),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_3),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_3),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_3),
.B(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_4),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g243 ( 
.A(n_4),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g425 ( 
.A(n_4),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_4),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_5),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_6),
.B(n_201),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_6),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g346 ( 
.A(n_6),
.B(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_6),
.B(n_39),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_6),
.B(n_408),
.Y(n_407)
);

AND2x2_ASAP7_75t_SL g424 ( 
.A(n_6),
.B(n_425),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_6),
.B(n_448),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_7),
.B(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_7),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_7),
.B(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_7),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_7),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_7),
.B(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_7),
.Y(n_454)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_8),
.Y(n_143)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_8),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_8),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_9),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_9),
.Y(n_126)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_9),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_9),
.Y(n_451)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_10),
.B(n_34),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_10),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_10),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_10),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_10),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_10),
.B(n_183),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_10),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_11),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_11),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_11),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_11),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_11),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_11),
.B(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_12),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_12),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_12),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_12),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_12),
.B(n_140),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_12),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_12),
.B(n_145),
.Y(n_144)
);

NAND2x1_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_159),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_13),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_13),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_14),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_14),
.B(n_223),
.Y(n_222)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_14),
.B(n_265),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_14),
.B(n_60),
.Y(n_322)
);

AND2x2_ASAP7_75t_SL g384 ( 
.A(n_14),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_14),
.B(n_412),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g418 ( 
.A(n_14),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_14),
.B(n_459),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_16),
.Y(n_185)
);

BUFx4f_ASAP7_75t_L g240 ( 
.A(n_16),
.Y(n_240)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_17),
.Y(n_147)
);

BUFx8_ASAP7_75t_L g166 ( 
.A(n_17),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_17),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_170),
.Y(n_19)
);

NAND2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_169),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_148),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_23),
.B(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_79),
.C(n_106),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_24),
.B(n_79),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_54),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_25),
.B(n_55),
.C(n_69),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_41),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_26),
.B(n_47),
.C(n_53),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_33),
.C(n_37),
.Y(n_26)
);

INVxp33_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_28),
.B(n_37),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_30),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_31),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_32),
.B(n_261),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_33),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_33),
.Y(n_133)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_35),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_36),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_37),
.B(n_197),
.C(n_198),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_37),
.A2(n_38),
.B1(n_198),
.B2(n_227),
.Y(n_226)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_40),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_41)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_48),
.B(n_137),
.C(n_144),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_48),
.B(n_144),
.Y(n_194)
);

MAJx2_ASAP7_75t_L g195 ( 
.A(n_48),
.B(n_196),
.C(n_199),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_48),
.A2(n_49),
.B1(n_199),
.B2(n_200),
.Y(n_230)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_52),
.Y(n_160)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_52),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_69),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_56),
.B(n_59),
.C(n_64),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_59),
.A2(n_68),
.B1(n_156),
.B2(n_157),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_59),
.B(n_100),
.C(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_59),
.A2(n_68),
.B1(n_221),
.B2(n_222),
.Y(n_332)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_62),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_64),
.B1(n_70),
.B2(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_63),
.B(n_118),
.Y(n_342)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.C(n_73),
.Y(n_69)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_64),
.B(n_119),
.C(n_280),
.Y(n_279)
);

OR2x2_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_70),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_84),
.C(n_89),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_70),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_111)
);

MAJx2_ASAP7_75t_L g321 ( 
.A(n_70),
.B(n_322),
.C(n_323),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_70),
.A2(n_82),
.B1(n_322),
.B2(n_377),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_72),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_77),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.C(n_96),
.Y(n_79)
);

XNOR2x2_ASAP7_75t_L g202 ( 
.A(n_80),
.B(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_83),
.B(n_96),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_139),
.C(n_142),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_84),
.A2(n_85),
.B1(n_142),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_85),
.B(n_234),
.Y(n_475)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_87),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_88),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_111),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.C(n_102),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_97),
.A2(n_98),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_98),
.B(n_129),
.Y(n_128)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_99),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_102),
.B1(n_103),
.B2(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_100),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_100),
.A2(n_130),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_101),
.Y(n_385)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_105),
.Y(n_457)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_107),
.B(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_131),
.C(n_136),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_109),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.C(n_127),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_110),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_112),
.B(n_128),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.C(n_123),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_113),
.A2(n_114),
.B1(n_123),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_122),
.Y(n_461)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_131),
.A2(n_132),
.B1(n_136),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_136),
.Y(n_207)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_139),
.B(n_191),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_182),
.B(n_186),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_182),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_142),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_142),
.A2(n_182),
.B1(n_192),
.B2(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_142),
.B(n_467),
.Y(n_466)
);

BUFx12f_ASAP7_75t_L g440 ( 
.A(n_143),
.Y(n_440)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_161),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_157),
.A2(n_158),
.B1(n_242),
.B2(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_158),
.Y(n_244)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_160),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_168),
.Y(n_161)
);

CKINVDCx12_ASAP7_75t_R g168 ( 
.A(n_162),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_163),
.Y(n_167)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_208),
.B(n_509),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_171),
.A2(n_511),
.B(n_512),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_172),
.B(n_174),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_202),
.C(n_204),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_175),
.B(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_193),
.C(n_195),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_212),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.C(n_190),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_177),
.B(n_180),
.Y(n_300)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_182),
.B(n_314),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_182),
.A2(n_219),
.B1(n_314),
.B2(n_315),
.Y(n_378)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_186),
.B(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_189),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_189),
.A2(n_345),
.B1(n_494),
.B2(n_495),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_190),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_192),
.B(n_467),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_195),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_196),
.B(n_230),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_SL g225 ( 
.A(n_197),
.B(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_198),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_202),
.A2(n_204),
.B1(n_205),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_248),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_245),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_210),
.B(n_245),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.C(n_215),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_211),
.B(n_213),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_215),
.B(n_394),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_228),
.C(n_231),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_216),
.B(n_298),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.C(n_225),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_217),
.B(n_220),
.Y(n_334)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2x2_ASAP7_75t_L g333 ( 
.A(n_225),
.B(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_298)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_242),
.C(n_244),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_233),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_241),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_237),
.Y(n_257)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_240),
.Y(n_410)
);

XNOR2x2_ASAP7_75t_SL g256 ( 
.A(n_241),
.B(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_243),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_396),
.Y(n_248)
);

A2O1A1O1Ixp25_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_335),
.B(n_388),
.C(n_389),
.D(n_395),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_251),
.B(n_390),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_303),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_252),
.B(n_303),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_296),
.Y(n_252)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_253),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_277),
.C(n_292),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_255),
.B(n_306),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_258),
.C(n_267),
.Y(n_255)
);

XNOR2x1_ASAP7_75t_SL g357 ( 
.A(n_256),
.B(n_358),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_258),
.A2(n_259),
.B1(n_267),
.B2(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_259),
.A2(n_260),
.B(n_264),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

INVx4_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_262),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_263),
.Y(n_413)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_267),
.Y(n_359)
);

MAJx3_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.C(n_275),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_268),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_271),
.B(n_477),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_272),
.B(n_275),
.Y(n_311)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_278),
.A2(n_292),
.B1(n_293),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_278),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_283),
.C(n_286),
.Y(n_278)
);

XNOR2x2_ASAP7_75t_SL g328 ( 
.A(n_279),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_280),
.B(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_286),
.Y(n_329)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_299),
.B1(n_301),
.B2(n_302),
.Y(n_296)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_297),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_299),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_299),
.B(n_301),
.C(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_333),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_304),
.A2(n_305),
.B1(n_333),
.B2(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_305),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_308),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_328),
.C(n_330),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_339),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.C(n_321),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_310),
.B(n_372),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_312),
.A2(n_313),
.B1(n_321),
.B2(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_317),
.Y(n_316)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g377 ( 
.A(n_322),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_323),
.B(n_376),
.Y(n_375)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_327),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_330),
.Y(n_339)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_333),
.Y(n_362)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_363),
.B(n_387),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_360),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_360),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_340),
.C(n_357),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_357),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.C(n_344),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_343),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_369),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.C(n_350),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_346),
.A2(n_350),
.B1(n_351),
.B2(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_346),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_366),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.C(n_374),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_367),
.A2(n_368),
.B1(n_504),
.B2(n_505),
.Y(n_503)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g505 ( 
.A1(n_370),
.A2(n_371),
.B1(n_374),
.B2(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_374),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_378),
.C(n_379),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_375),
.B(n_499),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_378),
.B(n_379),
.Y(n_499)
);

MAJx2_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_384),
.C(n_386),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_380),
.A2(n_381),
.B1(n_386),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_384),
.B(n_487),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_386),
.Y(n_488)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_387),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_393),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_393),
.Y(n_395)
);

NAND4xp25_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_398),
.C(n_399),
.D(n_400),
.Y(n_396)
);

OAI21x1_ASAP7_75t_SL g400 ( 
.A1(n_401),
.A2(n_502),
.B(n_508),
.Y(n_400)
);

AOI21x1_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_490),
.B(n_501),
.Y(n_401)
);

OAI21x1_ASAP7_75t_SL g402 ( 
.A1(n_403),
.A2(n_469),
.B(n_489),
.Y(n_402)
);

AOI21x1_ASAP7_75t_SL g403 ( 
.A1(n_404),
.A2(n_443),
.B(n_468),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_405),
.A2(n_430),
.B(n_442),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_414),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_406),
.B(n_414),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_411),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_407),
.B(n_411),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_407),
.B(n_439),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_422),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_415),
.B(n_424),
.C(n_426),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_418),
.Y(n_464)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_424),
.B1(n_426),
.B2(n_427),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_431),
.A2(n_438),
.B(n_441),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_437),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_432),
.B(n_437),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp67_ASAP7_75t_L g468 ( 
.A(n_444),
.B(n_445),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_462),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_464),
.C(n_465),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_452),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_447),
.B(n_458),
.C(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_458),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_453),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_463),
.A2(n_464),
.B1(n_465),
.B2(n_466),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_471),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_483),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_472),
.B(n_484),
.C(n_486),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_474),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_473),
.B(n_476),
.C(n_481),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_475),
.A2(n_476),
.B1(n_481),
.B2(n_482),
.Y(n_474)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_475),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_476),
.Y(n_482)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx8_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_486),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_500),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_SL g501 ( 
.A(n_491),
.B(n_500),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_498),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_497),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_493),
.B(n_497),
.C(n_498),
.Y(n_507)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_507),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_507),
.Y(n_508)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);


endmodule