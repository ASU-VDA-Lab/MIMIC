module real_jpeg_24794_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_1),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_38),
.B1(n_56),
.B2(n_57),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_1),
.A2(n_38),
.B1(n_72),
.B2(n_73),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_1),
.A2(n_28),
.B1(n_30),
.B2(n_38),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_26),
.B(n_197),
.C(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_1),
.B(n_27),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_30),
.B(n_54),
.C(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_1),
.B(n_71),
.C(n_72),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_1),
.B(n_52),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_1),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_1),
.B(n_69),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_3),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_6),
.A2(n_33),
.B1(n_56),
.B2(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_6),
.A2(n_33),
.B1(n_72),
.B2(n_73),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_7),
.A2(n_24),
.B1(n_39),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_127),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_127),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_7),
.A2(n_72),
.B1(n_73),
.B2(n_127),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_10),
.A2(n_28),
.B1(n_30),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_10),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_10),
.A2(n_32),
.B1(n_51),
.B2(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_10),
.A2(n_51),
.B1(n_72),
.B2(n_73),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_13),
.Y(n_96)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_13),
.Y(n_97)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_13),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_13),
.B(n_250),
.Y(n_255)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_13),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_323),
.Y(n_16)
);

OAI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_40),
.B1(n_44),
.B2(n_320),
.C(n_322),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_18),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_18),
.B(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_18),
.B(n_40),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_35),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_19),
.A2(n_27),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_20),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_21),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_24),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g197 ( 
.A1(n_25),
.A2(n_30),
.B(n_38),
.Y(n_197)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_37),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_27),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_27),
.B(n_126),
.Y(n_167)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_28),
.A2(n_30),
.B1(n_54),
.B2(n_59),
.Y(n_62)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVxp33_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_36),
.B(n_125),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_38),
.A2(n_56),
.B(n_59),
.Y(n_221)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_39),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_40),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_40),
.A2(n_94),
.B1(n_103),
.B2(n_108),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_41),
.A2(n_82),
.B(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_309),
.B(n_319),
.Y(n_44)
);

OAI211xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_128),
.B(n_145),
.C(n_308),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_104),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_47),
.B(n_104),
.Y(n_146)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_47),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_79),
.CI(n_93),
.CON(n_47),
.SN(n_47)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_48),
.A2(n_49),
.B(n_64),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_48),
.B(n_79),
.C(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_64),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_52),
.B(n_60),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_52),
.B(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_53),
.B(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_53),
.B(n_138),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_53),
.A2(n_61),
.B(n_138),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_53)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_57),
.B1(n_70),
.B2(n_71),
.Y(n_77)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_57),
.B(n_238),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_60),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_60),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_61),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_74),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_65),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_68),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_66),
.A2(n_68),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_67),
.B(n_76),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_75),
.B(n_101),
.Y(n_118)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_78),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_69),
.B(n_225),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_72),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_72),
.B(n_261),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_75),
.B(n_235),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_76),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_91),
.B2(n_92),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_80),
.A2(n_91),
.B1(n_133),
.B2(n_143),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_80),
.B(n_85),
.C(n_88),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_80),
.B(n_133),
.C(n_144),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_82),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_81),
.B(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_82),
.B(n_125),
.Y(n_192)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_88),
.B2(n_89),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_87),
.B(n_190),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_88),
.A2(n_89),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_88),
.B(n_179),
.C(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_88),
.A2(n_89),
.B1(n_181),
.B2(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_89),
.B(n_136),
.C(n_139),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_90),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_99),
.B(n_103),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_94),
.A2(n_100),
.B1(n_108),
.B2(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_94),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_94),
.A2(n_108),
.B1(n_220),
.B2(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B(n_98),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_95),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_95),
.B(n_98),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_95),
.B(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_100),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_102),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_102),
.B(n_224),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_109),
.C(n_110),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_105),
.A2(n_106),
.B1(n_109),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_109),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_110),
.B(n_169),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_119),
.C(n_123),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_118),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_112),
.B(n_118),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_113),
.B(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_116),
.A2(n_159),
.B(n_162),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_116),
.B(n_255),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_119),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_121),
.B(n_183),
.Y(n_276)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_SL g145 ( 
.A(n_129),
.B(n_146),
.C(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_130),
.B(n_131),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_144),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_133),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_137),
.B(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_140),
.Y(n_315)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_171),
.B(n_307),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_168),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_149),
.B(n_168),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_150),
.B(n_153),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_155),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_165),
.C(n_166),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_156),
.A2(n_157),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_163),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_158),
.B(n_163),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_161),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_161),
.B(n_248),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_164),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_165),
.A2(n_166),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_165),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_165),
.A2(n_296),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_165),
.B(n_311),
.C(n_316),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_166),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_302),
.B(n_306),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_213),
.B(n_288),
.C(n_301),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_201),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_174),
.B(n_201),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_187),
.B2(n_200),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_185),
.B2(n_186),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_177),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_177),
.B(n_186),
.C(n_200),
.Y(n_289)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_180),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_184),
.Y(n_191)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_189),
.B(n_194),
.C(n_195),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_199),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.C(n_208),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_202),
.A2(n_203),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_208),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.C(n_211),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_218),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_211),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_212),
.B(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_287),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_229),
.B(n_286),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_226),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_216),
.B(n_226),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.C(n_222),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_217),
.B(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_219),
.B(n_222),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_220),
.Y(n_279)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_228),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_281),
.B(n_285),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_272),
.B(n_280),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_252),
.B(n_271),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_239),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_233),
.B(n_239),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_251),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_242),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_245),
.C(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_246),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVxp33_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_258),
.B(n_270),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_256),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_254),
.B(n_256),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_266),
.B(n_269),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_267),
.B(n_268),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_274),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_289),
.B(n_290),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_298),
.B2(n_299),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_292),
.B(n_299),
.C(n_300),
.Y(n_303)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_303),
.B(n_304),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_318),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_318),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_317),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_313),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_314),
.Y(n_316)
);


endmodule