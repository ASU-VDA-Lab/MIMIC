module fake_jpeg_14161_n_167 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_167);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_167;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_18),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_20),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_16),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_45),
.Y(n_54)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

NOR2x1_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_26),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_60),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_32),
.B1(n_17),
.B2(n_42),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_45),
.B(n_37),
.C(n_36),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_30),
.A2(n_39),
.B1(n_41),
.B2(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_53),
.A2(n_56),
.B1(n_35),
.B2(n_1),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_17),
.B1(n_25),
.B2(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_32),
.B(n_28),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_28),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_14),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_68),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_18),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_72),
.Y(n_91)
);

OA22x2_ASAP7_75t_SL g71 ( 
.A1(n_64),
.A2(n_34),
.B1(n_45),
.B2(n_40),
.Y(n_71)
);

OAI32xp33_ASAP7_75t_L g98 ( 
.A1(n_71),
.A2(n_58),
.A3(n_49),
.B1(n_63),
.B2(n_3),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_15),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_76),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_74),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_75),
.A2(n_78),
.B1(n_85),
.B2(n_86),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_16),
.C(n_26),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_35),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_20),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_14),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_49),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_35),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_87),
.A2(n_52),
.B(n_51),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_63),
.B1(n_51),
.B2(n_58),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_99),
.B1(n_88),
.B2(n_79),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_98),
.B(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_99)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_93),
.B(n_67),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_106),
.B(n_114),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_112),
.B1(n_94),
.B2(n_103),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_66),
.C(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_116),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_96),
.B(n_103),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_110),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_78),
.B(n_71),
.Y(n_111)
);

OAI31xp33_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_98),
.A3(n_75),
.B(n_101),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_66),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_78),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_83),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_74),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_113),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_115),
.B(n_2),
.Y(n_140)
);

AOI322xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_99),
.A3(n_95),
.B1(n_77),
.B2(n_80),
.C1(n_75),
.C2(n_9),
.Y(n_125)
);

OAI321xp33_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_6),
.A3(n_11),
.B1(n_5),
.B2(n_9),
.C(n_100),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_109),
.B1(n_111),
.B2(n_107),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_127),
.A2(n_131),
.B1(n_108),
.B2(n_115),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_109),
.A2(n_95),
.B1(n_75),
.B2(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

NAND4xp25_ASAP7_75t_L g142 ( 
.A(n_137),
.B(n_140),
.C(n_141),
.D(n_124),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_128),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_139),
.Y(n_145)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_147),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_126),
.B(n_127),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_131),
.B(n_138),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_129),
.C(n_126),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_151),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_152),
.A2(n_155),
.B1(n_144),
.B2(n_146),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_153),
.B(n_154),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_121),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_123),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_147),
.C(n_146),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_140),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_159),
.A2(n_157),
.B1(n_156),
.B2(n_142),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_159),
.A2(n_154),
.B(n_6),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_161),
.A2(n_158),
.B(n_0),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_164),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_3),
.Y(n_167)
);


endmodule