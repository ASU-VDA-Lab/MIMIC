module fake_jpeg_15292_n_43 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx8_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

BUFx12_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_R g12 ( 
.A(n_6),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_22),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_13),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_21),
.B1(n_8),
.B2(n_20),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_19),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g18 ( 
.A1(n_13),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_18),
.A2(n_8),
.B1(n_17),
.B2(n_13),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_14),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

AO22x1_ASAP7_75t_L g21 ( 
.A1(n_12),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_28),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_11),
.C(n_14),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_34),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_33),
.B1(n_31),
.B2(n_25),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_32),
.A2(n_24),
.B(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_8),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_37),
.B(n_40),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_36),
.Y(n_43)
);


endmodule