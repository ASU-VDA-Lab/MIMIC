module real_jpeg_3655_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_1),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_70),
.B1(n_72),
.B2(n_133),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_47),
.B1(n_49),
.B2(n_133),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_1),
.A2(n_34),
.B1(n_42),
.B2(n_133),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_4),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_47),
.B1(n_49),
.B2(n_74),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_4),
.A2(n_34),
.B1(n_42),
.B2(n_74),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_47),
.B1(n_49),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_5),
.A2(n_56),
.B1(n_70),
.B2(n_72),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_5),
.A2(n_34),
.B1(n_42),
.B2(n_56),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_5),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_6),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_6),
.A2(n_70),
.B1(n_72),
.B2(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_6),
.A2(n_47),
.B1(n_49),
.B2(n_187),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_6),
.A2(n_34),
.B1(n_42),
.B2(n_187),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_7),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_7),
.A2(n_47),
.B1(n_49),
.B2(n_76),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_7),
.A2(n_34),
.B1(n_42),
.B2(n_76),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_8),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_8),
.A2(n_46),
.B1(n_70),
.B2(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_8),
.A2(n_46),
.B1(n_63),
.B2(n_64),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_8),
.A2(n_34),
.B1(n_42),
.B2(n_46),
.Y(n_162)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_9),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_10),
.B(n_63),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_168),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_10),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_10),
.A2(n_63),
.B(n_177),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_10),
.B(n_85),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_10),
.A2(n_72),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_10),
.B(n_34),
.C(n_52),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_10),
.A2(n_47),
.B1(n_49),
.B2(n_213),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_10),
.B(n_37),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_10),
.B(n_57),
.Y(n_269)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_14),
.A2(n_63),
.B1(n_64),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_14),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_14),
.A2(n_70),
.B1(n_72),
.B2(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_14),
.A2(n_47),
.B1(n_49),
.B2(n_167),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_14),
.A2(n_34),
.B1(n_42),
.B2(n_167),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_15),
.A2(n_21),
.B(n_334),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_15),
.B(n_335),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_16),
.A2(n_70),
.B1(n_72),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_16),
.A2(n_63),
.B1(n_64),
.B2(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_16),
.A2(n_47),
.B1(n_49),
.B2(n_82),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_16),
.A2(n_34),
.B1(n_42),
.B2(n_82),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_17),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_17),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_17),
.A2(n_41),
.B1(n_70),
.B2(n_72),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_17),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_323)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_329),
.B(n_332),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_321),
.B(n_325),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_308),
.B(n_320),
.Y(n_23)
);

AO21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_147),
.B(n_305),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_134),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_107),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_27),
.B(n_107),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_77),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_28),
.B(n_93),
.C(n_105),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_58),
.B(n_59),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_29),
.A2(n_30),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_43),
.Y(n_30)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_31),
.A2(n_58),
.B1(n_59),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_31),
.A2(n_43),
.B1(n_44),
.B2(n_58),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B(n_39),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_32),
.A2(n_36),
.B1(n_121),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_32),
.A2(n_36),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_32),
.A2(n_36),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_33),
.A2(n_37),
.B1(n_40),
.B2(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_33),
.A2(n_37),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_33),
.A2(n_37),
.B1(n_180),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_33),
.A2(n_37),
.B1(n_217),
.B2(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_33),
.A2(n_37),
.B1(n_213),
.B2(n_267),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_33),
.A2(n_37),
.B1(n_267),
.B2(n_271),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_34),
.B(n_265),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_50),
.B1(n_55),
.B2(n_57),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_45),
.A2(n_50),
.B1(n_57),
.B2(n_124),
.Y(n_123)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_49),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

AO22x2_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_49),
.B1(n_86),
.B2(n_88),
.Y(n_85)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_47),
.A2(n_72),
.A3(n_86),
.B1(n_212),
.B2(n_214),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_47),
.B(n_255),
.Y(n_254)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_49),
.B(n_88),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_50),
.A2(n_55),
.B1(n_57),
.B2(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_50),
.A2(n_57),
.B(n_92),
.Y(n_99)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_50),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_50),
.A2(n_57),
.B1(n_207),
.B2(n_209),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_50),
.A2(n_57),
.B1(n_209),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_50),
.A2(n_57),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_50),
.A2(n_57),
.B1(n_237),
.B2(n_258),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_54),
.A2(n_125),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_54),
.A2(n_160),
.B1(n_208),
.B2(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_69),
.B1(n_73),
.B2(n_75),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_60),
.A2(n_69),
.B1(n_75),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_60),
.A2(n_69),
.B1(n_73),
.B2(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_60),
.A2(n_69),
.B1(n_96),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_60),
.A2(n_69),
.B1(n_186),
.B2(n_188),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_60),
.A2(n_69),
.B1(n_186),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_132),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_61),
.A2(n_168),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_61),
.A2(n_168),
.B1(n_316),
.B2(n_323),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_61),
.A2(n_168),
.B(n_323),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AOI32xp33_ASAP7_75t_L g176 ( 
.A1(n_64),
.A2(n_67),
.A3(n_72),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_66),
.B(n_70),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_72),
.B1(n_86),
.B2(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_70),
.B(n_213),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_93),
.B1(n_105),
.B2(n_106),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_78),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_79),
.B(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_91),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_85),
.B2(n_90),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_84),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_83),
.A2(n_85),
.B1(n_90),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_83),
.A2(n_85),
.B1(n_128),
.B2(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_83),
.A2(n_85),
.B(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_84),
.A2(n_103),
.B1(n_129),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_84),
.A2(n_129),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_84),
.A2(n_129),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_84),
.A2(n_129),
.B1(n_183),
.B2(n_199),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_84),
.A2(n_129),
.B1(n_198),
.B2(n_246),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_85),
.Y(n_129)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_94),
.A2(n_95),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_99),
.C(n_101),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_95),
.B(n_138),
.C(n_145),
.Y(n_309)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_104),
.Y(n_98)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_99),
.A2(n_104),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_99),
.B(n_141),
.C(n_143),
.Y(n_319)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.C(n_115),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_108),
.A2(n_109),
.B1(n_113),
.B2(n_114),
.Y(n_150)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_126),
.C(n_130),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_117),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_123),
.Y(n_189)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_126),
.B(n_130),
.Y(n_153)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_134),
.A2(n_306),
.B(n_307),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_146),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_135),
.B(n_146),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_145),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_142),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_144),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_169),
.B(n_304),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_149),
.B(n_151),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.C(n_156),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_155),
.Y(n_191)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_153),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.C(n_165),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_158),
.B(n_161),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_162),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_192),
.B(n_303),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_190),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_171),
.B(n_190),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.C(n_189),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_172),
.B(n_189),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_174),
.B(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_182),
.C(n_185),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_175),
.B(n_293),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_176),
.B(n_179),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_182),
.B(n_185),
.Y(n_293)
);

AOI31xp33_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_287),
.A3(n_296),
.B(n_300),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_232),
.B(n_286),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_219),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_195),
.B(n_219),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_206),
.C(n_210),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_196),
.B(n_283),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_201),
.C(n_205),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_205),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_203),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_204),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_206),
.B(n_210),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_223),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_221),
.B(n_222),
.C(n_223),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_224),
.B(n_227),
.C(n_231),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_227),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_228),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_281),
.B(n_285),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_250),
.B(n_280),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_242),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_235),
.B(n_242),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_239),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_241),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_243),
.B(n_245),
.C(n_248),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_248),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_261),
.B(n_279),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_259),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_273),
.B(n_278),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_268),
.B(n_272),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_277),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_277),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_291),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_299),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_298),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_310),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_319),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_314),
.B1(n_317),
.B2(n_318),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_312),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_314),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_317),
.C(n_319),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_322),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_330),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_324),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_331),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule