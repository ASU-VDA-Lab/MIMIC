module fake_jpeg_27541_n_317 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_37),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_8),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_27),
.B(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_26),
.C(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_48),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_23),
.B1(n_27),
.B2(n_31),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_53),
.B1(n_33),
.B2(n_19),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_26),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_55),
.Y(n_72)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_51),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_42),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_23),
.B1(n_19),
.B2(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_32),
.B1(n_33),
.B2(n_19),
.Y(n_82)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_67),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_40),
.C(n_35),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_63),
.B(n_93),
.C(n_40),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_53),
.A2(n_28),
.B1(n_17),
.B2(n_25),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_52),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_70),
.B(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_39),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_98),
.Y(n_112)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_24),
.B1(n_25),
.B2(n_17),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_75),
.A2(n_83),
.B1(n_85),
.B2(n_90),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_32),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g126 ( 
.A(n_76),
.B(n_86),
.CI(n_88),
.CON(n_126),
.SN(n_126)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_24),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_52),
.B(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_20),
.B1(n_21),
.B2(n_36),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_57),
.A2(n_17),
.B1(n_24),
.B2(n_34),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_84),
.A2(n_87),
.B1(n_96),
.B2(n_36),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_32),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_21),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g89 ( 
.A(n_59),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_57),
.A2(n_34),
.B1(n_29),
.B2(n_28),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_91),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_59),
.A2(n_29),
.B(n_20),
.C(n_21),
.Y(n_92)
);

MAJx3_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_18),
.C(n_22),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_40),
.C(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_94),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_111),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_109),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_110),
.A2(n_120),
.B1(n_88),
.B2(n_86),
.Y(n_134)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_36),
.B1(n_42),
.B2(n_40),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_114),
.A2(n_123),
.B1(n_127),
.B2(n_68),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_77),
.A2(n_36),
.B1(n_11),
.B2(n_7),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_128),
.Y(n_138)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_118),
.B(n_73),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_96),
.A2(n_30),
.B1(n_18),
.B2(n_22),
.Y(n_120)
);

OR2x4_ASAP7_75t_L g152 ( 
.A(n_121),
.B(n_18),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_82),
.B1(n_71),
.B2(n_62),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_30),
.B1(n_18),
.B2(n_22),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_72),
.C(n_93),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_78),
.C(n_87),
.Y(n_137)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_85),
.B1(n_65),
.B2(n_64),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_123),
.B1(n_119),
.B2(n_105),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_134),
.B(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_138),
.C(n_156),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_157),
.Y(n_161)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_153),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_92),
.B(n_65),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g188 ( 
.A1(n_144),
.A2(n_150),
.B(n_0),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_SL g145 ( 
.A(n_121),
.B(n_80),
.Y(n_145)
);

NAND2xp33_ASAP7_75t_R g189 ( 
.A(n_145),
.B(n_7),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_107),
.A2(n_84),
.B(n_70),
.Y(n_146)
);

NAND2xp33_ASAP7_75t_SL g180 ( 
.A(n_146),
.B(n_152),
.Y(n_180)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_148),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_68),
.B(n_67),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_103),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_154),
.B(n_155),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_111),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_117),
.B(n_73),
.C(n_30),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_101),
.B(n_73),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_66),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_154),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_177),
.B1(n_149),
.B2(n_129),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_167),
.B(n_169),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_168),
.B(n_170),
.Y(n_197)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_152),
.B(n_110),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_173),
.B(n_175),
.Y(n_201)
);

AND2x6_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_126),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_104),
.B1(n_119),
.B2(n_126),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_129),
.B1(n_142),
.B2(n_10),
.Y(n_204)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_150),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_135),
.B(n_106),
.Y(n_183)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_9),
.C(n_15),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

AO22x1_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_66),
.B1(n_118),
.B2(n_18),
.Y(n_186)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_0),
.B(n_2),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_189),
.B(n_12),
.Y(n_198)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_212),
.B1(n_219),
.B2(n_171),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_138),
.C(n_137),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_196),
.B(n_203),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_198),
.A2(n_177),
.B1(n_174),
.B2(n_169),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_187),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_210),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_202),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_147),
.C(n_140),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_220),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_185),
.A2(n_188),
.B(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_206),
.A2(n_208),
.B(n_218),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_209),
.Y(n_230)
);

AO21x1_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_140),
.B(n_132),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_140),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_164),
.A2(n_132),
.B1(n_9),
.B2(n_10),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_159),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_217),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_176),
.A2(n_132),
.B(n_1),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_188),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_162),
.B1(n_161),
.B2(n_173),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_237),
.B1(n_241),
.B2(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_201),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_231),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_167),
.B(n_166),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_242),
.B(n_186),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_235),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_239),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_207),
.B(n_190),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_172),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_SL g242 ( 
.A1(n_220),
.A2(n_186),
.B(n_190),
.C(n_160),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_196),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_251),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_195),
.B1(n_197),
.B2(n_213),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_240),
.B1(n_242),
.B2(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_237),
.B1(n_192),
.B2(n_197),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_247),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_200),
.C(n_205),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_255),
.C(n_261),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_194),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_199),
.B1(n_219),
.B2(n_172),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_253),
.B1(n_256),
.B2(n_242),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_198),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_257),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_225),
.C(n_228),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_231),
.A2(n_202),
.B1(n_216),
.B2(n_191),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_175),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_163),
.C(n_217),
.Y(n_261)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_240),
.B(n_227),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_272),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_253),
.B1(n_258),
.B2(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_244),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_270),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_269),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_233),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_259),
.B(n_163),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_249),
.B(n_209),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_273),
.B(n_277),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_245),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_242),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_264),
.B(n_243),
.C(n_255),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_278),
.B(n_284),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_267),
.B1(n_259),
.B2(n_266),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_281),
.A2(n_282),
.B1(n_2),
.B2(n_3),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_251),
.C(n_254),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_277),
.B(n_271),
.C(n_268),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_287),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_222),
.C(n_242),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g290 ( 
.A(n_274),
.B(n_202),
.CI(n_12),
.CON(n_290),
.SN(n_290)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_290),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_274),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_295),
.Y(n_301)
);

OAI21x1_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_275),
.B(n_269),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_290),
.B(n_15),
.Y(n_296)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_296),
.A2(n_300),
.A3(n_280),
.B1(n_288),
.B2(n_14),
.C1(n_287),
.C2(n_6),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_14),
.B(n_13),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_281),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_14),
.B1(n_12),
.B2(n_4),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_302),
.A2(n_305),
.B1(n_298),
.B2(n_299),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_278),
.C(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_303),
.B(n_307),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_306),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_283),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_284),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_292),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_309),
.B(n_291),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_301),
.B(n_303),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_313),
.B(n_308),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_314),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_311),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_3),
.Y(n_317)
);


endmodule