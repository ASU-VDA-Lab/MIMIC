module real_jpeg_3279_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_332, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_332;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_1),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_31),
.B1(n_33),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_68),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_2),
.A2(n_50),
.B1(n_51),
.B2(n_68),
.Y(n_124)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_3),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_90),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_3),
.B(n_33),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_3),
.A2(n_25),
.B(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_3),
.B(n_42),
.C(n_44),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_3),
.A2(n_50),
.B1(n_51),
.B2(n_145),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_3),
.B(n_61),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_3),
.B(n_115),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_3),
.B(n_40),
.Y(n_247)
);

AOI21xp33_ASAP7_75t_L g262 ( 
.A1(n_3),
.A2(n_33),
.B(n_196),
.Y(n_262)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_4),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_5),
.A2(n_31),
.B1(n_33),
.B2(n_55),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_55),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_55),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_8),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_8),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_8),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_173)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_11),
.A2(n_31),
.B1(n_33),
.B2(n_107),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_50),
.B1(n_51),
.B2(n_107),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_107),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_12),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_105),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_105),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_105),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_152),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_14),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_152),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_14),
.A2(n_50),
.B1(n_51),
.B2(n_152),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_14),
.A2(n_43),
.B1(n_44),
.B2(n_152),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_15),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_15),
.A2(n_37),
.B1(n_43),
.B2(n_44),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_15),
.A2(n_37),
.B1(n_50),
.B2(n_51),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_92),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_19),
.B(n_83),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_77),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_20),
.A2(n_21),
.B1(n_73),
.B2(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_38),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_22),
.B(n_39),
.C(n_57),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_22)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_23),
.A2(n_36),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_23),
.A2(n_30),
.B1(n_104),
.B2(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_23),
.A2(n_30),
.B1(n_104),
.B2(n_151),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_23),
.A2(n_106),
.B(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_23),
.A2(n_30),
.B1(n_151),
.B2(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_23),
.A2(n_89),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_30),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_26),
.B(n_145),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_26),
.B(n_29),
.C(n_33),
.Y(n_146)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_28),
.Y(n_29)
);

OA22x2_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_29),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_28),
.A2(n_31),
.B(n_144),
.C(n_146),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_30),
.A2(n_34),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_31),
.A2(n_33),
.B1(n_63),
.B2(n_64),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g197 ( 
.A(n_31),
.B(n_50),
.C(n_63),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_56),
.B1(n_57),
.B2(n_72),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_39),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_73),
.C(n_78),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_39),
.A2(n_72),
.B1(n_78),
.B2(n_79),
.Y(n_321)
);

OAI21x1_ASAP7_75t_R g39 ( 
.A1(n_40),
.A2(n_48),
.B(n_53),
.Y(n_39)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_40),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_40),
.B(n_124),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_40),
.A2(n_48),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_40),
.A2(n_48),
.B1(n_229),
.B2(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_41),
.B(n_54),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_41)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_47),
.B1(n_50),
.B2(n_51),
.Y(n_49)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_44),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_44),
.B(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_48),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_48),
.A2(n_190),
.B(n_192),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_51),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx6p67_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g194 ( 
.A1(n_51),
.A2(n_64),
.B(n_195),
.C(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_51),
.B(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_54),
.A2(n_134),
.B(n_162),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_66),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_58),
.A2(n_70),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_62),
.B(n_70),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_60),
.A2(n_70),
.B(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_67),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_61),
.A2(n_69),
.B1(n_149),
.B2(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_61),
.A2(n_69),
.B1(n_81),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_62),
.A2(n_66),
.B(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_62),
.A2(n_70),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_62),
.A2(n_70),
.B1(n_182),
.B2(n_262),
.Y(n_261)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_80),
.B(n_82),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_73),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_73),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_77),
.B(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_90),
.B(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_314),
.B(n_327),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_292),
.B(n_313),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_176),
.B(n_291),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_153),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_99),
.B(n_153),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_125),
.C(n_136),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_100),
.B(n_125),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_109),
.B2(n_110),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_108),
.C(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_111),
.B(n_120),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_116),
.B(n_118),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_112),
.A2(n_114),
.B(n_129),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_112),
.A2(n_118),
.B(n_129),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_112),
.A2(n_114),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_113),
.B(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_115),
.B1(n_117),
.B2(n_141),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_113),
.A2(n_128),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_113),
.A2(n_115),
.B1(n_145),
.B2(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_113),
.A2(n_115),
.B1(n_243),
.B2(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_114),
.A2(n_131),
.B(n_142),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_115),
.B(n_119),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_121),
.A2(n_122),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_121),
.A2(n_134),
.B1(n_191),
.B2(n_264),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g308 ( 
.A(n_123),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_133),
.Y(n_166)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_134),
.A2(n_135),
.B(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_136),
.B(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_147),
.C(n_150),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_137),
.A2(n_138),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_139),
.A2(n_140),
.B1(n_143),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_143),
.Y(n_217)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_147),
.B(n_150),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_175),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_164),
.B2(n_165),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_157),
.B(n_165),
.C(n_175),
.Y(n_312)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_161),
.B2(n_163),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_159),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_159),
.B(n_161),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_159),
.A2(n_163),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

AOI21xp33_ASAP7_75t_L g318 ( 
.A1(n_159),
.A2(n_300),
.B(n_302),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_174),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_169),
.B(n_172),
.C(n_174),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_171),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_173),
.Y(n_310)
);

AOI321xp33_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_272),
.A3(n_283),
.B1(n_289),
.B2(n_290),
.C(n_332),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_218),
.B(n_271),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_199),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_179),
.B(n_199),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.C(n_193),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_180),
.B(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_185),
.C(n_188),
.Y(n_214)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_189),
.B(n_193),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_192),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_194),
.B(n_198),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_211),
.B2(n_212),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_200),
.B(n_213),
.C(n_216),
.Y(n_284)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_202),
.B(n_206),
.C(n_210),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_266),
.B(n_270),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_256),
.B(n_265),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_237),
.B(n_255),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_230),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_230),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_224),
.B1(n_226),
.B2(n_227),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_231),
.B(n_234),
.C(n_236),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_232),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_235),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_249),
.B(n_254),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_244),
.B(n_248),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_247),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_250),
.B(n_253),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_261),
.C(n_263),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_269),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_273),
.B(n_275),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_275),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_280),
.C(n_282),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_277),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_285),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_293),
.B(n_312),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_312),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_298),
.C(n_306),
.Y(n_316)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_305),
.B2(n_306),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_309),
.B(n_311),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_309),
.Y(n_311)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_318),
.CI(n_319),
.CON(n_317),
.SN(n_317)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_318),
.C(n_319),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_323),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_316),
.B(n_317),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g330 ( 
.A(n_317),
.Y(n_330)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI21xp33_ASAP7_75t_L g327 ( 
.A1(n_323),
.A2(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);


endmodule