module fake_jpeg_10764_n_63 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_15),
.B(n_7),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g26 ( 
.A(n_0),
.B(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_30),
.B(n_33),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_34),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_1),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_24),
.A2(n_2),
.B(n_3),
.C(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_42),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_31),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_25),
.B1(n_29),
.B2(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_40),
.B(n_31),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_48),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_39),
.B1(n_43),
.B2(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_3),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_29),
.B(n_25),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_4),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_43),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_53),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_54),
.B(n_49),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_57),
.C(n_56),
.Y(n_60)
);

AOI322xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_55),
.A3(n_46),
.B1(n_51),
.B2(n_6),
.C1(n_7),
.C2(n_13),
.Y(n_61)
);

AOI322xp5_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_17),
.C1(n_18),
.C2(n_19),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_51),
.B1(n_20),
.B2(n_21),
.Y(n_63)
);


endmodule