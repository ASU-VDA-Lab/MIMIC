module real_jpeg_19247_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_321, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;
input n_321;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_1),
.A2(n_22),
.B(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_1),
.B(n_22),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_34),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_54),
.Y(n_144)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_1),
.A2(n_10),
.B(n_48),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_1),
.B(n_62),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_1),
.A2(n_26),
.B(n_64),
.C(n_193),
.Y(n_192)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_3),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_58),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_58),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_58),
.Y(n_272)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_4),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_4),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_4),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_4),
.B(n_143),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_5),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_105),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_6),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_105),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_105),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_22),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_8),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_9),
.A2(n_22),
.B1(n_23),
.B2(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_9),
.A2(n_29),
.B1(n_48),
.B2(n_49),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_29),
.B1(n_42),
.B2(n_43),
.Y(n_99)
);

O2A1O1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_10),
.A2(n_42),
.B(n_46),
.C(n_47),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_10),
.B(n_42),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_11),
.Y(n_45)
);

MAJx2_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_16),
.C(n_277),
.Y(n_12)
);

OAI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_82),
.B(n_317),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_35),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_16),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_30),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_17),
.A2(n_25),
.B(n_57),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_18),
.B(n_103),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_19),
.B(n_32),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_19),
.A2(n_25),
.B(n_32),
.Y(n_278)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B(n_24),
.C(n_25),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_21),
.B(n_26),
.Y(n_128)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_24),
.Y(n_130)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_25),
.B(n_104),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_26),
.A2(n_63),
.B(n_64),
.C(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_64),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_27),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_30),
.B(n_115),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_34),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_36),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_74),
.C(n_76),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_37),
.A2(n_38),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_55),
.C(n_59),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_39),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_39),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_39),
.A2(n_107),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_39),
.A2(n_59),
.B1(n_60),
.B2(n_107),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_51),
.B(n_52),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_40),
.A2(n_98),
.B(n_235),
.Y(n_260)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_41),
.B(n_53),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_41),
.B(n_162),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_41),
.B(n_99),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_43),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

OAI21xp33_ASAP7_75t_L g193 ( 
.A1(n_42),
.A2(n_54),
.B(n_66),
.Y(n_193)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_43),
.A2(n_50),
.B(n_54),
.C(n_158),
.Y(n_157)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_47),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_47),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_47),
.B(n_53),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_49),
.B(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_51),
.B(n_54),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_51),
.A2(n_198),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_54),
.B(n_93),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_55),
.A2(n_56),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_57),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_68),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_61),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_70),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_63),
.B(n_73),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_63),
.A2(n_68),
.B(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_67),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_67),
.B(n_69),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_69),
.A2(n_138),
.B(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_70),
.B(n_120),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_74),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_74),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_74),
.A2(n_76),
.B1(n_241),
.B2(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_76),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_77),
.B(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_80),
.B(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_310),
.B(n_316),
.Y(n_82)
);

OAI321xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_286),
.A3(n_305),
.B1(n_308),
.B2(n_309),
.C(n_321),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_264),
.B(n_285),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_245),
.B(n_263),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_145),
.B(n_227),
.C(n_244),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_131),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_88),
.B(n_131),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_112),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_101),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_90),
.B(n_101),
.C(n_112),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_91),
.B(n_97),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B(n_95),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_92),
.A2(n_93),
.B(n_144),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_93),
.A2(n_94),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_98),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_107),
.C(n_108),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_104),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_106),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_107),
.B(n_290),
.C(n_295),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_110),
.B(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_113),
.Y(n_242)
);

FAx1_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_117),
.CI(n_121),
.CON(n_113),
.SN(n_113)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_122),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_124),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_124),
.B(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_125),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_154),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.C(n_135),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_132),
.B(n_223),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_224),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_134),
.Y(n_224)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.C(n_140),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_137),
.B(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_138),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_139),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_153),
.Y(n_169)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_226),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_220),
.B(n_225),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_205),
.B(n_219),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_186),
.B(n_204),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_174),
.B(n_185),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_163),
.B(n_173),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_155),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_157),
.B(n_159),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_168),
.B(n_172),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_165),
.B(n_166),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_176),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_183),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_181),
.C(n_183),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_182),
.B(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_188),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_195),
.B1(n_196),
.B2(n_203),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_189),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_194),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_190),
.A2(n_191),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_190),
.A2(n_191),
.B1(n_277),
.B2(n_278),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_190),
.A2(n_278),
.B(n_280),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_192),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_191),
.B(n_260),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_199),
.B1(n_200),
.B2(n_202),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_197),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_198),
.B(n_215),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_199),
.B(n_202),
.C(n_203),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_206),
.B(n_207),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_214),
.C(n_218),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_214),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_214),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_216),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_228),
.B(n_229),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_242),
.B2(n_243),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_236),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_236),
.C(n_243),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_234),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_242),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_246),
.B(n_247),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_262),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_258),
.B2(n_259),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_259),
.C(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_251),
.B(n_253),
.C(n_257),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_257),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_255),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_260),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_266),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_283),
.B2(n_284),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_274),
.B1(n_281),
.B2(n_282),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_269),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_282),
.C(n_284),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B(n_273),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_271),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_272),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_288),
.C(n_297),
.Y(n_287)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_273),
.B(n_288),
.CI(n_297),
.CON(n_307),
.SN(n_307)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_279),
.B2(n_280),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_275),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_276),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_298),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_298),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_289),
.A2(n_290),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_300),
.C(n_304),
.Y(n_311)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_304),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_312),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_313),
.Y(n_315)
);


endmodule