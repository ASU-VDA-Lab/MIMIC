module fake_netlist_1_8806_n_725 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_725);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_725;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_622;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_31), .Y(n_80) );
BUFx3_ASAP7_75t_L g81 ( .A(n_30), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_50), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_4), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_74), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVx2_ASAP7_75t_L g86 ( .A(n_39), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_27), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_1), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_72), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_11), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_79), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_53), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_26), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_70), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_25), .Y(n_96) );
NOR2xp33_ASAP7_75t_L g97 ( .A(n_49), .B(n_76), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_33), .Y(n_98) );
OR2x2_ASAP7_75t_L g99 ( .A(n_64), .B(n_36), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_22), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_0), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_54), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_55), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_32), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_47), .Y(n_105) );
CKINVDCx16_ASAP7_75t_R g106 ( .A(n_67), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_61), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_5), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_65), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_13), .Y(n_110) );
INVxp67_ASAP7_75t_SL g111 ( .A(n_21), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_51), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_57), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_41), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_6), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_10), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_17), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_8), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_7), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_40), .Y(n_122) );
INVxp67_ASAP7_75t_SL g123 ( .A(n_52), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_62), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_66), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_13), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_59), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_78), .Y(n_128) );
INVx1_ASAP7_75t_SL g129 ( .A(n_91), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_80), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_119), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_81), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g136 ( .A(n_82), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_84), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_91), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_90), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_88), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_88), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_106), .B(n_0), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_93), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_109), .B(n_1), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_108), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_92), .Y(n_149) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
HB1xp67_ASAP7_75t_L g151 ( .A(n_108), .Y(n_151) );
AND2x4_ASAP7_75t_L g152 ( .A(n_83), .B(n_2), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_83), .B(n_2), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_94), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_95), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_100), .B(n_3), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
INVxp67_ASAP7_75t_L g158 ( .A(n_85), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_96), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_96), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_98), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_98), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_107), .Y(n_163) );
INVxp67_ASAP7_75t_L g164 ( .A(n_85), .Y(n_164) );
AND2x4_ASAP7_75t_L g165 ( .A(n_87), .B(n_89), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_107), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_127), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_120), .Y(n_168) );
AND2x2_ASAP7_75t_L g169 ( .A(n_87), .B(n_3), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_89), .B(n_4), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_127), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_121), .B(n_5), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_102), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_93), .Y(n_174) );
BUFx10_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_168), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_168), .B(n_120), .Y(n_177) );
BUFx4f_ASAP7_75t_L g178 ( .A(n_152), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_148), .B(n_104), .Y(n_179) );
NOR2xp33_ASAP7_75t_SL g180 ( .A(n_148), .B(n_99), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
AND2x4_ASAP7_75t_L g182 ( .A(n_165), .B(n_121), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_151), .B(n_114), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_152), .Y(n_185) );
OR2x2_ASAP7_75t_SL g186 ( .A(n_151), .B(n_126), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_174), .B(n_128), .Y(n_187) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_173), .B(n_125), .Y(n_188) );
NAND2xp33_ASAP7_75t_L g189 ( .A(n_142), .B(n_99), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_132), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_132), .Y(n_191) );
INVx4_ASAP7_75t_L g192 ( .A(n_152), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_158), .B(n_124), .Y(n_193) );
BUFx10_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_158), .B(n_101), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_134), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_164), .B(n_113), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_132), .Y(n_198) );
AND2x6_ASAP7_75t_L g199 ( .A(n_152), .B(n_112), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_132), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_172), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_134), .Y(n_202) );
AND2x4_ASAP7_75t_L g203 ( .A(n_165), .B(n_110), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_129), .A2(n_140), .B1(n_144), .B2(n_172), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_172), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_132), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_141), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_172), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_165), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_165), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_164), .B(n_115), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_153), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_173), .B(n_122), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g214 ( .A(n_153), .B(n_103), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_129), .B(n_117), .Y(n_215) );
AND2x4_ASAP7_75t_L g216 ( .A(n_171), .B(n_116), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_142), .Y(n_217) );
AOI22x1_ASAP7_75t_L g218 ( .A1(n_138), .A2(n_105), .B1(n_111), .B2(n_123), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_153), .A2(n_118), .B1(n_97), .B2(n_9), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_130), .B(n_35), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_144), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_169), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_134), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_130), .B(n_6), .Y(n_224) );
AND2x4_ASAP7_75t_L g225 ( .A(n_137), .B(n_7), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_155), .Y(n_226) );
BUFx8_ASAP7_75t_SL g227 ( .A(n_131), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_169), .Y(n_228) );
INVx3_ASAP7_75t_L g229 ( .A(n_142), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_169), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_144), .B(n_10), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_155), .Y(n_232) );
BUFx10_ASAP7_75t_L g233 ( .A(n_147), .Y(n_233) );
AO22x2_ASAP7_75t_L g234 ( .A1(n_137), .A2(n_11), .B1(n_12), .B2(n_14), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_132), .Y(n_235) );
BUFx12f_ASAP7_75t_L g236 ( .A(n_194), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_180), .A2(n_156), .B1(n_171), .B2(n_167), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_195), .B(n_154), .Y(n_238) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_178), .A2(n_155), .B(n_157), .C(n_166), .Y(n_239) );
INVxp33_ASAP7_75t_L g240 ( .A(n_176), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_178), .A2(n_154), .B(n_167), .Y(n_241) );
BUFx12f_ASAP7_75t_L g242 ( .A(n_194), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_176), .Y(n_243) );
BUFx6f_ASAP7_75t_L g244 ( .A(n_225), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_178), .B(n_170), .Y(n_245) );
NOR3xp33_ASAP7_75t_SL g246 ( .A(n_207), .B(n_170), .C(n_166), .Y(n_246) );
OR2x6_ASAP7_75t_L g247 ( .A(n_214), .B(n_163), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_203), .B(n_163), .Y(n_248) );
AND2x4_ASAP7_75t_L g249 ( .A(n_212), .B(n_149), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_189), .A2(n_149), .B(n_161), .Y(n_250) );
INVx3_ASAP7_75t_L g251 ( .A(n_209), .Y(n_251) );
BUFx4f_ASAP7_75t_L g252 ( .A(n_214), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_209), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_221), .B(n_145), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_209), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g256 ( .A1(n_204), .A2(n_145), .B1(n_161), .B2(n_157), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_210), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_214), .B(n_157), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g259 ( .A1(n_222), .A2(n_143), .B(n_160), .C(n_159), .Y(n_259) );
INVx4_ASAP7_75t_L g260 ( .A(n_192), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_202), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_195), .B(n_157), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_225), .A2(n_143), .B1(n_160), .B2(n_159), .Y(n_263) );
NAND2x1p5_ASAP7_75t_L g264 ( .A(n_225), .B(n_155), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_202), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_192), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_182), .B(n_160), .Y(n_267) );
AO22x1_ASAP7_75t_L g268 ( .A1(n_207), .A2(n_159), .B1(n_143), .B2(n_138), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_182), .B(n_139), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_192), .B(n_139), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_194), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_182), .B(n_139), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_203), .B(n_138), .Y(n_273) );
BUFx3_ASAP7_75t_L g274 ( .A(n_175), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_203), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_179), .B(n_135), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_231), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g278 ( .A1(n_199), .A2(n_135), .B1(n_133), .B2(n_142), .Y(n_278) );
BUFx4f_ASAP7_75t_L g279 ( .A(n_199), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g280 ( .A1(n_234), .A2(n_162), .B1(n_150), .B2(n_142), .Y(n_280) );
NOR2x1p5_ASAP7_75t_L g281 ( .A(n_177), .B(n_135), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g282 ( .A(n_227), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_193), .B(n_133), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_175), .B(n_228), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_215), .B(n_133), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_199), .A2(n_162), .B1(n_150), .B2(n_142), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
INVx2_ASAP7_75t_L g288 ( .A(n_196), .Y(n_288) );
BUFx2_ASAP7_75t_L g289 ( .A(n_231), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_197), .B(n_162), .Y(n_290) );
AND2x6_ASAP7_75t_L g291 ( .A(n_185), .B(n_162), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_232), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_189), .A2(n_162), .B(n_150), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_186), .B(n_184), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_216), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_175), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_196), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_211), .B(n_162), .Y(n_298) );
BUFx6f_ASAP7_75t_L g299 ( .A(n_199), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g300 ( .A1(n_186), .A2(n_162), .B1(n_150), .B2(n_15), .Y(n_300) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_199), .A2(n_205), .B1(n_208), .B2(n_201), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_216), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_199), .A2(n_150), .B1(n_14), .B2(n_15), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g304 ( .A(n_252), .B(n_230), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_253), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_245), .A2(n_226), .B(n_223), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_247), .Y(n_307) );
AO21x2_ASAP7_75t_L g308 ( .A1(n_241), .A2(n_224), .B(n_220), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_255), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_247), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
OR2x6_ASAP7_75t_L g312 ( .A(n_247), .B(n_234), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_258), .Y(n_313) );
BUFx6f_ASAP7_75t_L g314 ( .A(n_299), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_251), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_277), .B(n_187), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_264), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_264), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g319 ( .A(n_240), .B(n_233), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_251), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_243), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_292), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_277), .B(n_226), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_287), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_258), .B(n_219), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_258), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_252), .B(n_233), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_257), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_300), .A2(n_188), .B(n_213), .C(n_183), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_243), .Y(n_331) );
AOI221x1_ASAP7_75t_L g332 ( .A1(n_293), .A2(n_234), .B1(n_150), .B2(n_235), .C(n_198), .Y(n_332) );
NOR2xp67_ASAP7_75t_L g333 ( .A(n_236), .B(n_12), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_244), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_244), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g336 ( .A1(n_284), .A2(n_233), .B1(n_234), .B2(n_223), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_275), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_274), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g339 ( .A1(n_241), .A2(n_248), .B(n_259), .C(n_285), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_289), .B(n_223), .Y(n_340) );
HB1xp67_ASAP7_75t_L g341 ( .A(n_271), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_268), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_293), .A2(n_259), .B(n_250), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_299), .Y(n_344) );
OR2x6_ASAP7_75t_SL g345 ( .A(n_282), .B(n_227), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_260), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_248), .A2(n_150), .B(n_229), .C(n_183), .Y(n_347) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_242), .Y(n_348) );
NAND2x1_ASAP7_75t_SL g349 ( .A(n_278), .B(n_229), .Y(n_349) );
A2O1A1Ixp33_ASAP7_75t_L g350 ( .A1(n_285), .A2(n_229), .B(n_235), .C(n_198), .Y(n_350) );
INVxp67_ASAP7_75t_L g351 ( .A(n_296), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_254), .B(n_16), .Y(n_352) );
O2A1O1Ixp5_ASAP7_75t_L g353 ( .A1(n_250), .A2(n_206), .B(n_200), .C(n_191), .Y(n_353) );
O2A1O1Ixp33_ASAP7_75t_L g354 ( .A1(n_294), .A2(n_206), .B(n_200), .C(n_191), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_238), .B(n_16), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_244), .Y(n_356) );
OR2x6_ASAP7_75t_L g357 ( .A(n_299), .B(n_218), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_260), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_249), .B(n_218), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_280), .A2(n_217), .B1(n_190), .B2(n_181), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g361 ( .A(n_307), .B(n_279), .Y(n_361) );
NOR2xp67_ASAP7_75t_L g362 ( .A(n_307), .B(n_266), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_321), .Y(n_363) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_319), .A2(n_301), .B(n_302), .Y(n_364) );
BUFx2_ASAP7_75t_L g365 ( .A(n_307), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_338), .Y(n_366) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_314), .Y(n_367) );
INVxp67_ASAP7_75t_SL g368 ( .A(n_310), .Y(n_368) );
AOI21x1_ASAP7_75t_L g369 ( .A1(n_332), .A2(n_190), .B(n_181), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_343), .A2(n_263), .B(n_286), .Y(n_370) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_350), .A2(n_263), .B(n_279), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_343), .A2(n_290), .B(n_298), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_329), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_332), .A2(n_301), .B(n_288), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
OAI22xp33_ASAP7_75t_SL g376 ( .A1(n_312), .A2(n_237), .B1(n_256), .B2(n_276), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_313), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_326), .A2(n_281), .B1(n_295), .B2(n_249), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_359), .A2(n_270), .B(n_262), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_353), .A2(n_297), .B(n_269), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_314), .Y(n_381) );
OAI21x1_ASAP7_75t_L g382 ( .A1(n_349), .A2(n_267), .B(n_272), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_322), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_322), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g385 ( .A1(n_312), .A2(n_273), .B1(n_283), .B2(n_266), .Y(n_385) );
AOI21x1_ASAP7_75t_L g386 ( .A1(n_312), .A2(n_261), .B(n_265), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_305), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_339), .A2(n_239), .B(n_246), .C(n_303), .Y(n_388) );
OAI21x1_ASAP7_75t_L g389 ( .A1(n_349), .A2(n_303), .B(n_280), .Y(n_389) );
OAI21x1_ASAP7_75t_SL g390 ( .A1(n_336), .A2(n_246), .B(n_291), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_331), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_305), .Y(n_392) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_313), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_309), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_352), .B(n_291), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_309), .Y(n_396) );
AOI221xp5_ASAP7_75t_L g397 ( .A1(n_376), .A2(n_316), .B1(n_326), .B2(n_352), .C(n_355), .Y(n_397) );
OR2x6_ASAP7_75t_L g398 ( .A(n_361), .B(n_327), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_378), .A2(n_326), .B1(n_355), .B2(n_330), .C(n_337), .Y(n_399) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_364), .A2(n_342), .B(n_312), .C(n_324), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g401 ( .A1(n_385), .A2(n_327), .B1(n_360), .B2(n_318), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_383), .Y(n_402) );
INVx4_ASAP7_75t_L g403 ( .A(n_365), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_373), .B(n_318), .Y(n_404) );
OAI33xp33_ASAP7_75t_L g405 ( .A1(n_373), .A2(n_354), .A3(n_304), .B1(n_328), .B2(n_311), .B3(n_325), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_383), .A2(n_333), .B1(n_357), .B2(n_345), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_384), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_365), .A2(n_317), .B1(n_341), .B2(n_358), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_375), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_375), .Y(n_411) );
AO21x2_ASAP7_75t_L g412 ( .A1(n_369), .A2(n_308), .B(n_347), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_388), .B(n_357), .C(n_317), .Y(n_413) );
INVx4_ASAP7_75t_SL g414 ( .A(n_384), .Y(n_414) );
OAI22xp33_ASAP7_75t_SL g415 ( .A1(n_363), .A2(n_345), .B1(n_351), .B2(n_357), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_392), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_387), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g418 ( .A1(n_391), .A2(n_340), .B1(n_348), .B2(n_358), .C(n_346), .Y(n_418) );
BUFx12f_ASAP7_75t_L g419 ( .A(n_377), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_362), .B(n_346), .Y(n_420) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_377), .B(n_346), .C(n_340), .Y(n_421) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_369), .A2(n_308), .B(n_306), .Y(n_422) );
AOI222xp33_ASAP7_75t_L g423 ( .A1(n_387), .A2(n_320), .B1(n_315), .B2(n_356), .C1(n_335), .C2(n_291), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_394), .Y(n_424) );
OAI21x1_ASAP7_75t_L g425 ( .A1(n_372), .A2(n_334), .B(n_356), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_392), .A2(n_357), .B1(n_335), .B2(n_320), .Y(n_426) );
OAI211xp5_ASAP7_75t_SL g427 ( .A1(n_418), .A2(n_366), .B(n_393), .C(n_368), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_409), .B(n_396), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_402), .B(n_396), .Y(n_429) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_402), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_407), .B(n_394), .Y(n_431) );
INVx2_ASAP7_75t_SL g432 ( .A(n_414), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_407), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_414), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_416), .B(n_372), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_416), .B(n_382), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_411), .B(n_382), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_414), .B(n_386), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_425), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_417), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_410), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_424), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_397), .A2(n_390), .B1(n_371), .B2(n_308), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_404), .Y(n_444) );
OA21x2_ASAP7_75t_L g445 ( .A1(n_413), .A2(n_389), .B(n_374), .Y(n_445) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_415), .A2(n_390), .B1(n_389), .B2(n_361), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_403), .B(n_370), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_399), .B(n_370), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_419), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_410), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_403), .B(n_374), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_398), .B(n_421), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_398), .B(n_395), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_398), .B(n_386), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_400), .B(n_379), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_426), .Y(n_456) );
INVx4_ASAP7_75t_SL g457 ( .A(n_420), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_410), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_421), .B(n_361), .Y(n_459) );
OR2x6_ASAP7_75t_L g460 ( .A(n_401), .B(n_381), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_422), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_440), .B(n_412), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_435), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_435), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g465 ( .A1(n_455), .A2(n_406), .B(n_408), .Y(n_465) );
NAND3xp33_ASAP7_75t_SL g466 ( .A(n_446), .B(n_408), .C(n_423), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_434), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_430), .B(n_412), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_437), .B(n_422), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_440), .B(n_406), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_433), .B(n_410), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_461), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_461), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_442), .B(n_420), .Y(n_474) );
AO21x2_ASAP7_75t_L g475 ( .A1(n_455), .A2(n_380), .B(n_405), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_427), .A2(n_315), .A3(n_334), .B(n_419), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_438), .Y(n_477) );
INVx2_ASAP7_75t_L g478 ( .A(n_439), .Y(n_478) );
NAND3xp33_ASAP7_75t_L g479 ( .A(n_427), .B(n_362), .C(n_217), .Y(n_479) );
NOR3xp33_ASAP7_75t_SL g480 ( .A(n_449), .B(n_405), .C(n_18), .Y(n_480) );
INVx4_ASAP7_75t_L g481 ( .A(n_434), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_439), .Y(n_482) );
BUFx2_ASAP7_75t_L g483 ( .A(n_438), .Y(n_483) );
NAND3xp33_ASAP7_75t_L g484 ( .A(n_446), .B(n_217), .C(n_367), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_437), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g486 ( .A(n_444), .B(n_17), .C(n_18), .D(n_19), .Y(n_486) );
AO21x2_ASAP7_75t_L g487 ( .A1(n_439), .A2(n_380), .B(n_381), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_442), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_444), .A2(n_381), .B1(n_367), .B2(n_323), .Y(n_489) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_447), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_429), .B(n_19), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_429), .B(n_20), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_436), .B(n_381), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_448), .A2(n_452), .B1(n_431), .B2(n_443), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_452), .B(n_20), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_431), .B(n_381), .Y(n_496) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_447), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_436), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_454), .Y(n_499) );
AOI322xp5_ASAP7_75t_L g500 ( .A1(n_428), .A2(n_344), .A3(n_217), .B1(n_28), .B2(n_29), .C1(n_34), .C2(n_37), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_441), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_451), .Y(n_502) );
INVx3_ASAP7_75t_L g503 ( .A(n_438), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_448), .B(n_367), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_428), .B(n_367), .Y(n_505) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_456), .A2(n_291), .B(n_217), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_454), .B(n_23), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_456), .B(n_24), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_453), .B(n_291), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_491), .B(n_459), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_491), .B(n_459), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_492), .B(n_453), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_488), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_492), .B(n_457), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_488), .B(n_457), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_486), .A2(n_432), .B(n_438), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_472), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_486), .A2(n_432), .B1(n_460), .B2(n_457), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_478), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_485), .B(n_457), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_485), .B(n_457), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_502), .B(n_445), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_472), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_473), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_495), .B(n_432), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_478), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_502), .B(n_445), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_466), .A2(n_460), .B1(n_445), .B2(n_450), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_495), .B(n_38), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_474), .B(n_458), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_508), .B(n_445), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_474), .B(n_458), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_508), .B(n_458), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_470), .B(n_450), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_498), .B(n_469), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_473), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_473), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_462), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_481), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_490), .B(n_460), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_490), .B(n_460), .Y(n_543) );
OAI33xp33_ASAP7_75t_L g544 ( .A1(n_470), .A2(n_450), .A3(n_441), .B1(n_44), .B2(n_45), .B3(n_46), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_498), .B(n_460), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_497), .B(n_441), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_478), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_462), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_499), .B(n_42), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_498), .B(n_43), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_463), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_466), .A2(n_344), .B1(n_323), .B2(n_314), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_494), .A2(n_323), .B1(n_314), .B2(n_58), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_469), .B(n_48), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_481), .Y(n_555) );
NOR2xp67_ASAP7_75t_L g556 ( .A(n_484), .B(n_56), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_482), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_469), .B(n_60), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_482), .Y(n_559) );
INVx2_ASAP7_75t_L g560 ( .A(n_482), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_497), .B(n_63), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_469), .B(n_68), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_504), .B(n_69), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_504), .B(n_71), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_499), .B(n_75), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_463), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_496), .B(n_314), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_463), .B(n_323), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_514), .B(n_494), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_514), .B(n_468), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_537), .B(n_468), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_518), .Y(n_572) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_541), .Y(n_573) );
OR2x6_ASAP7_75t_L g574 ( .A(n_541), .B(n_483), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_537), .B(n_503), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_518), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_555), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_540), .B(n_464), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_527), .B(n_481), .Y(n_579) );
NOR4xp25_ASAP7_75t_L g580 ( .A(n_517), .B(n_465), .C(n_479), .D(n_484), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_520), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_513), .B(n_464), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_545), .B(n_503), .Y(n_583) );
OR2x6_ASAP7_75t_L g584 ( .A(n_555), .B(n_483), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_520), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_526), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_545), .B(n_503), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_529), .B(n_503), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_525), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_529), .B(n_477), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_551), .B(n_464), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_533), .B(n_477), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_533), .B(n_501), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_551), .B(n_540), .Y(n_594) );
INVxp67_ASAP7_75t_L g595 ( .A(n_515), .Y(n_595) );
NOR3xp33_ASAP7_75t_L g596 ( .A(n_544), .B(n_479), .C(n_465), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_526), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_548), .B(n_481), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_548), .B(n_501), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_561), .Y(n_601) );
XNOR2x1_ASAP7_75t_L g602 ( .A(n_519), .B(n_507), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_566), .B(n_501), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_566), .B(n_493), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_536), .B(n_505), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_546), .B(n_505), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_511), .B(n_467), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_525), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_539), .B(n_493), .Y(n_609) );
NAND3xp33_ASAP7_75t_L g610 ( .A(n_530), .B(n_480), .C(n_476), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_538), .B(n_493), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_546), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_538), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_512), .B(n_467), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_532), .B(n_467), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_524), .B(n_493), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_524), .B(n_496), .Y(n_617) );
OR2x2_ASAP7_75t_L g618 ( .A(n_542), .B(n_475), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_534), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_535), .B(n_471), .Y(n_620) );
INVx2_ASAP7_75t_L g621 ( .A(n_521), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_561), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_580), .B(n_519), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_595), .B(n_619), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_577), .Y(n_625) );
NAND2xp5_ASAP7_75t_SL g626 ( .A(n_573), .B(n_476), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_610), .A2(n_531), .B1(n_480), .B2(n_516), .C(n_552), .Y(n_627) );
NOR5xp2_ASAP7_75t_L g628 ( .A(n_622), .B(n_556), .C(n_500), .D(n_553), .E(n_562), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_599), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_571), .B(n_554), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_602), .A2(n_556), .B1(n_553), .B2(n_523), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_594), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_599), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_569), .B(n_522), .Y(n_634) );
OA22x2_ASAP7_75t_L g635 ( .A1(n_574), .A2(n_562), .B1(n_558), .B2(n_554), .Y(n_635) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_602), .A2(n_579), .B1(n_607), .B2(n_614), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_594), .Y(n_637) );
NAND2x1p5_ASAP7_75t_L g638 ( .A(n_612), .B(n_558), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_620), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_572), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g641 ( .A1(n_596), .A2(n_565), .B1(n_543), .B2(n_542), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_576), .Y(n_642) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_574), .A2(n_543), .B(n_565), .Y(n_643) );
NAND2x1_ASAP7_75t_L g644 ( .A(n_574), .B(n_550), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_612), .B(n_528), .Y(n_645) );
AOI211xp5_ASAP7_75t_SL g646 ( .A1(n_601), .A2(n_563), .B(n_564), .C(n_507), .Y(n_646) );
AOI21xp33_ASAP7_75t_SL g647 ( .A1(n_574), .A2(n_563), .B(n_564), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_598), .B(n_550), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_584), .A2(n_489), .B1(n_509), .B2(n_549), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_581), .Y(n_650) );
OAI22xp33_ASAP7_75t_L g651 ( .A1(n_584), .A2(n_489), .B1(n_567), .B2(n_547), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_608), .Y(n_652) );
AOI322xp5_ASAP7_75t_L g653 ( .A1(n_571), .A2(n_509), .A3(n_521), .B1(n_560), .B2(n_559), .C1(n_547), .C2(n_557), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_584), .A2(n_506), .B(n_521), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_613), .Y(n_655) );
OAI221xp5_ASAP7_75t_SL g656 ( .A1(n_584), .A2(n_500), .B1(n_471), .B2(n_510), .C(n_559), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_617), .B(n_528), .Y(n_657) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_611), .A2(n_528), .B1(n_560), .B2(n_559), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_617), .B(n_560), .Y(n_659) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_606), .A2(n_557), .B1(n_547), .B2(n_510), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_585), .Y(n_661) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_623), .A2(n_582), .B(n_615), .C(n_570), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_636), .B(n_587), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_639), .B(n_592), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_661), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_629), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_624), .B(n_587), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_632), .B(n_592), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_637), .B(n_590), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_635), .A2(n_606), .B1(n_587), .B2(n_590), .Y(n_670) );
OAI321xp33_ASAP7_75t_L g671 ( .A1(n_656), .A2(n_618), .A3(n_605), .B1(n_616), .B2(n_588), .C(n_578), .Y(n_671) );
NAND4xp25_ASAP7_75t_L g672 ( .A(n_641), .B(n_618), .C(n_605), .D(n_611), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_658), .B(n_593), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_653), .B(n_593), .Y(n_674) );
INVxp67_ASAP7_75t_L g675 ( .A(n_625), .Y(n_675) );
AOI211xp5_ASAP7_75t_L g676 ( .A1(n_647), .A2(n_588), .B(n_575), .C(n_583), .Y(n_676) );
OAI32xp33_ASAP7_75t_L g677 ( .A1(n_638), .A2(n_575), .A3(n_578), .B1(n_599), .B2(n_583), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_634), .B(n_616), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_640), .B(n_589), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_642), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_650), .B(n_589), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_652), .Y(n_682) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_635), .A2(n_591), .B(n_604), .Y(n_683) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_645), .Y(n_684) );
AOI222xp33_ASAP7_75t_L g685 ( .A1(n_626), .A2(n_585), .B1(n_604), .B2(n_609), .C1(n_603), .C2(n_597), .Y(n_685) );
OA22x2_ASAP7_75t_L g686 ( .A1(n_683), .A2(n_631), .B1(n_644), .B2(n_630), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_671), .A2(n_670), .B1(n_662), .B2(n_663), .C(n_672), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_679), .Y(n_688) );
INVxp67_ASAP7_75t_L g689 ( .A(n_675), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_663), .A2(n_638), .B1(n_660), .B2(n_646), .Y(n_690) );
AOI31xp33_ASAP7_75t_L g691 ( .A1(n_676), .A2(n_627), .A3(n_649), .B(n_643), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_681), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_674), .B(n_655), .Y(n_693) );
AOI211xp5_ASAP7_75t_L g694 ( .A1(n_677), .A2(n_656), .B(n_651), .C(n_654), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_684), .A2(n_659), .B1(n_657), .B2(n_654), .C(n_648), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_684), .A2(n_633), .B1(n_649), .B2(n_609), .C(n_603), .Y(n_696) );
AOI221xp5_ASAP7_75t_L g697 ( .A1(n_667), .A2(n_597), .B1(n_586), .B2(n_621), .C(n_600), .Y(n_697) );
OAI21xp5_ASAP7_75t_L g698 ( .A1(n_685), .A2(n_628), .B(n_600), .Y(n_698) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_673), .Y(n_699) );
XNOR2x1_ASAP7_75t_L g700 ( .A(n_664), .B(n_628), .Y(n_700) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_691), .A2(n_667), .B1(n_682), .B2(n_680), .C(n_665), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_689), .B(n_678), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_687), .A2(n_669), .B1(n_668), .B2(n_666), .C(n_586), .Y(n_703) );
INVx2_ASAP7_75t_SL g704 ( .A(n_686), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_698), .A2(n_621), .B(n_568), .C(n_557), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_699), .A2(n_568), .B1(n_475), .B2(n_506), .C(n_487), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_688), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g708 ( .A1(n_695), .A2(n_475), .B1(n_506), .B2(n_487), .C(n_323), .Y(n_708) );
NAND5xp2_ASAP7_75t_SL g709 ( .A(n_696), .B(n_475), .C(n_487), .D(n_506), .E(n_700), .Y(n_709) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_704), .B(n_690), .Y(n_710) );
INVx1_ASAP7_75t_L g711 ( .A(n_707), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_702), .Y(n_712) );
NAND5xp2_ASAP7_75t_L g713 ( .A(n_701), .B(n_694), .C(n_697), .D(n_693), .E(n_692), .Y(n_713) );
INVx1_ASAP7_75t_L g714 ( .A(n_703), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_711), .Y(n_715) );
OAI21xp5_ASAP7_75t_L g716 ( .A1(n_710), .A2(n_705), .B(n_694), .Y(n_716) );
AND3x2_ASAP7_75t_L g717 ( .A(n_712), .B(n_708), .C(n_709), .Y(n_717) );
INVx2_ASAP7_75t_L g718 ( .A(n_715), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_716), .B(n_714), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
AND2x4_ASAP7_75t_L g721 ( .A(n_719), .B(n_712), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_721), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g723 ( .A1(n_722), .A2(n_720), .B(n_721), .Y(n_723) );
AOI22xp5_ASAP7_75t_SL g724 ( .A1(n_723), .A2(n_713), .B1(n_710), .B2(n_717), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_706), .B(n_487), .Y(n_725) );
endmodule