module real_jpeg_21841_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_150;
wire n_74;
wire n_41;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_0),
.A2(n_6),
.B1(n_23),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_0),
.A2(n_5),
.B1(n_38),
.B2(n_50),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_0),
.A2(n_4),
.B1(n_34),
.B2(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_1),
.A2(n_5),
.B1(n_38),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_1),
.A2(n_4),
.B1(n_34),
.B2(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_1),
.A2(n_6),
.B1(n_23),
.B2(n_40),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_2),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_20),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_2),
.A2(n_10),
.B1(n_25),
.B2(n_26),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_2),
.A2(n_20),
.B(n_25),
.C(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_4),
.A2(n_9),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_64),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_4),
.A2(n_10),
.B1(n_25),
.B2(n_34),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_4),
.A2(n_9),
.B(n_10),
.Y(n_150)
);

OAI22xp33_ASAP7_75t_L g37 ( 
.A1(n_5),
.A2(n_9),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_5),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_7),
.B1(n_38),
.B2(n_47),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_10),
.B1(n_25),
.B2(n_38),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_5),
.A2(n_25),
.B(n_35),
.C(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_6),
.A2(n_8),
.B1(n_20),
.B2(n_23),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_6),
.A2(n_10),
.B1(n_23),
.B2(n_25),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_6),
.A2(n_7),
.B1(n_23),
.B2(n_47),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_SL g126 ( 
.A1(n_6),
.A2(n_10),
.B(n_127),
.Y(n_126)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

O2A1O1Ixp33_ASAP7_75t_L g171 ( 
.A1(n_7),
.A2(n_10),
.B(n_23),
.C(n_172),
.Y(n_171)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_10),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_10),
.B(n_48),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_82),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_13),
.B(n_81),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_71),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_71),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_52),
.C(n_59),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_16),
.A2(n_52),
.B1(n_53),
.B2(n_102),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_16),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_27),
.B1(n_28),
.B2(n_51),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_17),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_17),
.A2(n_61),
.B(n_67),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_17),
.A2(n_51),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_17),
.A2(n_51),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_17),
.B(n_56),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_17),
.A2(n_51),
.B1(n_61),
.B2(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_17),
.A2(n_51),
.B1(n_56),
.B2(n_57),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_17),
.A2(n_51),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g209 ( 
.A1(n_17),
.A2(n_56),
.B(n_93),
.C(n_123),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_24),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_22),
.Y(n_18)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_20),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_22),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_25),
.B(n_33),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_25),
.B(n_90),
.Y(n_162)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_25),
.A2(n_38),
.B(n_47),
.Y(n_172)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_41),
.B2(n_42),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_29),
.A2(n_30),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_29),
.B(n_42),
.C(n_51),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_31),
.B(n_39),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_32),
.B(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_33),
.B(n_37),
.Y(n_36)
);

OA22x2_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_36),
.B1(n_39),
.B2(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_33),
.A2(n_36),
.B1(n_55),
.B2(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_34),
.B(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_48),
.B2(n_49),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_48),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_45),
.A2(n_48),
.B1(n_49),
.B2(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_57),
.Y(n_92)
);

AOI211xp5_ASAP7_75t_SL g111 ( 
.A1(n_51),
.A2(n_91),
.B(n_94),
.C(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_54),
.B(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_56),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_56),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_56),
.A2(n_57),
.B1(n_91),
.B2(n_113),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_56),
.A2(n_113),
.B(n_174),
.C(n_178),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_56),
.A2(n_57),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_57),
.B(n_128),
.C(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_60),
.B1(n_101),
.B2(n_103),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_61),
.A2(n_68),
.B1(n_99),
.B2(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_63),
.B(n_118),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_66),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_89),
.B1(n_90),
.B2(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_68),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_80),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_104),
.B(n_228),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_100),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_84),
.B(n_100),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_95),
.C(n_97),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_85),
.A2(n_86),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

OAI21xp33_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_92),
.B(n_93),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_87),
.A2(n_121),
.B1(n_122),
.B2(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_87),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_88),
.A2(n_91),
.B1(n_113),
.B2(n_203),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_91),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_113),
.B1(n_116),
.B2(n_119),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_91),
.A2(n_113),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_91),
.A2(n_113),
.B1(n_149),
.B2(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_91),
.B(n_128),
.C(n_153),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_91),
.A2(n_113),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_91),
.B(n_180),
.C(n_186),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_91),
.B(n_116),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_92),
.A2(n_93),
.B(n_205),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_95),
.A2(n_96),
.B1(n_97),
.B2(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_97),
.Y(n_226)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_101),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_222),
.B(n_227),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_212),
.B(n_221),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_142),
.B(n_197),
.C(n_211),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_130),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_108),
.B(n_130),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_120),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_115),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_110),
.B(n_115),
.C(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_112),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_113),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_116),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_129),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_121),
.A2(n_122),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_125),
.B1(n_128),
.B2(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_128),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_128),
.A2(n_137),
.B1(n_152),
.B2(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_128),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_137),
.B1(n_171),
.B2(n_173),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_128),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_183)
);

NAND2x1_ASAP7_75t_SL g187 ( 
.A(n_128),
.B(n_171),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.C(n_138),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_131),
.A2(n_132),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_133),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_134),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_193),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_138),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_196),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_189),
.B(n_195),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_176),
.B(n_188),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_167),
.B(n_175),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_156),
.B(n_166),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_151),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_149),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_152),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_169),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_170),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_171),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_179),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_190),
.B(n_191),
.Y(n_195)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_192),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_199),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_209),
.B2(n_210),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_204),
.B1(n_207),
.B2(n_208),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_208),
.C(n_210),
.Y(n_213)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_205),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g210 ( 
.A(n_209),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_213),
.B(n_214),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_215),
.B(n_223),
.Y(n_227)
);

FAx1_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_218),
.CI(n_220),
.CON(n_215),
.SN(n_215)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);


endmodule