module fake_jpeg_7264_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_39),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_9),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_46),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_43),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_21),
.B(n_16),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_56),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_21),
.B1(n_28),
.B2(n_27),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_55),
.A2(n_62),
.B1(n_27),
.B2(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_61),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_46),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_29),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_82),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_75),
.A2(n_86),
.B1(n_91),
.B2(n_30),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_41),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_81),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_41),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_51),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_84),
.B(n_95),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_37),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_85),
.B(n_90),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_23),
.B1(n_34),
.B2(n_17),
.Y(n_86)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_88),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_37),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_23),
.B1(n_17),
.B2(n_34),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_100),
.B(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_47),
.B1(n_17),
.B2(n_34),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_85),
.A2(n_64),
.B1(n_60),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_113),
.B1(n_124),
.B2(n_89),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_108),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_95),
.B(n_84),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_112),
.A2(n_125),
.B1(n_25),
.B2(n_30),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_81),
.A2(n_60),
.B1(n_40),
.B2(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_79),
.B(n_20),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_74),
.B(n_20),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_120),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_77),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_40),
.B1(n_50),
.B2(n_54),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_77),
.A2(n_52),
.B1(n_67),
.B2(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_126),
.Y(n_127)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_90),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_136),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_90),
.B(n_30),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_130),
.A2(n_149),
.B(n_153),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_131),
.A2(n_144),
.B1(n_35),
.B2(n_117),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_113),
.A2(n_38),
.B(n_76),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_140),
.B(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_78),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_19),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_151),
.Y(n_170)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_139),
.B(n_147),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_44),
.Y(n_140)
);

AO22x2_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_35),
.B1(n_66),
.B2(n_68),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_143),
.B1(n_83),
.B2(n_71),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_106),
.A2(n_83),
.B1(n_89),
.B2(n_71),
.Y(n_143)
);

INVx6_ASAP7_75t_SL g146 ( 
.A(n_102),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_146),
.Y(n_156)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_114),
.A2(n_25),
.B(n_33),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_19),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_111),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_128),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_159),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_158),
.A2(n_176),
.B1(n_177),
.B2(n_138),
.Y(n_201)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_122),
.C(n_45),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_178),
.C(n_127),
.Y(n_189)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_164),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_150),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_169),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_179),
.B(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_166),
.B(n_167),
.Y(n_207)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_99),
.Y(n_168)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_168),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_138),
.Y(n_169)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_127),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_172),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_140),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_174),
.Y(n_193)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_135),
.A2(n_103),
.B1(n_109),
.B2(n_126),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_175),
.A2(n_147),
.B1(n_141),
.B2(n_144),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_121),
.B1(n_111),
.B2(n_117),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_24),
.Y(n_178)
);

XOR2x2_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_129),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_135),
.A2(n_29),
.B(n_32),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_139),
.Y(n_199)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_186),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_184),
.A2(n_208),
.B(n_180),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_131),
.B1(n_130),
.B2(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_162),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_160),
.C(n_178),
.Y(n_214)
);

AND2x6_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_153),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_191),
.Y(n_229)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_162),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_206),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_156),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_199),
.B(n_205),
.Y(n_220)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_201),
.B(n_204),
.Y(n_234)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_148),
.Y(n_219)
);

OAI32xp33_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_149),
.A3(n_153),
.B1(n_22),
.B2(n_24),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_155),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_166),
.B(n_132),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_165),
.A2(n_133),
.B(n_152),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_133),
.B1(n_148),
.B2(n_102),
.Y(n_210)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_210),
.Y(n_225)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_173),
.B(n_159),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_181),
.B(n_174),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_217),
.C(n_223),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_170),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g221 ( 
.A(n_207),
.B(n_192),
.C(n_211),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_231),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_222),
.A2(n_235),
.B(n_236),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_186),
.B(n_157),
.C(n_161),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_224),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_192),
.C(n_208),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_238),
.C(n_188),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_227),
.A2(n_22),
.B(n_18),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_197),
.A2(n_31),
.B(n_102),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_233),
.B(n_220),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_31),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_18),
.Y(n_232)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_193),
.B(n_14),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_233),
.B(n_12),
.Y(n_259)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_187),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_237),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_148),
.C(n_68),
.Y(n_238)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_218),
.Y(n_240)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_229),
.A2(n_185),
.B1(n_200),
.B2(n_184),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_243),
.A2(n_259),
.B1(n_224),
.B2(n_215),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_202),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_244),
.B(n_252),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_248),
.C(n_251),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_203),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_229),
.A2(n_191),
.B1(n_195),
.B2(n_209),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_215),
.B1(n_225),
.B2(n_236),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_198),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_230),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_194),
.C(n_68),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_258),
.C(n_260),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_212),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_255),
.B(n_256),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_18),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_217),
.B(n_123),
.C(n_108),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_24),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_228),
.Y(n_270)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_243),
.A2(n_234),
.B1(n_213),
.B2(n_225),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_263),
.B(n_279),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_216),
.B(n_213),
.C(n_212),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_265),
.A2(n_259),
.B1(n_22),
.B2(n_2),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_247),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_265),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_22),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_277),
.C(n_22),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_235),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_254),
.B(n_261),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_222),
.C(n_232),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_276),
.C(n_253),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_257),
.A2(n_216),
.B1(n_237),
.B2(n_227),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_275),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_97),
.C(n_53),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_18),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_242),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_281),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_248),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_282),
.B(n_276),
.C(n_278),
.Y(n_299)
);

BUFx12_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_283),
.B(n_286),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_285),
.Y(n_305)
);

BUFx12_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_245),
.B(n_239),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_287),
.B(n_290),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_293),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_286),
.B(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_266),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_303),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_266),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_298),
.A2(n_308),
.B1(n_283),
.B2(n_1),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_283),
.C(n_1),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_288),
.A2(n_273),
.B1(n_270),
.B2(n_3),
.Y(n_302)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_302),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_280),
.B(n_22),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_284),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_8),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_10),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_288),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_317),
.C(n_312),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_311),
.A2(n_8),
.B1(n_3),
.B2(n_5),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_10),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_315),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_11),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_11),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_313),
.A2(n_298),
.B(n_300),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_320),
.A2(n_326),
.B(n_6),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_300),
.B1(n_308),
.B2(n_304),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_317),
.B1(n_5),
.B2(n_6),
.Y(n_327)
);

AO21x1_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_307),
.B(n_3),
.Y(n_323)
);

OAI321xp33_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_7),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C(n_16),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_324),
.B(n_325),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_12),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_327),
.Y(n_331)
);

XOR2x2_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_330),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_319),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_323),
.B(n_329),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_334),
.Y(n_335)
);

OAI32xp33_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_331),
.A3(n_322),
.B1(n_326),
.B2(n_15),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_7),
.B(n_14),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_0),
.Y(n_338)
);


endmodule