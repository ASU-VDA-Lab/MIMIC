module real_jpeg_3558_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_1),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_1),
.A2(n_36),
.B1(n_38),
.B2(n_144),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_1),
.A2(n_71),
.B1(n_73),
.B2(n_144),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_1),
.A2(n_59),
.B1(n_66),
.B2(n_144),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_3),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_4),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_4),
.A2(n_36),
.B1(n_38),
.B2(n_85),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_4),
.A2(n_71),
.B1(n_73),
.B2(n_85),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_4),
.A2(n_59),
.B1(n_66),
.B2(n_85),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_44),
.B1(n_71),
.B2(n_73),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_5),
.A2(n_36),
.B1(n_38),
.B2(n_44),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_5),
.A2(n_44),
.B1(n_59),
.B2(n_66),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_6),
.A2(n_36),
.B1(n_38),
.B2(n_197),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_6),
.A2(n_71),
.B1(n_73),
.B2(n_197),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_6),
.A2(n_59),
.B1(n_66),
.B2(n_197),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_7),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_7),
.A2(n_36),
.B1(n_38),
.B2(n_87),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_7),
.A2(n_71),
.B1(n_73),
.B2(n_87),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_7),
.A2(n_59),
.B1(n_66),
.B2(n_87),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_8),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_8),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_8),
.A2(n_36),
.B1(n_38),
.B2(n_70),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_70),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_8),
.A2(n_59),
.B1(n_66),
.B2(n_70),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_9),
.B(n_29),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_9),
.B(n_39),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_9),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_9),
.A2(n_29),
.B(n_187),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_9),
.B(n_96),
.Y(n_249)
);

AOI21xp33_ASAP7_75t_L g256 ( 
.A1(n_9),
.A2(n_38),
.B(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_9),
.B(n_59),
.C(n_76),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_9),
.A2(n_71),
.B1(n_73),
.B2(n_223),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_9),
.B(n_62),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_9),
.B(n_80),
.Y(n_279)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g76 ( 
.A(n_11),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_13),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_13),
.A2(n_36),
.B1(n_38),
.B2(n_178),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_13),
.A2(n_71),
.B1(n_73),
.B2(n_178),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_13),
.A2(n_59),
.B1(n_66),
.B2(n_178),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_20)
);

INVx4_ASAP7_75t_SL g21 ( 
.A(n_15),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_16),
.A2(n_36),
.B1(n_38),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_16),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_93),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_16),
.A2(n_71),
.B1(n_73),
.B2(n_93),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_16),
.A2(n_59),
.B1(n_66),
.B2(n_93),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_17),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_17),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_17),
.A2(n_41),
.B1(n_59),
.B2(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_17),
.A2(n_41),
.B1(n_71),
.B2(n_73),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_17),
.A2(n_36),
.B1(n_38),
.B2(n_41),
.Y(n_153)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_18),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_47),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_45),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_42),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_26),
.B(n_46),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_39),
.B(n_40),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_27),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_27),
.A2(n_39),
.B1(n_143),
.B2(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_27),
.A2(n_39),
.B1(n_43),
.B2(n_325),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_35),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g186 ( 
.A1(n_30),
.A2(n_33),
.A3(n_38),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OA22x2_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_33),
.B1(n_36),
.B2(n_38),
.Y(n_35)
);

NAND2xp33_ASAP7_75t_SL g188 ( 
.A(n_32),
.B(n_36),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_35),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_35),
.A2(n_83),
.B1(n_86),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_35),
.A2(n_83),
.B1(n_84),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_35),
.A2(n_83),
.B1(n_107),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_35),
.A2(n_83),
.B1(n_196),
.B2(n_198),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_35),
.A2(n_83),
.B1(n_196),
.B2(n_235),
.Y(n_234)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_36),
.A2(n_38),
.B1(n_97),
.B2(n_99),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_36),
.B(n_223),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g221 ( 
.A1(n_38),
.A2(n_71),
.A3(n_97),
.B1(n_222),
.B2(n_224),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_42),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_42),
.B(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_46),
.B(n_334),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_330),
.B(n_332),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_318),
.B(n_329),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_158),
.B(n_315),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_145),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_118),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_52),
.B(n_118),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_88),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_53),
.B(n_104),
.C(n_116),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_81),
.B(n_82),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_54),
.A2(n_55),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_67),
.Y(n_55)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_56),
.A2(n_81),
.B1(n_82),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_56),
.A2(n_67),
.B1(n_68),
.B2(n_81),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_61),
.B(n_64),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_57),
.A2(n_61),
.B1(n_132),
.B2(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_57),
.A2(n_61),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_57),
.A2(n_61),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_58),
.A2(n_62),
.B1(n_65),
.B2(n_131),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_58),
.A2(n_62),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_58),
.A2(n_62),
.B1(n_190),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_58),
.A2(n_62),
.B1(n_227),
.B2(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_58),
.A2(n_62),
.B1(n_223),
.B2(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_58),
.A2(n_62),
.B1(n_277),
.B2(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_66),
.B1(n_76),
.B2(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_59),
.B(n_275),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_74),
.B1(n_79),
.B2(n_80),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_69),
.A2(n_74),
.B1(n_80),
.B2(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_71),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_71),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

AO22x2_ASAP7_75t_SL g96 ( 
.A1(n_71),
.A2(n_73),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_71),
.B(n_265),
.Y(n_264)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_73),
.B(n_99),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_80),
.B(n_103),
.Y(n_110)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_74),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_74),
.A2(n_80),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_74),
.A2(n_80),
.B1(n_219),
.B2(n_239),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_74),
.A2(n_80),
.B1(n_247),
.B2(n_248),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_74),
.A2(n_80),
.B1(n_247),
.B2(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_78),
.A2(n_136),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_78),
.A2(n_171),
.B1(n_218),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_104),
.B1(n_116),
.B2(n_117),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_89),
.A2(n_90),
.B(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_102),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B1(n_96),
.B2(n_101),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_92),
.A2(n_95),
.B1(n_138),
.B2(n_140),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_94),
.A2(n_96),
.B1(n_101),
.B2(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_94),
.A2(n_96),
.B1(n_139),
.B2(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_94),
.A2(n_96),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_95),
.A2(n_114),
.B1(n_140),
.B2(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_95),
.A2(n_140),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_95),
.A2(n_140),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_95),
.A2(n_140),
.B1(n_193),
.B2(n_209),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_95),
.A2(n_140),
.B1(n_208),
.B2(n_256),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.Y(n_95)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_96),
.Y(n_140)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_104),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_105),
.A2(n_106),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_110),
.C(n_112),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_106),
.B(n_149),
.C(n_156),
.Y(n_319)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_111),
.B1(n_112),
.B2(n_115),
.Y(n_109)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_110),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_115),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_110),
.B(n_152),
.C(n_154),
.Y(n_328)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_124),
.C(n_126),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_120),
.B1(n_124),
.B2(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_161),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_137),
.C(n_141),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_128),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_129),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_199)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_141),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_145),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_157),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_146),
.B(n_157),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_156),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_154),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_153),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_155),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_179),
.B(n_314),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_160),
.B(n_162),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_166),
.Y(n_201)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_201),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_174),
.C(n_176),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_169),
.B(n_172),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_176),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_175),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_202),
.B(n_313),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_200),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_181),
.B(n_200),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_199),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_182),
.B(n_199),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_184),
.B(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.C(n_195),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_185),
.B(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_189),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_186),
.B(n_189),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_192),
.B(n_195),
.Y(n_303)
);

AOI31xp33_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_297),
.A3(n_306),
.B(n_310),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_242),
.B(n_296),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_229),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_205),
.B(n_229),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_216),
.C(n_220),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_206),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_211),
.C(n_215),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_214),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_216),
.B(n_220),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_225),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_231),
.B(n_232),
.C(n_233),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_234),
.B(n_237),
.C(n_241),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_236)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_237),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_238),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_291),
.B(n_295),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_260),
.B(n_290),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_252),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_252),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_249),
.C(n_250),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_249),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_248),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_270),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_255),
.C(n_258),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_271),
.B(n_289),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_269),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_266),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_283),
.B(n_288),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_278),
.B(n_282),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_287),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_294),
.Y(n_295)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_298),
.A2(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_301),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_301),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.C(n_305),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_305),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_328),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_324),
.B1(n_326),
.B2(n_327),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_324),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_326),
.C(n_328),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_331),
.Y(n_334)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);


endmodule