module real_jpeg_31646_n_20 (n_17, n_8, n_0, n_2, n_692, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_692;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_620;
wire n_328;
wire n_366;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_338;
wire n_175;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_314;
wire n_689;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_596;
wire n_617;
wire n_312;
wire n_325;
wire n_594;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_604;
wire n_420;
wire n_357;
wire n_431;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_616;
wire n_377;
wire n_109;
wire n_686;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_690;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g209 ( 
.A(n_0),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_0),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_0),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_1),
.A2(n_183),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_1),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_1),
.A2(n_292),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_1),
.A2(n_292),
.B1(n_530),
.B2(n_533),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_1),
.A2(n_292),
.B1(n_594),
.B2(n_595),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_2),
.Y(n_103)
);

OAI22x1_ASAP7_75t_SL g178 ( 
.A1(n_3),
.A2(n_179),
.B1(n_180),
.B2(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_3),
.Y(n_179)
);

AOI22x1_ASAP7_75t_SL g299 ( 
.A1(n_3),
.A2(n_179),
.B1(n_300),
.B2(n_304),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_3),
.A2(n_179),
.B1(n_339),
.B2(n_343),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_3),
.A2(n_179),
.B1(n_393),
.B2(n_398),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_4),
.A2(n_106),
.B1(n_109),
.B2(n_111),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_4),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_111),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_4),
.A2(n_111),
.B1(n_238),
.B2(n_240),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_4),
.A2(n_111),
.B1(n_430),
.B2(n_434),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_5),
.A2(n_73),
.B1(n_181),
.B2(n_373),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_5),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_5),
.A2(n_373),
.B1(n_378),
.B2(n_380),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g568 ( 
.A1(n_5),
.A2(n_373),
.B1(n_569),
.B2(n_571),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_SL g616 ( 
.A1(n_5),
.A2(n_373),
.B1(n_576),
.B2(n_617),
.Y(n_616)
);

AO22x1_ASAP7_75t_L g61 ( 
.A1(n_6),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_6),
.A2(n_64),
.B1(n_146),
.B2(n_149),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_64),
.B1(n_218),
.B2(n_221),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_7),
.A2(n_364),
.B(n_368),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_7),
.B(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g404 ( 
.A(n_7),
.Y(n_404)
);

OAI32xp33_ASAP7_75t_L g536 ( 
.A1(n_7),
.A2(n_408),
.A3(n_537),
.B1(n_540),
.B2(n_541),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_7),
.B(n_144),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g631 ( 
.A1(n_7),
.A2(n_210),
.B1(n_616),
.B2(n_632),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_7),
.A2(n_404),
.B1(n_657),
.B2(n_661),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_8),
.A2(n_134),
.B1(n_138),
.B2(n_142),
.Y(n_133)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_8),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_8),
.A2(n_142),
.B1(n_161),
.B2(n_167),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_8),
.A2(n_243),
.B(n_245),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_8),
.B(n_246),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_8),
.A2(n_142),
.B1(n_221),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_9),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_10),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_12),
.Y(n_433)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_13),
.Y(n_581)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_14),
.A2(n_73),
.B1(n_76),
.B2(n_77),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

OAI22x1_ASAP7_75t_SL g257 ( 
.A1(n_14),
.A2(n_76),
.B1(n_258),
.B2(n_264),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_14),
.A2(n_76),
.B1(n_274),
.B2(n_276),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_14),
.A2(n_76),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_15),
.A2(n_228),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_15),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_15),
.A2(n_231),
.B1(n_333),
.B2(n_336),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_15),
.A2(n_231),
.B1(n_454),
.B2(n_456),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_15),
.A2(n_231),
.B1(n_454),
.B2(n_456),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_15),
.A2(n_231),
.B1(n_545),
.B2(n_547),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g356 ( 
.A1(n_16),
.A2(n_354),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_16),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_16),
.A2(n_360),
.B1(n_463),
.B2(n_466),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_16),
.A2(n_360),
.B1(n_604),
.B2(n_607),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_SL g620 ( 
.A1(n_16),
.A2(n_360),
.B1(n_621),
.B2(n_624),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_17),
.A2(n_21),
.B(n_689),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_17),
.B(n_690),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_18),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_19),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_19),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_19),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_196),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_195),
.Y(n_22)
);

INVxp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_170),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_25),
.B(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_28),
.B1(n_154),
.B2(n_155),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_70),
.C(n_112),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_29),
.A2(n_113),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_29),
.A2(n_174),
.B1(n_189),
.B2(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_58),
.B(n_61),
.Y(n_29)
);

OA21x2_ASAP7_75t_L g174 ( 
.A1(n_30),
.A2(n_58),
.B(n_61),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_30),
.B(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_31),
.A2(n_59),
.B1(n_237),
.B2(n_242),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_31),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_31),
.A2(n_273),
.B1(n_338),
.B2(n_347),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_31),
.A2(n_347),
.B1(n_603),
.B2(n_609),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_40),
.B(n_48),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_37),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g608 ( 
.A(n_38),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_39),
.Y(n_131)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_39),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_39),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_39),
.Y(n_539)
);

INVxp33_ASAP7_75t_L g587 ( 
.A(n_40),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g345 ( 
.A(n_45),
.Y(n_345)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_46),
.Y(n_239)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_46),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_47),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_48),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_50),
.Y(n_390)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_50),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_50),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_50),
.Y(n_638)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_55),
.Y(n_215)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_55),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_55),
.Y(n_401)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_58),
.A2(n_61),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_58),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_58),
.B(n_280),
.Y(n_488)
);

AO22x1_ASAP7_75t_L g528 ( 
.A1(n_58),
.A2(n_331),
.B1(n_332),
.B2(n_529),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_58),
.A2(n_254),
.B1(n_529),
.B2(n_654),
.Y(n_653)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_59),
.B(n_404),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_60),
.Y(n_348)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_68),
.Y(n_241)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_69),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g567 ( 
.A(n_69),
.Y(n_567)
);

XOR2x2_ASAP7_75t_L g171 ( 
.A(n_70),
.B(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_83),
.B1(n_104),
.B2(n_105),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_72),
.A2(n_84),
.B1(n_178),
.B2(n_186),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_88),
.B1(n_91),
.B2(n_93),
.Y(n_87)
);

INVxp67_ASAP7_75t_SL g110 ( 
.A(n_74),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_75),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_75),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_75),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_75),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_75),
.Y(n_465)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_80),
.Y(n_182)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_81),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_82),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_83),
.A2(n_104),
.B1(n_105),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_84),
.A2(n_186),
.B1(n_461),
.B2(n_467),
.Y(n_460)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_85),
.A2(n_104),
.B1(n_363),
.B2(n_372),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_85),
.A2(n_104),
.B1(n_291),
.B2(n_462),
.Y(n_481)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_86),
.B(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_86),
.A2(n_186),
.B1(n_227),
.B2(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_95),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_90),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g412 ( 
.A(n_91),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_92),
.Y(n_418)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_99),
.B2(n_101),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_99),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_100),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_100),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_100),
.Y(n_422)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_104),
.Y(n_186)
);

NOR2x1_ASAP7_75t_L g403 ( 
.A(n_104),
.B(n_404),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_133),
.B1(n_143),
.B2(n_145),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_114),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_114),
.A2(n_133),
.B1(n_143),
.B2(n_190),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g349 ( 
.A1(n_114),
.A2(n_143),
.B1(n_350),
.B2(n_356),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_114),
.A2(n_143),
.B1(n_356),
.B2(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g452 ( 
.A1(n_114),
.A2(n_143),
.B1(n_350),
.B2(n_453),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_114),
.A2(n_143),
.B1(n_299),
.B2(n_483),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g655 ( 
.A1(n_114),
.A2(n_143),
.B1(n_377),
.B2(n_656),
.Y(n_655)
);

AO21x2_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_120),
.B(n_126),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_118),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_120),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_121),
.Y(n_304)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_122),
.Y(n_382)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_122),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_123),
.Y(n_267)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_126),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_126)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_127),
.Y(n_572)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_131),
.Y(n_244)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_137),
.Y(n_662)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_144),
.A2(n_157),
.B1(n_191),
.B2(n_257),
.Y(n_256)
);

AOI22x1_ASAP7_75t_L g297 ( 
.A1(n_144),
.A2(n_157),
.B1(n_257),
.B2(n_298),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_146),
.Y(n_192)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVx8_ASAP7_75t_L g353 ( 
.A(n_148),
.Y(n_353)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_153),
.Y(n_660)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_169),
.Y(n_442)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_175),
.C(n_187),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_171),
.B(n_320),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_175),
.C(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_175),
.Y(n_320)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_177),
.B(n_314),
.Y(n_313)
);

AOI21x1_ASAP7_75t_L g225 ( 
.A1(n_178),
.A2(n_186),
.B(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_187),
.B(n_319),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_189),
.Y(n_315)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

AO21x1_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_323),
.B(n_684),
.Y(n_196)
);

NOR2x1_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_316),
.Y(n_197)
);

NOR2xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_305),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_199),
.B(n_305),
.Y(n_686)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_251),
.C(n_269),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_201),
.A2(n_251),
.B1(n_252),
.B2(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_201),
.Y(n_511)
);

OAI22x1_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_235),
.B2(n_250),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_225),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_204),
.A2(n_307),
.B1(n_309),
.B2(n_692),
.Y(n_306)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_204),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_216),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_209),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_210),
.A2(n_217),
.B1(n_283),
.B2(n_286),
.Y(n_282)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_210),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_210),
.A2(n_286),
.B1(n_426),
.B2(n_429),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_210),
.A2(n_590),
.B1(n_592),
.B2(n_593),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_210),
.A2(n_616),
.B1(n_620),
.B2(n_627),
.Y(n_615)
);

OR2x6_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

BUFx2_ASAP7_75t_R g391 ( 
.A(n_211),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g644 ( 
.A(n_211),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_212),
.Y(n_628)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_212),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_221),
.Y(n_594)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_223),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx6_ASAP7_75t_L g397 ( 
.A(n_224),
.Y(n_397)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_224),
.Y(n_577)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_225),
.Y(n_310)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_230),
.Y(n_414)
);

INVx4_ASAP7_75t_SL g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_233),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_235),
.Y(n_308)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_236),
.Y(n_501)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_237),
.Y(n_280)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_238),
.Y(n_533)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_241),
.Y(n_275)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_SL g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_248),
.Y(n_570)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_256),
.B(n_268),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_256),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_254),
.A2(n_346),
.B1(n_560),
.B2(n_568),
.Y(n_559)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_267),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_269),
.B(n_510),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_288),
.C(n_296),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_270),
.B(n_505),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_279),
.B(n_281),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_271),
.B(n_488),
.Y(n_487)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx4f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_278),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_281),
.B(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_283),
.B(n_404),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g591 ( 
.A(n_285),
.Y(n_591)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_287),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_289),
.B(n_297),
.Y(n_505)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_312),
.C(n_322),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_310),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_317),
.B(n_686),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_SL g688 ( 
.A(n_318),
.B(n_321),
.Y(n_688)
);

AO21x2_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_512),
.B(n_677),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_491),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_471),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_444),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_327),
.B(n_444),
.Y(n_680)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_374),
.C(n_405),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_328),
.B(n_516),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_361),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_349),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_330),
.B(n_349),
.C(n_361),
.Y(n_449)
);

AOI22x1_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_337),
.B2(n_346),
.Y(n_330)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx5_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_343),
.B(n_404),
.Y(n_541)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx5_ASAP7_75t_L g359 ( 
.A(n_353),
.Y(n_359)
);

INVx5_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_353),
.Y(n_409)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g423 ( 
.A(n_368),
.Y(n_423)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_372),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_375),
.B(n_405),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_383),
.C(n_403),
.Y(n_375)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_376),
.Y(n_520)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_383),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_383),
.A2(n_521),
.B(n_522),
.Y(n_526)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_384),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_391),
.B1(n_392),
.B2(n_402),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_385),
.A2(n_402),
.B1(n_425),
.B2(n_428),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx4_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_392),
.A2(n_402),
.B1(n_544),
.B2(n_551),
.Y(n_543)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_397),
.Y(n_546)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_397),
.Y(n_586)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_397),
.Y(n_619)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_401),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_402),
.A2(n_642),
.B1(n_643),
.B2(n_644),
.Y(n_641)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_403),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_403),
.B(n_525),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_SL g560 ( 
.A1(n_404),
.A2(n_561),
.B(n_564),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_404),
.B(n_565),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_424),
.B1(n_438),
.B2(n_443),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_406),
.B(n_443),
.Y(n_470)
);

OAI32xp33_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_410),
.A3(n_413),
.B1(n_415),
.B2(n_423),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g439 ( 
.A1(n_407),
.A2(n_410),
.A3(n_415),
.B1(n_423),
.B2(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_419),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_424),
.Y(n_443)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_SL g426 ( 
.A(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_433),
.Y(n_599)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx4_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx4_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_437),
.Y(n_550)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_450),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_449),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_446),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_447),
.B(n_448),
.Y(n_478)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_449),
.Y(n_474)
);

MAJx2_ASAP7_75t_L g472 ( 
.A(n_450),
.B(n_473),
.C(n_474),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_470),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_460),
.B1(n_468),
.B2(n_469),
.Y(n_451)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_452),
.Y(n_468)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_460),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_468),
.C(n_470),
.Y(n_490)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx8_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

NAND2xp67_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_472),
.B(n_475),
.C(n_680),
.Y(n_679)
);

XOR2x2_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_490),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_477),
.A2(n_485),
.B1(n_486),
.B2(n_489),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_477),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g494 ( 
.A(n_477),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_480),
.C(n_497),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_480),
.A2(n_481),
.B1(n_482),
.B2(n_484),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_482),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_484),
.Y(n_497)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_490),
.C(n_494),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g677 ( 
.A1(n_491),
.A2(n_678),
.B(n_681),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_506),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_495),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_493),
.B(n_495),
.Y(n_682)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_496),
.B(n_499),
.C(n_508),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_504),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_503),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_502),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_504),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_506),
.A2(n_682),
.B(n_683),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_509),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_507),
.B(n_509),
.Y(n_683)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

AOI21x1_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_553),
.B(n_676),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_515),
.B(n_517),
.Y(n_514)
);

NOR2xp67_ASAP7_75t_SL g676 ( 
.A(n_515),
.B(n_517),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_528),
.C(n_534),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_518),
.B(n_671),
.Y(n_670)
);

AOI22x1_ASAP7_75t_L g518 ( 
.A1(n_519),
.A2(n_524),
.B1(n_526),
.B2(n_527),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_521),
.Y(n_519)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_520),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g671 ( 
.A1(n_528),
.A2(n_672),
.B(n_673),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_528),
.B(n_535),
.Y(n_673)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_534),
.Y(n_672)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_542),
.Y(n_535)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_536),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_536),
.B(n_543),
.Y(n_667)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_542),
.Y(n_666)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g592 ( 
.A(n_544),
.Y(n_592)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

BUFx4f_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g553 ( 
.A1(n_554),
.A2(n_669),
.B(n_675),
.Y(n_553)
);

AOI21x1_ASAP7_75t_L g554 ( 
.A1(n_555),
.A2(n_648),
.B(n_668),
.Y(n_554)
);

OAI21x1_ASAP7_75t_SL g555 ( 
.A1(n_556),
.A2(n_612),
.B(n_647),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_557),
.B(n_588),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_557),
.B(n_588),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_558),
.B(n_573),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_558),
.A2(n_559),
.B1(n_573),
.B2(n_574),
.Y(n_645)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_564),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_568),
.Y(n_609)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_570),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_572),
.Y(n_571)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_575),
.A2(n_582),
.B1(n_583),
.B2(n_587),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_576),
.B(n_578),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_589),
.B(n_600),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_589),
.B(n_602),
.C(n_610),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_593),
.Y(n_643)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_601),
.A2(n_602),
.B1(n_610),
.B2(n_611),
.Y(n_600)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_601),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_602),
.Y(n_611)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_603),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

AOI21x1_ASAP7_75t_SL g612 ( 
.A1(n_613),
.A2(n_640),
.B(n_646),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_614),
.A2(n_630),
.B(n_639),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_615),
.B(n_629),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_615),
.B(n_629),
.Y(n_639)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_620),
.Y(n_642)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_622),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_623),
.Y(n_622)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_626),
.Y(n_625)
);

INVx8_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_631),
.B(n_633),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_634),
.B(n_635),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

BUFx2_ASAP7_75t_SL g637 ( 
.A(n_638),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_641),
.B(n_645),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_L g646 ( 
.A(n_641),
.B(n_645),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_649),
.B(n_650),
.Y(n_648)
);

NOR2x1_ASAP7_75t_L g668 ( 
.A(n_649),
.B(n_650),
.Y(n_668)
);

XNOR2x1_ASAP7_75t_L g650 ( 
.A(n_651),
.B(n_664),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g651 ( 
.A1(n_652),
.A2(n_653),
.B1(n_655),
.B2(n_663),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_653),
.B(n_663),
.C(n_664),
.Y(n_674)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_655),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_658),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_662),
.Y(n_661)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_665),
.A2(n_666),
.B(n_667),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_SL g669 ( 
.A(n_670),
.B(n_674),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_670),
.B(n_674),
.Y(n_675)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_679),
.Y(n_678)
);

NAND2xp33_ASAP7_75t_SL g684 ( 
.A(n_685),
.B(n_687),
.Y(n_684)
);

INVxp33_ASAP7_75t_L g687 ( 
.A(n_688),
.Y(n_687)
);


endmodule