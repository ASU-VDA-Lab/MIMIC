module fake_jpeg_26325_n_130 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx8_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_3),
.B(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_35),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_26),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_24),
.Y(n_42)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_42),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_19),
.B1(n_13),
.B2(n_16),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_24),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_46),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_26),
.B(n_20),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_27),
.B(n_16),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_34),
.A2(n_19),
.B1(n_13),
.B2(n_20),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_35),
.B1(n_28),
.B2(n_33),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_45),
.B1(n_28),
.B2(n_33),
.Y(n_67)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_17),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_17),
.B(n_22),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_42),
.C(n_40),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_13),
.C(n_10),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_43),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_45),
.B1(n_35),
.B2(n_38),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_54),
.B1(n_49),
.B2(n_51),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_70),
.B(n_12),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_48),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_73),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_67),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_71),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_59),
.A2(n_31),
.B(n_29),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_61),
.C(n_59),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_76),
.C(n_73),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_88),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_21),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_63),
.A2(n_56),
.B1(n_45),
.B2(n_41),
.Y(n_82)
);

OAI21x1_ASAP7_75t_L g90 ( 
.A1(n_82),
.A2(n_87),
.B(n_56),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_47),
.B1(n_41),
.B2(n_69),
.Y(n_96)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_92),
.B(n_93),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_91),
.B(n_94),
.Y(n_106)
);

BUFx12f_ASAP7_75t_SL g92 ( 
.A(n_82),
.Y(n_92)
);

AOI322xp5_ASAP7_75t_SL g93 ( 
.A1(n_78),
.A2(n_65),
.A3(n_57),
.B1(n_76),
.B2(n_12),
.C1(n_10),
.C2(n_8),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_64),
.C(n_43),
.Y(n_94)
);

AOI322xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_9),
.A3(n_8),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_2),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_98),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_96),
.A2(n_97),
.B1(n_43),
.B2(n_69),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_85),
.A2(n_47),
.B1(n_41),
.B2(n_69),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_43),
.C(n_29),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_99),
.B(n_29),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_85),
.B(n_84),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

A2O1A1O1Ixp25_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_79),
.B(n_80),
.C(n_83),
.D(n_31),
.Y(n_101)
);

XOR2x1_ASAP7_75t_SL g114 ( 
.A(n_101),
.B(n_1),
.Y(n_114)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_105),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_97),
.B1(n_29),
.B2(n_14),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g108 ( 
.A1(n_94),
.A2(n_21),
.B1(n_25),
.B2(n_23),
.C(n_31),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_99),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_112),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_113),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_21),
.B1(n_23),
.B2(n_25),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_100),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_114),
.B(n_104),
.Y(n_117)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_119),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_117),
.B(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI321xp33_ASAP7_75t_L g126 ( 
.A1(n_122),
.A2(n_124),
.A3(n_117),
.B1(n_115),
.B2(n_106),
.C(n_6),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_1),
.Y(n_123)
);

BUFx24_ASAP7_75t_SL g125 ( 
.A(n_123),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_120),
.A2(n_115),
.B(n_103),
.C(n_106),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_126),
.B(n_127),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_1),
.B1(n_5),
.B2(n_124),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_128),
.Y(n_130)
);


endmodule