module fake_jpeg_3652_n_246 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_246);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_246;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g46 ( 
.A1(n_17),
.A2(n_0),
.B(n_2),
.Y(n_46)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_21),
.B(n_36),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx9p33_ASAP7_75t_R g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_54),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_23),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_25),
.B(n_22),
.C(n_35),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_32),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_74),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_51),
.A2(n_27),
.B1(n_36),
.B2(n_21),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_59),
.A2(n_61),
.B1(n_64),
.B2(n_77),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_27),
.B1(n_21),
.B2(n_19),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_44),
.A2(n_27),
.B1(n_19),
.B2(n_17),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_54),
.B1(n_53),
.B2(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_67),
.B1(n_84),
.B2(n_20),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_48),
.A2(n_28),
.B1(n_31),
.B2(n_33),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_68),
.B(n_73),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_23),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_50),
.B(n_29),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_76),
.B(n_0),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_40),
.A2(n_17),
.B1(n_36),
.B2(n_19),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_31),
.B1(n_33),
.B2(n_20),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_86),
.B1(n_20),
.B2(n_35),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_29),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_14),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_31),
.B1(n_33),
.B2(n_25),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_47),
.A2(n_31),
.B1(n_33),
.B2(n_20),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_87),
.A2(n_62),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_90),
.Y(n_119)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_103),
.B1(n_72),
.B2(n_62),
.Y(n_125)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_15),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_94),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_78),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_98),
.Y(n_131)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_22),
.B1(n_35),
.B2(n_37),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_99),
.A2(n_107),
.B1(n_111),
.B2(n_8),
.Y(n_141)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_78),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_106),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_35),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_102),
.A2(n_8),
.B(n_10),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_35),
.B1(n_22),
.B2(n_34),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_105),
.B(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_35),
.B1(n_37),
.B2(n_34),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_37),
.B(n_34),
.C(n_5),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_71),
.B(n_62),
.C(n_9),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_115),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_85),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_72),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_117),
.B1(n_83),
.B2(n_69),
.Y(n_134)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_79),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_75),
.B1(n_57),
.B2(n_69),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_69),
.B1(n_63),
.B2(n_75),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_121),
.A2(n_98),
.B1(n_101),
.B2(n_95),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_134),
.B1(n_102),
.B2(n_115),
.Y(n_155)
);

NOR3xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_132),
.C(n_110),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_87),
.A2(n_108),
.B(n_117),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_113),
.B(n_116),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_109),
.A2(n_79),
.B1(n_63),
.B2(n_83),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_103),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_83),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_139),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_104),
.B(n_6),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_110),
.B(n_10),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_143),
.B(n_113),
.Y(n_160)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_145),
.B(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_93),
.C(n_90),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_149),
.C(n_130),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_88),
.C(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_105),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_91),
.Y(n_152)
);

AO21x2_ASAP7_75t_L g176 ( 
.A1(n_153),
.A2(n_166),
.B(n_125),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_155),
.A2(n_131),
.B1(n_134),
.B2(n_121),
.Y(n_179)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_131),
.A2(n_114),
.A3(n_112),
.B1(n_89),
.B2(n_106),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_159),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_160),
.B(n_162),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_161),
.A2(n_167),
.B(n_133),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_100),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_164),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g164 ( 
.A(n_123),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_100),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_131),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_126),
.A2(n_96),
.B(n_12),
.C(n_13),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_126),
.A2(n_141),
.B(n_124),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_147),
.B(n_139),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_175),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_176),
.A2(n_179),
.B1(n_145),
.B2(n_137),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_128),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_182),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_150),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_160),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_177),
.C(n_182),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_128),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_140),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_183),
.B(n_156),
.Y(n_194)
);

OAI32xp33_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_131),
.A3(n_124),
.B1(n_119),
.B2(n_118),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_184),
.A2(n_166),
.B(n_145),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_185),
.A2(n_142),
.B(n_119),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_137),
.B1(n_136),
.B2(n_118),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

AOI221xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_148),
.B1(n_154),
.B2(n_147),
.C(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_187),
.A2(n_196),
.B1(n_135),
.B2(n_136),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_176),
.A2(n_165),
.B1(n_145),
.B2(n_161),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_198),
.B1(n_176),
.B2(n_168),
.Y(n_206)
);

INVxp33_ASAP7_75t_SL g203 ( 
.A(n_190),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_195),
.C(n_201),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_188),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_144),
.C(n_158),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_166),
.B(n_157),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_197),
.A2(n_202),
.B(n_168),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_151),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_209),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_206),
.B(n_214),
.Y(n_222)
);

AOI322xp5_ASAP7_75t_L g207 ( 
.A1(n_197),
.A2(n_172),
.A3(n_168),
.B1(n_176),
.B2(n_184),
.C1(n_173),
.C2(n_180),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_208),
.B(n_198),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_172),
.B(n_176),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_170),
.B(n_153),
.Y(n_209)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_142),
.C(n_135),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_210),
.B(n_202),
.Y(n_216)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_188),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_193),
.C(n_195),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_216),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_218),
.B(n_220),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_194),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_203),
.B(n_200),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_211),
.Y(n_228)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_222),
.A2(n_212),
.B1(n_208),
.B2(n_211),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_224),
.A2(n_229),
.B1(n_210),
.B2(n_206),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_228),
.Y(n_235)
);

INVx4_ASAP7_75t_SL g229 ( 
.A(n_217),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_222),
.A2(n_191),
.B1(n_199),
.B2(n_204),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_209),
.Y(n_233)
);

OAI21x1_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_219),
.B(n_220),
.Y(n_231)
);

AOI31xp33_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_234),
.A3(n_225),
.B(n_218),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_233),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_226),
.A2(n_213),
.B(n_201),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_235),
.B(n_226),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_238),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_229),
.Y(n_238)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_225),
.B(n_224),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g243 ( 
.A1(n_241),
.A2(n_237),
.B(n_12),
.C(n_13),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_237),
.B(n_135),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_242),
.A2(n_243),
.B(n_96),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_244),
.A2(n_10),
.B(n_12),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_13),
.Y(n_246)
);


endmodule