module fake_jpeg_18774_n_346 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_346);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_346;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx6_ASAP7_75t_SL g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_42),
.B(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_16),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_54),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_26),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_29),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_23),
.B1(n_37),
.B2(n_47),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_41),
.B1(n_23),
.B2(n_44),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_75),
.B1(n_86),
.B2(n_88),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_48),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_72),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_48),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_44),
.B1(n_43),
.B2(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_44),
.B1(n_45),
.B2(n_42),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_83),
.B1(n_84),
.B2(n_94),
.Y(n_111)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_96),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_45),
.B1(n_42),
.B2(n_23),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_37),
.B1(n_40),
.B2(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_47),
.B1(n_37),
.B2(n_46),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_19),
.B1(n_28),
.B2(n_34),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_87),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_59),
.B1(n_50),
.B2(n_55),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_55),
.B(n_49),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_100),
.C(n_25),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_59),
.A2(n_47),
.B1(n_46),
.B2(n_40),
.Y(n_94)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_21),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_21),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_66),
.B(n_39),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_54),
.A2(n_39),
.B1(n_38),
.B2(n_28),
.Y(n_97)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_99),
.B1(n_38),
.B2(n_36),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_19),
.B(n_28),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_25),
.C(n_34),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_39),
.B1(n_38),
.B2(n_19),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_39),
.C(n_38),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_61),
.A2(n_26),
.B1(n_27),
.B2(n_35),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_101),
.A2(n_27),
.B1(n_29),
.B2(n_35),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_76),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_104),
.B(n_114),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_108),
.B(n_75),
.Y(n_153)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_115),
.B(n_117),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_87),
.Y(n_116)
);

INVx5_ASAP7_75t_SL g159 ( 
.A(n_116),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_24),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_24),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_121),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_91),
.B(n_72),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_90),
.Y(n_122)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_125),
.B1(n_129),
.B2(n_132),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_21),
.Y(n_160)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_79),
.A2(n_31),
.B1(n_34),
.B2(n_17),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_74),
.A2(n_31),
.B1(n_17),
.B2(n_24),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_133),
.A2(n_95),
.B(n_86),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_73),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_138),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_106),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_137),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_100),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

BUFx24_ASAP7_75t_SL g141 ( 
.A(n_127),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_141),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_77),
.Y(n_142)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_142),
.Y(n_163)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_124),
.A2(n_128),
.B1(n_130),
.B2(n_133),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_144),
.A2(n_152),
.B1(n_154),
.B2(n_123),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_93),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_156),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_151),
.B(n_20),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_128),
.B1(n_126),
.B2(n_110),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_150),
.A2(n_160),
.B1(n_161),
.B2(n_131),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_107),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_126),
.A2(n_84),
.B1(n_83),
.B2(n_82),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_30),
.C(n_33),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_110),
.A2(n_85),
.B1(n_81),
.B2(n_94),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_111),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_81),
.Y(n_157)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_118),
.A2(n_67),
.B1(n_74),
.B2(n_80),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_162),
.A2(n_169),
.B1(n_143),
.B2(n_145),
.Y(n_202)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_131),
.B1(n_102),
.B2(n_120),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_3),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_18),
.B(n_114),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_185),
.B(n_187),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_150),
.A2(n_109),
.B1(n_122),
.B2(n_105),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_146),
.B(n_138),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_182),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_175),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_159),
.A2(n_160),
.B1(n_144),
.B2(n_147),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_210)
);

FAx1_ASAP7_75t_SL g175 ( 
.A(n_153),
.B(n_105),
.CI(n_109),
.CON(n_175),
.SN(n_175)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_147),
.A2(n_120),
.B1(n_68),
.B2(n_69),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_112),
.B1(n_92),
.B2(n_30),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_189),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_112),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_159),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_183),
.A2(n_188),
.B1(n_190),
.B2(n_2),
.Y(n_214)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_155),
.B(n_149),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_136),
.C(n_151),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_191),
.B(n_1),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_30),
.B1(n_33),
.B2(n_36),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_161),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_136),
.A2(n_36),
.B1(n_33),
.B2(n_20),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_192),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_193),
.B(n_203),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_197),
.B(n_205),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_185),
.A2(n_158),
.B1(n_137),
.B2(n_135),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_198),
.A2(n_211),
.B(n_191),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_200),
.A2(n_168),
.B1(n_186),
.B2(n_175),
.Y(n_232)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_178),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_202),
.A2(n_207),
.B1(n_209),
.B2(n_190),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_134),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_149),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_162),
.A2(n_139),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_163),
.A2(n_15),
.B(n_14),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_5),
.B(n_6),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_169),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_170),
.B(n_13),
.C(n_2),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_213),
.A2(n_216),
.B(n_218),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_217),
.B1(n_218),
.B2(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_215),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_172),
.A2(n_3),
.B(n_4),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_166),
.A2(n_3),
.B(n_4),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_3),
.C(n_4),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_184),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_220),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_181),
.Y(n_221)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_221),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_222),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_223),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_5),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_223),
.A2(n_217),
.B1(n_189),
.B2(n_167),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_227),
.A2(n_202),
.B1(n_207),
.B2(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_221),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_230),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_231),
.B(n_200),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_232),
.A2(n_231),
.B(n_233),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_193),
.Y(n_237)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_237),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_201),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_239),
.A2(n_242),
.B(n_244),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_210),
.A2(n_167),
.B1(n_177),
.B2(n_188),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_250),
.B1(n_214),
.B2(n_220),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_206),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_199),
.Y(n_245)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_245),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_199),
.Y(n_247)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_198),
.A2(n_180),
.B(n_192),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_248),
.A2(n_213),
.B(n_194),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_251),
.A2(n_235),
.B1(n_247),
.B2(n_245),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_194),
.B1(n_195),
.B2(n_208),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_238),
.B(n_173),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_254),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_255),
.A2(n_260),
.B1(n_250),
.B2(n_236),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_243),
.B(n_248),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_212),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_211),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_215),
.B1(n_196),
.B2(n_204),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_262),
.Y(n_286)
);

AOI221xp5_ASAP7_75t_L g264 ( 
.A1(n_233),
.A2(n_222),
.B1(n_211),
.B2(n_219),
.C(n_203),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_264),
.B(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_270),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_212),
.C(n_232),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_234),
.C(n_239),
.Y(n_273)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_226),
.Y(n_269)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_226),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_282),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_275),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_274),
.A2(n_271),
.B(n_265),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_276),
.A2(n_287),
.B1(n_288),
.B2(n_260),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_262),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_258),
.A2(n_235),
.B1(n_228),
.B2(n_242),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_258),
.A2(n_228),
.B1(n_249),
.B2(n_230),
.Y(n_283)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_283),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_259),
.Y(n_285)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_255),
.A2(n_249),
.B1(n_240),
.B2(n_244),
.Y(n_287)
);

AOI22x1_ASAP7_75t_L g288 ( 
.A1(n_256),
.A2(n_165),
.B1(n_209),
.B2(n_216),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_289),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_240),
.C(n_183),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_268),
.C(n_267),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_276),
.Y(n_291)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_291),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_294),
.B(n_286),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_295),
.B(n_301),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_271),
.C(n_263),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_274),
.A2(n_265),
.B1(n_266),
.B2(n_270),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_282),
.B1(n_283),
.B2(n_272),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_273),
.Y(n_302)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_302),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_263),
.C(n_261),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_286),
.C(n_275),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_288),
.B(n_287),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_307),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_299),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_310),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_317),
.C(n_288),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_284),
.B1(n_280),
.B2(n_269),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_316),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_292),
.B(n_252),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_279),
.C(n_252),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_323),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_297),
.B1(n_305),
.B2(n_294),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_320),
.A2(n_321),
.B1(n_315),
.B2(n_313),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_307),
.A2(n_305),
.B1(n_300),
.B2(n_301),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_303),
.B(n_293),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_325),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_165),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_7),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_322),
.B(n_317),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_327),
.B(n_329),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_318),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_330),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_326),
.B(n_173),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_333),
.A2(n_319),
.B(n_320),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_337),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_331),
.B(n_7),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g338 ( 
.A1(n_334),
.A2(n_332),
.B(n_8),
.Y(n_338)
);

OAI21xp33_ASAP7_75t_L g340 ( 
.A1(n_338),
.A2(n_7),
.B(n_8),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_339),
.C(n_9),
.Y(n_341)
);

NOR2xp67_ASAP7_75t_SL g342 ( 
.A(n_341),
.B(n_335),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_342),
.A2(n_7),
.B(n_9),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_9),
.C(n_10),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_10),
.Y(n_346)
);


endmodule