module fake_jpeg_9783_n_229 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_229);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_0),
.B(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_45),
.B(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_1),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx12_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_53),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_26),
.B1(n_17),
.B2(n_32),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_32),
.B1(n_22),
.B2(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_L g54 ( 
.A1(n_40),
.A2(n_23),
.B(n_29),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_21),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_61),
.Y(n_88)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_67),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_45),
.A2(n_26),
.B1(n_28),
.B2(n_17),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_60),
.A2(n_70),
.B1(n_22),
.B2(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_28),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_65),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_37),
.Y(n_65)
);

CKINVDCx12_ASAP7_75t_R g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_26),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_39),
.A2(n_1),
.B(n_2),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_18),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_19),
.C(n_34),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_77),
.Y(n_123)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_17),
.B1(n_18),
.B2(n_41),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_96),
.B1(n_71),
.B2(n_19),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_32),
.B1(n_30),
.B2(n_29),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_81),
.A2(n_103),
.B1(n_20),
.B2(n_31),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_84),
.B(n_85),
.Y(n_124)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_89),
.B(n_99),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_95),
.Y(n_110)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_55),
.B(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_27),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_73),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_65),
.A2(n_30),
.B1(n_21),
.B2(n_20),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_105),
.B(n_93),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_108),
.B1(n_122),
.B2(n_94),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_53),
.B(n_50),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_126),
.C(n_127),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_103),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_72),
.B1(n_62),
.B2(n_27),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_2),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_58),
.B(n_3),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_128),
.B(n_134),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_85),
.C(n_92),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_14),
.C(n_10),
.Y(n_165)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_89),
.Y(n_130)
);

AOI221xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_132),
.B1(n_126),
.B2(n_10),
.C(n_12),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_137),
.Y(n_169)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_91),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_139),
.Y(n_155)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_150),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_75),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_138),
.C(n_143),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_78),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_86),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_141),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_62),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_142),
.B(n_148),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_72),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_98),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g145 ( 
.A(n_120),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_145),
.A2(n_106),
.B1(n_121),
.B2(n_110),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_18),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_120),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_109),
.B(n_80),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_143),
.A2(n_113),
.B1(n_116),
.B2(n_109),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_151),
.A2(n_133),
.B1(n_146),
.B2(n_132),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_112),
.B(n_117),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_152),
.A2(n_154),
.B(n_157),
.Y(n_186)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_153),
.B(n_158),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_138),
.A2(n_112),
.B1(n_116),
.B2(n_104),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_126),
.B(n_83),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

OA21x2_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_165),
.B(n_130),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_166),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_118),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_170),
.B(n_2),
.C(n_3),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_154),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_146),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_183),
.C(n_185),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_173),
.Y(n_187)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_155),
.A2(n_160),
.A3(n_153),
.B1(n_151),
.B2(n_164),
.Y(n_174)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_174),
.Y(n_193)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_169),
.C(n_14),
.Y(n_196)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_166),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_178),
.B(n_179),
.Y(n_195)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_180),
.B(n_184),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_145),
.B(n_149),
.C(n_106),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_181),
.A2(n_177),
.B1(n_178),
.B2(n_175),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_118),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_159),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_192),
.Y(n_202)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_179),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_190),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_152),
.C(n_157),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_186),
.Y(n_204)
);

NAND3xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_5),
.C(n_6),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_164),
.B1(n_158),
.B2(n_156),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_181),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_198),
.B(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_199),
.B(n_206),
.Y(n_209)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_188),
.Y(n_203)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_203),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_204),
.B(n_189),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_205),
.B(n_5),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_192),
.A2(n_182),
.B(n_185),
.Y(n_206)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_207),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_202),
.C(n_191),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_210),
.B(n_214),
.Y(n_215)
);

AOI321xp33_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_193),
.A3(n_174),
.B1(n_194),
.B2(n_177),
.C(n_191),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_213),
.A2(n_195),
.B(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_187),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_216),
.A2(n_217),
.B(n_208),
.Y(n_220)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_190),
.A3(n_202),
.B1(n_175),
.B2(n_156),
.C1(n_205),
.C2(n_168),
.Y(n_218)
);

AOI211xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_9),
.B(n_7),
.C(n_8),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_5),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_6),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_220),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_211),
.B(n_213),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_221),
.B(n_222),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_224),
.B(n_225),
.C(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_226),
.B(n_227),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_7),
.C(n_8),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_8),
.Y(n_229)
);


endmodule