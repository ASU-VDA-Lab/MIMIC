module real_jpeg_30739_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_487;
wire n_493;
wire n_93;
wire n_242;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_0),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_0),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g366 ( 
.A(n_0),
.Y(n_366)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_0),
.Y(n_457)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_1),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_1),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_1),
.B(n_209),
.Y(n_368)
);

OAI32xp33_ASAP7_75t_L g470 ( 
.A1(n_1),
.A2(n_471),
.A3(n_476),
.B1(n_478),
.B2(n_483),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g499 ( 
.A1(n_1),
.A2(n_271),
.B1(n_500),
.B2(n_503),
.Y(n_499)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_1),
.A2(n_131),
.B(n_536),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_2),
.A2(n_203),
.B1(n_207),
.B2(n_208),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_2),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_2),
.A2(n_207),
.B1(n_288),
.B2(n_292),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_2),
.A2(n_207),
.B1(n_356),
.B2(n_358),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_2),
.A2(n_207),
.B1(n_461),
.B2(n_465),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_163),
.B1(n_166),
.B2(n_167),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_3),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_166),
.B1(n_224),
.B2(n_226),
.Y(n_223)
);

AOI22x1_ASAP7_75t_L g280 ( 
.A1(n_3),
.A2(n_166),
.B1(n_281),
.B2(n_286),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_3),
.A2(n_166),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_4),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_4),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_5),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_25)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_5),
.A2(n_31),
.B1(n_125),
.B2(n_128),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_31),
.B1(n_163),
.B2(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_6),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_6),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_7),
.A2(n_56),
.B1(n_61),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_173),
.B1(n_174),
.B2(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_8),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_8),
.A2(n_173),
.B1(n_303),
.B2(n_306),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g493 ( 
.A1(n_8),
.A2(n_32),
.B1(n_173),
.B2(n_494),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g527 ( 
.A1(n_8),
.A2(n_173),
.B1(n_528),
.B2(n_532),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_9),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_9),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_10),
.A2(n_296),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_10),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_10),
.A2(n_298),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g486 ( 
.A1(n_10),
.A2(n_298),
.B1(n_487),
.B2(n_490),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_L g580 ( 
.A1(n_10),
.A2(n_298),
.B1(n_361),
.B2(n_581),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_12),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_12),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_12),
.A2(n_76),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_12),
.A2(n_76),
.B1(n_240),
.B2(n_243),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_12),
.A2(n_76),
.B1(n_312),
.B2(n_317),
.Y(n_311)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_13),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_13),
.Y(n_192)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_14),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_15),
.A2(n_105),
.B1(n_109),
.B2(n_110),
.Y(n_104)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_15),
.A2(n_109),
.B1(n_145),
.B2(n_149),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_15),
.A2(n_109),
.B1(n_325),
.B2(n_329),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_16),
.Y(n_75)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_16),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_259),
.Y(n_17)
);

NAND2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_258),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2x1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_230),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_21),
.B(n_230),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_119),
.C(n_210),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_22),
.B(n_211),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_69),
.B(n_118),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_23),
.B(n_69),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_35),
.B1(n_57),
.B2(n_68),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_25),
.A2(n_36),
.B1(n_143),
.B2(n_144),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_30),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g39 ( 
.A(n_34),
.Y(n_39)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_35),
.A2(n_57),
.B(n_68),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_35),
.A2(n_68),
.B1(n_279),
.B2(n_287),
.Y(n_278)
);

AO22x2_ASAP7_75t_SL g523 ( 
.A1(n_35),
.A2(n_68),
.B1(n_287),
.B2(n_524),
.Y(n_523)
);

OAI211xp5_ASAP7_75t_L g565 ( 
.A1(n_35),
.A2(n_566),
.B(n_567),
.C(n_568),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_36),
.A2(n_143),
.B1(n_144),
.B2(n_152),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_36),
.A2(n_143),
.B1(n_152),
.B2(n_280),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_36),
.A2(n_143),
.B1(n_486),
.B2(n_493),
.Y(n_485)
);

OAI21xp33_ASAP7_75t_SL g508 ( 
.A1(n_36),
.A2(n_493),
.B(n_509),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_48),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_37)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_38),
.Y(n_286)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_39),
.Y(n_293)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22x1_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_49),
.B1(n_52),
.B2(n_55),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_44),
.Y(n_563)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_47),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_47),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_51),
.Y(n_584)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_68),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_68),
.B(n_287),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_81),
.B1(n_104),
.B2(n_115),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_70),
.A2(n_81),
.B1(n_117),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g168 ( 
.A(n_75),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_75),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_75),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_79),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_80),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_80),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_81),
.A2(n_104),
.B1(n_115),
.B2(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_81),
.A2(n_115),
.B1(n_295),
.B2(n_301),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g354 ( 
.A(n_81),
.B(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_81),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_91),
.Y(n_81)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_87),
.Y(n_559)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_95),
.B(n_98),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_97),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_101),
.Y(n_108)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_101),
.Y(n_307)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_102),
.Y(n_357)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_102),
.Y(n_505)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_114),
.Y(n_300)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_114),
.Y(n_358)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI21xp33_ASAP7_75t_SL g352 ( 
.A1(n_116),
.A2(n_353),
.B(n_354),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_116),
.A2(n_384),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

NOR2x1_ASAP7_75t_L g525 ( 
.A(n_116),
.B(n_271),
.Y(n_525)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_117),
.B(n_355),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_118),
.Y(n_235)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2x2_ASAP7_75t_L g417 ( 
.A(n_120),
.B(n_418),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_160),
.C(n_169),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_122),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_142),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_123),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.Y(n_411)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_123),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_131),
.B1(n_138),
.B2(n_140),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_124),
.A2(n_131),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g330 ( 
.A(n_130),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_131),
.A2(n_138),
.B(n_214),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_131),
.A2(n_311),
.B1(n_360),
.B2(n_365),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_131),
.A2(n_527),
.B(n_536),
.Y(n_526)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_132),
.A2(n_310),
.B1(n_321),
.B2(n_324),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_132),
.B(n_460),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_132),
.A2(n_596),
.B1(n_597),
.B2(n_598),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_136),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_137),
.Y(n_538)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_142),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_143),
.B(n_271),
.Y(n_578)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_149),
.Y(n_567)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_151),
.Y(n_291)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_151),
.Y(n_497)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_159),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_161),
.B(n_170),
.Y(n_424)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_162),
.Y(n_408)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_168),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_201),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_182),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g409 ( 
.A1(n_172),
.A2(n_182),
.B1(n_209),
.B2(n_389),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_175),
.Y(n_208)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_177),
.Y(n_270)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx4f_ASAP7_75t_SL g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g242 ( 
.A(n_180),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_181),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_181),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_202),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_182),
.Y(n_238)
);

NAND2xp33_ASAP7_75t_SL g268 ( 
.A(n_182),
.B(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_183),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B1(n_189),
.B2(n_190),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_185),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_192),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_198),
.Y(n_391)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_201),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.Y(n_201)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_209),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_209),
.B(n_389),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g232 ( 
.A(n_212),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_213),
.A2(n_217),
.B1(n_219),
.B2(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

BUFx4f_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_217),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B(n_228),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_219),
.A2(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_229),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_220),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_221),
.B(n_388),
.Y(n_387)
);

AOI22x1_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_238),
.B1(n_239),
.B2(n_246),
.Y(n_237)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_224),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_226),
.Y(n_390)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_248),
.Y(n_236)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_256),
.B2(n_257),
.Y(n_248)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2x1_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_441),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_415),
.B(n_436),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_397),
.C(n_398),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_369),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_265),
.B(n_370),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_308),
.C(n_350),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_266),
.B(n_607),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_277),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_267),
.B(n_278),
.C(n_294),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B(n_272),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_271),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_271),
.B(n_555),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_271),
.B(n_554),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_271),
.B(n_593),
.Y(n_592)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_273),
.A2(n_332),
.B1(n_337),
.B2(n_343),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx6_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_294),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g489 ( 
.A(n_285),
.Y(n_489)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_295),
.Y(n_353)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx4f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_300),
.Y(n_479)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_302),
.A2(n_384),
.B(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g502 ( 
.A(n_305),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g607 ( 
.A1(n_308),
.A2(n_350),
.B1(n_351),
.B2(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_308),
.Y(n_608)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_331),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g393 ( 
.A(n_309),
.B(n_331),
.Y(n_393)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_316),
.Y(n_464)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_319),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx6_ASAP7_75t_L g328 ( 
.A(n_320),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_320),
.Y(n_468)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_320),
.Y(n_535)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_324),
.Y(n_377)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_328),
.Y(n_364)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx2_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp33_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_359),
.C(n_367),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_352),
.B(n_514),
.Y(n_513)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_355),
.Y(n_407)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_359),
.A2(n_367),
.B1(n_368),
.B2(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_359),
.Y(n_515)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_360),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx4_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

INVx8_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_380),
.B1(n_395),
.B2(n_396),
.Y(n_370)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_371),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B1(n_378),
.B2(n_379),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_378),
.C(n_396),
.Y(n_397)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_375),
.Y(n_404)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_376),
.Y(n_597)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_381),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_380)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_381),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_386),
.B2(n_387),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_386),
.C(n_392),
.Y(n_400)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_384),
.A2(n_385),
.B(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_397),
.Y(n_444)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_399),
.A2(n_444),
.B(n_445),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_411),
.C(n_432),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_410),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_402),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_405),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_404),
.B(n_409),
.C(n_427),
.Y(n_426)
);

XNOR2x1_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_406),
.Y(n_427)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_416),
.B(n_443),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_419),
.B(n_430),
.Y(n_416)
);

NOR2x1_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_419),
.Y(n_440)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_420),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_425),
.C(n_428),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_422),
.A2(n_423),
.B1(n_428),
.B2(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_434),
.Y(n_433)
);

INVxp33_ASAP7_75t_SL g435 ( 
.A(n_428),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_433),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_438),
.B(n_440),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_446),
.Y(n_441)
);

OAI21x1_ASAP7_75t_SL g446 ( 
.A1(n_447),
.A2(n_602),
.B(n_609),
.Y(n_446)
);

AOI21x1_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_516),
.B(n_601),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_506),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_L g601 ( 
.A(n_449),
.B(n_506),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_485),
.C(n_498),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_451),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_451),
.B(n_520),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_469),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_452),
.B(n_470),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_459),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_458),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_457),
.Y(n_588)
);

OAI21xp33_ASAP7_75t_L g579 ( 
.A1(n_459),
.A2(n_580),
.B(n_585),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g536 ( 
.A(n_460),
.B(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx3_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_476),
.Y(n_484)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_498),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_486),
.Y(n_524)
);

BUFx4f_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx3_ASAP7_75t_SL g504 ( 
.A(n_505),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_513),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_508),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.Y(n_507)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_508),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_509),
.B(n_565),
.Y(n_564)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_510),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_510),
.B(n_511),
.C(n_605),
.Y(n_604)
);

INVxp67_ASAP7_75t_L g605 ( 
.A(n_513),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_539),
.B(n_571),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_518),
.B(n_572),
.C(n_575),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_521),
.Y(n_518)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_519),
.Y(n_541)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_521),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.C(n_526),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

XNOR2x1_ASAP7_75t_L g570 ( 
.A(n_523),
.B(n_525),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g569 ( 
.A(n_526),
.B(n_570),
.Y(n_569)
);

INVxp33_ASAP7_75t_SL g598 ( 
.A(n_527),
.Y(n_598)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

BUFx2_ASAP7_75t_SL g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_532),
.B(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_532),
.Y(n_556)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_540),
.A2(n_541),
.B1(n_542),
.B2(n_569),
.Y(n_539)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_542),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_564),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g600 ( 
.A(n_543),
.B(n_564),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_544),
.A2(n_552),
.B1(n_556),
.B2(n_557),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx6_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

CKINVDCx14_ASAP7_75t_R g552 ( 
.A(n_553),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVxp67_ASAP7_75t_SL g566 ( 
.A(n_554),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_558),
.B(n_560),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_569),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_574),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_576),
.B(n_595),
.C(n_599),
.Y(n_575)
);

OA21x2_ASAP7_75t_SL g576 ( 
.A1(n_577),
.A2(n_589),
.B(n_594),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_578),
.B(n_579),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_578),
.B(n_579),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g596 ( 
.A(n_580),
.Y(n_596)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_582),
.B(n_592),
.Y(n_591)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_586),
.Y(n_585)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_586),
.Y(n_593)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVx2_ASAP7_75t_SL g587 ( 
.A(n_588),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_590),
.B(n_591),
.Y(n_589)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_600),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_606),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_604),
.B(n_610),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_606),
.Y(n_610)
);


endmodule