module real_jpeg_18745_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_14;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_0),
.A2(n_305),
.B1(n_309),
.B2(n_310),
.Y(n_304)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_0),
.Y(n_311)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_2),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_2),
.Y(n_75)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_51),
.B1(n_120),
.B2(n_123),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_3),
.A2(n_51),
.B1(n_141),
.B2(n_144),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_3),
.A2(n_51),
.B1(n_193),
.B2(n_195),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_4),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_4),
.A2(n_27),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_4),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_4),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_4),
.A2(n_27),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_125),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_4),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_4),
.B(n_228),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_5),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_5),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_6),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_6),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_6),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_7),
.A2(n_320),
.B1(n_325),
.B2(n_326),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_7),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_9),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_10),
.Y(n_153)
);

BUFx4f_ASAP7_75t_L g324 ( 
.A(n_10),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_345),
.Y(n_12)
);

AOI21xp5_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_289),
.B(n_341),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_219),
.B(n_288),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_182),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_17),
.B(n_182),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_18),
.B(n_127),
.C(n_160),
.Y(n_337)
);

XOR2x1_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_55),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_20),
.B(n_352),
.C(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_21),
.A2(n_22),
.B1(n_300),
.B2(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_21),
.B(n_57),
.C(n_82),
.Y(n_335)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_31),
.B1(n_41),
.B2(n_49),
.Y(n_22)
);

OA22x2_ASAP7_75t_L g294 ( 
.A1(n_23),
.A2(n_31),
.B1(n_41),
.B2(n_49),
.Y(n_294)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_25),
.B(n_39),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_27),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_27),
.B(n_54),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_27),
.B(n_251),
.Y(n_250)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21x1_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_38),
.B(n_41),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_32),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_41),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_42),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_42),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_52),
.B2(n_54),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_82),
.B2(n_83),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_76),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_58),
.A2(n_67),
.B1(n_76),
.B2(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_58),
.Y(n_227)
);

NAND2x1p5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_67),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_65),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_62),
.Y(n_212)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_66),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_67),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_67),
.A2(n_357),
.B(n_367),
.Y(n_356)
);

OA22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_70),
.Y(n_265)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_74),
.Y(n_247)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_76),
.Y(n_226)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_82),
.A2(n_83),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_82),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_82),
.A2(n_83),
.B1(n_294),
.B2(n_331),
.Y(n_373)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_107),
.B1(n_119),
.B2(n_125),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_84),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_84),
.A2(n_107),
.B(n_125),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_100),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_91),
.B1(n_95),
.B2(n_99),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_90),
.Y(n_106)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_96),
.Y(n_205)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_100),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

OA22x2_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_105),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_102),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g241 ( 
.A(n_102),
.Y(n_241)
);

INVx4_ASAP7_75t_L g365 ( 
.A(n_102),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_113),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

OAI32xp33_ASAP7_75t_L g199 ( 
.A1(n_113),
.A2(n_200),
.A3(n_202),
.B1(n_203),
.B2(n_206),
.Y(n_199)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_160),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_132),
.C(n_134),
.Y(n_127)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_128),
.A2(n_190),
.B1(n_294),
.B2(n_331),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_132),
.A2(n_134),
.B1(n_187),
.B2(n_188),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_SL g255 ( 
.A(n_134),
.B(n_256),
.Y(n_255)
);

OA21x2_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_139),
.B(n_147),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_148),
.B1(n_154),
.B2(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_143),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_143),
.Y(n_326)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_147),
.A2(n_304),
.B(n_312),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_148),
.B(n_216),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_148),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_150),
.Y(n_313)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_152),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g214 ( 
.A(n_154),
.Y(n_214)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_176),
.B2(n_177),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_162),
.B(n_176),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_173),
.B2(n_175),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_176),
.A2(n_177),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_177),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_177),
.B(n_267),
.Y(n_268)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_191),
.C(n_198),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_183),
.A2(n_184),
.B1(n_284),
.B2(n_286),
.Y(n_283)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_190),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_SL g236 ( 
.A(n_188),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_188),
.B(n_237),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_189),
.B(n_294),
.C(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_191),
.B(n_232),
.C(n_233),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_191),
.A2(n_233),
.B1(n_275),
.B2(n_276),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_191),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_191),
.A2(n_198),
.B1(n_275),
.B2(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_191),
.A2(n_275),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_198),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_213),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NOR2xp67_ASAP7_75t_SL g369 ( 
.A(n_215),
.B(n_319),
.Y(n_369)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_218),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_279),
.B(n_287),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_234),
.B(n_278),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_231),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_222),
.B(n_231),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_230),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_225),
.B1(n_238),
.B2(n_239),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_224),
.A2(n_225),
.B1(n_303),
.B2(n_333),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

NAND2xp33_ASAP7_75t_R g271 ( 
.A(n_225),
.B(n_239),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_225),
.B(n_303),
.Y(n_302)
);

AO22x2_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_226),
.B(n_227),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_230),
.B(n_281),
.C(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_233),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_270),
.B(n_277),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_254),
.B(n_269),
.Y(n_235)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI32xp33_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_242),
.A3(n_246),
.B1(n_248),
.B2(n_250),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_266),
.B(n_268),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_261),
.Y(n_256)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_264),
.Y(n_309)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_265),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_272),
.Y(n_277)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_275),
.B(n_317),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_283),
.Y(n_287)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_284),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_336),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_291),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_328),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_328),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_315),
.C(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

XNOR2x1_ASAP7_75t_L g329 ( 
.A(n_295),
.B(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_314),
.B2(n_315),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_297),
.Y(n_349)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2x1_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_300),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_303),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_318),
.B1(n_319),
.B2(n_327),
.Y(n_317)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_310),
.A2(n_359),
.B1(n_363),
.B2(n_366),
.Y(n_358)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_310),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_332),
.C(n_334),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_332),
.A2(n_334),
.B1(n_335),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_332),
.Y(n_340)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_337),
.B(n_338),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_344),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_374),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_350),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_371),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_368),
.B1(n_369),
.B2(n_370),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_356),
.Y(n_370)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2x1_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);


endmodule