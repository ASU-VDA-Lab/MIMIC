module real_jpeg_3588_n_16 (n_5, n_4, n_8, n_0, n_12, n_337, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_337;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_1),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_35),
.B1(n_37),
.B2(n_115),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_1),
.A2(n_51),
.B1(n_53),
.B2(n_115),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_1),
.A2(n_63),
.B1(n_64),
.B2(n_115),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_3),
.A2(n_35),
.B1(n_37),
.B2(n_39),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_3),
.A2(n_39),
.B1(n_51),
.B2(n_53),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_3),
.A2(n_39),
.B1(n_63),
.B2(n_64),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_4),
.A2(n_35),
.B1(n_37),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_4),
.A2(n_44),
.B1(n_63),
.B2(n_64),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_44),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_4),
.A2(n_44),
.B1(n_51),
.B2(n_53),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_5),
.A2(n_63),
.B1(n_64),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_5),
.A2(n_51),
.B1(n_53),
.B2(n_71),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_5),
.A2(n_35),
.B1(n_37),
.B2(n_71),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_6),
.A2(n_35),
.B1(n_37),
.B2(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_6),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_56),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_7),
.A2(n_51),
.B1(n_53),
.B2(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_7),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_63),
.B1(n_64),
.B2(n_81),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_7),
.A2(n_35),
.B1(n_37),
.B2(n_81),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_81),
.Y(n_299)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g78 ( 
.A(n_10),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_12),
.B(n_134),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_12),
.B(n_37),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_12),
.A2(n_29),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_12),
.B(n_63),
.C(n_78),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_12),
.A2(n_51),
.B1(n_53),
.B2(n_106),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_12),
.B(n_57),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_12),
.B(n_67),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_12),
.B(n_76),
.Y(n_214)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_12),
.A2(n_37),
.B(n_163),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_14),
.A2(n_35),
.B1(n_37),
.B2(n_41),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_14),
.A2(n_41),
.B1(n_51),
.B2(n_53),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_14),
.A2(n_41),
.B1(n_63),
.B2(n_64),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_328),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_318),
.B(n_327),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_284),
.B(n_315),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_259),
.B(n_283),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_142),
.B(n_258),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_116),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_22),
.B(n_116),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_86),
.C(n_97),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_23),
.B(n_86),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_58),
.B2(n_59),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_42),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_26),
.B(n_42),
.C(n_58),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_34),
.B1(n_38),
.B2(n_40),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_27),
.A2(n_34),
.B1(n_38),
.B2(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_27),
.A2(n_40),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_27),
.A2(n_34),
.B1(n_114),
.B2(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_27),
.A2(n_271),
.B(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_27),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_27),
.A2(n_34),
.B1(n_299),
.B2(n_311),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_27),
.A2(n_272),
.B(n_311),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_30),
.B(n_106),
.Y(n_105)
);

NAND3xp33_ASAP7_75t_L g107 ( 
.A(n_30),
.B(n_33),
.C(n_37),
.Y(n_107)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_32),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_37),
.Y(n_34)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_32),
.A2(n_35),
.B(n_105),
.C(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_34),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_34),
.A2(n_299),
.B(n_300),
.Y(n_298)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_37),
.B1(n_47),
.B2(n_49),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g164 ( 
.A(n_35),
.B(n_49),
.C(n_53),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_54),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_43),
.A2(n_45),
.B(n_50),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_45),
.A2(n_109),
.B(n_111),
.Y(n_108)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_45),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_45),
.A2(n_50),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_45),
.A2(n_50),
.B1(n_148),
.B2(n_229),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_45),
.A2(n_54),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_47),
.A2(n_51),
.B(n_162),
.C(n_164),
.Y(n_161)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_50),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_50),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g85 ( 
.A1(n_51),
.A2(n_53),
.B1(n_78),
.B2(n_79),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_51),
.B(n_192),
.Y(n_191)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_55),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_57),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_57),
.A2(n_110),
.B1(n_139),
.B2(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_57),
.A2(n_139),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_74),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_60),
.B(n_74),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_69),
.B(n_72),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_66),
.B(n_90),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_61),
.A2(n_72),
.B(n_90),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_61),
.A2(n_66),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_73),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_67),
.B1(n_70),
.B2(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_62),
.A2(n_89),
.B(n_199),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_62),
.A2(n_67),
.B1(n_106),
.B2(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_62),
.A2(n_67),
.B1(n_210),
.B2(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_64),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_63),
.B(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_66),
.A2(n_92),
.B(n_103),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_67),
.B(n_73),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_80),
.B(n_82),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_75),
.A2(n_80),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_75),
.A2(n_95),
.B1(n_157),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_76),
.B(n_83),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_76),
.A2(n_84),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_76),
.A2(n_84),
.B1(n_196),
.B2(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_76),
.A2(n_84),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_77),
.B(n_159),
.Y(n_158)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_78),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_82),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_84),
.A2(n_156),
.B(n_158),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_96),
.B(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_95),
.A2(n_125),
.B(n_159),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_97),
.B(n_241),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_108),
.C(n_113),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_98),
.A2(n_99),
.B1(n_245),
.B2(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_104),
.Y(n_184)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_108),
.B(n_113),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_111),
.B(n_138),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_141),
.Y(n_116)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_127),
.B2(n_128),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_120),
.B(n_128),
.C(n_141),
.Y(n_282)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_122),
.B(n_124),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_122),
.A2(n_126),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g288 ( 
.A1(n_122),
.A2(n_267),
.B(n_269),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_140),
.Y(n_128)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_129),
.Y(n_140)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_132),
.B(n_136),
.C(n_140),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_133),
.B(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_134),
.B(n_273),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_135),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_137),
.Y(n_279)
);

AOI321xp33_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_239),
.A3(n_250),
.B1(n_256),
.B2(n_257),
.C(n_337),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_185),
.B(n_238),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_166),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_145),
.B(n_166),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_155),
.C(n_160),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_146),
.B(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_147),
.B(n_151),
.C(n_154),
.Y(n_181)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_155),
.B(n_160),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_158),
.B(n_277),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_159),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_161),
.B(n_165),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_178),
.B2(n_179),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_167),
.B(n_180),
.C(n_183),
.Y(n_251)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_169),
.B(n_173),
.C(n_177),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_176),
.B2(n_177),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_233),
.B(n_237),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_223),
.B(n_232),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_204),
.B(n_222),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_197),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_197),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_190),
.A2(n_191),
.B1(n_193),
.B2(n_194),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_201),
.C(n_203),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_216),
.B(n_221),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_215),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_212),
.B(n_214),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_220),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_224),
.B(n_225),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_228),
.C(n_230),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_234),
.B(n_236),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_242),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_242),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.C(n_249),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_243),
.A2(n_244),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_252),
.Y(n_256)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_282),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_282),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_265),
.C(n_275),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_273),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_278),
.B(n_281),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_278),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_280),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g287 ( 
.A(n_281),
.B(n_288),
.CI(n_289),
.CON(n_287),
.SN(n_287)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_288),
.C(n_289),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_303),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_287),
.Y(n_316)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_287),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_298),
.B2(n_302),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_295),
.B2(n_296),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_296),
.C(n_298),
.Y(n_306)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_296),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_296),
.B(n_310),
.C(n_314),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_298),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_298),
.A2(n_302),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_306),
.C(n_308),
.Y(n_319)
);

AOI21xp33_ASAP7_75t_L g315 ( 
.A1(n_303),
.A2(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_304),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_312),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_320),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_323),
.B(n_324),
.C(n_326),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_333),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_334),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);


endmodule