module fake_jpeg_690_n_581 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_581);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_581;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_4),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_56),
.B(n_59),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_58),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_62),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_23),
.B(n_22),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_69),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_66),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_65),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_67),
.Y(n_158)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_68),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_22),
.B(n_19),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g162 ( 
.A(n_70),
.Y(n_162)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_74),
.B(n_89),
.Y(n_134)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_34),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_79),
.Y(n_110)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_36),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_80),
.Y(n_122)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_82),
.Y(n_161)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_90),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_88),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_17),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_50),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_25),
.Y(n_91)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_100),
.Y(n_137)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_97),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_98),
.Y(n_151)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_52),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_103),
.Y(n_150)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_52),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_26),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_104),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_165)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_20),
.Y(n_105)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_33),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_106),
.B(n_38),
.Y(n_148)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_53),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_74),
.A2(n_26),
.B1(n_40),
.B2(n_39),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_113),
.A2(n_120),
.B1(n_165),
.B2(n_60),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_72),
.B(n_40),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_119),
.B(n_129),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_104),
.A2(n_20),
.B1(n_39),
.B2(n_24),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_94),
.B1(n_97),
.B2(n_99),
.Y(n_126)
);

AO22x1_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_149),
.B1(n_91),
.B2(n_116),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_128),
.B(n_138),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_40),
.B1(n_81),
.B2(n_71),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_136),
.B(n_28),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_70),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_68),
.B(n_35),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_153),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_61),
.A2(n_42),
.B1(n_41),
.B2(n_48),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_143),
.A2(n_145),
.B1(n_152),
.B2(n_42),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_56),
.A2(n_66),
.B1(n_64),
.B2(n_59),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_148),
.B(n_163),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_53),
.B1(n_38),
.B2(n_48),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_77),
.A2(n_42),
.B1(n_41),
.B2(n_46),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_82),
.B(n_51),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_88),
.A2(n_51),
.B(n_47),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_95),
.B(n_47),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_164),
.B(n_168),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_78),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_45),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_171),
.B(n_173),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_73),
.B(n_44),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_119),
.A2(n_86),
.B1(n_103),
.B2(n_79),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_174),
.A2(n_215),
.B1(n_216),
.B2(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_175),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_113),
.A2(n_101),
.B1(n_100),
.B2(n_87),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_176),
.A2(n_234),
.B1(n_235),
.B2(n_183),
.Y(n_242)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_127),
.Y(n_177)
);

BUFx2_ASAP7_75t_L g256 ( 
.A(n_177),
.Y(n_256)
);

INVxp33_ASAP7_75t_L g283 ( 
.A(n_178),
.Y(n_283)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_127),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_179),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_180),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_115),
.Y(n_181)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_182),
.Y(n_252)
);

INVx11_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_185),
.Y(n_254)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_125),
.Y(n_186)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_186),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_187),
.B(n_197),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_188),
.Y(n_288)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_189),
.Y(n_291)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_190),
.Y(n_240)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_110),
.Y(n_191)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_191),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_114),
.B(n_91),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_192),
.B(n_194),
.Y(n_278)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_134),
.B(n_91),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_133),
.Y(n_196)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_196),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_140),
.B(n_28),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_150),
.Y(n_198)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_199),
.Y(n_266)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_111),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_202),
.B(n_203),
.Y(n_243)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_111),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_21),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_204),
.B(n_219),
.Y(n_263)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_123),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_205),
.B(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_83),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_207),
.B(n_208),
.Y(n_261)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_147),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_210),
.Y(n_253)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_212),
.B(n_213),
.Y(n_264)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_118),
.Y(n_213)
);

INVx11_ASAP7_75t_L g214 ( 
.A(n_145),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_214),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_119),
.A2(n_90),
.B1(n_96),
.B2(n_98),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_129),
.A2(n_67),
.B1(n_57),
.B2(n_93),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_112),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_217),
.B(n_218),
.Y(n_275)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_109),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_122),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_160),
.B(n_148),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_220),
.B(n_222),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_152),
.A2(n_65),
.B1(n_85),
.B2(n_55),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_121),
.B(n_62),
.C(n_58),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_155),
.C(n_133),
.Y(n_251)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_144),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_224),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_146),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_226),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g226 ( 
.A(n_126),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_159),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_230),
.Y(n_248)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_141),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_149),
.B(n_21),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_232),
.Y(n_255)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_146),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_233),
.B(n_236),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_149),
.B(n_84),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_143),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_126),
.B(n_18),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_242),
.A2(n_247),
.B1(n_258),
.B2(n_276),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_246),
.B(n_265),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_234),
.A2(n_131),
.B1(n_112),
.B2(n_157),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_251),
.B(n_196),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_226),
.A2(n_131),
.B1(n_158),
.B2(n_157),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_211),
.B(n_228),
.C(n_174),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_271),
.C(n_272),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_211),
.B(n_141),
.C(n_142),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_142),
.C(n_155),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_158),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_273),
.B(n_277),
.C(n_292),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_175),
.A2(n_156),
.B1(n_154),
.B2(n_169),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_223),
.B(n_185),
.C(n_186),
.Y(n_277)
);

AO21x2_ASAP7_75t_L g280 ( 
.A1(n_221),
.A2(n_169),
.B(n_102),
.Y(n_280)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_280),
.A2(n_217),
.B(n_203),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_216),
.A2(n_156),
.B1(n_154),
.B2(n_107),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_284),
.A2(n_286),
.B1(n_290),
.B2(n_6),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_175),
.A2(n_80),
.B1(n_75),
.B2(n_54),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_215),
.A2(n_117),
.B1(n_76),
.B2(n_3),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_201),
.B(n_117),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_230),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_214),
.A2(n_162),
.B(n_2),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_245),
.B(n_267),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_199),
.A2(n_18),
.B1(n_2),
.B2(n_3),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_189),
.B(n_162),
.C(n_2),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_248),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_314),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_294),
.B(n_304),
.Y(n_347)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_296),
.B(n_306),
.C(n_311),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_SL g354 ( 
.A1(n_297),
.A2(n_322),
.B(n_286),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_250),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_298),
.B(n_301),
.Y(n_351)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_248),
.Y(n_299)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_299),
.Y(n_369)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_279),
.Y(n_300)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_300),
.Y(n_382)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_243),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_303),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_212),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_264),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_200),
.C(n_205),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_249),
.B(n_190),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_307),
.B(n_309),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_308),
.B(n_320),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_249),
.B(n_208),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_257),
.B(n_202),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_310),
.B(n_312),
.Y(n_387)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_213),
.C(n_182),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_257),
.B(n_268),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_237),
.Y(n_314)
);

NOR2x1_ASAP7_75t_L g315 ( 
.A(n_255),
.B(n_179),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_315),
.B(n_317),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_268),
.B(n_222),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_245),
.A2(n_219),
.B(n_184),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_319),
.A2(n_280),
.B(n_285),
.Y(n_346)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_267),
.A2(n_210),
.B1(n_209),
.B2(n_188),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_321),
.A2(n_329),
.B1(n_333),
.B2(n_334),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_289),
.A2(n_177),
.B(n_162),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_181),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_324),
.C(n_292),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g324 ( 
.A(n_274),
.B(n_180),
.C(n_3),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_281),
.B(n_1),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_325),
.B(n_327),
.Y(n_349)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_326),
.B(n_328),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_275),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_255),
.B(n_1),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_4),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_338),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_244),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_332),
.Y(n_353)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_288),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_265),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_260),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_281),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_339),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_276),
.A2(n_15),
.B1(n_8),
.B2(n_9),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_336),
.A2(n_329),
.B1(n_318),
.B2(n_280),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_SL g372 ( 
.A1(n_337),
.A2(n_340),
.B(n_343),
.Y(n_372)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_261),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_288),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_341),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_239),
.B(n_8),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_342),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_263),
.B(n_8),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_346),
.A2(n_354),
.B(n_365),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_358),
.B(n_324),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_297),
.A2(n_283),
.B(n_287),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_360),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_296),
.B(n_302),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_363),
.B(n_367),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_251),
.C(n_271),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_364),
.B(n_370),
.C(n_371),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_283),
.B(n_246),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_316),
.B(n_270),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_316),
.B(n_270),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_311),
.B(n_240),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_323),
.B(n_269),
.C(n_240),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_374),
.C(n_375),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_304),
.B(n_247),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_291),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_313),
.A2(n_284),
.B(n_280),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_376),
.B(n_308),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_313),
.B(n_291),
.C(n_252),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_379),
.C(n_381),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_330),
.B(n_252),
.C(n_259),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_294),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_383),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_299),
.B(n_259),
.C(n_256),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_305),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_385),
.A2(n_386),
.B1(n_333),
.B2(n_319),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_318),
.A2(n_280),
.B1(n_266),
.B2(n_258),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_256),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_388),
.B(n_320),
.C(n_341),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_344),
.B(n_293),
.Y(n_389)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_389),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_351),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_391),
.B(n_396),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_380),
.B(n_357),
.Y(n_392)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_392),
.Y(n_442)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_382),
.Y(n_393)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_393),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_394),
.Y(n_444)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_382),
.Y(n_395)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_395),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_315),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_364),
.C(n_367),
.Y(n_437)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_384),
.Y(n_400)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_400),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_363),
.B(n_328),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_401),
.B(n_420),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_365),
.A2(n_352),
.B1(n_346),
.B2(n_369),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_402),
.A2(n_419),
.B1(n_366),
.B2(n_385),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_353),
.Y(n_403)
);

BUFx24_ASAP7_75t_L g439 ( 
.A(n_403),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_386),
.A2(n_321),
.B1(n_331),
.B2(n_334),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_412),
.B1(n_418),
.B2(n_422),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_362),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_406),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_303),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_387),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_407),
.Y(n_434)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_369),
.Y(n_408)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_357),
.B(n_300),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_414),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_368),
.B(n_340),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g415 ( 
.A(n_388),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_415),
.B(n_416),
.Y(n_446)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_368),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_377),
.B(n_338),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_352),
.A2(n_336),
.B1(n_266),
.B2(n_253),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_370),
.B(n_326),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_421),
.B(n_373),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_377),
.B(n_332),
.Y(n_422)
);

OA22x2_ASAP7_75t_L g423 ( 
.A1(n_354),
.A2(n_314),
.B1(n_295),
.B2(n_238),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_423),
.B(n_426),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_348),
.B(n_238),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_425),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g426 ( 
.A1(n_359),
.A2(n_241),
.B1(n_10),
.B2(n_11),
.Y(n_426)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_427),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_424),
.A2(n_360),
.B(n_350),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_428),
.A2(n_432),
.B(n_456),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_355),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_429),
.B(n_460),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_350),
.B(n_366),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_449),
.C(n_450),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_412),
.A2(n_366),
.B1(n_374),
.B2(n_372),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_438),
.A2(n_447),
.B1(n_455),
.B2(n_415),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_402),
.A2(n_347),
.B1(n_375),
.B2(n_359),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_371),
.C(n_355),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_417),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_451),
.B(n_442),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_390),
.B(n_358),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_452),
.B(n_454),
.C(n_356),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_399),
.B(n_347),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_417),
.A2(n_378),
.B1(n_376),
.B2(n_381),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_410),
.A2(n_424),
.B(n_417),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_389),
.A2(n_349),
.B(n_345),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_458),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_420),
.B(n_379),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_403),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_461),
.B(n_440),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_458),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_463),
.B(n_464),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_431),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_430),
.B(n_413),
.Y(n_467)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_467),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_414),
.Y(n_468)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_468),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_448),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_469),
.B(n_475),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_437),
.B(n_411),
.C(n_409),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_472),
.C(n_476),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_411),
.C(n_409),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_473),
.A2(n_483),
.B1(n_484),
.B2(n_485),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_439),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_398),
.C(n_421),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_445),
.Y(n_477)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_478),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_450),
.B(n_401),
.C(n_416),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_486),
.C(n_423),
.Y(n_510)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_433),
.Y(n_480)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_480),
.Y(n_506)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_433),
.Y(n_481)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_481),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_442),
.B(n_392),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_482),
.Y(n_508)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_436),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_443),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_408),
.C(n_423),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_441),
.A2(n_419),
.B1(n_423),
.B2(n_400),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_487),
.A2(n_488),
.B1(n_444),
.B2(n_455),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_427),
.A2(n_438),
.B1(n_444),
.B2(n_447),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_429),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_492),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_474),
.A2(n_456),
.B(n_432),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_494),
.A2(n_495),
.B(n_498),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_474),
.A2(n_428),
.B(n_446),
.Y(n_495)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_496),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_486),
.A2(n_446),
.B(n_439),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_502),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_480),
.B1(n_481),
.B2(n_487),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_503),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_460),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_466),
.A2(n_453),
.B1(n_439),
.B2(n_435),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_472),
.B(n_435),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_510),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_465),
.B(n_393),
.C(n_397),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_511),
.B(n_470),
.C(n_465),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_471),
.B(n_459),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_512),
.B(n_508),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_515),
.B(n_522),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_490),
.C(n_504),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_517),
.B(n_518),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_513),
.B(n_471),
.Y(n_518)
);

XOR2x1_ASAP7_75t_L g521 ( 
.A(n_503),
.B(n_473),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_521),
.B(n_491),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_490),
.B(n_462),
.C(n_476),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_479),
.Y(n_524)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_524),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_525),
.B(n_527),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_502),
.B(n_462),
.C(n_488),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_482),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_528),
.B(n_531),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_500),
.B(n_468),
.C(n_467),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_529),
.B(n_530),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_498),
.A2(n_478),
.B(n_477),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_493),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_492),
.B(n_495),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_532),
.B(n_484),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g534 ( 
.A1(n_514),
.A2(n_494),
.B(n_501),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_534),
.B(n_538),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_517),
.B(n_499),
.C(n_491),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_536),
.B(n_539),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_523),
.A2(n_507),
.B1(n_509),
.B2(n_506),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g550 ( 
.A1(n_537),
.A2(n_540),
.B1(n_520),
.B2(n_532),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_515),
.B(n_509),
.C(n_506),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_520),
.A2(n_526),
.B1(n_453),
.B2(n_521),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_505),
.C(n_493),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_543),
.B(n_527),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_505),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_544),
.B(n_546),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_483),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_547),
.B(n_542),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_548),
.B(n_516),
.Y(n_549)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_549),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_550),
.B(n_554),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_516),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_551),
.B(n_553),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_535),
.B(n_519),
.C(n_457),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_556),
.B(n_559),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_538),
.A2(n_395),
.B1(n_361),
.B2(n_345),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_557),
.A2(n_540),
.B1(n_539),
.B2(n_536),
.Y(n_562)
);

AOI21xp33_ASAP7_75t_L g558 ( 
.A1(n_545),
.A2(n_361),
.B(n_10),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g561 ( 
.A1(n_558),
.A2(n_534),
.B(n_544),
.Y(n_561)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_543),
.Y(n_559)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_561),
.Y(n_572)
);

CKINVDCx20_ASAP7_75t_R g573 ( 
.A(n_562),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_549),
.B(n_541),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_556),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g566 ( 
.A1(n_555),
.A2(n_9),
.B(n_10),
.Y(n_566)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_566),
.B(n_552),
.C(n_560),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_570),
.Y(n_576)
);

AOI21x1_ASAP7_75t_L g570 ( 
.A1(n_567),
.A2(n_552),
.B(n_560),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_571),
.B(n_563),
.Y(n_574)
);

AOI21xp5_ASAP7_75t_SL g577 ( 
.A1(n_574),
.A2(n_572),
.B(n_568),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_573),
.B(n_564),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_575),
.A2(n_568),
.B(n_11),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_577),
.A2(n_578),
.B1(n_576),
.B2(n_9),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_9),
.B1(n_13),
.B2(n_475),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_13),
.Y(n_581)
);


endmodule