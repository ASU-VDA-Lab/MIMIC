module fake_jpeg_22496_n_171 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_171);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_171;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx8_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_36),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx16f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g34 ( 
.A(n_23),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_35),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g35 ( 
.A1(n_26),
.A2(n_2),
.B(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_54),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_27),
.B1(n_26),
.B2(n_28),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_51),
.B1(n_27),
.B2(n_37),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_19),
.B1(n_28),
.B2(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_30),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_55),
.B(n_30),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_20),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_27),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_52),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_50),
.B1(n_49),
.B2(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_20),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_53),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_68),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_17),
.B1(n_18),
.B2(n_24),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_54),
.B(n_17),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_42),
.B(n_18),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_69),
.B(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_51),
.A2(n_18),
.B1(n_24),
.B2(n_16),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_25),
.B1(n_16),
.B2(n_21),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_21),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_55),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_91),
.C(n_88),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_80),
.B1(n_86),
.B2(n_72),
.Y(n_105)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_63),
.A2(n_55),
.B(n_48),
.C(n_56),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_15),
.B1(n_21),
.B2(n_22),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_50),
.B1(n_49),
.B2(n_41),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_88),
.B1(n_67),
.B2(n_72),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_62),
.A2(n_47),
.B1(n_16),
.B2(n_25),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_56),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_69),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_58),
.A2(n_47),
.B1(n_19),
.B2(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_92),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_52),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_90),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_98),
.B1(n_105),
.B2(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_103),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_64),
.B1(n_60),
.B2(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_102),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_100),
.B(n_79),
.C(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_101),
.A2(n_106),
.B1(n_78),
.B2(n_73),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_60),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_104),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_82),
.Y(n_117)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_115),
.C(n_96),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_100),
.A2(n_80),
.B(n_76),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_111),
.A2(n_121),
.B(n_122),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_105),
.A2(n_84),
.B1(n_80),
.B2(n_77),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_118),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_102),
.C(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_119),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_94),
.A2(n_73),
.B1(n_15),
.B2(n_25),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_120),
.B(n_98),
.C(n_5),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_82),
.B(n_86),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_24),
.B(n_22),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_4),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_132),
.B(n_117),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.C(n_134),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_101),
.Y(n_127)
);

AOI322xp5_ASAP7_75t_L g128 ( 
.A1(n_121),
.A2(n_93),
.A3(n_15),
.B1(n_9),
.B2(n_12),
.C1(n_13),
.C2(n_10),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_112),
.B(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_131),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_5),
.B(n_6),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_9),
.C(n_10),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_135),
.A2(n_113),
.B1(n_114),
.B2(n_112),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_126),
.B1(n_129),
.B2(n_134),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_143),
.Y(n_153)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_141),
.B(n_142),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_132),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_116),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_144),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_127),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_123),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_150),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_140),
.B(n_122),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_151),
.B(n_147),
.C(n_148),
.Y(n_157)
);

XNOR2x1_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_119),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_152),
.B(n_136),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_146),
.A2(n_137),
.B1(n_140),
.B2(n_138),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_154),
.A2(n_149),
.B1(n_7),
.B2(n_8),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_139),
.C(n_12),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_149),
.B(n_6),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_158),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_160),
.Y(n_166)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_6),
.B(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_156),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_163),
.C(n_155),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_162),
.B(n_160),
.Y(n_168)
);

AOI31xp33_ASAP7_75t_L g170 ( 
.A1(n_168),
.A2(n_169),
.A3(n_167),
.B(n_7),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_8),
.Y(n_171)
);


endmodule