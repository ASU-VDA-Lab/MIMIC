module fake_jpeg_7399_n_334 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_334);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_334;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_25),
.Y(n_54)
);

INVx11_ASAP7_75t_SL g40 ( 
.A(n_35),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_32),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_0),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_23),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_60),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_57),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_54),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_24),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_28),
.B1(n_33),
.B2(n_19),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_68),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_38),
.B(n_23),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_20),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_30),
.B(n_20),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_21),
.C(n_32),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_26),
.B1(n_21),
.B2(n_36),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_75),
.Y(n_111)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_76),
.B(n_81),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_90),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_65),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_83),
.B(n_86),
.Y(n_117)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_84),
.Y(n_122)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_65),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_37),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_19),
.B1(n_28),
.B2(n_33),
.Y(n_105)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_60),
.B(n_27),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_112),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_64),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_91),
.C(n_88),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_105),
.A2(n_107),
.B1(n_124),
.B2(n_26),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_108),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_73),
.A2(n_45),
.B1(n_52),
.B2(n_65),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_82),
.B(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_71),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_70),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_0),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_114),
.A2(n_125),
.B(n_110),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_118),
.Y(n_153)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_126),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_86),
.A2(n_46),
.B1(n_41),
.B2(n_61),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_11),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_76),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_71),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_131),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_52),
.B1(n_78),
.B2(n_56),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_140),
.B1(n_146),
.B2(n_152),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_71),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_136),
.C(n_137),
.Y(n_165)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_132),
.Y(n_162)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_133),
.B(n_150),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_122),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_77),
.C(n_93),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_144),
.B(n_154),
.Y(n_176)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_139),
.B(n_143),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_75),
.B1(n_46),
.B2(n_45),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_95),
.Y(n_144)
);

XOR2x2_ASAP7_75t_SL g186 ( 
.A(n_147),
.B(n_8),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_148),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_105),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_93),
.C(n_44),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_44),
.C(n_119),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_99),
.A2(n_45),
.B1(n_96),
.B2(n_84),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_115),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_111),
.B(n_34),
.Y(n_155)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_113),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_99),
.A2(n_67),
.B1(n_62),
.B2(n_36),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_157),
.A2(n_108),
.B1(n_101),
.B2(n_98),
.Y(n_160)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_163),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_164),
.B1(n_174),
.B2(n_182),
.Y(n_193)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_139),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_62),
.B1(n_55),
.B2(n_36),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_111),
.B(n_44),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_166),
.A2(n_168),
.B(n_171),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_167),
.B(n_169),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_36),
.B1(n_74),
.B2(n_101),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

HB1xp67_ASAP7_75t_SL g218 ( 
.A(n_170),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_153),
.B1(n_128),
.B2(n_141),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_98),
.B1(n_74),
.B2(n_59),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_149),
.A2(n_44),
.B(n_87),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_177),
.A2(n_181),
.B(n_134),
.Y(n_192)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_185),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_147),
.A2(n_98),
.B1(n_18),
.B2(n_31),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_180),
.A2(n_100),
.B1(n_29),
.B2(n_25),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_154),
.A2(n_18),
.B(n_31),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_127),
.A2(n_131),
.B1(n_137),
.B2(n_146),
.Y(n_182)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_184),
.Y(n_197)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_8),
.C(n_16),
.Y(n_210)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_157),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_187),
.B(n_191),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_133),
.A2(n_38),
.A3(n_18),
.B1(n_31),
.B2(n_29),
.Y(n_188)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_188),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_129),
.C(n_147),
.Y(n_203)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_192),
.A2(n_196),
.B(n_204),
.Y(n_233)
);

XOR2x2_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_138),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_135),
.B(n_130),
.C(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

NAND2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_136),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_202),
.B(n_214),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_206),
.C(n_211),
.Y(n_232)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_44),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_205),
.A2(n_181),
.B(n_173),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_182),
.B(n_44),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_100),
.Y(n_207)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_207),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_81),
.B1(n_120),
.B2(n_59),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_209),
.B1(n_213),
.B2(n_220),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_162),
.A2(n_92),
.B1(n_25),
.B2(n_34),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_216),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_165),
.B(n_22),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_168),
.A2(n_22),
.B1(n_10),
.B2(n_12),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_212),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_170),
.A2(n_22),
.B1(n_2),
.B2(n_3),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_174),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_166),
.A2(n_7),
.B1(n_15),
.B2(n_14),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_219),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_164),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_222),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_223),
.B(n_224),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_194),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_167),
.B(n_169),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_228),
.A2(n_216),
.B1(n_193),
.B2(n_199),
.Y(n_259)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_230),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_201),
.B(n_159),
.Y(n_231)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_165),
.C(n_190),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_241),
.C(n_243),
.Y(n_253)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_198),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_240),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_192),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_218),
.B(n_185),
.Y(n_239)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_161),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_161),
.C(n_183),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_207),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_244),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_177),
.C(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_195),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_196),
.B(n_188),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_245),
.B(n_246),
.C(n_200),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_180),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_237),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_244),
.A2(n_217),
.B1(n_199),
.B2(n_195),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_252),
.A2(n_262),
.B1(n_264),
.B2(n_247),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_255),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_208),
.C(n_193),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_265),
.C(n_267),
.Y(n_274)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_204),
.B1(n_220),
.B2(n_197),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_260),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_197),
.B1(n_158),
.B2(n_189),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_240),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_263),
.B(n_226),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_230),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_232),
.B(n_186),
.C(n_179),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_227),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_215),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_256),
.A2(n_228),
.B(n_249),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_268),
.A2(n_278),
.B(n_281),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_250),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_270),
.B(n_277),
.Y(n_292)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_272),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_266),
.A2(n_225),
.B1(n_234),
.B2(n_224),
.Y(n_273)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_250),
.B(n_238),
.CI(n_233),
.CON(n_275),
.SN(n_275)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_7),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_255),
.B(n_245),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_246),
.C(n_248),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_251),
.A2(n_234),
.B1(n_233),
.B2(n_239),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_279),
.A2(n_252),
.B1(n_258),
.B2(n_254),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_258),
.A2(n_235),
.B(n_229),
.Y(n_281)
);

AO221x1_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_235),
.B1(n_213),
.B2(n_229),
.C(n_243),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_257),
.C(n_265),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_226),
.Y(n_291)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_285),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_253),
.C(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_288),
.C(n_294),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_291),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_253),
.C(n_241),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_290),
.B(n_280),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_271),
.B(n_275),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_7),
.C(n_14),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_276),
.B(n_6),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_299),
.C(n_10),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_5),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_1),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_5),
.C(n_13),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_302),
.B(n_304),
.C(n_305),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_280),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_268),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_295),
.A2(n_269),
.B1(n_271),
.B2(n_282),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_306),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_277),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_307),
.B(n_275),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_309),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_281),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_310),
.B(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_311),
.B(n_12),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_312),
.B(n_315),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_317),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_300),
.B(n_299),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_SL g318 ( 
.A(n_304),
.B(n_288),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_305),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_302),
.C(n_5),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_303),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_322),
.B(n_4),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_320),
.B(n_307),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_326),
.Y(n_328)
);

AOI21x1_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_314),
.B(n_312),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_329),
.C(n_323),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_328),
.C(n_325),
.Y(n_331)
);

AOI321xp33_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_4),
.A3(n_12),
.B1(n_13),
.B2(n_16),
.C(n_2),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_1),
.Y(n_333)
);

HAxp5_ASAP7_75t_SL g334 ( 
.A(n_333),
.B(n_3),
.CON(n_334),
.SN(n_334)
);


endmodule