module real_jpeg_30991_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_0),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_0),
.B(n_86),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_0),
.B(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_1),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_1),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_1),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_205),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_1),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_1),
.B(n_284),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_2),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_2),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_3),
.B(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_3),
.B(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_5),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_5),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_5),
.B(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_5),
.B(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_5),
.B(n_245),
.Y(n_244)
);

NAND2x1p5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_6),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_6),
.B(n_107),
.Y(n_106)
);

NAND2x1_ASAP7_75t_L g155 ( 
.A(n_6),
.B(n_122),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_6),
.B(n_237),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_7),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_7),
.B(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_7),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_7),
.B(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_7),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_9),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_9),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_9),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_9),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_9),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_9),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_9),
.B(n_293),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_10),
.Y(n_238)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_11),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_14),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_15),
.B(n_73),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_15),
.B(n_174),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_189),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_188),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_145),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_20),
.B(n_145),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_101),
.C(n_132),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_21),
.B(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_23),
.B(n_63),
.C(n_147),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_24)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_29),
.B(n_35),
.C(n_36),
.Y(n_151)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_33),
.Y(n_293)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_34),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.C(n_44),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g131 ( 
.A(n_37),
.Y(n_131)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_40),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_41),
.A2(n_44),
.B1(n_45),
.B2(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_41),
.Y(n_130)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_43),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_43),
.Y(n_310)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_48),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_60),
.B2(n_61),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_51),
.B(n_55),
.C(n_61),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_54),
.Y(n_112)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_54),
.Y(n_171)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_59),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_59),
.Y(n_259)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_78),
.C(n_87),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_64),
.B(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_65),
.B(n_72),
.C(n_76),
.Y(n_142)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_76),
.B2(n_77),
.Y(n_69)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_78),
.A2(n_79),
.B1(n_87),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_80),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_80),
.A2(n_83),
.B1(n_187),
.B2(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_82),
.Y(n_246)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_82),
.Y(n_299)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_83),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_86),
.Y(n_285)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_87),
.Y(n_196)
);

MAJx2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_90),
.C(n_95),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_88),
.A2(n_95),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_88),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_89),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_90),
.B(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_99),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2x1_ASAP7_75t_SL g192 ( 
.A(n_102),
.B(n_132),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_119),
.C(n_127),
.Y(n_102)
);

XNOR2x1_ASAP7_75t_L g222 ( 
.A(n_103),
.B(n_223),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.C(n_113),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_104),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_106),
.A2(n_182),
.B1(n_183),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g182 ( 
.A(n_106),
.Y(n_182)
);

AO22x1_ASAP7_75t_SL g327 ( 
.A1(n_106),
.A2(n_182),
.B1(n_244),
.B2(n_328),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_107),
.Y(n_317)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_109),
.B(n_114),
.Y(n_249)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_120),
.B(n_128),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_123),
.B(n_126),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_123),
.Y(n_126)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_126),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.Y(n_128)
);

XOR2x2_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

MAJx2_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_142),
.C(n_143),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_139),
.C(n_140),
.Y(n_153)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_140),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_162),
.Y(n_148)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_161),
.Y(n_149)
);

AO22x2_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_159),
.B2(n_160),
.Y(n_150)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

XOR2x2_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_176),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_173),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_165),
.A2(n_166),
.B1(n_169),
.B2(n_172),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_169),
.Y(n_172)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_175),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_182),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_183),
.Y(n_186)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_224),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NOR2xp67_ASAP7_75t_SL g226 ( 
.A(n_191),
.B(n_193),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_197),
.C(n_221),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_222),
.Y(n_230)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.C(n_218),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_199),
.B(n_233),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_203),
.B(n_218),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_208),
.C(n_215),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_204),
.B(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_207),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_208),
.A2(n_209),
.B1(n_215),
.B2(n_216),
.Y(n_268)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_210),
.B(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2x1p5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_250),
.B(n_338),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_229),
.B(n_231),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.C(n_247),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_239),
.C(n_243),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_239),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_238),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_240),
.B(n_285),
.Y(n_296)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_244),
.Y(n_328)
);

BUFx4f_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_271),
.B(n_337),
.Y(n_250)
);

NOR2x1_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_269),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_252),
.B(n_269),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_265),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_254),
.B(n_334),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_256),
.A2(n_266),
.B1(n_267),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_256),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_262),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_257),
.B(n_260),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_262),
.B(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_298),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_331),
.B(n_336),
.Y(n_271)
);

OAI21x1_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_319),
.B(n_330),
.Y(n_272)
);

OA21x2_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_300),
.B(n_318),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_286),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_286),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_282),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_277),
.A2(n_278),
.B1(n_282),
.B2(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_277),
.B(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_294),
.B2(n_295),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_292),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_292),
.C(n_294),
.Y(n_329)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_297),
.Y(n_325)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_312),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_311),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_303),
.A2(n_311),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_316),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx8_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_329),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_320),
.B(n_329),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_321),
.B(n_324),
.C(n_327),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_324),
.A2(n_325),
.B1(n_326),
.B2(n_327),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);


endmodule