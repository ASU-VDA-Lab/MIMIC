module real_jpeg_24939_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_348, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_348;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_1),
.A2(n_42),
.B1(n_44),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_1),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_131),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_131),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_1),
.A2(n_58),
.B1(n_65),
.B2(n_131),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_4),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_5),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_5),
.A2(n_26),
.B1(n_27),
.B2(n_59),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_59),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_5),
.A2(n_42),
.B1(n_44),
.B2(n_59),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_6),
.A2(n_37),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_6),
.A2(n_37),
.B1(n_57),
.B2(n_66),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_7),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_7),
.B(n_67),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_7),
.B(n_29),
.C(n_33),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_7),
.B(n_45),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_7),
.A2(n_108),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_10),
.A2(n_65),
.B1(n_70),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_10),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_10),
.A2(n_42),
.B1(n_44),
.B2(n_138),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_138),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_138),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_11),
.A2(n_42),
.B1(n_44),
.B2(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_11),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_129),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_11),
.A2(n_26),
.B1(n_27),
.B2(n_129),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_129),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_13),
.A2(n_42),
.B1(n_44),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_13),
.A2(n_51),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_13),
.A2(n_33),
.B1(n_34),
.B2(n_51),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_51),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_14),
.A2(n_69),
.B1(n_70),
.B2(n_73),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_14),
.A2(n_42),
.B1(n_44),
.B2(n_69),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_69),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_69),
.Y(n_279)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_15),
.Y(n_152)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_15),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_98),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_96),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_85),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_85),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_74),
.C(n_79),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_20),
.A2(n_74),
.B1(n_332),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_20),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_38),
.B2(n_39),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_74),
.C(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_22),
.A2(n_23),
.B1(n_80),
.B2(n_81),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_23),
.B(n_38),
.C(n_54),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_32),
.B(n_35),
.Y(n_23)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_24),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_24),
.A2(n_35),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_24),
.A2(n_32),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_24),
.A2(n_32),
.B1(n_184),
.B2(n_191),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_24),
.A2(n_249),
.B(n_250),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_24),
.A2(n_32),
.B1(n_117),
.B2(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_24),
.A2(n_125),
.B(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_32),
.Y(n_24)
);

OAI22xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_26),
.A2(n_27),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

NAND3xp33_ASAP7_75t_L g228 ( 
.A(n_26),
.B(n_42),
.C(n_48),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_27),
.B(n_180),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_47),
.B(n_227),
.C(n_228),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_31),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_32),
.A2(n_117),
.B(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_32),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_32),
.B(n_134),
.Y(n_218)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_33),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_34),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_36),
.B(n_126),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_49),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_40),
.A2(n_83),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_41),
.A2(n_45),
.B(n_52),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_41),
.Y(n_272)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_44),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_42),
.A2(n_62),
.B(n_135),
.C(n_154),
.Y(n_153)
);

HAxp5_ASAP7_75t_SL g227 ( 
.A(n_42),
.B(n_134),
.CON(n_227),
.SN(n_227)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND3xp33_ASAP7_75t_L g154 ( 
.A(n_44),
.B(n_58),
.C(n_63),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_45),
.B(n_50),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_45),
.A2(n_52),
.B1(n_128),
.B2(n_130),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_45),
.A2(n_52),
.B1(n_164),
.B2(n_227),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_45),
.A2(n_52),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_46),
.A2(n_83),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_46),
.A2(n_49),
.B(n_302),
.Y(n_301)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_52),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_67),
.B2(n_68),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_56),
.A2(n_61),
.B(n_75),
.Y(n_74)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_60),
.A2(n_68),
.B(n_90),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_60),
.A2(n_67),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_60),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_60),
.A2(n_67),
.B1(n_145),
.B2(n_269),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_61),
.A2(n_137),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_66),
.B(n_134),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_67),
.B(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_67),
.B(n_300),
.Y(n_299)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_70),
.A2(n_134),
.B(n_135),
.Y(n_133)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_74),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_74),
.Y(n_332)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_79),
.B(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_82),
.Y(n_325)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_83),
.A2(n_84),
.B(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_94),
.B2(n_95),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_88),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_89),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_91),
.A2(n_143),
.B(n_318),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI321xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_329),
.A3(n_340),
.B1(n_345),
.B2(n_346),
.C(n_348),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_307),
.B(n_328),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_284),
.B(n_306),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_172),
.B(n_260),
.C(n_283),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_156),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_103),
.B(n_156),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_139),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B1(n_121),
.B2(n_122),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_105),
.B(n_122),
.C(n_139),
.Y(n_261)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_116),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_107),
.B(n_116),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_110),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_108),
.B(n_115),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_108),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_108),
.A2(n_202),
.B1(n_209),
.B2(n_215),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_108),
.A2(n_113),
.B(n_291),
.Y(n_290)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx3_ASAP7_75t_SL g170 ( 
.A(n_109),
.Y(n_170)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_109),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_112),
.A2(n_196),
.B(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_113),
.Y(n_195)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_118),
.B(n_250),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_120),
.A2(n_126),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_127),
.C(n_132),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_130),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_132),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_134),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_148),
.B2(n_155),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_142),
.B(n_146),
.C(n_155),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_143),
.A2(n_298),
.B(n_299),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_148),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_153),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_151),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_160),
.C(n_161),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_157),
.B(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_160),
.B(n_161),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.C(n_168),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_162),
.B(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_244)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_171),
.B(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_259),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_254),
.B(n_258),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_239),
.B(n_253),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_223),
.B(n_238),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_197),
.B(n_222),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_185),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_178),
.B(n_185),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_179),
.Y(n_205)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_193),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_196),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_206),
.B(n_221),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_204),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_217),
.B(n_220),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_213),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_219),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_237),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_237),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_232),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_233),
.C(n_236),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_229),
.B1(n_230),
.B2(n_231),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_226),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_231),
.Y(n_247)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_229),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_235),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_243),
.B1(n_245),
.B2(n_246),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_242),
.B(n_248),
.C(n_251),
.Y(n_257)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_251),
.B2(n_252),
.Y(n_246)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_247),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_257),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_262),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_282),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_273),
.B1(n_280),
.B2(n_281),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_268),
.C(n_270),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_271),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_273),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_280),
.C(n_282),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_274),
.B(n_278),
.Y(n_303)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_285),
.B(n_286),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_305),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_294),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_288),
.B(n_294),
.C(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_289),
.A2(n_290),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_313),
.B(n_317),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_292),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_292),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_301),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_297),
.B(n_301),
.C(n_304),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_300),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_302),
.Y(n_324)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_308),
.B(n_309),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_327),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_320),
.B2(n_321),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_312),
.B(n_320),
.C(n_327),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_315),
.B2(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B(n_326),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_326),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_326),
.A2(n_331),
.B1(n_335),
.B2(n_344),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_337),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_330),
.B(n_337),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.C(n_336),
.Y(n_330)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_331),
.Y(n_344)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_343),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_341),
.B(n_342),
.Y(n_345)
);


endmodule