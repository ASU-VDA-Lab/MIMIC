module fake_jpeg_28650_n_479 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_479);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_479;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_288;
wire n_21;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_52),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_68),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_58),
.Y(n_129)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_36),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx13_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_63),
.Y(n_112)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_64),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_15),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_69),
.B(n_85),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_71),
.Y(n_139)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_76),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_77),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_78),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_80),
.B(n_83),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_81),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_13),
.Y(n_85)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_16),
.Y(n_86)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_91),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_89),
.Y(n_131)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_92),
.Y(n_145)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_33),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_19),
.Y(n_143)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_26),
.Y(n_94)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_94),
.Y(n_138)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_97),
.Y(n_120)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_82),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_89),
.B(n_49),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_48),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_137),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_61),
.B(n_38),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_38),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_53),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_127),
.B(n_140),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_49),
.C(n_16),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_143),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_42),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_93),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_51),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_141),
.B(n_142),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_42),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_31),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_146),
.B(n_31),
.Y(n_183)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_150),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_153),
.Y(n_231)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

CKINVDCx12_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_156),
.B(n_157),
.Y(n_216)
);

CKINVDCx12_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_118),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_158),
.Y(n_205)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_160),
.Y(n_232)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_118),
.Y(n_162)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

INVx2_ASAP7_75t_R g166 ( 
.A(n_116),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_166),
.A2(n_183),
.B(n_32),
.Y(n_208)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_167),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_168),
.B(n_179),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_132),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_173),
.B1(n_180),
.B2(n_103),
.Y(n_201)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

INVx13_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_55),
.B1(n_50),
.B2(n_74),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_143),
.A2(n_88),
.B1(n_67),
.B2(n_73),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_175),
.A2(n_177),
.B1(n_194),
.B2(n_107),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_52),
.B1(n_60),
.B2(n_65),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_130),
.Y(n_178)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_178),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_101),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_108),
.A2(n_70),
.B1(n_95),
.B2(n_33),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_182),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_124),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

INVx13_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_186),
.B(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_187),
.B(n_199),
.Y(n_228)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_196),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_111),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_190),
.B(n_81),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_124),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_191),
.A2(n_198),
.B1(n_134),
.B2(n_102),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_125),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_144),
.A2(n_105),
.B1(n_110),
.B2(n_107),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_129),
.Y(n_196)
);

CKINVDCx9p33_ASAP7_75t_R g197 ( 
.A(n_111),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_197),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_138),
.B(n_32),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_200),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_201),
.A2(n_152),
.B1(n_133),
.B2(n_102),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_120),
.B(n_103),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_202),
.A2(n_224),
.B(n_228),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_195),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_206),
.B(n_219),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_208),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_138),
.C(n_109),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_175),
.C(n_188),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_161),
.B(n_110),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g224 ( 
.A1(n_166),
.A2(n_47),
.B(n_43),
.C(n_37),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_180),
.A2(n_152),
.B1(n_105),
.B2(n_134),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

INVx13_ASAP7_75t_L g241 ( 
.A(n_227),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_139),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_237),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_202),
.A2(n_164),
.B(n_153),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_240),
.A2(n_205),
.B(n_204),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_233),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_242),
.B(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_190),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_253),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_246),
.B(n_254),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_212),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_248),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_249),
.A2(n_258),
.B1(n_273),
.B2(n_209),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_206),
.B(n_48),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_250),
.B(n_266),
.Y(n_302)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_251),
.Y(n_282)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_231),
.B(n_171),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_234),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_255),
.Y(n_304)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_261),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_201),
.A2(n_215),
.B1(n_210),
.B2(n_231),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_178),
.C(n_162),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_260),
.C(n_205),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_181),
.C(n_200),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_158),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_263),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_155),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_230),
.B(n_172),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_264),
.B(n_265),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_155),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_224),
.B(n_41),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_222),
.B(n_47),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_41),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_197),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_268),
.B(n_205),
.Y(n_280)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_272),
.Y(n_291)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_213),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_211),
.A2(n_117),
.B1(n_114),
.B2(n_163),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_257),
.A2(n_177),
.B1(n_194),
.B2(n_117),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_274),
.A2(n_276),
.B1(n_284),
.B2(n_285),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_246),
.A2(n_114),
.B1(n_211),
.B2(n_207),
.Y(n_276)
);

AND2x4_ASAP7_75t_SL g278 ( 
.A(n_246),
.B(n_245),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_278),
.A2(n_283),
.B(n_287),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_280),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_258),
.A2(n_266),
.B(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_248),
.A2(n_191),
.B1(n_198),
.B2(n_174),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_176),
.B1(n_185),
.B2(n_207),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_247),
.A2(n_236),
.B1(n_213),
.B2(n_214),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_286),
.A2(n_298),
.B1(n_255),
.B2(n_241),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_240),
.B(n_204),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_294),
.C(n_289),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_270),
.A2(n_236),
.B1(n_218),
.B2(n_232),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_273),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_209),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_263),
.A2(n_253),
.B(n_265),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_295),
.A2(n_277),
.B(n_239),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_296),
.A2(n_299),
.B1(n_305),
.B2(n_306),
.Y(n_333)
);

AOI22x1_ASAP7_75t_SL g298 ( 
.A1(n_241),
.A2(n_186),
.B1(n_145),
.B2(n_131),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_249),
.A2(n_232),
.B1(n_218),
.B2(n_234),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_303),
.B(n_250),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_268),
.A2(n_217),
.B1(n_238),
.B2(n_100),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_242),
.A2(n_217),
.B1(n_104),
.B2(n_147),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_300),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_307),
.B(n_311),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_308),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_306),
.Y(n_347)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_313),
.B(n_325),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_281),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_327),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_289),
.B(n_260),
.C(n_259),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_321),
.C(n_292),
.Y(n_343)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_320),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_279),
.B(n_244),
.C(n_239),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_322),
.Y(n_340)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_323),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_324),
.B(n_334),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_290),
.B(n_256),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_269),
.Y(n_326)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_326),
.Y(n_365)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_261),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_328),
.B(n_329),
.Y(n_366)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_300),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_277),
.B(n_267),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_330),
.B(n_331),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_283),
.B(n_295),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_271),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_332),
.B(n_23),
.Y(n_363)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_301),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_296),
.A2(n_241),
.B1(n_251),
.B2(n_243),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_335),
.A2(n_336),
.B1(n_293),
.B2(n_272),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_287),
.A2(n_262),
.B1(n_252),
.B2(n_104),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_301),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_337),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_294),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_341),
.B(n_347),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_343),
.B(n_346),
.C(n_349),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_316),
.A2(n_278),
.B1(n_276),
.B2(n_305),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_344),
.A2(n_354),
.B1(n_335),
.B2(n_333),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_317),
.B(n_280),
.C(n_278),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_321),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_309),
.B(n_304),
.C(n_288),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_352),
.B(n_360),
.C(n_362),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_316),
.A2(n_299),
.B1(n_274),
.B2(n_288),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_325),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_357),
.B(n_323),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_318),
.A2(n_320),
.B(n_337),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_358),
.A2(n_336),
.B(n_318),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_291),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_361),
.A2(n_356),
.B1(n_355),
.B2(n_362),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_315),
.B(n_145),
.C(n_147),
.Y(n_362)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_363),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_329),
.B(n_193),
.C(n_272),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_364),
.B(n_308),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_327),
.Y(n_367)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_365),
.A2(n_307),
.B1(n_324),
.B2(n_334),
.Y(n_368)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_368),
.Y(n_397)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_358),
.Y(n_369)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_369),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_319),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_370),
.B(n_374),
.Y(n_403)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_338),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_372),
.Y(n_396)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_338),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_364),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_375),
.B(n_376),
.Y(n_399)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_339),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_359),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_377),
.B(n_386),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_378),
.A2(n_347),
.B(n_341),
.Y(n_398)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_350),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_379),
.B(n_384),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_380),
.A2(n_390),
.B1(n_345),
.B2(n_356),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_381),
.A2(n_388),
.B1(n_39),
.B2(n_21),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_351),
.A2(n_308),
.B1(n_313),
.B2(n_333),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_382),
.A2(n_43),
.B1(n_37),
.B2(n_30),
.Y(n_405)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_346),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_344),
.A2(n_345),
.B1(n_354),
.B2(n_353),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_345),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_389),
.B(n_271),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_373),
.B(n_349),
.C(n_352),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_392),
.B(n_407),
.C(n_383),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_393),
.B(n_406),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_369),
.A2(n_361),
.B(n_343),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_395),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_400),
.B(n_378),
.Y(n_422)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_404),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_405),
.A2(n_409),
.B1(n_372),
.B2(n_371),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_391),
.B(n_30),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_373),
.B(n_23),
.C(n_22),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_384),
.A2(n_22),
.B1(n_21),
.B2(n_13),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_410),
.A2(n_390),
.B1(n_379),
.B2(n_376),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_383),
.B(n_39),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_411),
.B(n_391),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_385),
.Y(n_412)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_428),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_422),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_375),
.C(n_380),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_417),
.B(n_425),
.C(n_426),
.Y(n_431)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_408),
.Y(n_418)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_418),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_419),
.A2(n_393),
.B1(n_394),
.B2(n_402),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_398),
.A2(n_367),
.B(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_420),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_423),
.Y(n_442)
);

INVx13_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_424),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_388),
.C(n_381),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_11),
.C(n_10),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_10),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_397),
.C(n_411),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_440),
.C(n_5),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_435),
.B(n_439),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_421),
.A2(n_396),
.B1(n_403),
.B2(n_410),
.Y(n_436)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_436),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_413),
.A2(n_408),
.B1(n_406),
.B2(n_396),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_437),
.A2(n_427),
.B1(n_426),
.B2(n_416),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_419),
.A2(n_407),
.B1(n_3),
.B2(n_4),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_2),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_427),
.A2(n_2),
.B(n_3),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_443),
.B(n_424),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_430),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_445),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_415),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_448),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_417),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_454),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_413),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_452),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_441),
.A2(n_2),
.B(n_4),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_453),
.B(n_440),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_438),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_434),
.A2(n_5),
.B(n_6),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_455),
.A2(n_443),
.B(n_439),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_429),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_459),
.A2(n_437),
.B(n_6),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_460),
.B(n_461),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_433),
.C(n_429),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_435),
.Y(n_463)
);

AOI32xp33_ASAP7_75t_L g465 ( 
.A1(n_463),
.A2(n_457),
.A3(n_462),
.B1(n_450),
.B2(n_442),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_464),
.B(n_448),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_465),
.A2(n_468),
.B(n_457),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_467),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_5),
.C(n_6),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_469),
.A2(n_458),
.B(n_8),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_SL g474 ( 
.A(n_470),
.B(n_472),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_471),
.B(n_469),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_473),
.A2(n_474),
.B(n_466),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_475),
.B(n_7),
.Y(n_476)
);

AO21x1_ASAP7_75t_L g477 ( 
.A1(n_476),
.A2(n_7),
.B(n_9),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g478 ( 
.A(n_477),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_478),
.B(n_9),
.Y(n_479)
);


endmodule