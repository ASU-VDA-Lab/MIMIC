module fake_netlist_5_960_n_24 (n_8, n_4, n_5, n_7, n_0, n_9, n_2, n_3, n_6, n_1, n_24);

input n_8;
input n_4;
input n_5;
input n_7;
input n_0;
input n_9;
input n_2;
input n_3;
input n_6;
input n_1;

output n_24;

wire n_16;
wire n_12;
wire n_18;
wire n_22;
wire n_10;
wire n_21;
wire n_11;
wire n_17;
wire n_19;
wire n_15;
wire n_14;
wire n_23;
wire n_13;
wire n_20;

INVx4_ASAP7_75t_SL g10 ( 
.A(n_6),
.Y(n_10)
);

AND2x4_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_3),
.B(n_0),
.Y(n_12)
);

OR2x6_ASAP7_75t_L g13 ( 
.A(n_1),
.B(n_3),
.Y(n_13)
);

BUFx6f_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

AO21x2_ASAP7_75t_L g16 ( 
.A1(n_12),
.A2(n_1),
.B(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_17),
.B(n_11),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_11),
.B(n_12),
.C(n_15),
.Y(n_19)
);

NAND3xp33_ASAP7_75t_L g20 ( 
.A(n_19),
.B(n_13),
.C(n_14),
.Y(n_20)
);

AOI222xp33_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.C1(n_16),
.C2(n_4),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_8),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_21),
.B(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g24 ( 
.A1(n_23),
.A2(n_9),
.B1(n_10),
.B2(n_22),
.Y(n_24)
);


endmodule