module fake_jpeg_1002_n_100 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_24),
.B(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_3),
.Y(n_27)
);

INVxp33_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_11),
.B(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_30),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_7),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_31),
.B(n_17),
.Y(n_38)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_14),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_38),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_16),
.B1(n_12),
.B2(n_17),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_14),
.B1(n_21),
.B2(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_12),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_12),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_11),
.Y(n_52)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_47),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_32),
.B(n_16),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_56),
.C(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2x1_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_21),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_44),
.B(n_41),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_43),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_20),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_46),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_34),
.B1(n_43),
.B2(n_41),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g75 ( 
.A1(n_63),
.A2(n_53),
.B(n_49),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_50),
.B(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_66),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_76),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_56),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_73),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_67),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_65),
.B1(n_54),
.B2(n_55),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_77),
.B(n_62),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_78),
.A2(n_13),
.B1(n_15),
.B2(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_80),
.B(n_82),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_67),
.C(n_63),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_71),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_70),
.B1(n_59),
.B2(n_58),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_78),
.A2(n_75),
.B1(n_69),
.B2(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_86),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_88),
.C(n_79),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

AOI321xp33_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_45),
.A3(n_9),
.B1(n_10),
.B2(n_15),
.C(n_13),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_94),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_85),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_93),
.B(n_88),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_95),
.A2(n_13),
.B(n_15),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

OAI321xp33_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_0),
.A3(n_1),
.B1(n_15),
.B2(n_96),
.C(n_78),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_0),
.Y(n_100)
);


endmodule