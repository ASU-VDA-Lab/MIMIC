module real_jpeg_18961_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_556;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_78;
wire n_83;
wire n_288;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_487;
wire n_93;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_602;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_0),
.A2(n_21),
.B(n_642),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_0),
.B(n_643),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_1),
.Y(n_243)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_1),
.Y(n_411)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_2),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_4),
.A2(n_182),
.B1(n_184),
.B2(n_186),
.Y(n_181)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_4),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_4),
.A2(n_186),
.B1(n_310),
.B2(n_314),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_4),
.A2(n_186),
.B1(n_330),
.B2(n_333),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_4),
.A2(n_186),
.B1(n_377),
.B2(n_382),
.Y(n_376)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_5),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g143 ( 
.A(n_5),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_5),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_208),
.B1(n_213),
.B2(n_214),
.Y(n_207)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_6),
.A2(n_213),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_6),
.A2(n_213),
.B1(n_491),
.B2(n_494),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_6),
.A2(n_213),
.B1(n_487),
.B2(n_589),
.Y(n_588)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_7),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_7),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_7),
.A2(n_215),
.B1(n_269),
.B2(n_370),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_7),
.A2(n_269),
.B1(n_483),
.B2(n_487),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_7),
.A2(n_269),
.B1(n_505),
.B2(n_549),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_8),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_8),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_8),
.A2(n_222),
.B1(n_355),
.B2(n_358),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_8),
.A2(n_222),
.B1(n_417),
.B2(n_419),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_8),
.A2(n_222),
.B1(n_500),
.B2(n_505),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_9),
.A2(n_59),
.B1(n_61),
.B2(n_62),
.Y(n_58)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_9),
.A2(n_62),
.B1(n_106),
.B2(n_110),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_9),
.A2(n_62),
.B1(n_158),
.B2(n_162),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_9),
.A2(n_62),
.B1(n_244),
.B2(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_10),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g141 ( 
.A(n_10),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g246 ( 
.A(n_10),
.Y(n_246)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_10),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_11),
.A2(n_126),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_11),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_11),
.A2(n_271),
.B1(n_343),
.B2(n_345),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_11),
.A2(n_271),
.B1(n_514),
.B2(n_518),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_11),
.A2(n_271),
.B1(n_525),
.B2(n_527),
.Y(n_524)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_12),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_12),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_12),
.A2(n_125),
.B1(n_192),
.B2(n_194),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_12),
.A2(n_125),
.B1(n_257),
.B2(n_261),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_12),
.A2(n_125),
.B1(n_279),
.B2(n_283),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_13),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_13),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_52),
.B2(n_56),
.Y(n_46)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_56),
.B1(n_68),
.B2(n_73),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_14),
.A2(n_56),
.B1(n_292),
.B2(n_294),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_14),
.A2(n_56),
.B1(n_399),
.B2(n_402),
.Y(n_398)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_15),
.Y(n_104)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_15),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_15),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_15),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g486 ( 
.A(n_15),
.Y(n_486)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_16),
.A2(n_116),
.B1(n_119),
.B2(n_121),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_16),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_16),
.A2(n_121),
.B1(n_249),
.B2(n_251),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_16),
.A2(n_121),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g421 ( 
.A1(n_16),
.A2(n_121),
.B1(n_422),
.B2(n_426),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_17),
.B(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_17),
.A2(n_237),
.B(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_17),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_17),
.B(n_167),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_17),
.A2(n_241),
.B1(n_548),
.B2(n_551),
.Y(n_547)
);

OAI32xp33_ASAP7_75t_L g565 ( 
.A1(n_17),
.A2(n_280),
.A3(n_566),
.B1(n_570),
.B2(n_572),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_17),
.A2(n_389),
.B1(n_581),
.B2(n_583),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g239 ( 
.A(n_19),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_171),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_169),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_63),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_24),
.B(n_63),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_46),
.B1(n_57),
.B2(n_58),
.Y(n_24)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_25),
.A2(n_46),
.B1(n_57),
.B2(n_165),
.Y(n_164)
);

OAI22x1_ASAP7_75t_L g180 ( 
.A1(n_25),
.A2(n_57),
.B1(n_115),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_25),
.A2(n_57),
.B1(n_265),
.B2(n_270),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_25),
.A2(n_57),
.B1(n_270),
.B2(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_25),
.A2(n_57),
.B1(n_265),
.B2(n_349),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_25),
.A2(n_57),
.B1(n_321),
.B2(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_25),
.A2(n_57),
.B1(n_181),
.B2(n_416),
.Y(n_449)
);

AO21x2_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B(n_39),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_30),
.Y(n_326)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_32),
.A2(n_208),
.B1(n_229),
.B2(n_236),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_34),
.Y(n_183)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_34),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_38),
.Y(n_233)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_39),
.A2(n_114),
.B1(n_122),
.B2(n_123),
.Y(n_113)
);

AO22x2_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_41),
.Y(n_217)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_42),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_42),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_51),
.Y(n_185)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_55),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_55),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_55),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_57),
.B(n_389),
.Y(n_388)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g351 ( 
.A(n_60),
.Y(n_351)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_61),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_164),
.C(n_166),
.Y(n_63)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_64),
.B(n_164),
.CI(n_166),
.CON(n_174),
.SN(n_174)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_113),
.C(n_128),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_65),
.A2(n_66),
.B1(n_128),
.B2(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI22x1_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_78),
.B1(n_105),
.B2(n_112),
.Y(n_66)
);

OAI22x1_ASAP7_75t_L g190 ( 
.A1(n_67),
.A2(n_78),
.B1(n_112),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_69),
.Y(n_585)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_71),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_71),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

BUFx5_ASAP7_75t_L g212 ( 
.A(n_72),
.Y(n_212)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_77),
.Y(n_221)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_77),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_78),
.A2(n_112),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_78),
.A2(n_112),
.B1(n_342),
.B2(n_347),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_78),
.A2(n_112),
.B1(n_342),
.B2(n_369),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_78),
.A2(n_112),
.B1(n_328),
.B2(n_329),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_78),
.A2(n_112),
.B1(n_329),
.B2(n_421),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_R g435 ( 
.A1(n_78),
.A2(n_112),
.B1(n_329),
.B2(n_421),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_78),
.A2(n_112),
.B1(n_369),
.B2(n_580),
.Y(n_579)
);

INVx3_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_79),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_79),
.A2(n_167),
.B1(n_207),
.B2(n_218),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_79),
.A2(n_167),
.B1(n_439),
.B2(n_440),
.Y(n_438)
);

OA21x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_88),
.B(n_95),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_85),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_85),
.Y(n_344)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_87),
.Y(n_569)
);

INVxp33_ASAP7_75t_L g572 ( 
.A(n_88),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_96),
.B1(n_99),
.B2(n_102),
.Y(n_95)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_93),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_94),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_101),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_102),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g589 ( 
.A(n_102),
.Y(n_589)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g161 ( 
.A(n_104),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

BUFx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g582 ( 
.A(n_108),
.Y(n_582)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_109),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_128),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_128),
.B(n_189),
.C(n_190),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_128),
.B(n_190),
.Y(n_625)
);

OA21x2_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_144),
.B(n_157),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_129),
.B(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_129),
.A2(n_144),
.B1(n_285),
.B2(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_129),
.A2(n_144),
.B1(n_157),
.B2(n_442),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_129),
.A2(n_144),
.B1(n_478),
.B2(n_482),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_129),
.A2(n_144),
.B1(n_482),
.B2(n_513),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_129),
.A2(n_144),
.B1(n_513),
.B2(n_588),
.Y(n_587)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_130),
.A2(n_353),
.B1(n_354),
.B2(n_359),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_130),
.A2(n_278),
.B1(n_353),
.B2(n_398),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_130),
.B(n_389),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g601 ( 
.A1(n_130),
.A2(n_353),
.B1(n_354),
.B2(n_602),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_131),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_135),
.B1(n_139),
.B2(n_142),
.Y(n_131)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_134),
.Y(n_474)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_137),
.Y(n_254)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_137),
.Y(n_293)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_138),
.Y(n_304)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_140),
.Y(n_462)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_141),
.Y(n_295)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_141),
.Y(n_504)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_141),
.Y(n_526)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_144),
.B(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_144),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_150),
.B1(n_153),
.B2(n_155),
.Y(n_145)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_146),
.Y(n_286)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_149),
.Y(n_316)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_149),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_149),
.Y(n_517)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_154),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_156),
.Y(n_313)
);

BUFx12f_ASAP7_75t_L g481 ( 
.A(n_156),
.Y(n_481)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_160),
.Y(n_461)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_162),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_163),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_199),
.B(n_640),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_174),
.B(n_175),
.Y(n_641)
);

BUFx24_ASAP7_75t_SL g644 ( 
.A(n_174),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_180),
.C(n_187),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_177),
.A2(n_180),
.B1(n_189),
.B2(n_622),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_177),
.Y(n_622)
);

INVxp67_ASAP7_75t_SL g189 ( 
.A(n_180),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_180),
.A2(n_189),
.B1(n_625),
.B2(n_626),
.Y(n_624)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_188),
.B(n_621),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_191),
.Y(n_440)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_192),
.Y(n_333)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_616),
.B(n_636),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_453),
.B(n_611),
.Y(n_200)
);

NAND3xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_390),
.C(n_432),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_334),
.B(n_360),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_203),
.B(n_334),
.C(n_613),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_273),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_204),
.B(n_274),
.C(n_305),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_227),
.C(n_263),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_206),
.A2(n_263),
.B1(n_264),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_206),
.Y(n_337)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_207),
.Y(n_347)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_212),
.Y(n_235)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_218),
.Y(n_328)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_225),
.Y(n_427)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_227),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_240),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_228),
.B(n_240),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_238),
.Y(n_272)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_247),
.B1(n_255),
.B2(n_256),
.Y(n_240)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_241),
.A2(n_256),
.B1(n_291),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_241),
.A2(n_302),
.B(n_406),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_241),
.A2(n_255),
.B1(n_490),
.B2(n_498),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_241),
.A2(n_524),
.B1(n_548),
.B2(n_556),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_242),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_243),
.Y(n_300)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_246),
.Y(n_384)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_246),
.Y(n_475)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_246),
.Y(n_493)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_246),
.Y(n_497)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_246),
.Y(n_529)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_246),
.Y(n_545)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_248),
.A2(n_296),
.B1(n_376),
.B2(n_385),
.Y(n_375)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_255),
.Y(n_574)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_259),
.Y(n_508)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_259),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_260),
.Y(n_381)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_305),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_289),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_284),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_276),
.A2(n_284),
.B(n_289),
.Y(n_428)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_282),
.Y(n_401)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_296),
.B1(n_297),
.B2(n_301),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_296),
.A2(n_523),
.B1(n_530),
.B2(n_534),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g573 ( 
.A1(n_296),
.A2(n_376),
.B1(n_499),
.B2(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_297),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_300),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_319),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_306),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_317),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_307),
.A2(n_308),
.B1(n_317),
.B2(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_327),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_320),
.B(n_393),
.C(n_394),
.Y(n_392)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_338),
.C(n_340),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g361 ( 
.A(n_335),
.B(n_362),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_340),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_348),
.C(n_352),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_341),
.B(n_352),
.Y(n_365)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_348),
.B(n_365),
.Y(n_364)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_361),
.B(n_363),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.C(n_367),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_364),
.B(n_608),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_366),
.B(n_367),
.Y(n_608)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_374),
.C(n_388),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_SL g595 ( 
.A(n_368),
.B(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_374),
.A2(n_375),
.B1(n_388),
.B2(n_597),
.Y(n_596)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_388),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_389),
.B(n_467),
.Y(n_466)
);

OAI21xp33_ASAP7_75t_SL g478 ( 
.A1(n_389),
.A2(n_466),
.B(n_479),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_389),
.B(n_531),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_389),
.B(n_571),
.Y(n_570)
);

A2O1A1O1Ixp25_ASAP7_75t_L g611 ( 
.A1(n_390),
.A2(n_432),
.B(n_612),
.C(n_614),
.D(n_615),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_431),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_SL g614 ( 
.A(n_391),
.B(n_431),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_392),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_396),
.A2(n_413),
.B1(n_429),
.B2(n_430),
.Y(n_395)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_396),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_396),
.B(n_429),
.C(n_452),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_397),
.A2(n_404),
.B1(n_405),
.B2(n_412),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_397),
.B(n_405),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_398),
.Y(n_442)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_402),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_404),
.A2(n_405),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_404),
.A2(n_449),
.B(n_450),
.Y(n_628)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_411),
.Y(n_533)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_413),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_428),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_420),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_415),
.B(n_428),
.C(n_435),
.Y(n_434)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_421),
.Y(n_439)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_451),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_433),
.B(n_451),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_436),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_434),
.B(n_631),
.C(n_632),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_444),
.Y(n_436)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_437),
.Y(n_632)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_441),
.B(n_443),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_438),
.B(n_441),
.Y(n_443)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_443),
.Y(n_627)
);

AOI22xp5_ASAP7_75t_L g634 ( 
.A1(n_443),
.A2(n_624),
.B1(n_627),
.B2(n_635),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g631 ( 
.A(n_444),
.Y(n_631)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_445),
.A2(n_446),
.B1(n_447),
.B2(n_450),
.Y(n_444)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_445),
.Y(n_450)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

AOI21x1_ASAP7_75t_L g453 ( 
.A1(n_454),
.A2(n_606),
.B(n_610),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_591),
.B(n_605),
.Y(n_454)
);

AOI21x1_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_561),
.B(n_590),
.Y(n_455)
);

OAI21x1_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_520),
.B(n_560),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_488),
.Y(n_457)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_458),
.B(n_488),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_476),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_459),
.A2(n_476),
.B1(n_477),
.B2(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_459),
.Y(n_536)
);

OAI32xp33_ASAP7_75t_L g459 ( 
.A1(n_460),
.A2(n_462),
.A3(n_463),
.B1(n_466),
.B2(n_470),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_475),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_481),
.Y(n_571)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_483),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_509),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_489),
.B(n_511),
.C(n_519),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_490),
.Y(n_534)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_508),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_510),
.A2(n_511),
.B1(n_512),
.B2(n_519),
.Y(n_509)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_510),
.Y(n_519)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_521),
.A2(n_537),
.B(n_559),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_535),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_522),
.B(n_535),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx6_ASAP7_75t_L g556 ( 
.A(n_533),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_538),
.A2(n_554),
.B(n_558),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_547),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_546),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_557),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_555),
.B(n_557),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_562),
.B(n_563),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_SL g590 ( 
.A(n_562),
.B(n_563),
.Y(n_590)
);

XOR2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_577),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_564),
.B(n_578),
.C(n_587),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_565),
.A2(n_573),
.B1(n_575),
.B2(n_576),
.Y(n_564)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_565),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_565),
.B(n_576),
.Y(n_600)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_567),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_573),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_578),
.A2(n_579),
.B1(n_586),
.B2(n_587),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_588),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_593),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_592),
.B(n_593),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_594),
.A2(n_595),
.B1(n_598),
.B2(n_599),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g609 ( 
.A(n_594),
.B(n_601),
.C(n_603),
.Y(n_609)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_600),
.A2(n_601),
.B1(n_603),
.B2(n_604),
.Y(n_599)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_600),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_601),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_607),
.B(n_609),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_607),
.B(n_609),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_629),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_619),
.A2(n_638),
.B(n_639),
.Y(n_637)
);

NOR2xp67_ASAP7_75t_SL g619 ( 
.A(n_620),
.B(n_623),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_620),
.B(n_623),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_627),
.C(n_628),
.Y(n_623)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_624),
.Y(n_635)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_625),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g633 ( 
.A(n_628),
.B(n_634),
.Y(n_633)
);

OR2x2_ASAP7_75t_L g629 ( 
.A(n_630),
.B(n_633),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_630),
.B(n_633),
.Y(n_638)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);


endmodule