module real_jpeg_11203_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_205;
wire n_110;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_244;
wire n_179;
wire n_213;
wire n_202;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_206;
wire n_127;
wire n_53;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx24_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_1),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_1),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_1),
.A2(n_54),
.B1(n_56),
.B2(n_73),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_1),
.A2(n_28),
.B1(n_32),
.B2(n_73),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_73),
.Y(n_220)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_66),
.B1(n_72),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_54),
.B1(n_56),
.B2(n_77),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_77),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_77),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_4),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_4),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_4),
.A2(n_206),
.B(n_230),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_7),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_7),
.A2(n_33),
.B1(n_38),
.B2(n_39),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_9),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_55),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_9),
.A2(n_28),
.B1(n_32),
.B2(n_55),
.Y(n_164)
);

BUFx6f_ASAP7_75t_SL g59 ( 
.A(n_10),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_11),
.A2(n_66),
.B1(n_72),
.B2(n_94),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_11),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_11),
.A2(n_54),
.B1(n_56),
.B2(n_94),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_11),
.A2(n_38),
.B1(n_39),
.B2(n_94),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_11),
.A2(n_28),
.B1(n_32),
.B2(n_94),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_13),
.A2(n_40),
.B1(n_54),
.B2(n_56),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_28),
.B1(n_32),
.B2(n_40),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_15),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_28),
.B1(n_32),
.B2(n_48),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_16),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_16),
.A2(n_54),
.B(n_68),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_16),
.A2(n_66),
.B1(n_72),
.B2(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_16),
.B(n_75),
.Y(n_161)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_16),
.A2(n_38),
.B(n_42),
.C(n_174),
.D(n_175),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_16),
.B(n_38),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_16),
.B(n_61),
.Y(n_183)
);

OAI21xp33_ASAP7_75t_L g208 ( 
.A1(n_16),
.A2(n_26),
.B(n_189),
.Y(n_208)
);

A2O1A1O1Ixp25_ASAP7_75t_L g221 ( 
.A1(n_16),
.A2(n_56),
.B(n_57),
.C(n_124),
.D(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_16),
.B(n_56),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_20),
.B(n_102),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_78),
.B2(n_79),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_25),
.B(n_36),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_34),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_26),
.A2(n_27),
.B(n_34),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_26),
.A2(n_27),
.B1(n_88),
.B2(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_26),
.A2(n_27),
.B1(n_118),
.B2(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_26),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_26),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_26),
.B(n_191),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_28),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_27),
.A2(n_196),
.B(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_27),
.B(n_115),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_28),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_28),
.A2(n_45),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_32),
.B(n_43),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_32),
.B(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_90),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_39),
.B1(n_58),
.B2(n_59),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_38),
.A2(n_222),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_39),
.B(n_59),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_41),
.A2(n_49),
.B1(n_186),
.B2(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_41),
.A2(n_220),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_42),
.B(n_137),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_46),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_49),
.A2(n_90),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_49),
.B(n_138),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_49),
.A2(n_136),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_49),
.B(n_115),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_53),
.Y(n_97)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

O2A1O1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_54),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_58),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_56),
.B1(n_67),
.B2(n_68),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_57),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_60),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_61),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_71),
.B(n_74),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_66),
.A2(n_67),
.B(n_69),
.C(n_70),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_66),
.B(n_67),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_66),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_67),
.B(n_115),
.C(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_70),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g109 ( 
.A1(n_70),
.A2(n_93),
.B(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_74),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_84),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_82),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.C(n_95),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_87),
.B(n_89),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_91),
.A2(n_92),
.B1(n_95),
.B2(n_96),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_101),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_98),
.A2(n_121),
.B1(n_122),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_98),
.A2(n_99),
.B(n_144),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.C(n_106),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_103),
.B(n_105),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_106),
.A2(n_107),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_112),
.C(n_119),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_108),
.A2(n_109),
.B1(n_119),
.B2(n_120),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_113),
.A2(n_114),
.B1(n_117),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_117),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B(n_123),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_166),
.Y(n_127)
);

INVxp33_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_150),
.B(n_165),
.Y(n_129)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_130),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_147),
.Y(n_130)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_147),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_133),
.CI(n_145),
.CON(n_131),
.SN(n_131)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_139),
.C(n_142),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_135),
.B1(n_142),
.B2(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_151),
.B(n_152),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.C(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_153),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_155),
.A2(n_157),
.B1(n_158),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_162),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_159),
.A2(n_160),
.B1(n_237),
.B2(n_239),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_161),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_164),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_251),
.C(n_252),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_245),
.B(n_250),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_233),
.B(n_244),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_214),
.B(n_232),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_171),
.A2(n_192),
.B(n_213),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_180),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_172),
.B(n_180),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_173),
.A2(n_176),
.B1(n_177),
.B2(n_200),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_174),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_188),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_201),
.B(n_212),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_194),
.B(n_199),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_207),
.B(n_211),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_203),
.B(n_204),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_215),
.B(n_216),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_225),
.B2(n_231),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_221),
.B1(n_223),
.B2(n_224),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_219),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_221),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_224),
.C(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_225),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_229),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_235),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_240),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_236),
.B(n_241),
.C(n_242),
.Y(n_246)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_237),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_246),
.B(n_247),
.Y(n_250)
);


endmodule