module real_aes_7946_n_239 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_239);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_239;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_766;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_763;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_693;
wire n_496;
wire n_281;
wire n_468;
wire n_755;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_417;
wire n_363;
wire n_754;
wire n_607;
wire n_449;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_733;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_751;
wire n_490;
wire n_261;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_392;
wire n_562;
wire n_288;
wire n_756;
wire n_404;
wire n_598;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_749;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_712;
wire n_266;
wire n_312;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_762;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_554;
wire n_475;
wire n_264;
wire n_668;
CKINVDCx20_ASAP7_75t_R g295 ( .A(n_0), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_1), .A2(n_182), .B1(n_426), .B2(n_526), .Y(n_525) );
XOR2x2_ASAP7_75t_L g348 ( .A(n_2), .B(n_349), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_3), .A2(n_202), .B1(n_439), .B2(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_4), .A2(n_154), .B1(n_360), .B2(n_384), .Y(n_440) );
INVx1_ASAP7_75t_L g433 ( .A(n_5), .Y(n_433) );
AOI222xp33_ASAP7_75t_L g378 ( .A1(n_6), .A2(n_25), .B1(n_192), .B2(n_379), .C1(n_380), .C2(n_383), .Y(n_378) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_7), .A2(n_207), .B1(n_358), .B2(n_359), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_8), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_9), .B(n_355), .Y(n_437) );
INVx1_ASAP7_75t_L g757 ( .A(n_10), .Y(n_757) );
OA22x2_ASAP7_75t_L g761 ( .A1(n_11), .A2(n_733), .B1(n_734), .B2(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_11), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_12), .A2(n_139), .B1(n_307), .B2(n_478), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_13), .A2(n_69), .B1(n_368), .B2(n_370), .Y(n_367) );
AOI22xp33_ASAP7_75t_SL g505 ( .A1(n_14), .A2(n_91), .B1(n_359), .B2(n_384), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_15), .A2(n_58), .B1(n_416), .B2(n_418), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_16), .A2(n_18), .B1(n_616), .B2(n_617), .C(n_619), .Y(n_615) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_17), .A2(n_195), .B1(n_711), .B2(n_712), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g290 ( .A(n_19), .Y(n_290) );
XOR2x2_ASAP7_75t_L g458 ( .A(n_20), .B(n_459), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_21), .A2(n_174), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_22), .A2(n_83), .B1(n_383), .B2(n_570), .Y(n_638) );
AO22x2_ASAP7_75t_L g270 ( .A1(n_23), .A2(n_75), .B1(n_262), .B2(n_267), .Y(n_270) );
INVx1_ASAP7_75t_L g729 ( .A(n_23), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_24), .Y(n_544) );
AOI222xp33_ASAP7_75t_L g511 ( .A1(n_26), .A2(n_90), .B1(n_110), .B2(n_380), .C1(n_393), .C2(n_512), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_27), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_28), .A2(n_138), .B1(n_417), .B2(n_647), .Y(n_679) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_29), .A2(n_31), .B1(n_375), .B2(n_582), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_30), .A2(n_203), .B1(n_257), .B2(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g667 ( .A(n_32), .Y(n_667) );
AOI222xp33_ASAP7_75t_L g688 ( .A1(n_33), .A2(n_81), .B1(n_219), .B2(n_382), .C1(n_432), .C2(n_572), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_34), .Y(n_542) );
AOI22xp33_ASAP7_75t_SL g701 ( .A1(n_35), .A2(n_59), .B1(n_408), .B2(n_702), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_36), .A2(n_37), .B1(n_352), .B2(n_355), .Y(n_351) );
INVx1_ASAP7_75t_L g755 ( .A(n_38), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_39), .A2(n_141), .B1(n_495), .B2(n_496), .Y(n_494) );
AO22x2_ASAP7_75t_L g272 ( .A1(n_40), .A2(n_78), .B1(n_262), .B2(n_263), .Y(n_272) );
INVx1_ASAP7_75t_L g730 ( .A(n_40), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_41), .A2(n_116), .B1(n_451), .B2(n_453), .Y(n_450) );
AOI22xp33_ASAP7_75t_SL g644 ( .A1(n_42), .A2(n_45), .B1(n_307), .B2(n_479), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g640 ( .A1(n_43), .A2(n_102), .B1(n_257), .B2(n_368), .Y(n_640) );
INVx1_ASAP7_75t_L g749 ( .A(n_44), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g606 ( .A1(n_46), .A2(n_237), .B1(n_482), .B2(n_607), .C(n_608), .Y(n_606) );
INVx1_ASAP7_75t_L g743 ( .A(n_47), .Y(n_743) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_48), .A2(n_229), .B1(n_380), .B2(n_512), .Y(n_634) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_49), .Y(n_327) );
INVx1_ASAP7_75t_L g748 ( .A(n_50), .Y(n_748) );
AOI22xp33_ASAP7_75t_SL g581 ( .A1(n_51), .A2(n_128), .B1(n_526), .B2(n_582), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_52), .B(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_53), .A2(n_204), .B1(n_489), .B2(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g620 ( .A(n_54), .Y(n_620) );
AOI22xp33_ASAP7_75t_SL g641 ( .A1(n_55), .A2(n_173), .B1(n_418), .B2(n_642), .Y(n_641) );
XOR2x2_ASAP7_75t_L g628 ( .A(n_56), .B(n_629), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_57), .A2(n_184), .B1(n_279), .B2(n_285), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_60), .B(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_SL g434 ( .A1(n_61), .A2(n_227), .B1(n_382), .B2(n_435), .Y(n_434) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_62), .A2(n_180), .B1(n_279), .B2(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_63), .B(n_439), .Y(n_438) );
OA22x2_ASAP7_75t_L g561 ( .A1(n_64), .A2(n_562), .B1(n_563), .B2(n_586), .Y(n_561) );
CKINVDCx20_ASAP7_75t_R g562 ( .A(n_64), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_65), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_66), .B(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_67), .A2(n_145), .B1(n_413), .B2(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g347 ( .A(n_68), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_70), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g599 ( .A(n_71), .Y(n_599) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_72), .A2(n_101), .B1(n_302), .B2(n_411), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g703 ( .A1(n_73), .A2(n_223), .B1(n_439), .B2(n_704), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_74), .A2(n_230), .B1(n_356), .B2(n_471), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_76), .A2(n_80), .B1(n_384), .B2(n_751), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_77), .A2(n_196), .B1(n_570), .B2(n_572), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_79), .A2(n_225), .B1(n_302), .B2(n_447), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g603 ( .A(n_82), .Y(n_603) );
INVx1_ASAP7_75t_L g246 ( .A(n_84), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_85), .A2(n_112), .B1(n_257), .B2(n_273), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_86), .B(n_470), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_87), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_88), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g243 ( .A(n_89), .Y(n_243) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_92), .A2(n_228), .B1(n_273), .B2(n_686), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_93), .A2(n_130), .B1(n_292), .B2(n_374), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_94), .A2(n_205), .B1(n_364), .B2(n_366), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_95), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_96), .A2(n_167), .B1(n_413), .B2(n_478), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_97), .A2(n_153), .B1(n_275), .B2(n_377), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_98), .A2(n_103), .B1(n_364), .B2(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g669 ( .A(n_99), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g612 ( .A(n_100), .Y(n_612) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_104), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g357 ( .A1(n_105), .A2(n_113), .B1(n_358), .B2(n_359), .Y(n_357) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_106), .A2(n_190), .B1(n_510), .B2(n_523), .Y(n_576) );
INVx1_ASAP7_75t_L g663 ( .A(n_107), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g312 ( .A(n_108), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_109), .A2(n_157), .B1(n_579), .B2(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_111), .A2(n_183), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_114), .A2(n_234), .B1(n_374), .B2(n_375), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_115), .Y(n_604) );
INVx1_ASAP7_75t_L g736 ( .A(n_117), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_118), .A2(n_121), .B1(n_616), .B2(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g665 ( .A(n_119), .Y(n_665) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_120), .A2(n_217), .B1(n_532), .B2(n_579), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_122), .Y(n_696) );
AOI222xp33_ASAP7_75t_L g670 ( .A1(n_123), .A2(n_159), .B1(n_163), .B2(n_326), .C1(n_358), .C2(n_399), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_124), .B(n_335), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_125), .A2(n_215), .B1(n_335), .B2(n_407), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_126), .A2(n_171), .B1(n_481), .B2(n_482), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_127), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_129), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g424 ( .A1(n_131), .A2(n_162), .B1(n_425), .B2(n_426), .Y(n_424) );
INVx2_ASAP7_75t_L g247 ( .A(n_132), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_133), .A2(n_208), .B1(n_329), .B2(n_465), .Y(n_464) );
AO22x1_ASAP7_75t_L g588 ( .A1(n_134), .A2(n_589), .B1(n_624), .B2(n_625), .Y(n_588) );
INVx1_ASAP7_75t_L g624 ( .A(n_134), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g594 ( .A(n_135), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_136), .A2(n_238), .B1(n_435), .B2(n_546), .Y(n_567) );
AOI22xp33_ASAP7_75t_SL g583 ( .A1(n_137), .A2(n_143), .B1(n_481), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_140), .A2(n_220), .B1(n_498), .B2(n_499), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_142), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g484 ( .A1(n_144), .A2(n_191), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI22xp33_ASAP7_75t_SL g577 ( .A1(n_146), .A2(n_235), .B1(n_578), .B2(n_579), .Y(n_577) );
AND2x6_ASAP7_75t_L g242 ( .A(n_147), .B(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_147), .Y(n_723) );
AO22x2_ASAP7_75t_L g261 ( .A1(n_148), .A2(n_200), .B1(n_262), .B2(n_263), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g655 ( .A1(n_149), .A2(n_226), .B1(n_486), .B2(n_490), .Y(n_655) );
AOI22xp33_ASAP7_75t_SL g395 ( .A1(n_150), .A2(n_178), .B1(n_396), .B2(n_399), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_151), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_152), .B(n_471), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g420 ( .A1(n_155), .A2(n_236), .B1(n_421), .B2(n_422), .Y(n_420) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_156), .Y(n_343) );
INVx1_ASAP7_75t_L g657 ( .A(n_158), .Y(n_657) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_160), .Y(n_513) );
INVx1_ASAP7_75t_L g671 ( .A(n_161), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g732 ( .A1(n_164), .A2(n_733), .B1(n_734), .B2(n_758), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g758 ( .A(n_164), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_165), .B(n_601), .Y(n_600) );
AO22x2_ASAP7_75t_L g266 ( .A1(n_166), .A2(n_210), .B1(n_262), .B2(n_267), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_168), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g443 ( .A1(n_169), .A2(n_213), .B1(n_444), .B2(n_445), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_170), .B(n_402), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g446 ( .A1(n_172), .A2(n_177), .B1(n_279), .B2(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g622 ( .A(n_175), .Y(n_622) );
INVx1_ASAP7_75t_L g754 ( .A(n_176), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_179), .A2(n_216), .B1(n_570), .B2(n_572), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_181), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_185), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_186), .B(n_659), .Y(n_658) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_187), .Y(n_524) );
INVx1_ASAP7_75t_L g737 ( .A(n_188), .Y(n_737) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_189), .A2(n_232), .B1(n_646), .B2(n_647), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g300 ( .A(n_193), .Y(n_300) );
AOI211xp5_ASAP7_75t_L g239 ( .A1(n_194), .A2(n_240), .B(n_248), .C(n_731), .Y(n_239) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_197), .Y(n_339) );
XOR2x2_ASAP7_75t_L g388 ( .A(n_198), .B(n_389), .Y(n_388) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_199), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_200), .B(n_728), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_201), .Y(n_548) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_206), .Y(n_501) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_209), .Y(n_566) );
INVx1_ASAP7_75t_L g726 ( .A(n_210), .Y(n_726) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_211), .Y(n_609) );
INVx1_ASAP7_75t_L g394 ( .A(n_212), .Y(n_394) );
OA22x2_ASAP7_75t_L g691 ( .A1(n_214), .A2(n_692), .B1(n_693), .B2(n_714), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_214), .Y(n_692) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_218), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_221), .B(n_471), .Y(n_637) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_222), .Y(n_697) );
INVx1_ASAP7_75t_L g262 ( .A(n_224), .Y(n_262) );
INVx1_ASAP7_75t_L g264 ( .A(n_224), .Y(n_264) );
INVx1_ASAP7_75t_L g744 ( .A(n_231), .Y(n_744) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_233), .A2(n_517), .B1(n_553), .B2(n_554), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_233), .Y(n_553) );
INVx2_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_242), .B(n_244), .Y(n_241) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_243), .Y(n_722) );
OA21x2_ASAP7_75t_L g768 ( .A1(n_244), .A2(n_721), .B(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
HB1xp67_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AOI221xp5_ASAP7_75t_L g248 ( .A1(n_249), .A2(n_556), .B1(n_716), .B2(n_717), .C(n_718), .Y(n_248) );
INVx1_ASAP7_75t_L g716 ( .A(n_249), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B1(n_385), .B2(n_555), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
XOR2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_348), .Y(n_251) );
XOR2xp5_ASAP7_75t_SL g252 ( .A(n_253), .B(n_347), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_310), .Y(n_253) );
NOR3xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_289), .C(n_299), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_256), .B(n_278), .Y(n_255) );
BUFx2_ASAP7_75t_SL g257 ( .A(n_258), .Y(n_257) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_258), .Y(n_377) );
INVx2_ASAP7_75t_L g452 ( .A(n_258), .Y(n_452) );
BUFx2_ASAP7_75t_SL g616 ( .A(n_258), .Y(n_616) );
AND2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_268), .Y(n_258) );
AND2x6_ASAP7_75t_L g275 ( .A(n_259), .B(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g294 ( .A(n_259), .B(n_284), .Y(n_294) );
AND2x6_ASAP7_75t_L g326 ( .A(n_259), .B(n_321), .Y(n_326) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_265), .Y(n_259) );
AND2x2_ASAP7_75t_L g304 ( .A(n_260), .B(n_266), .Y(n_304) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g282 ( .A(n_261), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_261), .B(n_266), .Y(n_288) );
AND2x2_ASAP7_75t_L g316 ( .A(n_261), .B(n_270), .Y(n_316) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g267 ( .A(n_264), .Y(n_267) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g283 ( .A(n_266), .Y(n_283) );
INVx1_ASAP7_75t_L g332 ( .A(n_266), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_268), .B(n_282), .Y(n_298) );
AND2x4_ASAP7_75t_L g303 ( .A(n_268), .B(n_304), .Y(n_303) );
AND2x4_ASAP7_75t_L g308 ( .A(n_268), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g365 ( .A(n_268), .B(n_282), .Y(n_365) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
OR2x2_ASAP7_75t_L g277 ( .A(n_269), .B(n_272), .Y(n_277) );
AND2x2_ASAP7_75t_L g284 ( .A(n_269), .B(n_272), .Y(n_284) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g321 ( .A(n_270), .B(n_272), .Y(n_321) );
INVx1_ASAP7_75t_L g317 ( .A(n_271), .Y(n_317) );
AND2x2_ASAP7_75t_L g337 ( .A(n_271), .B(n_332), .Y(n_337) );
INVx2_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g287 ( .A(n_272), .Y(n_287) );
INVx1_ASAP7_75t_L g668 ( .A(n_273), .Y(n_668) );
INVx3_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx4_ASAP7_75t_L g374 ( .A(n_274), .Y(n_374) );
INVx4_ASAP7_75t_L g526 ( .A(n_274), .Y(n_526) );
INVx2_ASAP7_75t_SL g646 ( .A(n_274), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_274), .A2(n_623), .B1(n_743), .B2(n_744), .C(n_745), .Y(n_742) );
INVx11_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx11_ASAP7_75t_L g414 ( .A(n_275), .Y(n_414) );
AND2x4_ASAP7_75t_L g354 ( .A(n_276), .B(n_304), .Y(n_354) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g341 ( .A(n_277), .B(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_279), .Y(n_578) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx5_ASAP7_75t_L g417 ( .A(n_280), .Y(n_417) );
BUFx3_ASAP7_75t_L g487 ( .A(n_280), .Y(n_487) );
INVx3_ASAP7_75t_L g498 ( .A(n_280), .Y(n_498) );
INVx1_ASAP7_75t_L g533 ( .A(n_280), .Y(n_533) );
INVx4_ASAP7_75t_L g741 ( .A(n_280), .Y(n_741) );
INVx8_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_282), .B(n_284), .Y(n_611) );
INVx1_ASAP7_75t_L g323 ( .A(n_283), .Y(n_323) );
NAND2x1p5_ASAP7_75t_L g346 ( .A(n_284), .B(n_304), .Y(n_346) );
AND2x6_ASAP7_75t_L g356 ( .A(n_284), .B(n_304), .Y(n_356) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx6_ASAP7_75t_SL g366 ( .A(n_286), .Y(n_366) );
INVx1_ASAP7_75t_SL g534 ( .A(n_286), .Y(n_534) );
OR2x6_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx1_ASAP7_75t_L g361 ( .A(n_287), .Y(n_361) );
INVx1_ASAP7_75t_L g309 ( .A(n_288), .Y(n_309) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_295), .B2(n_296), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_291), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_666) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g425 ( .A(n_293), .Y(n_425) );
INVx2_ASAP7_75t_L g485 ( .A(n_293), .Y(n_485) );
INVx6_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx3_ASAP7_75t_L g375 ( .A(n_294), .Y(n_375) );
BUFx3_ASAP7_75t_L g510 ( .A(n_294), .Y(n_510) );
BUFx3_ASAP7_75t_L g647 ( .A(n_294), .Y(n_647) );
OAI221xp5_ASAP7_75t_SL g527 ( .A1(n_296), .A2(n_528), .B1(n_529), .B2(n_530), .C(n_531), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_296), .A2(n_663), .B1(n_664), .B2(n_665), .Y(n_662) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_305), .B2(n_306), .Y(n_299) );
INVx4_ASAP7_75t_L g607 ( .A(n_301), .Y(n_607) );
INVx3_ASAP7_75t_L g654 ( .A(n_301), .Y(n_654) );
OAI221xp5_ASAP7_75t_SL g735 ( .A1(n_301), .A2(n_520), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_735) );
INVx4_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
BUFx3_ASAP7_75t_L g453 ( .A(n_303), .Y(n_453) );
BUFx3_ASAP7_75t_L g489 ( .A(n_303), .Y(n_489) );
BUFx3_ASAP7_75t_L g508 ( .A(n_303), .Y(n_508) );
INVx1_ASAP7_75t_L g342 ( .A(n_304), .Y(n_342) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g371 ( .A(n_308), .Y(n_371) );
BUFx2_ASAP7_75t_SL g426 ( .A(n_308), .Y(n_426) );
BUFx2_ASAP7_75t_L g445 ( .A(n_308), .Y(n_445) );
BUFx3_ASAP7_75t_L g482 ( .A(n_308), .Y(n_482) );
BUFx3_ASAP7_75t_L g496 ( .A(n_308), .Y(n_496) );
BUFx3_ASAP7_75t_L g585 ( .A(n_308), .Y(n_585) );
BUFx3_ASAP7_75t_L g686 ( .A(n_308), .Y(n_686) );
AND2x2_ASAP7_75t_L g447 ( .A(n_309), .B(n_317), .Y(n_447) );
NOR3xp33_ASAP7_75t_L g310 ( .A(n_311), .B(n_324), .C(n_338), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B1(n_318), .B2(n_319), .Y(n_311) );
INVx3_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g549 ( .A(n_314), .Y(n_549) );
INVx4_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
AND2x4_ASAP7_75t_L g330 ( .A(n_316), .B(n_331), .Y(n_330) );
AND2x4_ASAP7_75t_L g336 ( .A(n_316), .B(n_337), .Y(n_336) );
AND2x4_ASAP7_75t_L g360 ( .A(n_316), .B(n_361), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g552 ( .A(n_319), .Y(n_552) );
OR2x6_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x4_ASAP7_75t_L g384 ( .A(n_321), .B(n_323), .Y(n_384) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
OAI221xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_327), .B1(n_328), .B2(n_333), .C(n_334), .Y(n_324) );
INVx4_ASAP7_75t_L g393 ( .A(n_325), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g752 ( .A1(n_325), .A2(n_753), .B1(n_754), .B2(n_755), .C1(n_756), .C2(n_757), .Y(n_752) );
INVx4_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
BUFx6f_ASAP7_75t_L g379 ( .A(n_326), .Y(n_379) );
BUFx3_ASAP7_75t_L g432 ( .A(n_326), .Y(n_432) );
INVx2_ASAP7_75t_SL g462 ( .A(n_326), .Y(n_462) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g546 ( .A(n_329), .Y(n_546) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_330), .Y(n_382) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_330), .Y(n_399) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_L g358 ( .A(n_336), .Y(n_358) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_336), .Y(n_398) );
BUFx4f_ASAP7_75t_SL g435 ( .A(n_336), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_343), .B2(n_344), .Y(n_338) );
BUFx3_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVx2_ASAP7_75t_L g539 ( .A(n_341), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_344), .A2(n_537), .B1(n_538), .B2(n_540), .Y(n_536) );
OAI221xp5_ASAP7_75t_L g746 ( .A1(n_344), .A2(n_747), .B1(n_748), .B2(n_749), .C(n_750), .Y(n_746) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_SL g595 ( .A(n_345), .Y(n_595) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g503 ( .A(n_346), .Y(n_503) );
NAND4xp75_ASAP7_75t_L g349 ( .A(n_350), .B(n_362), .C(n_372), .D(n_378), .Y(n_349) );
AND2x2_ASAP7_75t_SL g350 ( .A(n_351), .B(n_357), .Y(n_350) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g405 ( .A(n_353), .Y(n_405) );
INVx2_ASAP7_75t_L g439 ( .A(n_353), .Y(n_439) );
INVx5_ASAP7_75t_L g471 ( .A(n_353), .Y(n_471) );
INVx4_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
BUFx4f_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g403 ( .A(n_356), .Y(n_403) );
BUFx2_ASAP7_75t_L g473 ( .A(n_356), .Y(n_473) );
BUFx2_ASAP7_75t_L g704 ( .A(n_356), .Y(n_704) );
BUFx6f_ASAP7_75t_L g512 ( .A(n_358), .Y(n_512) );
BUFx3_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
BUFx2_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
INVx1_ASAP7_75t_L g571 ( .A(n_360), .Y(n_571) );
BUFx2_ASAP7_75t_L g702 ( .A(n_360), .Y(n_702) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_367), .Y(n_362) );
INVx1_ASAP7_75t_L g423 ( .A(n_364), .Y(n_423) );
BUFx3_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx3_ASAP7_75t_L g444 ( .A(n_365), .Y(n_444) );
BUFx3_ASAP7_75t_L g479 ( .A(n_365), .Y(n_479) );
BUFx3_ASAP7_75t_L g495 ( .A(n_365), .Y(n_495) );
BUFx2_ASAP7_75t_L g418 ( .A(n_366), .Y(n_418) );
BUFx2_ASAP7_75t_L g490 ( .A(n_366), .Y(n_490) );
BUFx2_ASAP7_75t_L g499 ( .A(n_366), .Y(n_499) );
BUFx2_ASAP7_75t_L g579 ( .A(n_366), .Y(n_579) );
BUFx4f_ASAP7_75t_SL g614 ( .A(n_366), .Y(n_614) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_376), .Y(n_372) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_377), .Y(n_421) );
INVx3_ASAP7_75t_L g520 ( .A(n_377), .Y(n_520) );
BUFx3_ASAP7_75t_L g711 ( .A(n_377), .Y(n_711) );
INVx2_ASAP7_75t_SL g632 ( .A(n_379), .Y(n_632) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx4f_ASAP7_75t_SL g601 ( .A(n_382), .Y(n_601) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
BUFx2_ASAP7_75t_SL g408 ( .A(n_384), .Y(n_408) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_384), .Y(n_467) );
BUFx3_ASAP7_75t_L g572 ( .A(n_384), .Y(n_572) );
INVx1_ASAP7_75t_L g555 ( .A(n_385), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_455), .B2(n_456), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
XNOR2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_427), .Y(n_387) );
NAND3x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_409), .C(n_419), .Y(n_389) );
NOR2x1_ASAP7_75t_SL g390 ( .A(n_391), .B(n_400), .Y(n_390) );
OAI21xp5_ASAP7_75t_SL g391 ( .A1(n_392), .A2(n_394), .B(n_395), .Y(n_391) );
OAI222xp33_ASAP7_75t_L g695 ( .A1(n_392), .A2(n_543), .B1(n_696), .B2(n_697), .C1(n_698), .C2(n_699), .Y(n_695) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g753 ( .A(n_396), .Y(n_753) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx4_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g698 ( .A(n_399), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g400 ( .A(n_401), .B(n_404), .C(n_406), .Y(n_400) );
INVx1_ASAP7_75t_SL g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_SL g574 ( .A(n_403), .Y(n_574) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_415), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
BUFx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_417), .Y(n_642) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_424), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g623 ( .A(n_425), .Y(n_623) );
XOR2x2_ASAP7_75t_L g427 ( .A(n_428), .B(n_454), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g428 ( .A(n_429), .B(n_441), .Y(n_428) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_430), .B(n_436), .Y(n_429) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_433), .B(n_434), .Y(n_430) );
OAI21xp5_ASAP7_75t_SL g565 ( .A1(n_431), .A2(n_566), .B(n_567), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g596 ( .A1(n_431), .A2(n_597), .B1(n_598), .B2(n_599), .C(n_600), .Y(n_596) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g543 ( .A(n_435), .Y(n_543) );
NAND3xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .C(n_440), .Y(n_436) );
BUFx2_ASAP7_75t_L g659 ( .A(n_439), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_448), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_446), .Y(n_442) );
INVx1_ASAP7_75t_L g618 ( .A(n_444), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx3_ASAP7_75t_L g481 ( .A(n_452), .Y(n_481) );
INVx1_ASAP7_75t_L g713 ( .A(n_453), .Y(n_713) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_516), .Y(n_456) );
AO22x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_491), .B1(n_514), .B2(n_515), .Y(n_457) );
INVx2_ASAP7_75t_L g514 ( .A(n_458), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_460), .B(n_475), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_468), .Y(n_460) );
OAI21xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_463), .B(n_464), .Y(n_461) );
OAI221xp5_ASAP7_75t_L g541 ( .A1(n_462), .A2(n_542), .B1(n_543), .B2(n_544), .C(n_545), .Y(n_541) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_472), .C(n_474), .Y(n_468) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_476), .B(n_483), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_477), .B(n_480), .Y(n_476) );
BUFx4f_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_488), .Y(n_483) );
INVx3_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx3_ASAP7_75t_SL g515 ( .A(n_491), .Y(n_515) );
XOR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_513), .Y(n_491) );
NAND4xp75_ASAP7_75t_L g492 ( .A(n_493), .B(n_500), .C(n_506), .D(n_511), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_497), .Y(n_493) );
BUFx3_ASAP7_75t_L g582 ( .A(n_495), .Y(n_582) );
INVxp67_ASAP7_75t_L g664 ( .A(n_496), .Y(n_664) );
OA211x2_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B(n_504), .C(n_505), .Y(n_500) );
OA211x2_ASAP7_75t_L g656 ( .A1(n_502), .A2(n_657), .B(n_658), .C(n_660), .Y(n_656) );
BUFx3_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
BUFx2_ASAP7_75t_L g523 ( .A(n_508), .Y(n_523) );
INVx1_ASAP7_75t_L g528 ( .A(n_510), .Y(n_528) );
INVx2_ASAP7_75t_SL g598 ( .A(n_512), .Y(n_598) );
INVx2_ASAP7_75t_L g554 ( .A(n_517), .Y(n_554) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_518), .B(n_535), .Y(n_517) );
NOR2xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_527), .Y(n_518) );
OAI221xp5_ASAP7_75t_SL g519 ( .A1(n_520), .A2(n_521), .B1(n_522), .B2(n_524), .C(n_525), .Y(n_519) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g621 ( .A(n_526), .Y(n_621) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NOR3xp33_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .C(n_547), .Y(n_535) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_SL g593 ( .A(n_539), .Y(n_593) );
INVx2_ASAP7_75t_L g747 ( .A(n_539), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B1(n_550), .B2(n_551), .Y(n_547) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_549), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g605 ( .A(n_552), .Y(n_605) );
INVx1_ASAP7_75t_L g717 ( .A(n_556), .Y(n_717) );
AOI22xp5_ASAP7_75t_SL g556 ( .A1(n_557), .A2(n_558), .B1(n_674), .B2(n_675), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_560), .B1(n_627), .B2(n_673), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_587), .B1(n_588), .B2(n_626), .Y(n_560) );
INVx1_ASAP7_75t_L g626 ( .A(n_561), .Y(n_626) );
INVx1_ASAP7_75t_SL g586 ( .A(n_563), .Y(n_586) );
NAND3x1_ASAP7_75t_L g563 ( .A(n_564), .B(n_575), .C(n_580), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_573), .Y(n_568) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g751 ( .A(n_571), .Y(n_751) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
BUFx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g625 ( .A(n_589), .Y(n_625) );
AND3x1_ASAP7_75t_L g589 ( .A(n_590), .B(n_606), .C(n_615), .Y(n_589) );
NOR3xp33_ASAP7_75t_L g590 ( .A(n_591), .B(n_596), .C(n_602), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B1(n_594), .B2(n_595), .Y(n_591) );
INVx1_ASAP7_75t_L g756 ( .A(n_601), .Y(n_756) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_612), .B2(n_613), .Y(n_608) );
BUFx2_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_619) );
INVx1_ASAP7_75t_L g673 ( .A(n_627), .Y(n_673) );
OAI22xp5_ASAP7_75t_SL g627 ( .A1(n_628), .A2(n_648), .B1(n_649), .B2(n_672), .Y(n_627) );
INVx1_ASAP7_75t_L g672 ( .A(n_628), .Y(n_672) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_639), .C(n_643), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_635), .Y(n_630) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_633), .B(n_634), .Y(n_631) );
NAND3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .C(n_638), .Y(n_635) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
AND2x2_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
XOR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_671), .Y(n_650) );
NAND4xp75_ASAP7_75t_L g651 ( .A(n_652), .B(n_656), .C(n_661), .D(n_670), .Y(n_651) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_666), .Y(n_661) );
CKINVDCx16_ASAP7_75t_R g674 ( .A(n_675), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_690), .B1(n_691), .B2(n_715), .Y(n_675) );
INVx2_ASAP7_75t_SL g715 ( .A(n_676), .Y(n_715) );
XOR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_689), .Y(n_676) );
NAND4xp75_ASAP7_75t_L g677 ( .A(n_678), .B(n_681), .C(n_684), .D(n_688), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
AND2x2_ASAP7_75t_SL g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g714 ( .A(n_693), .Y(n_714) );
NAND3x1_ASAP7_75t_L g693 ( .A(n_694), .B(n_705), .C(n_708), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_700), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
AND2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .Y(n_719) );
OR2x2_ASAP7_75t_SL g765 ( .A(n_720), .B(n_725), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_721), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_722), .B(n_760), .Y(n_769) );
CKINVDCx16_ASAP7_75t_R g760 ( .A(n_723), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_727), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_730), .Y(n_728) );
OAI222xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_759), .B1(n_761), .B2(n_762), .C1(n_763), .C2(n_766), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OR4x1_ASAP7_75t_L g734 ( .A(n_735), .B(n_742), .C(n_746), .D(n_752), .Y(n_734) );
INVx3_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
endmodule