module fake_jpeg_24837_n_265 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_239;
wire n_72;
wire n_107;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_91;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_29),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_44),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_18),
.B(n_0),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_53),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_38),
.B(n_25),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_56),
.C(n_30),
.Y(n_98)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_33),
.C(n_28),
.Y(n_56)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g58 ( 
.A(n_38),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_60),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_82),
.B1(n_83),
.B2(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_64),
.B(n_78),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_46),
.B(n_23),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_66),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_43),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_67),
.B(n_68),
.Y(n_114)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_26),
.B1(n_22),
.B2(n_24),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_69),
.A2(n_21),
.B1(n_30),
.B2(n_27),
.Y(n_93)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_37),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_72),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_23),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_42),
.B(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_75),
.B(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_47),
.B(n_32),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_32),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_81),
.Y(n_91)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_45),
.A2(n_26),
.B1(n_35),
.B2(n_34),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_38),
.A2(n_22),
.B1(n_17),
.B2(n_34),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_46),
.A2(n_17),
.B1(n_35),
.B2(n_31),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_30),
.B1(n_21),
.B2(n_27),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_27),
.B1(n_28),
.B2(n_36),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_90),
.B(n_94),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_93),
.A2(n_106),
.B1(n_113),
.B2(n_2),
.Y(n_137)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_33),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_2),
.Y(n_138)
);

OAI211xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_36),
.B(n_31),
.C(n_20),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_96),
.A2(n_97),
.A3(n_117),
.B1(n_101),
.B2(n_102),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_95),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_100),
.A2(n_86),
.B1(n_59),
.B2(n_84),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_20),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_109),
.Y(n_133)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_105),
.Y(n_126)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_80),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_1),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_80),
.A2(n_19),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_86),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_91),
.A2(n_81),
.B1(n_87),
.B2(n_65),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_119),
.A2(n_121),
.B1(n_123),
.B2(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_130),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_91),
.A2(n_65),
.B1(n_52),
.B2(n_71),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_122),
.B(n_138),
.C(n_147),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_52),
.B1(n_54),
.B2(n_56),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_98),
.B(n_57),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_124),
.A2(n_125),
.B(n_128),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_111),
.A2(n_61),
.B(n_63),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_83),
.B1(n_82),
.B2(n_61),
.Y(n_127)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_127),
.A2(n_142),
.B1(n_90),
.B2(n_8),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_68),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_97),
.A2(n_60),
.B1(n_83),
.B2(n_53),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_134),
.B1(n_125),
.B2(n_89),
.Y(n_170)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_131),
.Y(n_156)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_83),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_136),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_77),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_143),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_103),
.B(n_16),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_141),
.Y(n_159)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_4),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_117),
.B(n_4),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_114),
.B(n_16),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

NOR3xp33_ASAP7_75t_SL g148 ( 
.A(n_112),
.B(n_5),
.C(n_6),
.Y(n_148)
);

INVx13_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_149),
.B(n_153),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_136),
.B(n_101),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_171),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_152),
.B(n_160),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_104),
.C(n_88),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_161),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_104),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_146),
.B1(n_121),
.B2(n_119),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_162),
.A2(n_167),
.B1(n_134),
.B2(n_115),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_108),
.B1(n_115),
.B2(n_90),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_170),
.A2(n_173),
.B1(n_142),
.B2(n_148),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_126),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_122),
.B(n_88),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_122),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_120),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_175),
.B(n_133),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_177),
.B(n_194),
.Y(n_201)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_183),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_182),
.B(n_188),
.Y(n_199)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_167),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_133),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_162),
.A2(n_172),
.B1(n_149),
.B2(n_155),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_186),
.A2(n_197),
.B1(n_170),
.B2(n_173),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_128),
.Y(n_187)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_135),
.B(n_129),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_189),
.B(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_132),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_172),
.B(n_175),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_128),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_193),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_173),
.B(n_124),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_195),
.B(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_166),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_198),
.B(n_205),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_207),
.B1(n_210),
.B2(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_204),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_168),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_158),
.B1(n_156),
.B2(n_164),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_197),
.A2(n_164),
.B1(n_143),
.B2(n_153),
.Y(n_210)
);

AO32x1_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_157),
.A3(n_89),
.B1(n_141),
.B2(n_139),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_213),
.B(n_177),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_182),
.C(n_190),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_218),
.C(n_224),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_211),
.A2(n_194),
.B(n_188),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_217),
.B(n_225),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_196),
.C(n_181),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_219),
.A2(n_228),
.B1(n_202),
.B2(n_210),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_220),
.A2(n_214),
.B(n_209),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_212),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_189),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_222),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_196),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_181),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_157),
.C(n_193),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_225),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_201),
.A2(n_184),
.B1(n_178),
.B2(n_195),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_223),
.B(n_200),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_229),
.B(n_203),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_232),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_226),
.A2(n_209),
.B1(n_201),
.B2(n_200),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_231),
.A2(n_237),
.B1(n_221),
.B2(n_213),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g236 ( 
.A1(n_224),
.A2(n_204),
.B(n_213),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_236),
.A2(n_238),
.B(n_239),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_215),
.A2(n_207),
.B1(n_204),
.B2(n_214),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_240),
.A2(n_218),
.B(n_227),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_242),
.A2(n_233),
.B(n_236),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_245),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_206),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_5),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_216),
.B(n_180),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g249 ( 
.A1(n_247),
.A2(n_232),
.A3(n_236),
.B1(n_239),
.B2(n_237),
.C1(n_240),
.C2(n_234),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_165),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_248),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_245),
.C(n_241),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_252),
.B(n_243),
.Y(n_257)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_247),
.A2(n_238),
.B(n_234),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_163),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_255),
.B(n_253),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_253),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_258),
.B(n_107),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_251),
.A2(n_233),
.B(n_163),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_259),
.Y(n_263)
);

AOI322xp5_ASAP7_75t_L g262 ( 
.A1(n_260),
.A2(n_261),
.A3(n_107),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_8),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_10),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_264),
.B(n_263),
.Y(n_265)
);


endmodule