module fake_jpeg_15746_n_88 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_88);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_88;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx11_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_25),
.B(n_18),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_2),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_0),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_33),
.B1(n_29),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.Y(n_65)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_54),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_52),
.B(n_55),
.Y(n_59)
);

A2O1A1Ixp33_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_39),
.B(n_55),
.C(n_51),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_56),
.B(n_57),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_61),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_60),
.A2(n_65),
.B1(n_6),
.B2(n_7),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_63),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_71),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_8),
.B(n_9),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_70),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_10),
.Y(n_71)
);

NOR3xp33_ASAP7_75t_SL g74 ( 
.A(n_58),
.B(n_11),
.C(n_12),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_16),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_61),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_75),
.B(n_19),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_79),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_69),
.C(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_81),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_67),
.C(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_72),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_80),
.B(n_72),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_85),
.A2(n_77),
.B1(n_79),
.B2(n_24),
.Y(n_86)
);

AOI21x1_ASAP7_75t_SL g87 ( 
.A1(n_86),
.A2(n_27),
.B(n_23),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_21),
.Y(n_88)
);


endmodule