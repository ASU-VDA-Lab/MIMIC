module real_aes_6515_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_769;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g187 ( .A1(n_0), .A2(n_188), .B(n_191), .C(n_195), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_1), .B(n_179), .Y(n_198) );
INVx1_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_3), .B(n_189), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_4), .A2(n_152), .B(n_155), .C(n_545), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_5), .A2(n_147), .B(n_569), .Y(n_568) );
AOI21xp5_ASAP7_75t_L g243 ( .A1(n_6), .A2(n_147), .B(n_244), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_7), .B(n_179), .Y(n_575) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_8), .A2(n_181), .B(n_253), .Y(n_252) );
AND2x6_ASAP7_75t_L g152 ( .A(n_9), .B(n_153), .Y(n_152) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_10), .A2(n_152), .B(n_155), .C(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g536 ( .A(n_11), .Y(n_536) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g462 ( .A(n_12), .B(n_39), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g547 ( .A(n_13), .B(n_194), .Y(n_547) );
INVx1_ASAP7_75t_L g173 ( .A(n_14), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_15), .B(n_189), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g554 ( .A1(n_16), .A2(n_190), .B(n_555), .C(n_557), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_17), .B(n_179), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_18), .B(n_167), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_19), .A2(n_155), .B(n_158), .C(n_166), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g584 ( .A1(n_20), .A2(n_193), .B(n_261), .C(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_21), .B(n_194), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_22), .B(n_194), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_23), .Y(n_517) );
INVx1_ASAP7_75t_L g497 ( .A(n_24), .Y(n_497) );
A2O1A1Ixp33_ASAP7_75t_L g255 ( .A1(n_25), .A2(n_155), .B(n_166), .C(n_256), .Y(n_255) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_26), .Y(n_151) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_27), .Y(n_543) );
INVx1_ASAP7_75t_L g511 ( .A(n_28), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_29), .A2(n_147), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g150 ( .A(n_30), .Y(n_150) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_31), .A2(n_205), .B(n_206), .C(n_210), .Y(n_204) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_32), .A2(n_33), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_32), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_33), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g571 ( .A1(n_34), .A2(n_193), .B(n_572), .C(n_574), .Y(n_571) );
INVxp67_ASAP7_75t_L g512 ( .A(n_35), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_36), .B(n_258), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_37), .A2(n_155), .B(n_166), .C(n_496), .Y(n_495) );
CKINVDCx14_ASAP7_75t_R g570 ( .A(n_38), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_40), .A2(n_195), .B(n_534), .C(n_535), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_41), .B(n_146), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g274 ( .A(n_42), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_43), .B(n_189), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_44), .B(n_147), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_45), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_46), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_47), .A2(n_205), .B(n_210), .C(n_235), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_48), .A2(n_105), .B1(n_116), .B2(n_771), .Y(n_104) );
INVx1_ASAP7_75t_L g192 ( .A(n_49), .Y(n_192) );
INVx1_ASAP7_75t_L g236 ( .A(n_50), .Y(n_236) );
INVx1_ASAP7_75t_L g583 ( .A(n_51), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_52), .B(n_147), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g175 ( .A(n_53), .Y(n_175) );
CKINVDCx14_ASAP7_75t_R g532 ( .A(n_54), .Y(n_532) );
AOI22xp5_ASAP7_75t_SL g468 ( .A1(n_55), .A2(n_460), .B1(n_469), .B2(n_766), .Y(n_468) );
INVx1_ASAP7_75t_L g153 ( .A(n_56), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_57), .B(n_147), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_58), .B(n_179), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_59), .A2(n_165), .B(n_221), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g172 ( .A(n_60), .Y(n_172) );
INVx1_ASAP7_75t_SL g573 ( .A(n_61), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_62), .Y(n_121) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_63), .B(n_189), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_64), .B(n_179), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_65), .B(n_190), .Y(n_271) );
INVx1_ASAP7_75t_L g520 ( .A(n_66), .Y(n_520) );
CKINVDCx16_ASAP7_75t_R g185 ( .A(n_67), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_68), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_69), .A2(n_155), .B(n_210), .C(n_219), .Y(n_218) );
CKINVDCx16_ASAP7_75t_R g245 ( .A(n_70), .Y(n_245) );
INVx1_ASAP7_75t_L g115 ( .A(n_71), .Y(n_115) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_72), .A2(n_147), .B(n_531), .Y(n_530) );
AOI22xp5_ASAP7_75t_L g131 ( .A1(n_73), .A2(n_95), .B1(n_132), .B2(n_133), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_73), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g524 ( .A(n_74), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g478 ( .A1(n_75), .A2(n_103), .B1(n_479), .B2(n_480), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_75), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_76), .A2(n_147), .B(n_552), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_77), .A2(n_146), .B(n_507), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_78), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_79), .A2(n_476), .B1(n_477), .B2(n_478), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_79), .Y(n_476) );
INVx1_ASAP7_75t_L g553 ( .A(n_80), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_81), .B(n_163), .Y(n_162) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_82), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_83), .A2(n_147), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g556 ( .A(n_84), .Y(n_556) );
INVx2_ASAP7_75t_L g170 ( .A(n_85), .Y(n_170) );
INVx1_ASAP7_75t_L g546 ( .A(n_86), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_87), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_88), .B(n_194), .Y(n_272) );
NAND3xp33_ASAP7_75t_SL g111 ( .A(n_89), .B(n_112), .C(n_113), .Y(n_111) );
OR2x2_ASAP7_75t_L g459 ( .A(n_89), .B(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g471 ( .A(n_89), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_90), .A2(n_155), .B(n_210), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_91), .B(n_147), .Y(n_203) );
INVx1_ASAP7_75t_L g207 ( .A(n_92), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_93), .B(n_464), .Y(n_463) );
INVxp67_ASAP7_75t_L g248 ( .A(n_94), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_95), .Y(n_132) );
AOI22xp5_ASAP7_75t_L g474 ( .A1(n_96), .A2(n_475), .B1(n_481), .B2(n_482), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_96), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_97), .B(n_181), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_98), .B(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g220 ( .A(n_99), .Y(n_220) );
INVx1_ASAP7_75t_L g267 ( .A(n_100), .Y(n_267) );
INVx2_ASAP7_75t_L g586 ( .A(n_101), .Y(n_586) );
AND2x2_ASAP7_75t_L g238 ( .A(n_102), .B(n_169), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_103), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
INVx5_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
CKINVDCx9p33_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx4f_ASAP7_75t_SL g771 ( .A(n_108), .Y(n_771) );
OR2x4_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND2x2_ASAP7_75t_L g461 ( .A(n_112), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AO21x2_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_122), .B(n_467), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g770 ( .A(n_121), .Y(n_770) );
OAI21xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_457), .B(n_463), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_125), .B1(n_128), .B2(n_129), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g548 ( .A(n_126), .B(n_180), .Y(n_548) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_131), .B1(n_134), .B2(n_135), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_134), .A2(n_135), .B1(n_473), .B2(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_412), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_347), .Y(n_136) );
NAND4xp25_ASAP7_75t_SL g137 ( .A(n_138), .B(n_292), .C(n_316), .D(n_339), .Y(n_137) );
AOI221xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_229), .B1(n_263), .B2(n_276), .C(n_279), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_199), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_141), .A2(n_177), .B1(n_230), .B2(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_141), .B(n_200), .Y(n_350) );
AND2x2_ASAP7_75t_L g369 ( .A(n_141), .B(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_141), .B(n_353), .Y(n_439) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_177), .Y(n_141) );
AND2x2_ASAP7_75t_L g307 ( .A(n_142), .B(n_200), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_142), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g330 ( .A(n_142), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g335 ( .A(n_142), .B(n_178), .Y(n_335) );
INVx2_ASAP7_75t_L g367 ( .A(n_142), .Y(n_367) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_142), .Y(n_411) );
AND2x2_ASAP7_75t_L g428 ( .A(n_142), .B(n_305), .Y(n_428) );
INVx5_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g346 ( .A(n_143), .B(n_305), .Y(n_346) );
AND2x4_ASAP7_75t_L g360 ( .A(n_143), .B(n_177), .Y(n_360) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_143), .Y(n_364) );
AND2x2_ASAP7_75t_L g384 ( .A(n_143), .B(n_299), .Y(n_384) );
AND2x2_ASAP7_75t_L g434 ( .A(n_143), .B(n_201), .Y(n_434) );
AND2x2_ASAP7_75t_L g444 ( .A(n_143), .B(n_178), .Y(n_444) );
OR2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_174), .Y(n_143) );
AOI21xp5_ASAP7_75t_SL g144 ( .A1(n_145), .A2(n_154), .B(n_167), .Y(n_144) );
BUFx2_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_152), .Y(n_147) );
NAND2x1p5_ASAP7_75t_L g268 ( .A(n_148), .B(n_152), .Y(n_268) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx1_ASAP7_75t_L g165 ( .A(n_149), .Y(n_165) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
INVx1_ASAP7_75t_L g262 ( .A(n_150), .Y(n_262) );
INVx1_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
INVx3_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_151), .Y(n_194) );
INVx1_ASAP7_75t_L g258 ( .A(n_151), .Y(n_258) );
BUFx3_ASAP7_75t_L g166 ( .A(n_152), .Y(n_166) );
INVx4_ASAP7_75t_SL g197 ( .A(n_152), .Y(n_197) );
INVx5_ASAP7_75t_L g186 ( .A(n_155), .Y(n_186) );
AND2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
BUFx3_ASAP7_75t_L g196 ( .A(n_156), .Y(n_196) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_156), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_162), .B(n_164), .Y(n_158) );
INVx2_ASAP7_75t_L g163 ( .A(n_160), .Y(n_163) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx4_ASAP7_75t_L g222 ( .A(n_161), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_163), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_163), .A2(n_209), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_163), .A2(n_520), .B(n_521), .C(n_522), .Y(n_519) );
O2A1O1Ixp5_ASAP7_75t_L g545 ( .A1(n_163), .A2(n_522), .B(n_546), .C(n_547), .Y(n_545) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_164), .A2(n_189), .B(n_497), .C(n_498), .Y(n_496) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_165), .B(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_168), .B(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_169), .A2(n_203), .B(n_204), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_169), .A2(n_233), .B(n_234), .Y(n_232) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_169), .A2(n_268), .B(n_494), .C(n_495), .Y(n_493) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_169), .A2(n_530), .B(n_537), .Y(n_529) );
AND2x2_ASAP7_75t_SL g169 ( .A(n_170), .B(n_171), .Y(n_169) );
AND2x2_ASAP7_75t_L g182 ( .A(n_170), .B(n_171), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
AO21x2_ASAP7_75t_L g541 ( .A1(n_176), .A2(n_542), .B(n_548), .Y(n_541) );
AND2x2_ASAP7_75t_L g300 ( .A(n_177), .B(n_200), .Y(n_300) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_177), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_177), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g390 ( .A(n_177), .Y(n_390) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g278 ( .A(n_178), .B(n_215), .Y(n_278) );
AND2x2_ASAP7_75t_L g305 ( .A(n_178), .B(n_216), .Y(n_305) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_183), .B(n_198), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_180), .B(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_180), .A2(n_217), .B(n_227), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_180), .B(n_228), .Y(n_227) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_180), .A2(n_266), .B(n_273), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_180), .B(n_500), .Y(n_499) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_180), .A2(n_516), .B(n_523), .Y(n_515) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_181), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_181), .A2(n_254), .B(n_255), .Y(n_253) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g275 ( .A(n_182), .Y(n_275) );
O2A1O1Ixp33_ASAP7_75t_SL g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_197), .Y(n_184) );
INVx2_ASAP7_75t_L g205 ( .A(n_186), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_186), .A2(n_197), .B(n_245), .C(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_186), .A2(n_197), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_186), .A2(n_197), .B(n_532), .C(n_533), .Y(n_531) );
O2A1O1Ixp33_ASAP7_75t_SL g552 ( .A1(n_186), .A2(n_197), .B(n_553), .C(n_554), .Y(n_552) );
O2A1O1Ixp33_ASAP7_75t_L g569 ( .A1(n_186), .A2(n_197), .B(n_570), .C(n_571), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_SL g582 ( .A1(n_186), .A2(n_197), .B(n_583), .C(n_584), .Y(n_582) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_189), .B(n_248), .Y(n_247) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_189), .A2(n_222), .B1(n_511), .B2(n_512), .Y(n_510) );
INVx5_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_190), .B(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_192), .B(n_193), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_193), .B(n_573), .Y(n_572) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g534 ( .A(n_194), .Y(n_534) );
INVx2_ASAP7_75t_L g522 ( .A(n_195), .Y(n_522) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
HB1xp67_ASAP7_75t_L g209 ( .A(n_196), .Y(n_209) );
INVx1_ASAP7_75t_L g557 ( .A(n_196), .Y(n_557) );
INVx1_ASAP7_75t_L g210 ( .A(n_197), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_199), .B(n_364), .Y(n_363) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_213), .Y(n_199) );
OR2x2_ASAP7_75t_L g331 ( .A(n_200), .B(n_214), .Y(n_331) );
AND2x2_ASAP7_75t_L g368 ( .A(n_200), .B(n_278), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_200), .B(n_299), .Y(n_379) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_200), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_200), .B(n_335), .Y(n_452) );
INVx5_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
BUFx2_ASAP7_75t_L g277 ( .A(n_201), .Y(n_277) );
AND2x2_ASAP7_75t_L g286 ( .A(n_201), .B(n_214), .Y(n_286) );
AND2x2_ASAP7_75t_L g402 ( .A(n_201), .B(n_297), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_201), .B(n_335), .Y(n_424) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_211), .Y(n_201) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_214), .Y(n_370) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_215), .Y(n_322) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
BUFx2_ASAP7_75t_L g299 ( .A(n_216), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_226), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_223), .C(n_224), .Y(n_219) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_222), .B(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_222), .B(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx3_ASAP7_75t_L g574 ( .A(n_225), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_230), .B(n_239), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_230), .B(n_312), .Y(n_431) );
HB1xp67_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_231), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g283 ( .A(n_231), .B(n_284), .Y(n_283) );
INVx5_ASAP7_75t_SL g291 ( .A(n_231), .Y(n_291) );
OR2x2_ASAP7_75t_L g314 ( .A(n_231), .B(n_284), .Y(n_314) );
OR2x2_ASAP7_75t_L g324 ( .A(n_231), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g387 ( .A(n_231), .B(n_241), .Y(n_387) );
AND2x2_ASAP7_75t_SL g425 ( .A(n_231), .B(n_240), .Y(n_425) );
NOR4xp25_ASAP7_75t_L g446 ( .A(n_231), .B(n_367), .C(n_447), .D(n_448), .Y(n_446) );
AND2x2_ASAP7_75t_L g456 ( .A(n_231), .B(n_288), .Y(n_456) );
OR2x6_ASAP7_75t_L g231 ( .A(n_232), .B(n_238), .Y(n_231) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g281 ( .A(n_240), .B(n_277), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_240), .B(n_283), .Y(n_450) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_250), .Y(n_240) );
OR2x2_ASAP7_75t_L g290 ( .A(n_241), .B(n_291), .Y(n_290) );
INVx3_ASAP7_75t_L g297 ( .A(n_241), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_241), .B(n_265), .Y(n_309) );
INVxp67_ASAP7_75t_L g312 ( .A(n_241), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_241), .B(n_284), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_241), .B(n_251), .Y(n_378) );
AND2x2_ASAP7_75t_L g393 ( .A(n_241), .B(n_288), .Y(n_393) );
OR2x2_ASAP7_75t_L g422 ( .A(n_241), .B(n_251), .Y(n_422) );
OA21x2_ASAP7_75t_L g241 ( .A1(n_242), .A2(n_243), .B(n_249), .Y(n_241) );
OA21x2_ASAP7_75t_L g550 ( .A1(n_242), .A2(n_551), .B(n_558), .Y(n_550) );
OA21x2_ASAP7_75t_L g567 ( .A1(n_242), .A2(n_568), .B(n_575), .Y(n_567) );
OA21x2_ASAP7_75t_L g580 ( .A1(n_242), .A2(n_581), .B(n_587), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_250), .B(n_327), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_250), .B(n_291), .Y(n_430) );
OR2x2_ASAP7_75t_L g451 ( .A(n_250), .B(n_328), .Y(n_451) );
INVx1_ASAP7_75t_SL g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g264 ( .A(n_251), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g288 ( .A(n_251), .B(n_284), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_251), .B(n_265), .Y(n_303) );
AND2x2_ASAP7_75t_L g373 ( .A(n_251), .B(n_297), .Y(n_373) );
AND2x2_ASAP7_75t_L g407 ( .A(n_251), .B(n_291), .Y(n_407) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_252), .B(n_291), .Y(n_310) );
AND2x2_ASAP7_75t_L g338 ( .A(n_252), .B(n_265), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_259), .B(n_260), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_260), .A2(n_271), .B(n_272), .Y(n_270) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_263), .B(n_346), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g405 ( .A1(n_264), .A2(n_353), .B1(n_389), .B2(n_406), .C(n_408), .Y(n_405) );
INVx5_ASAP7_75t_SL g284 ( .A(n_265), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_269), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_268), .A2(n_517), .B(n_518), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g542 ( .A1(n_268), .A2(n_543), .B(n_544), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
INVx2_ASAP7_75t_L g505 ( .A(n_275), .Y(n_505) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
OAI33xp33_ASAP7_75t_L g304 ( .A1(n_277), .A2(n_305), .A3(n_306), .B1(n_308), .B2(n_311), .B3(n_315), .Y(n_304) );
OR2x2_ASAP7_75t_L g320 ( .A(n_277), .B(n_321), .Y(n_320) );
AOI322xp5_ASAP7_75t_L g429 ( .A1(n_277), .A2(n_346), .A3(n_353), .B1(n_430), .B2(n_431), .C1(n_432), .C2(n_435), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_277), .B(n_305), .Y(n_447) );
A2O1A1Ixp33_ASAP7_75t_SL g453 ( .A1(n_277), .A2(n_305), .B(n_454), .C(n_456), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g292 ( .A1(n_278), .A2(n_293), .B1(n_298), .B2(n_301), .C(n_304), .Y(n_292) );
INVx1_ASAP7_75t_L g385 ( .A(n_278), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_278), .B(n_434), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_282), .B1(n_285), .B2(n_287), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g362 ( .A(n_283), .B(n_297), .Y(n_362) );
AND2x2_ASAP7_75t_L g420 ( .A(n_283), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g328 ( .A(n_284), .B(n_291), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_284), .B(n_297), .Y(n_356) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_286), .B(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_286), .B(n_364), .Y(n_418) );
OAI321xp33_ASAP7_75t_L g437 ( .A1(n_286), .A2(n_359), .A3(n_438), .B1(n_439), .B2(n_440), .C(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g404 ( .A(n_287), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_288), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g343 ( .A(n_288), .B(n_291), .Y(n_343) );
AOI321xp33_ASAP7_75t_L g401 ( .A1(n_288), .A2(n_305), .A3(n_402), .B1(n_403), .B2(n_404), .C(n_405), .Y(n_401) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g318 ( .A(n_290), .B(n_303), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_291), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_291), .B(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_291), .B(n_377), .Y(n_414) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x4_ASAP7_75t_L g337 ( .A(n_295), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OR2x2_ASAP7_75t_L g302 ( .A(n_296), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g410 ( .A(n_297), .Y(n_410) );
AND2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_300), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_307), .B(n_342), .Y(n_391) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
OR2x2_ASAP7_75t_L g355 ( .A(n_310), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g400 ( .A(n_310), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_311), .A2(n_358), .B1(n_361), .B2(n_363), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g455 ( .A(n_314), .B(n_378), .Y(n_455) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_319), .B1(n_323), .B2(n_329), .C(n_332), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx2_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
INVx1_ASAP7_75t_SL g399 ( .A(n_325), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_327), .B(n_377), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_327), .A2(n_395), .B(n_397), .Y(n_394) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g440 ( .A(n_328), .B(n_422), .Y(n_440) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_SL g342 ( .A(n_331), .Y(n_342) );
AOI21xp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B(n_336), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g386 ( .A(n_338), .B(n_387), .Y(n_386) );
INVxp67_ASAP7_75t_L g448 ( .A(n_338), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_343), .B(n_344), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_342), .B(n_360), .Y(n_396) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g417 ( .A(n_346), .Y(n_417) );
NAND5xp2_ASAP7_75t_L g347 ( .A(n_348), .B(n_365), .C(n_374), .D(n_394), .E(n_401), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_351), .B(n_354), .C(n_357), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g389 ( .A(n_353), .Y(n_389) );
CKINVDCx16_ASAP7_75t_R g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_361), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g403 ( .A(n_363), .Y(n_403) );
OAI21xp5_ASAP7_75t_SL g365 ( .A1(n_366), .A2(n_369), .B(n_371), .Y(n_365) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_366), .A2(n_420), .B1(n_423), .B2(n_425), .C(n_426), .Y(n_419) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AOI321xp33_ASAP7_75t_L g374 ( .A1(n_367), .A2(n_375), .A3(n_379), .B1(n_380), .B2(n_386), .C(n_388), .Y(n_374) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g445 ( .A(n_379), .Y(n_445) );
NAND2xp5_ASAP7_75t_SL g380 ( .A(n_381), .B(n_385), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g397 ( .A(n_382), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NOR2xp67_ASAP7_75t_SL g409 ( .A(n_383), .B(n_390), .Y(n_409) );
AOI321xp33_ASAP7_75t_SL g441 ( .A1(n_386), .A2(n_442), .A3(n_443), .B1(n_444), .B2(n_445), .C(n_446), .Y(n_441) );
O2A1O1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B(n_391), .C(n_392), .Y(n_388) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_399), .B(n_407), .Y(n_436) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NAND3xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .C(n_411), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_437), .C(n_449), .Y(n_412) );
OAI211xp5_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_415), .B(n_419), .C(n_429), .Y(n_413) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_SL g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OAI221xp5_ASAP7_75t_L g449 ( .A1(n_418), .A2(n_450), .B1(n_451), .B2(n_452), .C(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g438 ( .A(n_420), .Y(n_438) );
INVx1_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_SL g442 ( .A(n_440), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
CKINVDCx14_ASAP7_75t_R g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g466 ( .A(n_459), .Y(n_466) );
NOR2x2_ASAP7_75t_L g768 ( .A(n_460), .B(n_471), .Y(n_768) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_463), .A2(n_468), .B(n_769), .Y(n_467) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B1(n_483), .B2(n_485), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g484 ( .A(n_471), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_473), .A2(n_474), .B1(n_486), .B2(n_487), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g482 ( .A(n_475), .Y(n_482) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR4x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_656), .C(n_703), .D(n_743), .Y(n_487) );
NAND3xp33_ASAP7_75t_SL g488 ( .A(n_489), .B(n_602), .C(n_631), .Y(n_488) );
AOI211xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_525), .B(n_559), .C(n_595), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_L g631 ( .A1(n_490), .A2(n_615), .B(n_632), .C(n_636), .Y(n_631) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_492), .B(n_594), .Y(n_593) );
INVx3_ASAP7_75t_SL g598 ( .A(n_492), .Y(n_598) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_492), .Y(n_610) );
AND2x4_ASAP7_75t_L g614 ( .A(n_492), .B(n_566), .Y(n_614) );
AND2x2_ASAP7_75t_L g625 ( .A(n_492), .B(n_515), .Y(n_625) );
OR2x2_ASAP7_75t_L g649 ( .A(n_492), .B(n_562), .Y(n_649) );
AND2x2_ASAP7_75t_L g662 ( .A(n_492), .B(n_567), .Y(n_662) );
AND2x2_ASAP7_75t_L g702 ( .A(n_492), .B(n_688), .Y(n_702) );
AND2x2_ASAP7_75t_L g709 ( .A(n_492), .B(n_672), .Y(n_709) );
AND2x2_ASAP7_75t_L g739 ( .A(n_492), .B(n_502), .Y(n_739) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_499), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_501), .B(n_666), .Y(n_678) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_514), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_502), .B(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g616 ( .A(n_502), .B(n_514), .Y(n_616) );
BUFx3_ASAP7_75t_L g624 ( .A(n_502), .Y(n_624) );
OR2x2_ASAP7_75t_L g645 ( .A(n_502), .B(n_528), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_502), .B(n_666), .Y(n_756) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_506), .B(n_513), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g562 ( .A1(n_504), .A2(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g563 ( .A(n_506), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_513), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_514), .B(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g609 ( .A(n_514), .Y(n_609) );
AND2x2_ASAP7_75t_L g672 ( .A(n_514), .B(n_567), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_514), .A2(n_675), .B1(n_677), .B2(n_679), .C(n_680), .Y(n_674) );
AND2x2_ASAP7_75t_L g688 ( .A(n_514), .B(n_562), .Y(n_688) );
AND2x2_ASAP7_75t_L g714 ( .A(n_514), .B(n_598), .Y(n_714) );
INVx2_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g594 ( .A(n_515), .B(n_567), .Y(n_594) );
BUFx2_ASAP7_75t_L g728 ( .A(n_515), .Y(n_728) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
OAI32xp33_ASAP7_75t_L g694 ( .A1(n_526), .A2(n_655), .A3(n_669), .B1(n_695), .B2(n_696), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_538), .Y(n_526) );
AND2x2_ASAP7_75t_L g635 ( .A(n_527), .B(n_579), .Y(n_635) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g617 ( .A(n_528), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_528), .B(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g689 ( .A(n_528), .B(n_579), .Y(n_689) );
AND2x2_ASAP7_75t_L g700 ( .A(n_528), .B(n_592), .Y(n_700) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g601 ( .A(n_529), .B(n_580), .Y(n_601) );
AND2x2_ASAP7_75t_L g605 ( .A(n_529), .B(n_580), .Y(n_605) );
AND2x2_ASAP7_75t_L g640 ( .A(n_529), .B(n_591), .Y(n_640) );
AND2x2_ASAP7_75t_L g647 ( .A(n_529), .B(n_549), .Y(n_647) );
OAI211xp5_ASAP7_75t_L g652 ( .A1(n_529), .A2(n_598), .B(n_609), .C(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g706 ( .A(n_529), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_529), .B(n_540), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_538), .B(n_589), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_538), .B(n_605), .Y(n_695) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g600 ( .A(n_539), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_549), .Y(n_539) );
AND2x2_ASAP7_75t_L g592 ( .A(n_540), .B(n_550), .Y(n_592) );
OR2x2_ASAP7_75t_L g607 ( .A(n_540), .B(n_550), .Y(n_607) );
AND2x2_ASAP7_75t_L g630 ( .A(n_540), .B(n_591), .Y(n_630) );
INVx1_ASAP7_75t_L g634 ( .A(n_540), .Y(n_634) );
AND2x2_ASAP7_75t_L g653 ( .A(n_540), .B(n_590), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g663 ( .A1(n_540), .A2(n_618), .B1(n_664), .B2(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_540), .B(n_706), .Y(n_730) );
AND2x2_ASAP7_75t_L g745 ( .A(n_540), .B(n_605), .Y(n_745) );
INVx4_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx3_ASAP7_75t_L g577 ( .A(n_541), .Y(n_577) );
AND2x2_ASAP7_75t_L g619 ( .A(n_541), .B(n_550), .Y(n_619) );
AND2x2_ASAP7_75t_L g621 ( .A(n_541), .B(n_579), .Y(n_621) );
AND3x2_ASAP7_75t_L g683 ( .A(n_541), .B(n_647), .C(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g718 ( .A(n_549), .B(n_590), .Y(n_718) );
INVx1_ASAP7_75t_SL g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g579 ( .A(n_550), .B(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_550), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_550), .B(n_589), .Y(n_651) );
NAND3xp33_ASAP7_75t_L g758 ( .A(n_550), .B(n_630), .C(n_706), .Y(n_758) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_576), .B1(n_588), .B2(n_593), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_562), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g670 ( .A(n_562), .Y(n_670) );
OAI31xp33_ASAP7_75t_L g686 ( .A1(n_565), .A2(n_687), .A3(n_688), .B(n_689), .Y(n_686) );
AND2x2_ASAP7_75t_L g711 ( .A(n_565), .B(n_598), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_565), .B(n_624), .Y(n_757) );
AND2x2_ASAP7_75t_L g666 ( .A(n_566), .B(n_598), .Y(n_666) );
AND2x2_ASAP7_75t_L g727 ( .A(n_566), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g597 ( .A(n_567), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g655 ( .A(n_567), .Y(n_655) );
OR2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
CKINVDCx16_ASAP7_75t_R g676 ( .A(n_577), .Y(n_676) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_578), .B(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AOI221x1_ASAP7_75t_SL g643 ( .A1(n_579), .A2(n_644), .B1(n_646), .B2(n_648), .C(n_650), .Y(n_643) );
INVx2_ASAP7_75t_L g591 ( .A(n_580), .Y(n_591) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_580), .Y(n_685) );
INVx1_ASAP7_75t_L g673 ( .A(n_588), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_592), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_589), .B(n_606), .Y(n_698) );
INVx1_ASAP7_75t_SL g761 ( .A(n_589), .Y(n_761) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g679 ( .A(n_592), .B(n_605), .Y(n_679) );
INVx1_ASAP7_75t_L g747 ( .A(n_593), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_593), .B(n_676), .Y(n_760) );
INVx2_ASAP7_75t_SL g599 ( .A(n_594), .Y(n_599) );
AND2x2_ASAP7_75t_L g642 ( .A(n_594), .B(n_598), .Y(n_642) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_594), .B(n_649), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_594), .B(n_669), .Y(n_696) );
AOI21xp33_ASAP7_75t_SL g595 ( .A1(n_596), .A2(n_599), .B(n_600), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_597), .B(n_669), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_597), .B(n_624), .Y(n_765) );
OR2x2_ASAP7_75t_L g637 ( .A(n_598), .B(n_616), .Y(n_637) );
AND2x2_ASAP7_75t_L g736 ( .A(n_598), .B(n_727), .Y(n_736) );
OAI22xp5_ASAP7_75t_SL g611 ( .A1(n_599), .A2(n_612), .B1(n_617), .B2(n_620), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g644 ( .A(n_599), .B(n_645), .Y(n_644) );
OR2x2_ASAP7_75t_L g659 ( .A(n_601), .B(n_607), .Y(n_659) );
INVx1_ASAP7_75t_L g723 ( .A(n_601), .Y(n_723) );
AOI311xp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_608), .A3(n_610), .B(n_611), .C(n_622), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
AOI221xp5_ASAP7_75t_L g749 ( .A1(n_606), .A2(n_738), .B1(n_750), .B2(n_753), .C(n_755), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_606), .B(n_761), .Y(n_763) );
INVx2_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g660 ( .A(n_608), .Y(n_660) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_609), .A2(n_651), .B(n_652), .C(n_654), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
O2A1O1Ixp33_ASAP7_75t_SL g719 ( .A1(n_613), .A2(n_615), .B(n_720), .C(n_721), .Y(n_719) );
INVx3_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_614), .B(n_688), .Y(n_754) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_617), .A2(n_637), .B1(n_638), .B2(n_641), .C(n_643), .Y(n_636) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g639 ( .A(n_619), .B(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g722 ( .A(n_619), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
NOR2xp33_ASAP7_75t_L g622 ( .A(n_623), .B(n_626), .Y(n_622) );
A2O1A1Ixp33_ASAP7_75t_L g680 ( .A1(n_623), .A2(n_681), .B(n_682), .C(n_686), .Y(n_680) );
NAND2xp5_ASAP7_75t_SL g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_624), .B(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_624), .B(n_727), .Y(n_726) );
OR2x2_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
INVxp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g646 ( .A(n_630), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_634), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g748 ( .A(n_637), .Y(n_748) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_640), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g675 ( .A(n_640), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g752 ( .A(n_640), .Y(n_752) );
INVx1_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g693 ( .A(n_642), .B(n_669), .Y(n_693) );
INVx1_ASAP7_75t_SL g687 ( .A(n_649), .Y(n_687) );
INVx1_ASAP7_75t_L g664 ( .A(n_655), .Y(n_664) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_674), .C(n_690), .Y(n_656) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_660), .A3(n_661), .B1(n_663), .B2(n_667), .C1(n_671), .C2(n_673), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g710 ( .A1(n_658), .A2(n_711), .B(n_712), .C(n_719), .Y(n_710) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_661), .A2(n_682), .B1(n_713), .B2(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g671 ( .A(n_669), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g708 ( .A(n_669), .B(n_709), .Y(n_708) );
AOI32xp33_ASAP7_75t_L g759 ( .A1(n_669), .A2(n_760), .A3(n_761), .B1(n_762), .B2(n_764), .Y(n_759) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g681 ( .A(n_672), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_672), .A2(n_725), .B1(n_729), .B2(n_731), .C(n_734), .Y(n_724) );
AND2x2_ASAP7_75t_L g738 ( .A(n_672), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g741 ( .A(n_676), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g751 ( .A(n_676), .B(n_752), .Y(n_751) );
INVxp67_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVxp67_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g742 ( .A(n_685), .B(n_706), .Y(n_742) );
AOI211xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B(n_694), .C(n_697), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B(n_701), .Y(n_697) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g703 ( .A1(n_704), .A2(n_707), .B(n_710), .C(n_724), .Y(n_703) );
INVxp67_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_718), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g733 ( .A(n_730), .Y(n_733) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B(n_740), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
OAI211xp5_ASAP7_75t_SL g743 ( .A1(n_744), .A2(n_746), .B(n_749), .C(n_759), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_747), .B(n_748), .Y(n_746) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AOI21xp33_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_758), .Y(n_755) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
INVx3_ASAP7_75t_SL g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
endmodule