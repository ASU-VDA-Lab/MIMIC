module fake_jpeg_26759_n_333 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_333);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_333;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_14),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_33),
.Y(n_48)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_39),
.B(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_47),
.B(n_63),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_48),
.B(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_40),
.A2(n_17),
.B(n_29),
.C(n_35),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_19),
.B(n_30),
.C(n_25),
.Y(n_80)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_58),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_33),
.B1(n_17),
.B2(n_35),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_60),
.Y(n_94)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_40),
.B(n_19),
.Y(n_66)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_44),
.B1(n_38),
.B2(n_46),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_54),
.B1(n_61),
.B2(n_53),
.Y(n_102)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_74),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_18),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_80),
.Y(n_118)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_96),
.Y(n_101)
);

NAND2x1_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_40),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_41),
.C(n_20),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_81),
.B(n_89),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_85),
.B(n_87),
.Y(n_100)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_30),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_95),
.B1(n_51),
.B2(n_55),
.Y(n_107)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_93),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_61),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_94),
.A2(n_28),
.B1(n_27),
.B2(n_58),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_111),
.B1(n_74),
.B2(n_73),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_56),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_105),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_94),
.A2(n_68),
.B1(n_55),
.B2(n_56),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_106),
.A2(n_79),
.B(n_84),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_107),
.B(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_45),
.B1(n_41),
.B2(n_37),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_87),
.B(n_36),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_88),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_80),
.A2(n_41),
.B1(n_37),
.B2(n_23),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_114),
.A2(n_120),
.B1(n_123),
.B2(n_125),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_83),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_84),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_121),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_88),
.A2(n_24),
.B1(n_22),
.B2(n_34),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_32),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_76),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g123 ( 
.A1(n_78),
.A2(n_42),
.B1(n_34),
.B2(n_21),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_88),
.A2(n_24),
.B1(n_22),
.B2(n_34),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_100),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_126),
.B(n_129),
.Y(n_169)
);

OA21x2_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_82),
.B(n_83),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_123),
.B(n_109),
.Y(n_157)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_128),
.B(n_131),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_134),
.B1(n_136),
.B2(n_152),
.Y(n_160)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_90),
.B1(n_96),
.B2(n_91),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_90),
.B1(n_86),
.B2(n_71),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_113),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_138),
.B(n_140),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_139),
.A2(n_145),
.B(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_72),
.Y(n_140)
);

AOI22x1_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_42),
.B1(n_77),
.B2(n_71),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_141),
.A2(n_110),
.B1(n_124),
.B2(n_104),
.Y(n_173)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_124),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_98),
.A2(n_72),
.B(n_32),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_148),
.Y(n_156)
);

INVxp33_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_108),
.A2(n_106),
.B(n_114),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_115),
.B(n_32),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_124),
.C(n_104),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_111),
.A2(n_76),
.B1(n_79),
.B2(n_21),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_140),
.B(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_155),
.B(n_163),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_178),
.B1(n_171),
.B2(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_149),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_158),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_161),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_164),
.B(n_175),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_102),
.B1(n_107),
.B2(n_123),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_165),
.A2(n_153),
.B1(n_150),
.B2(n_130),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_182),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_142),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_168),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_120),
.B1(n_119),
.B2(n_116),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_170),
.A2(n_152),
.B1(n_137),
.B2(n_151),
.Y(n_203)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_171),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_139),
.A2(n_0),
.B(n_1),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_172),
.A2(n_179),
.B(n_180),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_173),
.A2(n_178),
.B1(n_134),
.B2(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_131),
.C(n_97),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_128),
.B(n_104),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_177),
.B(n_97),
.Y(n_191)
);

OAI22x1_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_97),
.B1(n_21),
.B2(n_20),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_127),
.A2(n_0),
.B(n_2),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_143),
.A2(n_0),
.B(n_2),
.Y(n_180)
);

XOR2x1_ASAP7_75t_L g181 ( 
.A(n_126),
.B(n_15),
.Y(n_181)
);

XNOR2x1_ASAP7_75t_SL g189 ( 
.A(n_181),
.B(n_145),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_133),
.Y(n_182)
);

NAND2x1p5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_127),
.Y(n_183)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_183),
.B(n_161),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_129),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_10),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_190),
.B1(n_192),
.B2(n_197),
.Y(n_212)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_155),
.B(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_153),
.B1(n_132),
.B2(n_146),
.Y(n_192)
);

OAI32xp33_ASAP7_75t_L g193 ( 
.A1(n_167),
.A2(n_168),
.A3(n_175),
.B1(n_159),
.B2(n_181),
.Y(n_193)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_193),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_194),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_233)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_195),
.B(n_198),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_162),
.A2(n_132),
.B(n_127),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_196),
.A2(n_180),
.B(n_158),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_178),
.A2(n_176),
.B1(n_179),
.B2(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_138),
.Y(n_200)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_204),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_203),
.A2(n_177),
.B1(n_172),
.B2(n_160),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_207),
.C(n_210),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_169),
.B(n_20),
.C(n_15),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_162),
.B(n_14),
.C(n_13),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_211),
.B(n_236),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_216),
.A2(n_221),
.B(n_187),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_208),
.B(n_156),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_218),
.B(n_227),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_220),
.A2(n_230),
.B1(n_233),
.B2(n_197),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_222),
.Y(n_237)
);

NAND3xp33_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_193),
.C(n_185),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_182),
.C(n_174),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_225),
.C(n_226),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_174),
.C(n_14),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_13),
.C(n_11),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_209),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_209),
.B1(n_198),
.B2(n_195),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_192),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_13),
.B(n_11),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_231),
.B(n_232),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_200),
.B(n_11),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_10),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_234),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_207),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_208),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_248),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_252),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_244),
.B1(n_245),
.B2(n_230),
.Y(n_275)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_242),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_220),
.A2(n_188),
.B1(n_183),
.B2(n_201),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_216),
.A2(n_183),
.B1(n_199),
.B2(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_251),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_205),
.Y(n_250)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_222),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_196),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_253),
.A2(n_250),
.B(n_254),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_205),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_255),
.A2(n_246),
.B(n_249),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_203),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_212),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_185),
.C(n_210),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_225),
.C(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_265),
.Y(n_283)
);

BUFx24_ASAP7_75t_SL g261 ( 
.A(n_241),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_261),
.B(n_263),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_238),
.A2(n_214),
.B1(n_211),
.B2(n_216),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

AOI21x1_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_221),
.B(n_214),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_267),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_217),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_247),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_226),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_270),
.A2(n_237),
.B(n_255),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_213),
.C(n_212),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_243),
.C(n_258),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_275),
.A2(n_245),
.B(n_229),
.Y(n_287)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_276),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_252),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_285),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_285),
.C(n_277),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_279),
.B(n_287),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_264),
.A2(n_244),
.B1(n_240),
.B2(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_290),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_263),
.A2(n_248),
.B1(n_213),
.B2(n_229),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_282),
.A2(n_288),
.B1(n_280),
.B2(n_276),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_267),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_239),
.C(n_228),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_289),
.B(n_278),
.C(n_283),
.Y(n_293)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_269),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_291),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_281),
.B(n_268),
.Y(n_292)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_292),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_287),
.C(n_286),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_300),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_209),
.Y(n_298)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_289),
.B(n_265),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_301),
.B(n_256),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_259),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_5),
.B(n_6),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_306),
.C(n_311),
.Y(n_319)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_274),
.B(n_4),
.Y(n_309)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_3),
.C(n_4),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_297),
.B(n_4),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_313),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_303),
.Y(n_315)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_315),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_305),
.B(n_294),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_320),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_302),
.C(n_295),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_308),
.B(n_294),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_321),
.A2(n_322),
.B(n_6),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_311),
.B(n_5),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_319),
.A2(n_314),
.B1(n_7),
.B2(n_8),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_325),
.A2(n_326),
.B(n_316),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_327),
.A2(n_328),
.B(n_318),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_SL g328 ( 
.A1(n_324),
.A2(n_318),
.B(n_7),
.C(n_8),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_323),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_6),
.C(n_8),
.Y(n_331)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_9),
.B(n_309),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_9),
.Y(n_333)
);


endmodule