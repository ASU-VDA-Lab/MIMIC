module real_aes_17820_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_831, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_831;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_449;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_617;
wire n_552;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g115 ( .A(n_0), .B(n_116), .Y(n_115) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_1), .A2(n_4), .B1(n_157), .B2(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g199 ( .A1(n_2), .A2(n_40), .B1(n_164), .B2(n_200), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_3), .A2(n_23), .B1(n_200), .B2(n_242), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_5), .A2(n_15), .B1(n_154), .B2(n_231), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_6), .A2(n_58), .B1(n_214), .B2(n_244), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g600 ( .A1(n_7), .A2(n_16), .B1(n_164), .B2(n_185), .Y(n_600) );
INVx1_ASAP7_75t_L g116 ( .A(n_8), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g513 ( .A(n_9), .Y(n_513) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_10), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_11), .A2(n_17), .B1(n_213), .B2(n_216), .Y(n_212) );
BUFx2_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
OR2x2_ASAP7_75t_L g126 ( .A(n_12), .B(n_36), .Y(n_126) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_13), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g235 ( .A(n_14), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g153 ( .A1(n_18), .A2(n_99), .B1(n_154), .B2(n_157), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_19), .A2(n_37), .B1(n_189), .B2(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_20), .B(n_155), .Y(n_186) );
OAI21x1_ASAP7_75t_L g172 ( .A1(n_21), .A2(n_54), .B(n_173), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_22), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_24), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_25), .B(n_161), .Y(n_520) );
INVx4_ASAP7_75t_R g568 ( .A(n_26), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g201 ( .A1(n_27), .A2(n_45), .B1(n_202), .B2(n_203), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g282 ( .A1(n_28), .A2(n_51), .B1(n_154), .B2(n_203), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_29), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_30), .B(n_189), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_31), .Y(n_265) );
INVx1_ASAP7_75t_L g499 ( .A(n_32), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_33), .B(n_200), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_SL g511 ( .A1(n_34), .A2(n_160), .B(n_164), .C(n_512), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_35), .A2(n_52), .B1(n_164), .B2(n_203), .Y(n_488) );
HB1xp67_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
AOI22xp5_ASAP7_75t_L g240 ( .A1(n_38), .A2(n_85), .B1(n_164), .B2(n_241), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_39), .A2(n_44), .B1(n_164), .B2(n_185), .Y(n_217) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_41), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_42), .A2(n_56), .B1(n_154), .B2(n_163), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_43), .A2(n_70), .B1(n_129), .B2(n_130), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_43), .Y(n_130) );
INVx1_ASAP7_75t_L g523 ( .A(n_46), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_47), .B(n_164), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_48), .Y(n_540) );
INVx2_ASAP7_75t_L g121 ( .A(n_49), .Y(n_121) );
INVx1_ASAP7_75t_L g110 ( .A(n_50), .Y(n_110) );
BUFx3_ASAP7_75t_L g124 ( .A(n_50), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_53), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_55), .A2(n_86), .B1(n_164), .B2(n_203), .Y(n_601) );
OAI22xp5_ASAP7_75t_L g804 ( .A1(n_57), .A2(n_66), .B1(n_805), .B2(n_806), .Y(n_804) );
INVx1_ASAP7_75t_L g806 ( .A(n_57), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_59), .A2(n_74), .B1(n_163), .B2(n_202), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_60), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_61), .A2(n_76), .B1(n_164), .B2(n_185), .Y(n_263) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_62), .Y(n_828) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_63), .A2(n_98), .B1(n_154), .B2(n_216), .Y(n_262) );
AND2x4_ASAP7_75t_L g150 ( .A(n_64), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g173 ( .A(n_65), .Y(n_173) );
INVx1_ASAP7_75t_L g805 ( .A(n_66), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_67), .A2(n_89), .B1(n_202), .B2(n_203), .Y(n_495) );
AO22x1_ASAP7_75t_L g557 ( .A1(n_68), .A2(n_75), .B1(n_228), .B2(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g151 ( .A(n_69), .Y(n_151) );
INVx1_ASAP7_75t_L g129 ( .A(n_70), .Y(n_129) );
AND2x2_ASAP7_75t_L g515 ( .A(n_71), .B(n_195), .Y(n_515) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_72), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_73), .B(n_244), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_77), .B(n_200), .Y(n_541) );
INVx2_ASAP7_75t_L g161 ( .A(n_78), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_79), .B(n_195), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_80), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_81), .A2(n_97), .B1(n_203), .B2(n_244), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_82), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_83), .B(n_171), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_84), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g826 ( .A(n_87), .Y(n_826) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_88), .B(n_195), .Y(n_194) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_90), .Y(n_223) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_91), .B(n_195), .Y(n_537) );
INVx1_ASAP7_75t_L g114 ( .A(n_92), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_92), .B(n_811), .Y(n_810) );
AOI21xp5_ASAP7_75t_L g814 ( .A1(n_93), .A2(n_815), .B(n_822), .Y(n_814) );
NAND2xp33_ASAP7_75t_L g191 ( .A(n_94), .B(n_155), .Y(n_191) );
A2O1A1Ixp33_ASAP7_75t_L g563 ( .A1(n_95), .A2(n_219), .B(n_244), .C(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g570 ( .A(n_96), .B(n_571), .Y(n_570) );
NAND2xp33_ASAP7_75t_L g545 ( .A(n_100), .B(n_190), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_117), .B(n_827), .Y(n_101) );
BUFx8_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
BUFx12f_ASAP7_75t_L g829 ( .A(n_103), .Y(n_829) );
BUFx12f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NOR2x1p5_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_107), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
AND3x2_ASAP7_75t_L g825 ( .A(n_109), .B(n_113), .C(n_125), .Y(n_825) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g811 ( .A(n_110), .Y(n_811) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g136 ( .A(n_114), .Y(n_136) );
AO21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_127), .B(n_801), .Y(n_117) );
BUFx12f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x6_ASAP7_75t_SL g119 ( .A(n_120), .B(n_122), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g813 ( .A(n_121), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g818 ( .A(n_121), .B(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_125), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NOR2x1_ASAP7_75t_L g821 ( .A(n_124), .B(n_126), .Y(n_821) );
AND2x6_ASAP7_75t_SL g809 ( .A(n_125), .B(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
XNOR2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_131), .Y(n_127) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
OAI22xp5_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_137), .B1(n_477), .B2(n_478), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_135), .Y(n_477) );
BUFx8_ASAP7_75t_SL g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g820 ( .A(n_136), .B(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
XOR2xp5_ASAP7_75t_L g803 ( .A(n_138), .B(n_804), .Y(n_803) );
OR2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_380), .Y(n_138) );
NAND4xp25_ASAP7_75t_L g139 ( .A(n_140), .B(n_304), .C(n_335), .D(n_364), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_141), .B(n_271), .Y(n_140) );
OAI322xp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_207), .A3(n_236), .B1(n_249), .B2(n_257), .C1(n_266), .C2(n_268), .Y(n_141) );
INVxp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_143), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g143 ( .A(n_144), .B(n_177), .Y(n_143) );
AND2x2_ASAP7_75t_L g301 ( .A(n_144), .B(n_302), .Y(n_301) );
INVx4_ASAP7_75t_L g337 ( .A(n_144), .Y(n_337) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g312 ( .A(n_145), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g315 ( .A(n_145), .B(n_209), .Y(n_315) );
AND2x2_ASAP7_75t_L g332 ( .A(n_145), .B(n_225), .Y(n_332) );
AND2x2_ASAP7_75t_L g430 ( .A(n_145), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g253 ( .A(n_146), .Y(n_253) );
AND2x4_ASAP7_75t_L g436 ( .A(n_146), .B(n_431), .Y(n_436) );
AO31x2_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_152), .A3(n_168), .B(n_174), .Y(n_146) );
AO31x2_ASAP7_75t_L g260 ( .A1(n_147), .A2(n_220), .A3(n_261), .B(n_264), .Y(n_260) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_148), .A2(n_563), .B(n_566), .Y(n_562) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
AO31x2_ASAP7_75t_L g197 ( .A1(n_149), .A2(n_198), .A3(n_204), .B(n_205), .Y(n_197) );
AO31x2_ASAP7_75t_L g210 ( .A1(n_149), .A2(n_211), .A3(n_220), .B(n_222), .Y(n_210) );
AO31x2_ASAP7_75t_L g225 ( .A1(n_149), .A2(n_226), .A3(n_233), .B(n_234), .Y(n_225) );
AO31x2_ASAP7_75t_L g598 ( .A1(n_149), .A2(n_176), .A3(n_599), .B(n_602), .Y(n_598) );
BUFx10_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
BUFx10_ASAP7_75t_L g490 ( .A(n_150), .Y(n_490) );
INVx1_ASAP7_75t_L g514 ( .A(n_150), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_159), .B1(n_162), .B2(n_165), .Y(n_152) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_155), .Y(n_558) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g158 ( .A(n_156), .Y(n_158) );
INVx3_ASAP7_75t_L g164 ( .A(n_156), .Y(n_164) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_156), .Y(n_200) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_156), .Y(n_203) );
INVx1_ASAP7_75t_L g215 ( .A(n_156), .Y(n_215) );
INVx1_ASAP7_75t_L g229 ( .A(n_156), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_156), .Y(n_232) );
INVx2_ASAP7_75t_L g242 ( .A(n_156), .Y(n_242) );
INVx1_ASAP7_75t_L g244 ( .A(n_156), .Y(n_244) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_158), .B(n_508), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_159), .A2(n_188), .B(n_191), .Y(n_187) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_159), .A2(n_165), .B1(n_199), .B2(n_201), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g211 ( .A1(n_159), .A2(n_212), .B1(n_217), .B2(n_218), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g226 ( .A1(n_159), .A2(n_165), .B1(n_227), .B2(n_230), .Y(n_226) );
OAI22xp5_ASAP7_75t_L g239 ( .A1(n_159), .A2(n_240), .B1(n_243), .B2(n_245), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g261 ( .A1(n_159), .A2(n_218), .B1(n_262), .B2(n_263), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_159), .A2(n_165), .B1(n_281), .B2(n_282), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_159), .A2(n_487), .B1(n_488), .B2(n_489), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_159), .A2(n_245), .B1(n_495), .B2(n_496), .Y(n_494) );
OAI22x1_ASAP7_75t_L g599 ( .A1(n_159), .A2(n_245), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx6_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
O2A1O1Ixp5_ASAP7_75t_L g183 ( .A1(n_160), .A2(n_184), .B(n_185), .C(n_186), .Y(n_183) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_160), .A2(n_545), .B(n_546), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_160), .B(n_557), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g614 ( .A1(n_160), .A2(n_553), .B(n_557), .C(n_560), .Y(n_614) );
BUFx8_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g167 ( .A(n_161), .Y(n_167) );
INVx1_ASAP7_75t_L g219 ( .A(n_161), .Y(n_219) );
INVx1_ASAP7_75t_L g510 ( .A(n_161), .Y(n_510) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx4_ASAP7_75t_L g185 ( .A(n_164), .Y(n_185) );
INVx1_ASAP7_75t_L g216 ( .A(n_164), .Y(n_216) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g489 ( .A(n_166), .Y(n_489) );
BUFx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g543 ( .A(n_167), .Y(n_543) );
AO31x2_ASAP7_75t_L g279 ( .A1(n_168), .A2(n_246), .A3(n_280), .B(n_283), .Y(n_279) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_168), .A2(n_562), .B(n_570), .Y(n_561) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
NOR2xp33_ASAP7_75t_SL g222 ( .A(n_170), .B(n_223), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_170), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g176 ( .A(n_171), .Y(n_176) );
INVx2_ASAP7_75t_L g221 ( .A(n_171), .Y(n_221) );
OAI21xp33_ASAP7_75t_L g560 ( .A1(n_171), .A2(n_514), .B(n_555), .Y(n_560) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_172), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_176), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g441 ( .A(n_177), .B(n_342), .Y(n_441) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g270 ( .A(n_178), .Y(n_270) );
INVxp67_ASAP7_75t_SL g428 ( .A(n_178), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_179), .B(n_196), .Y(n_178) );
AND2x2_ASAP7_75t_L g258 ( .A(n_179), .B(n_197), .Y(n_258) );
INVx1_ASAP7_75t_L g299 ( .A(n_179), .Y(n_299) );
OAI21x1_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_182), .B(n_194), .Y(n_179) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_180), .A2(n_182), .B(n_194), .Y(n_294) );
INVx2_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
INVx4_ASAP7_75t_L g195 ( .A(n_181), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_181), .B(n_206), .Y(n_205) );
BUFx3_ASAP7_75t_L g233 ( .A(n_181), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_181), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_181), .B(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g527 ( .A(n_181), .B(n_490), .Y(n_527) );
OAI21x1_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_187), .B(n_192), .Y(n_182) );
O2A1O1Ixp33_ASAP7_75t_L g539 ( .A1(n_185), .A2(n_540), .B(n_541), .C(n_542), .Y(n_539) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g202 ( .A(n_190), .Y(n_202) );
OAI22xp33_ASAP7_75t_L g567 ( .A1(n_190), .A2(n_232), .B1(n_568), .B2(n_569), .Y(n_567) );
INVx2_ASAP7_75t_SL g192 ( .A(n_193), .Y(n_192) );
INVx2_ASAP7_75t_SL g246 ( .A(n_193), .Y(n_246) );
INVx2_ASAP7_75t_L g204 ( .A(n_195), .Y(n_204) );
NOR2x1_ASAP7_75t_L g547 ( .A(n_195), .B(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g290 ( .A(n_196), .Y(n_290) );
AND2x2_ASAP7_75t_L g354 ( .A(n_196), .B(n_293), .Y(n_354) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g308 ( .A(n_197), .Y(n_308) );
HB1xp67_ASAP7_75t_L g361 ( .A(n_197), .Y(n_361) );
OR2x2_ASAP7_75t_L g432 ( .A(n_197), .B(n_238), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_200), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g497 ( .A(n_203), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_203), .B(n_522), .Y(n_521) );
AO31x2_ASAP7_75t_L g485 ( .A1(n_204), .A2(n_486), .A3(n_490), .B(n_491), .Y(n_485) );
NAND4xp25_ASAP7_75t_L g310 ( .A(n_207), .B(n_311), .C(n_314), .D(n_316), .Y(n_310) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
AND2x2_ASAP7_75t_L g448 ( .A(n_208), .B(n_436), .Y(n_448) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_224), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_209), .B(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g302 ( .A(n_209), .B(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g322 ( .A(n_209), .Y(n_322) );
INVx1_ASAP7_75t_L g339 ( .A(n_209), .Y(n_339) );
INVx1_ASAP7_75t_L g347 ( .A(n_209), .Y(n_347) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_209), .Y(n_461) );
INVx4_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_210), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g379 ( .A(n_210), .B(n_279), .Y(n_379) );
AND2x2_ASAP7_75t_L g387 ( .A(n_210), .B(n_225), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_210), .B(n_410), .Y(n_409) );
BUFx2_ASAP7_75t_L g452 ( .A(n_210), .Y(n_452) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_215), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g245 ( .A(n_219), .Y(n_245) );
AO31x2_ASAP7_75t_L g493 ( .A1(n_220), .A2(n_246), .A3(n_494), .B(n_498), .Y(n_493) );
AOI21x1_ASAP7_75t_L g502 ( .A1(n_220), .A2(n_503), .B(n_515), .Y(n_502) );
BUFx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_221), .B(n_492), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_221), .B(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g571 ( .A(n_221), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_221), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g256 ( .A(n_225), .Y(n_256) );
OR2x2_ASAP7_75t_L g317 ( .A(n_225), .B(n_279), .Y(n_317) );
INVx2_ASAP7_75t_L g324 ( .A(n_225), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_225), .B(n_277), .Y(n_348) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_225), .Y(n_435) );
OAI21xp33_ASAP7_75t_SL g519 ( .A1(n_228), .A2(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AO31x2_ASAP7_75t_L g238 ( .A1(n_233), .A2(n_239), .A3(n_246), .B(n_247), .Y(n_238) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_236), .B(n_407), .Y(n_406) );
BUFx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g259 ( .A(n_238), .B(n_260), .Y(n_259) );
BUFx2_ASAP7_75t_L g269 ( .A(n_238), .Y(n_269) );
INVx2_ASAP7_75t_L g287 ( .A(n_238), .Y(n_287) );
AND2x4_ASAP7_75t_L g319 ( .A(n_238), .B(n_291), .Y(n_319) );
OR2x2_ASAP7_75t_L g399 ( .A(n_238), .B(n_299), .Y(n_399) );
INVx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_242), .B(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_245), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_250), .B(n_254), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_251), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g316 ( .A(n_251), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_251), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_252), .B(n_322), .Y(n_330) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g275 ( .A(n_253), .Y(n_275) );
OR2x2_ASAP7_75t_L g368 ( .A(n_253), .B(n_278), .Y(n_368) );
INVx1_ASAP7_75t_L g295 ( .A(n_254), .Y(n_295) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g267 ( .A(n_255), .Y(n_267) );
INVx1_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
OAI322xp33_ASAP7_75t_L g271 ( .A1(n_258), .A2(n_272), .A3(n_285), .B1(n_288), .B2(n_295), .C1(n_296), .C2(n_300), .Y(n_271) );
AND2x4_ASAP7_75t_L g318 ( .A(n_258), .B(n_319), .Y(n_318) );
AOI211xp5_ASAP7_75t_SL g349 ( .A1(n_258), .A2(n_350), .B(n_351), .C(n_355), .Y(n_349) );
AND2x2_ASAP7_75t_L g369 ( .A(n_258), .B(n_259), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_258), .B(n_286), .Y(n_375) );
AND2x4_ASAP7_75t_SL g297 ( .A(n_259), .B(n_298), .Y(n_297) );
NAND3xp33_ASAP7_75t_L g388 ( .A(n_259), .B(n_315), .C(n_343), .Y(n_388) );
AND2x2_ASAP7_75t_L g419 ( .A(n_259), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g286 ( .A(n_260), .B(n_287), .Y(n_286) );
INVx3_ASAP7_75t_L g291 ( .A(n_260), .Y(n_291) );
BUFx2_ASAP7_75t_L g359 ( .A(n_260), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_269), .B(n_293), .Y(n_292) );
NAND2x1_ASAP7_75t_L g333 ( .A(n_269), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g352 ( .A(n_269), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_270), .B(n_286), .Y(n_417) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_276), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g360 ( .A(n_275), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
AND2x4_ASAP7_75t_L g323 ( .A(n_279), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g410 ( .A(n_279), .Y(n_410) );
INVx2_ASAP7_75t_L g431 ( .A(n_279), .Y(n_431) );
OAI22xp33_ASAP7_75t_L g443 ( .A1(n_285), .A2(n_444), .B1(n_446), .B2(n_447), .Y(n_443) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g355 ( .A(n_286), .B(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_L g309 ( .A(n_287), .B(n_293), .Y(n_309) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
INVx1_ASAP7_75t_L g328 ( .A(n_289), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x4_ASAP7_75t_L g298 ( .A(n_290), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g420 ( .A(n_290), .Y(n_420) );
INVx2_ASAP7_75t_L g306 ( .A(n_291), .Y(n_306) );
AND2x2_ASAP7_75t_L g334 ( .A(n_291), .B(n_293), .Y(n_334) );
INVx3_ASAP7_75t_L g342 ( .A(n_291), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_291), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g327 ( .A(n_292), .Y(n_327) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g343 ( .A(n_294), .Y(n_343) );
OAI222xp33_ASAP7_75t_L g466 ( .A1(n_296), .A2(n_456), .B1(n_467), .B2(n_470), .C1(n_472), .C2(n_474), .Y(n_466) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g407 ( .A(n_298), .Y(n_407) );
AND2x2_ASAP7_75t_L g471 ( .A(n_298), .B(n_341), .Y(n_471) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_301), .B(n_392), .Y(n_391) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_310), .B1(n_318), .B2(n_320), .C(n_325), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_307), .Y(n_305) );
INVx1_ASAP7_75t_L g393 ( .A(n_306), .Y(n_393) );
INVx2_ASAP7_75t_L g455 ( .A(n_307), .Y(n_455) );
AND2x4_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx2_ASAP7_75t_L g356 ( .A(n_308), .Y(n_356) );
AND2x2_ASAP7_75t_L g392 ( .A(n_308), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g358 ( .A(n_309), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g384 ( .A(n_309), .B(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g473 ( .A(n_309), .Y(n_473) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g422 ( .A(n_313), .Y(n_422) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g445 ( .A(n_315), .B(n_323), .Y(n_445) );
AND2x2_ASAP7_75t_L g468 ( .A(n_315), .B(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g329 ( .A(n_317), .B(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g464 ( .A(n_317), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_318), .A2(n_372), .B1(n_406), .B2(n_408), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g433 ( .A1(n_318), .A2(n_434), .B(n_437), .Y(n_433) );
INVxp67_ASAP7_75t_L g350 ( .A(n_319), .Y(n_350) );
INVx2_ASAP7_75t_SL g454 ( .A(n_319), .Y(n_454) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_323), .Y(n_320) );
OR2x2_ASAP7_75t_L g367 ( .A(n_321), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g465 ( .A(n_321), .B(n_464), .Y(n_465) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g338 ( .A(n_323), .B(n_339), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_323), .B(n_347), .Y(n_363) );
INVx2_ASAP7_75t_L g390 ( .A(n_323), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B1(n_331), .B2(n_333), .Y(n_325) );
NOR2xp33_ASAP7_75t_SL g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g413 ( .A1(n_327), .A2(n_401), .B1(n_414), .B2(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g423 ( .A(n_332), .B(n_424), .Y(n_423) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_340), .B(n_344), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g404 ( .A(n_337), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_337), .B(n_387), .Y(n_415) );
INVx1_ASAP7_75t_L g373 ( .A(n_339), .Y(n_373) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_341), .B(n_354), .Y(n_446) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
OAI21xp33_ASAP7_75t_L g459 ( .A1(n_342), .A2(n_460), .B(n_462), .Y(n_459) );
OAI21xp5_ASAP7_75t_SL g344 ( .A1(n_345), .A2(n_349), .B(n_357), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g403 ( .A(n_348), .Y(n_403) );
INVx1_ASAP7_75t_L g469 ( .A(n_348), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
INVx1_ASAP7_75t_L g442 ( .A(n_352), .Y(n_442) );
OR2x2_ASAP7_75t_L g453 ( .A(n_353), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_358), .B(n_360), .C(n_362), .Y(n_357) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_358), .A2(n_419), .B1(n_421), .B2(n_423), .Y(n_418) );
INVx1_ASAP7_75t_L g385 ( .A(n_359), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_360), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_363), .B(n_367), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g425 ( .A1(n_363), .A2(n_426), .B1(n_429), .B2(n_432), .C(n_433), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B(n_370), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g374 ( .A(n_368), .Y(n_374) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B1(n_376), .B2(n_831), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g457 ( .A(n_379), .B(n_435), .Y(n_457) );
NAND4xp25_ASAP7_75t_L g380 ( .A(n_381), .B(n_411), .C(n_438), .D(n_458), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_382), .B(n_394), .Y(n_381) );
OAI221xp5_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_386), .B1(n_388), .B2(n_389), .C(n_391), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_384), .A2(n_441), .B1(n_463), .B2(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g437 ( .A(n_386), .Y(n_437) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g421 ( .A(n_387), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_387), .B(n_430), .Y(n_429) );
NAND2x1_ASAP7_75t_L g474 ( .A(n_387), .B(n_475), .Y(n_474) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_389), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g396 ( .A(n_393), .B(n_397), .Y(n_396) );
OAI21xp33_ASAP7_75t_SL g394 ( .A1(n_395), .A2(n_400), .B(n_405), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g424 ( .A(n_410), .Y(n_424) );
AOI211xp5_ASAP7_75t_L g438 ( .A1(n_410), .A2(n_439), .B(n_443), .C(n_449), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_425), .Y(n_411) );
NAND2xp5_ASAP7_75t_SL g412 ( .A(n_413), .B(n_418), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g472 ( .A(n_420), .B(n_473), .Y(n_472) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx3_ASAP7_75t_L g476 ( .A(n_436), .Y(n_476) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp33_ASAP7_75t_R g449 ( .A1(n_450), .A2(n_453), .B1(n_455), .B2(n_456), .Y(n_449) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g463 ( .A(n_452), .B(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_459), .B(n_466), .Y(n_458) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g478 ( .A(n_479), .B(n_693), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_480), .B(n_635), .Y(n_479) );
NAND3xp33_ASAP7_75t_SL g480 ( .A(n_481), .B(n_572), .C(n_617), .Y(n_480) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_528), .B(n_549), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_482), .A2(n_573), .B1(n_592), .B2(n_604), .Y(n_572) );
AOI22x1_ASAP7_75t_L g697 ( .A1(n_482), .A2(n_698), .B1(n_702), .B2(n_703), .Y(n_697) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_500), .Y(n_483) );
OR2x2_ASAP7_75t_L g658 ( .A(n_484), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_493), .Y(n_484) );
OR2x2_ASAP7_75t_L g533 ( .A(n_485), .B(n_493), .Y(n_533) );
AND2x2_ASAP7_75t_L g576 ( .A(n_485), .B(n_577), .Y(n_576) );
INVx2_ASAP7_75t_SL g584 ( .A(n_485), .Y(n_584) );
BUFx2_ASAP7_75t_L g634 ( .A(n_485), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_489), .A2(n_525), .B(n_526), .Y(n_524) );
OAI21x1_ASAP7_75t_L g553 ( .A1(n_489), .A2(n_554), .B(n_555), .Y(n_553) );
INVx1_ASAP7_75t_L g548 ( .A(n_490), .Y(n_548) );
AND2x2_ASAP7_75t_L g579 ( .A(n_493), .B(n_516), .Y(n_579) );
INVx1_ASAP7_75t_L g586 ( .A(n_493), .Y(n_586) );
INVx1_ASAP7_75t_L g591 ( .A(n_493), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_493), .B(n_584), .Y(n_653) );
INVx1_ASAP7_75t_L g674 ( .A(n_493), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g744 ( .A(n_493), .B(n_577), .Y(n_744) );
INVx1_ASAP7_75t_L g637 ( .A(n_500), .Y(n_637) );
OR2x2_ASAP7_75t_L g689 ( .A(n_500), .B(n_653), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_516), .Y(n_500) );
AND2x2_ASAP7_75t_L g534 ( .A(n_501), .B(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g582 ( .A(n_501), .B(n_583), .Y(n_582) );
INVxp67_ASAP7_75t_L g588 ( .A(n_501), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_501), .B(n_531), .Y(n_665) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g577 ( .A(n_502), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_511), .B(n_514), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_507), .B(n_509), .Y(n_504) );
BUFx4f_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_510), .B(n_523), .Y(n_522) );
INVx3_ASAP7_75t_L g531 ( .A(n_516), .Y(n_531) );
INVx1_ASAP7_75t_L g631 ( .A(n_516), .Y(n_631) );
AND2x2_ASAP7_75t_L g633 ( .A(n_516), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g651 ( .A(n_516), .B(n_652), .Y(n_651) );
OR2x2_ASAP7_75t_L g673 ( .A(n_516), .B(n_674), .Y(n_673) );
NAND2x1p5_ASAP7_75t_SL g684 ( .A(n_516), .B(n_660), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_516), .B(n_591), .Y(n_774) );
AND2x4_ASAP7_75t_L g516 ( .A(n_517), .B(n_518), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_524), .B(n_527), .Y(n_518) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_534), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_529), .A2(n_713), .B1(n_714), .B2(n_716), .Y(n_712) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_530), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_530), .B(n_769), .Y(n_768) );
OR2x2_ASAP7_75t_L g791 ( .A(n_530), .B(n_649), .Y(n_791) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
AND2x4_ASAP7_75t_L g590 ( .A(n_531), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_531), .B(n_660), .Y(n_659) );
OR2x2_ASAP7_75t_L g679 ( .A(n_531), .B(n_680), .Y(n_679) );
AND2x4_ASAP7_75t_L g630 ( .A(n_532), .B(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_L g720 ( .A(n_533), .Y(n_720) );
OR2x2_ASAP7_75t_L g794 ( .A(n_533), .B(n_721), .Y(n_794) );
INVx1_ASAP7_75t_L g625 ( .A(n_534), .Y(n_625) );
INVx3_ASAP7_75t_L g629 ( .A(n_535), .Y(n_629) );
BUFx2_ASAP7_75t_L g640 ( .A(n_535), .Y(n_640) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g610 ( .A(n_536), .B(n_561), .Y(n_610) );
INVx2_ASAP7_75t_L g656 ( .A(n_536), .Y(n_656) );
INVx1_ASAP7_75t_L g688 ( .A(n_536), .Y(n_688) );
AND2x2_ASAP7_75t_L g701 ( .A(n_536), .B(n_598), .Y(n_701) );
AND2x2_ASAP7_75t_L g723 ( .A(n_536), .B(n_622), .Y(n_723) );
NAND2x1p5_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
OAI21x1_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_544), .B(n_547), .Y(n_538) );
INVx2_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g714 ( .A(n_550), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_550), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g739 ( .A(n_550), .B(n_607), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_550), .B(n_741), .Y(n_740) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_561), .Y(n_550) );
INVx2_ASAP7_75t_L g596 ( .A(n_551), .Y(n_596) );
AND2x2_ASAP7_75t_L g623 ( .A(n_551), .B(n_624), .Y(n_623) );
AOI21x1_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_556), .B(n_559), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g597 ( .A(n_561), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g616 ( .A(n_561), .Y(n_616) );
INVx2_ASAP7_75t_L g624 ( .A(n_561), .Y(n_624) );
OR2x2_ASAP7_75t_L g644 ( .A(n_561), .B(n_598), .Y(n_644) );
AND2x2_ASAP7_75t_L g655 ( .A(n_561), .B(n_656), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_578), .B1(n_580), .B2(n_585), .C(n_587), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI32xp33_ASAP7_75t_L g685 ( .A1(n_575), .A2(n_589), .A3(n_686), .B1(n_689), .B2(n_690), .Y(n_685) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g675 ( .A(n_576), .Y(n_675) );
AND2x2_ASAP7_75t_L g711 ( .A(n_576), .B(n_590), .Y(n_711) );
INVx1_ASAP7_75t_L g775 ( .A(n_576), .Y(n_775) );
OR2x2_ASAP7_75t_L g649 ( .A(n_577), .B(n_584), .Y(n_649) );
INVx2_ASAP7_75t_L g660 ( .A(n_577), .Y(n_660) );
BUFx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g799 ( .A(n_579), .B(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g786 ( .A(n_582), .Y(n_786) );
INVx1_ASAP7_75t_L g800 ( .A(n_582), .Y(n_800) );
OR2x2_ASAP7_75t_L g680 ( .A(n_583), .B(n_660), .Y(n_680) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_585), .B(n_680), .Y(n_702) );
INVx1_ASAP7_75t_L g733 ( .A(n_585), .Y(n_733) );
BUFx3_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g767 ( .A(n_586), .Y(n_767) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2x1_ASAP7_75t_L g736 ( .A(n_588), .B(n_737), .Y(n_736) );
OAI21xp5_ASAP7_75t_SL g758 ( .A1(n_589), .A2(n_759), .B(n_764), .Y(n_758) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx2_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_597), .Y(n_593) );
AND2x2_ASAP7_75t_L g668 ( .A(n_594), .B(n_610), .Y(n_668) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_594), .Y(n_798) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g700 ( .A(n_595), .Y(n_700) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g682 ( .A(n_596), .B(n_656), .Y(n_682) );
AND2x2_ASAP7_75t_L g753 ( .A(n_596), .B(n_624), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_597), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g681 ( .A(n_597), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g760 ( .A(n_597), .B(n_761), .Y(n_760) );
INVx2_ASAP7_75t_L g609 ( .A(n_598), .Y(n_609) );
INVx2_ASAP7_75t_L g622 ( .A(n_598), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_598), .B(n_613), .Y(n_670) );
AND2x2_ASAP7_75t_L g730 ( .A(n_598), .B(n_624), .Y(n_730) );
NAND2xp33_ASAP7_75t_SL g604 ( .A(n_605), .B(n_611), .Y(n_604) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g705 ( .A(n_608), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_608), .B(n_688), .Y(n_780) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OR2x2_ASAP7_75t_L g612 ( .A(n_609), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g741 ( .A(n_609), .B(n_656), .Y(n_741) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_615), .Y(n_611) );
OR2x2_ASAP7_75t_L g686 ( .A(n_612), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g643 ( .A(n_613), .Y(n_643) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g669 ( .A(n_616), .B(n_670), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_630), .B1(n_632), .B2(n_633), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_625), .B(n_626), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g632 ( .A(n_620), .B(n_629), .Y(n_632) );
BUFx2_ASAP7_75t_L g650 ( .A(n_620), .Y(n_650) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g661 ( .A(n_621), .Y(n_661) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g676 ( .A(n_623), .B(n_640), .Y(n_676) );
INVx2_ASAP7_75t_L g692 ( .A(n_623), .Y(n_692) );
AND2x2_ASAP7_75t_L g734 ( .A(n_623), .B(n_656), .Y(n_734) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g709 ( .A(n_629), .B(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g756 ( .A(n_630), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g787 ( .A(n_631), .Y(n_787) );
INVx2_ASAP7_75t_L g726 ( .A(n_634), .Y(n_726) );
NAND4xp25_ASAP7_75t_L g635 ( .A(n_636), .B(n_645), .C(n_662), .D(n_677), .Y(n_635) );
NAND2xp33_ASAP7_75t_SL g636 ( .A(n_637), .B(n_638), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g731 ( .A1(n_638), .A2(n_716), .B1(n_732), .B2(n_734), .C(n_735), .Y(n_731) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2x1_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g713 ( .A(n_642), .Y(n_713) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_644), .Y(n_642) );
INVx2_ASAP7_75t_L g706 ( .A(n_643), .Y(n_706) );
INVx2_ASAP7_75t_L g778 ( .A(n_644), .Y(n_778) );
AOI222xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B1(n_651), .B2(n_654), .C1(n_657), .C2(n_661), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g732 ( .A(n_648), .B(n_733), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g759 ( .A1(n_648), .A2(n_760), .B(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g771 ( .A(n_649), .B(n_715), .Y(n_771) );
OAI21xp33_ASAP7_75t_SL g745 ( .A1(n_650), .A2(n_671), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g664 ( .A(n_653), .B(n_665), .Y(n_664) );
INVxp67_ASAP7_75t_SL g716 ( .A(n_653), .Y(n_716) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
BUFx2_ASAP7_75t_L g715 ( .A(n_656), .Y(n_715) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g721 ( .A(n_660), .Y(n_721) );
AOI22xp33_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_666), .B1(n_671), .B2(n_676), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_668), .A2(n_678), .B1(n_681), .B2(n_683), .C(n_685), .Y(n_677) );
INVx3_ASAP7_75t_R g792 ( .A(n_669), .Y(n_792) );
INVx1_ASAP7_75t_L g710 ( .A(n_670), .Y(n_710) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
OR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_675), .Y(n_672) );
INVxp67_ASAP7_75t_SL g727 ( .A(n_673), .Y(n_727) );
INVx1_ASAP7_75t_L g737 ( .A(n_673), .Y(n_737) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_682), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g755 ( .A(n_682), .Y(n_755) );
AND2x2_ASAP7_75t_L g783 ( .A(n_682), .B(n_730), .Y(n_783) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g777 ( .A(n_687), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NOR2x1_ASAP7_75t_L g693 ( .A(n_694), .B(n_749), .Y(n_693) );
NAND3xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_731), .C(n_745), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_707), .C(n_717), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_698), .A2(n_709), .B(n_711), .Y(n_708) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g748 ( .A(n_700), .Y(n_748) );
AND2x2_ASAP7_75t_L g789 ( .A(n_700), .B(n_778), .Y(n_789) );
NAND2x1_ASAP7_75t_L g747 ( .A(n_701), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
INVx1_ASAP7_75t_L g769 ( .A(n_706), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_708), .B(n_712), .Y(n_707) );
INVx1_ASAP7_75t_L g761 ( .A(n_715), .Y(n_761) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_722), .B1(n_724), .B2(n_728), .Y(n_717) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g757 ( .A(n_721), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_723), .B(n_753), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_727), .Y(n_724) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g796 ( .A(n_729), .Y(n_796) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OAI22xp33_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_738), .B1(n_740), .B2(n_742), .Y(n_735) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx2_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_776), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_754), .B(n_756), .C(n_758), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
OAI21xp33_ASAP7_75t_L g765 ( .A1(n_752), .A2(n_766), .B(n_768), .Y(n_765) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
O2A1O1Ixp5_ASAP7_75t_SL g776 ( .A1(n_756), .A2(n_777), .B(n_779), .C(n_781), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_760), .A2(n_765), .B1(n_770), .B2(n_772), .Y(n_764) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI211xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .B(n_788), .C(n_795), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g788 ( .A1(n_789), .A2(n_790), .B1(n_792), .B2(n_793), .Y(n_788) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI21xp5_ASAP7_75t_SL g795 ( .A1(n_796), .A2(n_797), .B(n_799), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_802), .A2(n_812), .B(n_814), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_803), .B(n_807), .Y(n_802) );
BUFx2_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
BUFx8_ASAP7_75t_SL g812 ( .A(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
BUFx10_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_823), .B(n_826), .Y(n_822) );
BUFx2_ASAP7_75t_SL g823 ( .A(n_824), .Y(n_823) );
INVx4_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
NOR2xp33_ASAP7_75t_R g827 ( .A(n_828), .B(n_829), .Y(n_827) );
endmodule