module fake_jpeg_27346_n_68 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_66;

INVx3_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_SL g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_35),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_0),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_40),
.B(n_41),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_1),
.B(n_2),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_13),
.B1(n_24),
.B2(n_23),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_50),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_12),
.B1(n_22),
.B2(n_21),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_49),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_9),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_4),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_3),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_35),
.A2(n_10),
.B1(n_20),
.B2(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx24_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_4),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_5),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_53),
.C(n_60),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_58),
.C(n_62),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_64),
.A2(n_62),
.B(n_52),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_SL g66 ( 
.A(n_65),
.B(n_52),
.C(n_49),
.Y(n_66)
);

AOI322xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_5),
.A3(n_7),
.B1(n_8),
.B2(n_14),
.C1(n_15),
.C2(n_16),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_25),
.Y(n_68)
);


endmodule