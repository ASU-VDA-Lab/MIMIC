module fake_ibex_1075_n_2420 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_338, n_173, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_463, n_624, n_411, n_135, n_520, n_658, n_512, n_615, n_283, n_366, n_397, n_111, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_563, n_132, n_277, n_555, n_337, n_522, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_501, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_260, n_620, n_462, n_302, n_450, n_443, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_489, n_399, n_254, n_213, n_424, n_565, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_2420);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_338;
input n_173;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_658;
input n_512;
input n_615;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_501;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_2420;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_992;
wire n_1582;
wire n_2201;
wire n_766;
wire n_2175;
wire n_2071;
wire n_1110;
wire n_1382;
wire n_1998;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_1234;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_773;
wire n_2038;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_2074;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_802;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_2276;
wire n_1045;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2139;
wire n_1308;
wire n_1138;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_667;
wire n_884;
wire n_2396;
wire n_850;
wire n_1971;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_876;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_2343;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_2192;
wire n_1766;
wire n_1922;
wire n_2032;
wire n_1937;
wire n_2311;
wire n_893;
wire n_1654;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_824;
wire n_1945;
wire n_694;
wire n_787;
wire n_2015;
wire n_1130;
wire n_1228;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_2363;
wire n_2003;
wire n_1970;
wire n_1778;
wire n_2347;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2333;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_1955;
wire n_917;
wire n_2249;
wire n_2413;
wire n_2362;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_2090;
wire n_666;
wire n_2260;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_793;
wire n_937;
wire n_2116;
wire n_1645;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_2393;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_1445;
wire n_2283;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_2022;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_2275;
wire n_1853;
wire n_2189;
wire n_745;
wire n_2112;
wire n_1753;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2171;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_906;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_978;
wire n_899;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_2166;
wire n_2150;
wire n_695;
wire n_1549;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_2292;
wire n_2334;
wire n_1424;
wire n_2350;
wire n_1742;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_1040;
wire n_2203;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2397;
wire n_1121;
wire n_693;
wire n_2256;
wire n_737;
wire n_1571;
wire n_1980;
wire n_2019;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2355;
wire n_1543;
wire n_823;
wire n_2233;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_1441;
wire n_2028;
wire n_1924;
wire n_1921;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_2033;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1964;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_2052;
wire n_981;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_2377;
wire n_1591;
wire n_2289;
wire n_2288;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_2101;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2390;
wire n_859;
wire n_1109;
wire n_965;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_1884;
wire n_2176;
wire n_1825;
wire n_1589;
wire n_2204;
wire n_1210;
wire n_2319;
wire n_1933;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2132;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_2297;
wire n_1792;
wire n_1712;
wire n_1984;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_2006;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_669;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_938;
wire n_1178;
wire n_878;
wire n_2358;
wire n_2361;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2252;
wire n_1982;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_1695;
wire n_1418;
wire n_2402;
wire n_1137;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_1602;
wire n_1776;
wire n_2372;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_2287;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_1146;
wire n_705;
wire n_2142;
wire n_1548;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2234;
wire n_847;
wire n_1436;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_2332;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_1545;
wire n_2369;
wire n_1471;
wire n_1738;
wire n_998;
wire n_1115;
wire n_1395;
wire n_1729;
wire n_801;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2241;
wire n_1470;
wire n_2109;
wire n_2098;
wire n_1761;
wire n_1836;
wire n_2398;
wire n_1593;
wire n_986;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_927;
wire n_1563;
wire n_803;
wire n_1875;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1599;
wire n_1539;
wire n_1806;
wire n_1575;
wire n_2209;
wire n_1448;
wire n_2077;
wire n_817;
wire n_2193;
wire n_2095;
wire n_2395;
wire n_951;
wire n_2053;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2352;
wire n_863;
wire n_2185;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_1405;
wire n_997;
wire n_2308;
wire n_1428;
wire n_2243;
wire n_2400;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_2270;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_903;
wire n_1967;
wire n_2340;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_2042;
wire n_1048;
wire n_774;
wire n_1925;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_1247;
wire n_836;
wire n_1475;
wire n_1263;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_2298;
wire n_895;
wire n_687;
wire n_1035;
wire n_2045;
wire n_1535;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_1437;
wire n_1707;
wire n_1941;
wire n_2064;
wire n_1679;
wire n_2342;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_1578;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_972;
wire n_1815;
wire n_1917;
wire n_1444;
wire n_920;
wire n_1067;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_1920;
wire n_887;
wire n_1162;
wire n_1997;
wire n_1894;
wire n_2110;
wire n_961;
wire n_991;
wire n_1331;
wire n_1223;
wire n_1349;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_1777;
wire n_1353;
wire n_2386;
wire n_1429;
wire n_2029;
wire n_2026;
wire n_1546;
wire n_1432;
wire n_2103;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_2271;
wire n_2356;
wire n_1830;
wire n_2261;
wire n_1629;
wire n_2011;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_1626;
wire n_674;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_2344;
wire n_2317;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_1099;
wire n_2141;
wire n_1422;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2210;
wire n_1517;
wire n_690;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_1952;
wire n_2180;
wire n_2087;
wire n_1598;
wire n_977;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2075;
wire n_1625;
wire n_2380;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_2309;
wire n_842;
wire n_2274;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_1259;
wire n_2108;
wire n_1001;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_2196;
wire n_1538;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2351;
wire n_2049;
wire n_1456;
wire n_1889;
wire n_2113;
wire n_1124;
wire n_1690;
wire n_1673;
wire n_2018;
wire n_922;
wire n_1790;
wire n_993;
wire n_851;
wire n_2085;
wire n_1725;
wire n_2149;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_1938;
wire n_830;
wire n_1241;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_839;
wire n_768;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_2153;
wire n_1270;
wire n_834;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_2027;
wire n_2072;
wire n_2012;
wire n_722;
wire n_2251;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_1057;
wire n_1473;
wire n_2125;
wire n_1403;
wire n_2181;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_2159;
wire n_975;
wire n_675;
wire n_934;
wire n_775;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_2286;
wire n_1879;
wire n_1959;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_1261;
wire n_2299;
wire n_2078;
wire n_2265;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_2315;
wire n_2157;
wire n_1282;
wire n_2067;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_681;
wire n_1718;
wire n_2225;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2348;
wire n_786;
wire n_2417;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_1085;
wire n_2388;
wire n_2222;
wire n_1907;
wire n_885;
wire n_1530;
wire n_877;
wire n_2135;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_2232;
wire n_2121;
wire n_1893;
wire n_1570;
wire n_2231;
wire n_701;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_1256;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_1961;
wire n_1050;
wire n_2218;
wire n_1769;
wire n_2130;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1542;
wire n_1097;
wire n_1909;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_1872;
wire n_1940;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_2020;
wire n_1978;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_1585;
wire n_2316;
wire n_1861;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_1131;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_828;
wire n_1438;
wire n_1973;
wire n_2314;
wire n_2156;
wire n_753;
wire n_2126;
wire n_1147;
wire n_747;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_698;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_2266;
wire n_682;
wire n_2061;
wire n_1373;
wire n_1686;
wire n_2131;
wire n_1302;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_755;
wire n_2091;
wire n_1029;
wire n_2394;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_854;
wire n_2405;
wire n_1369;
wire n_714;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_2323;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2371;
wire n_914;
wire n_1986;
wire n_1024;
wire n_1141;
wire n_1949;
wire n_1197;
wire n_2408;
wire n_1168;
wire n_865;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2305;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_2048;
wire n_987;
wire n_1299;
wire n_750;
wire n_2096;
wire n_2129;
wire n_1101;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_1911;
wire n_2293;
wire n_731;
wire n_1336;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_2227;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2111;
wire n_2169;
wire n_1262;
wire n_1904;
wire n_1692;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_1092;
wire n_1808;
wire n_1658;
wire n_1386;
wire n_910;
wire n_2291;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_1142;
wire n_783;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2357;
wire n_924;
wire n_2331;
wire n_1600;
wire n_1661;
wire n_1965;
wire n_1757;
wire n_699;
wire n_2136;
wire n_2403;
wire n_918;
wire n_2056;
wire n_1913;
wire n_672;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2092;
wire n_1365;
wire n_1472;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_1974;
wire n_2066;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2378;
wire n_888;
wire n_1325;
wire n_2014;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_1837;
wire n_1744;
wire n_1975;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_2202;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_1468;
wire n_2327;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_1354;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_866;
wire n_1559;
wire n_2321;
wire n_1579;
wire n_1280;
wire n_1335;
wire n_2285;
wire n_1934;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_1843;
wire n_2186;
wire n_2030;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_1194;
wire n_1150;
wire n_683;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_867;
wire n_983;
wire n_1417;
wire n_2282;
wire n_970;
wire n_921;
wire n_1534;
wire n_908;
wire n_1346;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_2368;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_2065;
wire n_1743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_200),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_48),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_587),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_651),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_641),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_190),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_591),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_600),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_660),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_656),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_472),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_621),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_17),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_520),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_208),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_249),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_557),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_599),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_369),
.Y(n_684)
);

CKINVDCx20_ASAP7_75t_R g685 ( 
.A(n_100),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_585),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_620),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_609),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_414),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_69),
.Y(n_690)
);

BUFx2_ASAP7_75t_L g691 ( 
.A(n_151),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_213),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_193),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_528),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_598),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_258),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_315),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_374),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_430),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_438),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_580),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_201),
.Y(n_702)
);

BUFx5_ASAP7_75t_L g703 ( 
.A(n_435),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_306),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_596),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_64),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_647),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_646),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_369),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_623),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_515),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_586),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_289),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_583),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_96),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_187),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_440),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_237),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_336),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_296),
.Y(n_720)
);

CKINVDCx14_ASAP7_75t_R g721 ( 
.A(n_398),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_133),
.Y(n_722)
);

BUFx5_ASAP7_75t_L g723 ( 
.A(n_635),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_539),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_188),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_41),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_447),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_305),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_171),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_303),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_644),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_280),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_626),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_589),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_214),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_115),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_436),
.Y(n_737)
);

INVx2_ASAP7_75t_SL g738 ( 
.A(n_524),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_50),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_167),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_160),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_605),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_89),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_251),
.Y(n_744)
);

INVx1_ASAP7_75t_SL g745 ( 
.A(n_303),
.Y(n_745)
);

CKINVDCx20_ASAP7_75t_R g746 ( 
.A(n_202),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_631),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_401),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_657),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_596),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_161),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_628),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_582),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_649),
.Y(n_754)
);

CKINVDCx20_ASAP7_75t_R g755 ( 
.A(n_394),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_399),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_615),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_636),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_544),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_404),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_662),
.Y(n_761)
);

BUFx5_ASAP7_75t_L g762 ( 
.A(n_205),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_259),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_203),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_418),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_630),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_338),
.Y(n_767)
);

INVx4_ASAP7_75t_R g768 ( 
.A(n_648),
.Y(n_768)
);

CKINVDCx16_ASAP7_75t_R g769 ( 
.A(n_591),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_359),
.Y(n_770)
);

CKINVDCx14_ASAP7_75t_R g771 ( 
.A(n_570),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_414),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_610),
.Y(n_773)
);

HB1xp67_ASAP7_75t_L g774 ( 
.A(n_451),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_292),
.Y(n_775)
);

CKINVDCx16_ASAP7_75t_R g776 ( 
.A(n_389),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_661),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_243),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_373),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_551),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_618),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_330),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_604),
.Y(n_783)
);

BUFx10_ASAP7_75t_L g784 ( 
.A(n_496),
.Y(n_784)
);

BUFx5_ASAP7_75t_L g785 ( 
.A(n_212),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_629),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_593),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_329),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_637),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_483),
.Y(n_790)
);

BUFx5_ASAP7_75t_L g791 ( 
.A(n_193),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_588),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_655),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_636),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_361),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_622),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_471),
.Y(n_797)
);

INVx2_ASAP7_75t_SL g798 ( 
.A(n_0),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_437),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_595),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_590),
.Y(n_801)
);

INVx1_ASAP7_75t_SL g802 ( 
.A(n_209),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_348),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_483),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_320),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_639),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_567),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_605),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_479),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_237),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_619),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_519),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_568),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_581),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_477),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_625),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_584),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_453),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_148),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_634),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_597),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_25),
.Y(n_822)
);

INVx1_ASAP7_75t_SL g823 ( 
.A(n_171),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_61),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_173),
.Y(n_825)
);

INVx3_ASAP7_75t_L g826 ( 
.A(n_28),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_385),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_352),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_659),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_612),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_415),
.Y(n_831)
);

BUFx10_ASAP7_75t_L g832 ( 
.A(n_1),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_226),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_142),
.Y(n_834)
);

CKINVDCx16_ASAP7_75t_R g835 ( 
.A(n_56),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_355),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_213),
.Y(n_837)
);

CKINVDCx16_ASAP7_75t_R g838 ( 
.A(n_543),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_108),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_83),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_175),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_190),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_220),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_221),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_470),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_608),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_424),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_107),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_311),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_632),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_606),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_616),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_257),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_631),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_164),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_150),
.Y(n_856)
);

BUFx10_ASAP7_75t_L g857 ( 
.A(n_484),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_499),
.Y(n_858)
);

BUFx10_ASAP7_75t_L g859 ( 
.A(n_650),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_169),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_81),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_601),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_195),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_100),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_144),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_471),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_633),
.Y(n_867)
);

CKINVDCx20_ASAP7_75t_R g868 ( 
.A(n_59),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_623),
.Y(n_869)
);

CKINVDCx6p67_ASAP7_75t_R g870 ( 
.A(n_355),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_388),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_120),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_72),
.Y(n_873)
);

BUFx6f_ASAP7_75t_L g874 ( 
.A(n_614),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_287),
.Y(n_875)
);

CKINVDCx20_ASAP7_75t_R g876 ( 
.A(n_307),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_153),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_273),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_617),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_166),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_402),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_462),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_248),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_274),
.Y(n_884)
);

BUFx6f_ASAP7_75t_L g885 ( 
.A(n_17),
.Y(n_885)
);

CKINVDCx5p33_ASAP7_75t_R g886 ( 
.A(n_651),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_451),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_293),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_473),
.Y(n_889)
);

INVxp67_ASAP7_75t_L g890 ( 
.A(n_515),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_444),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_217),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_162),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_643),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_126),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_317),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_309),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_4),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_640),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_433),
.Y(n_900)
);

CKINVDCx16_ASAP7_75t_R g901 ( 
.A(n_624),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_77),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_481),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_642),
.Y(n_904)
);

INVx1_ASAP7_75t_SL g905 ( 
.A(n_55),
.Y(n_905)
);

HB1xp67_ASAP7_75t_L g906 ( 
.A(n_183),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_173),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_181),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_48),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_390),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_116),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_592),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_283),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_395),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_157),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_173),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_228),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_328),
.Y(n_918)
);

BUFx2_ASAP7_75t_L g919 ( 
.A(n_44),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_84),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_197),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_559),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_540),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_164),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_400),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_300),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_423),
.Y(n_927)
);

BUFx2_ASAP7_75t_SL g928 ( 
.A(n_521),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_405),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_383),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_400),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_283),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_22),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_23),
.Y(n_934)
);

CKINVDCx20_ASAP7_75t_R g935 ( 
.A(n_594),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_278),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_531),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_179),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_532),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_233),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_187),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_282),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_652),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_416),
.Y(n_944)
);

CKINVDCx20_ASAP7_75t_R g945 ( 
.A(n_613),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_611),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_607),
.Y(n_947)
);

INVx1_ASAP7_75t_SL g948 ( 
.A(n_633),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_627),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_39),
.Y(n_950)
);

INVxp33_ASAP7_75t_R g951 ( 
.A(n_602),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_377),
.Y(n_952)
);

CKINVDCx16_ASAP7_75t_R g953 ( 
.A(n_368),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_425),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_89),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_479),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_558),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_23),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_561),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_393),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_270),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_277),
.Y(n_962)
);

INVxp33_ASAP7_75t_L g963 ( 
.A(n_413),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_654),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_485),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_157),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_120),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_653),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_658),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_563),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_198),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_163),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_523),
.Y(n_973)
);

BUFx10_ASAP7_75t_L g974 ( 
.A(n_443),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_R g975 ( 
.A(n_523),
.Y(n_975)
);

CKINVDCx5p33_ASAP7_75t_R g976 ( 
.A(n_250),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_12),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_21),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_127),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_68),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_172),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_645),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_638),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_302),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_603),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_374),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_369),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_262),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_721),
.Y(n_989)
);

INVxp67_ASAP7_75t_SL g990 ( 
.A(n_963),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_670),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_776),
.B(n_0),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_721),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_870),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_774),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_771),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_670),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_771),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_685),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_798),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_896),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_907),
.Y(n_1002)
);

INVxp67_ASAP7_75t_SL g1003 ( 
.A(n_826),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_746),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_835),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_953),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_723),
.Y(n_1007)
);

INVxp67_ASAP7_75t_SL g1008 ( 
.A(n_826),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_748),
.Y(n_1009)
);

CKINVDCx20_ASAP7_75t_R g1010 ( 
.A(n_755),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_691),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_984),
.B(n_763),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_831),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_666),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_919),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_894),
.B(n_0),
.Y(n_1016)
);

CKINVDCx20_ASAP7_75t_R g1017 ( 
.A(n_834),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_855),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_667),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_707),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_679),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_L g1022 ( 
.A(n_738),
.B(n_1),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_906),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_678),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_680),
.Y(n_1025)
);

CKINVDCx20_ASAP7_75t_R g1026 ( 
.A(n_853),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_681),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_696),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_868),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_684),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_690),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_871),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_692),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_876),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_693),
.Y(n_1035)
);

INVxp67_ASAP7_75t_SL g1036 ( 
.A(n_698),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_713),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_881),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_793),
.B(n_2),
.Y(n_1039)
);

INVxp33_ASAP7_75t_SL g1040 ( 
.A(n_964),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_720),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_973),
.B(n_2),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_890),
.B(n_2),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_735),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_888),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_697),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_740),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_743),
.Y(n_1048)
);

INVxp33_ASAP7_75t_SL g1049 ( 
.A(n_700),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_914),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_R g1051 ( 
.A(n_702),
.B(n_704),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_706),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_709),
.Y(n_1053)
);

NOR2xp67_ASAP7_75t_L g1054 ( 
.A(n_744),
.B(n_3),
.Y(n_1054)
);

INVxp67_ASAP7_75t_SL g1055 ( 
.A(n_751),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_756),
.Y(n_1056)
);

HB1xp67_ASAP7_75t_L g1057 ( 
.A(n_909),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_SL g1058 ( 
.A(n_689),
.Y(n_1058)
);

CKINVDCx20_ASAP7_75t_R g1059 ( 
.A(n_958),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_765),
.Y(n_1060)
);

CKINVDCx14_ASAP7_75t_R g1061 ( 
.A(n_689),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_772),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_775),
.Y(n_1063)
);

HB1xp67_ASAP7_75t_L g1064 ( 
.A(n_909),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_961),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_778),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_779),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_799),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_715),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_717),
.Y(n_1070)
);

HB1xp67_ASAP7_75t_L g1071 ( 
.A(n_913),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_719),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_722),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_818),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_723),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_1061),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_994),
.B(n_769),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_990),
.B(n_832),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_1049),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1014),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_1019),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1057),
.Y(n_1082)
);

BUFx2_ASAP7_75t_SL g1083 ( 
.A(n_1058),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_1007),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1064),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_1075),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1071),
.Y(n_1087)
);

CKINVDCx20_ASAP7_75t_R g1088 ( 
.A(n_999),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_991),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_995),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_995),
.B(n_974),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_1024),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_1004),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1003),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1008),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_997),
.Y(n_1096)
);

OR2x6_ASAP7_75t_L g1097 ( 
.A(n_1012),
.B(n_928),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1036),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_1009),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_1011),
.B(n_707),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_1025),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_R g1102 ( 
.A(n_993),
.B(n_1005),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1055),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1001),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_1027),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1018),
.B(n_838),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1002),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1030),
.Y(n_1108)
);

CKINVDCx20_ASAP7_75t_R g1109 ( 
.A(n_1010),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_1028),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_1031),
.Y(n_1111)
);

OR2x2_ASAP7_75t_L g1112 ( 
.A(n_1023),
.B(n_901),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1037),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_1033),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1035),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_R g1116 ( 
.A(n_1006),
.B(n_727),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1041),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1046),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_1044),
.A2(n_1048),
.B(n_1047),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1013),
.B(n_913),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_1074),
.Y(n_1121)
);

OA21x2_ASAP7_75t_L g1122 ( 
.A1(n_1056),
.A2(n_716),
.B(n_671),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1015),
.B(n_986),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1060),
.Y(n_1124)
);

OA21x2_ASAP7_75t_L g1125 ( 
.A1(n_1062),
.A2(n_716),
.B(n_671),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1063),
.B(n_728),
.Y(n_1126)
);

BUFx2_ASAP7_75t_L g1127 ( 
.A(n_1052),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1066),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1067),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_1053),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1068),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_996),
.B(n_730),
.Y(n_1132)
);

AND2x6_ASAP7_75t_L g1133 ( 
.A(n_1022),
.B(n_950),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_998),
.B(n_732),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1073),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1042),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_1016),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_1072),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_1069),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1039),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1054),
.Y(n_1141)
);

CKINVDCx20_ASAP7_75t_R g1142 ( 
.A(n_1017),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_1070),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1026),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1043),
.Y(n_1145)
);

AND3x2_ASAP7_75t_L g1146 ( 
.A(n_992),
.B(n_749),
.C(n_951),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1040),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1021),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_1029),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1032),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_1065),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1034),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1038),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_1045),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1059),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1050),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1020),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_1061),
.Y(n_1158)
);

BUFx6f_ASAP7_75t_L g1159 ( 
.A(n_1007),
.Y(n_1159)
);

NOR2xp33_ASAP7_75t_L g1160 ( 
.A(n_1000),
.B(n_736),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_990),
.B(n_737),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_989),
.B(n_703),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_999),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1020),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1020),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1057),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1057),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_995),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1000),
.B(n_739),
.Y(n_1169)
);

AND3x1_ASAP7_75t_L g1170 ( 
.A(n_992),
.B(n_676),
.C(n_672),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_R g1171 ( 
.A(n_1061),
.B(n_741),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_999),
.Y(n_1172)
);

OA21x2_ASAP7_75t_L g1173 ( 
.A1(n_1007),
.A2(n_839),
.B(n_822),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_990),
.B(n_714),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1061),
.Y(n_1175)
);

INVxp67_ASAP7_75t_L g1176 ( 
.A(n_995),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_1061),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1057),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1007),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1057),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1020),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1057),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1057),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_999),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1007),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1061),
.Y(n_1186)
);

BUFx8_ASAP7_75t_L g1187 ( 
.A(n_1058),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_L g1188 ( 
.A(n_1012),
.B(n_714),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1000),
.B(n_760),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1020),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1057),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1057),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1057),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_1007),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1057),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1057),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_990),
.B(n_950),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1057),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1057),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1051),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1057),
.Y(n_1201)
);

BUFx10_ASAP7_75t_L g1202 ( 
.A(n_1076),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1137),
.A2(n_827),
.B1(n_833),
.B2(n_819),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1091),
.Y(n_1204)
);

CKINVDCx14_ASAP7_75t_R g1205 ( 
.A(n_1171),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1168),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_SL g1207 ( 
.A(n_1176),
.B(n_840),
.Y(n_1207)
);

AND2x4_ASAP7_75t_L g1208 ( 
.A(n_1097),
.B(n_987),
.Y(n_1208)
);

INVx4_ASAP7_75t_L g1209 ( 
.A(n_1158),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1080),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1112),
.B(n_699),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1122),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1181),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1106),
.B(n_669),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_L g1215 ( 
.A(n_1133),
.B(n_762),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1104),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1145),
.B(n_843),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1089),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1096),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1083),
.B(n_695),
.Y(n_1220)
);

OR2x2_ASAP7_75t_L g1221 ( 
.A(n_1081),
.B(n_718),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1136),
.A2(n_841),
.B1(n_847),
.B2(n_837),
.Y(n_1222)
);

NAND2xp33_ASAP7_75t_L g1223 ( 
.A(n_1133),
.B(n_762),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1161),
.B(n_762),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1078),
.A2(n_767),
.B1(n_770),
.B2(n_764),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1105),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1125),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_1175),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_SL g1229 ( 
.A(n_1174),
.B(n_877),
.Y(n_1229)
);

INVx4_ASAP7_75t_L g1230 ( 
.A(n_1177),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1126),
.B(n_785),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1173),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1173),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1098),
.B(n_785),
.Y(n_1234)
);

NOR2xp33_ASAP7_75t_L g1235 ( 
.A(n_1094),
.B(n_782),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1131),
.Y(n_1236)
);

BUFx10_ASAP7_75t_L g1237 ( 
.A(n_1186),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1095),
.B(n_1134),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_SL g1239 ( 
.A(n_1079),
.B(n_788),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1103),
.Y(n_1240)
);

AND3x2_ASAP7_75t_L g1241 ( 
.A(n_1156),
.B(n_892),
.C(n_668),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1119),
.Y(n_1242)
);

AOI22xp33_ASAP7_75t_L g1243 ( 
.A1(n_1082),
.A2(n_856),
.B1(n_865),
.B2(n_863),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1085),
.A2(n_872),
.B1(n_880),
.B2(n_878),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

BUFx2_ASAP7_75t_L g1246 ( 
.A(n_1127),
.Y(n_1246)
);

AOI22xp33_ASAP7_75t_L g1247 ( 
.A1(n_1087),
.A2(n_882),
.B1(n_898),
.B2(n_897),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1119),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1084),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1120),
.Y(n_1250)
);

INVx5_ASAP7_75t_L g1251 ( 
.A(n_1086),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1166),
.A2(n_805),
.B1(n_810),
.B2(n_803),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1167),
.A2(n_900),
.B1(n_911),
.B2(n_910),
.Y(n_1253)
);

OR2x2_ASAP7_75t_L g1254 ( 
.A(n_1147),
.B(n_745),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1113),
.B(n_791),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1110),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1117),
.B(n_791),
.Y(n_1257)
);

BUFx6f_ASAP7_75t_L g1258 ( 
.A(n_1200),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1086),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1124),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1159),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1128),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1178),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1180),
.Y(n_1264)
);

AND2x6_ASAP7_75t_L g1265 ( 
.A(n_1182),
.B(n_966),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1183),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1092),
.Y(n_1267)
);

AND2x6_ASAP7_75t_L g1268 ( 
.A(n_1191),
.B(n_967),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1192),
.Y(n_1269)
);

AND2x6_ASAP7_75t_L g1270 ( 
.A(n_1193),
.B(n_967),
.Y(n_1270)
);

AND2x6_ASAP7_75t_L g1271 ( 
.A(n_1195),
.B(n_1196),
.Y(n_1271)
);

AND2x6_ASAP7_75t_L g1272 ( 
.A(n_1198),
.B(n_979),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1199),
.Y(n_1273)
);

AND2x6_ASAP7_75t_L g1274 ( 
.A(n_1201),
.B(n_979),
.Y(n_1274)
);

BUFx10_ASAP7_75t_L g1275 ( 
.A(n_1101),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_1188),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1132),
.B(n_824),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1140),
.B(n_825),
.Y(n_1278)
);

INVxp67_ASAP7_75t_SL g1279 ( 
.A(n_1129),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1108),
.Y(n_1280)
);

INVx4_ASAP7_75t_L g1281 ( 
.A(n_1111),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1115),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1157),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1164),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1118),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1170),
.B(n_802),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1144),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1165),
.Y(n_1288)
);

INVxp67_ASAP7_75t_SL g1289 ( 
.A(n_1116),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1141),
.B(n_1123),
.Y(n_1290)
);

INVx5_ASAP7_75t_L g1291 ( 
.A(n_1179),
.Y(n_1291)
);

AND2x6_ASAP7_75t_L g1292 ( 
.A(n_1160),
.B(n_725),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1190),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1179),
.Y(n_1294)
);

INVx4_ASAP7_75t_SL g1295 ( 
.A(n_1151),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1169),
.A2(n_915),
.B1(n_918),
.B2(n_916),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1130),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1189),
.Y(n_1298)
);

AND2x2_ASAP7_75t_SL g1299 ( 
.A(n_1154),
.B(n_920),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1154),
.B(n_695),
.Y(n_1300)
);

INVx2_ASAP7_75t_SL g1301 ( 
.A(n_1135),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1162),
.B(n_828),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1138),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1139),
.B(n_1143),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1102),
.B(n_784),
.Y(n_1305)
);

OR2x6_ASAP7_75t_L g1306 ( 
.A(n_1152),
.B(n_712),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1077),
.Y(n_1307)
);

AND2x2_ASAP7_75t_SL g1308 ( 
.A(n_1153),
.B(n_925),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1185),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1149),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_SL g1311 ( 
.A(n_1194),
.B(n_836),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1088),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1146),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1150),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1155),
.Y(n_1315)
);

AND2x6_ASAP7_75t_L g1316 ( 
.A(n_1093),
.B(n_725),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1099),
.B(n_842),
.Y(n_1317)
);

AND2x2_ASAP7_75t_SL g1318 ( 
.A(n_1109),
.B(n_927),
.Y(n_1318)
);

NAND2xp33_ASAP7_75t_SL g1319 ( 
.A(n_1142),
.B(n_988),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1163),
.A2(n_929),
.B1(n_933),
.B2(n_931),
.Y(n_1320)
);

AND2x2_ASAP7_75t_SL g1321 ( 
.A(n_1172),
.B(n_954),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1184),
.Y(n_1322)
);

INVx5_ASAP7_75t_L g1323 ( 
.A(n_1121),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1187),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1137),
.A2(n_971),
.B1(n_980),
.B2(n_978),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_SL g1326 ( 
.A(n_1081),
.B(n_844),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1197),
.B(n_791),
.Y(n_1327)
);

INVx4_ASAP7_75t_L g1328 ( 
.A(n_1076),
.Y(n_1328)
);

BUFx10_ASAP7_75t_L g1329 ( 
.A(n_1076),
.Y(n_1329)
);

INVx1_ASAP7_75t_SL g1330 ( 
.A(n_1090),
.Y(n_1330)
);

OR2x2_ASAP7_75t_SL g1331 ( 
.A(n_1114),
.B(n_761),
.Y(n_1331)
);

INVx5_ASAP7_75t_L g1332 ( 
.A(n_1121),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1107),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1107),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1107),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1187),
.Y(n_1336)
);

AND2x6_ASAP7_75t_L g1337 ( 
.A(n_1136),
.B(n_725),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1136),
.B(n_849),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1107),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1187),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1137),
.A2(n_981),
.B1(n_861),
.B2(n_864),
.Y(n_1341)
);

AND3x1_ASAP7_75t_L g1342 ( 
.A(n_1148),
.B(n_686),
.C(n_677),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1122),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1090),
.B(n_823),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1176),
.B(n_857),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1176),
.B(n_873),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1122),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1137),
.A2(n_726),
.B1(n_729),
.B2(n_725),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1212),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1279),
.B(n_875),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1263),
.B(n_694),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1264),
.B(n_883),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1266),
.B(n_884),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1224),
.A2(n_710),
.B(n_705),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1210),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1269),
.B(n_724),
.Y(n_1356)
);

OAI221xp5_ASAP7_75t_L g1357 ( 
.A1(n_1320),
.A2(n_1211),
.B1(n_1225),
.B2(n_1244),
.C(n_1243),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1273),
.B(n_887),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1227),
.Y(n_1359)
);

OAI22xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1331),
.A2(n_945),
.B1(n_969),
.B2(n_935),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_SL g1361 ( 
.A(n_1281),
.B(n_975),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1338),
.B(n_891),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_SL g1363 ( 
.A(n_1206),
.B(n_908),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1250),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1298),
.B(n_895),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1216),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1341),
.B(n_902),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1235),
.B(n_977),
.Y(n_1368)
);

AND2x4_ASAP7_75t_SL g1369 ( 
.A(n_1275),
.B(n_857),
.Y(n_1369)
);

NAND3xp33_ASAP7_75t_L g1370 ( 
.A(n_1239),
.B(n_924),
.C(n_921),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_SL g1371 ( 
.A(n_1326),
.B(n_926),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_1204),
.B(n_1214),
.Y(n_1372)
);

BUFx8_ASAP7_75t_L g1373 ( 
.A(n_1324),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_1347),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1221),
.B(n_938),
.Y(n_1375)
);

AND2x6_ASAP7_75t_L g1376 ( 
.A(n_1242),
.B(n_726),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_SL g1377 ( 
.A(n_1344),
.B(n_930),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1265),
.B(n_932),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1268),
.B(n_976),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1254),
.B(n_934),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_L g1381 ( 
.A(n_1345),
.B(n_936),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1268),
.B(n_940),
.Y(n_1382)
);

NAND2xp33_ASAP7_75t_L g1383 ( 
.A(n_1347),
.B(n_942),
.Y(n_1383)
);

CKINVDCx20_ASAP7_75t_R g1384 ( 
.A(n_1226),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1343),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_L g1386 ( 
.A(n_1317),
.B(n_944),
.C(n_905),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1246),
.B(n_962),
.Y(n_1387)
);

NOR2xp33_ASAP7_75t_SL g1388 ( 
.A(n_1282),
.B(n_952),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1270),
.B(n_955),
.Y(n_1389)
);

BUFx8_ASAP7_75t_L g1390 ( 
.A(n_1340),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1272),
.B(n_960),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1274),
.B(n_1203),
.Y(n_1392)
);

NAND2xp33_ASAP7_75t_L g1393 ( 
.A(n_1274),
.B(n_723),
.Y(n_1393)
);

BUFx5_ASAP7_75t_L g1394 ( 
.A(n_1248),
.Y(n_1394)
);

NOR2xp33_ASAP7_75t_L g1395 ( 
.A(n_1346),
.B(n_673),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1333),
.Y(n_1396)
);

INVx8_ASAP7_75t_L g1397 ( 
.A(n_1220),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1334),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1325),
.B(n_674),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1232),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1222),
.B(n_675),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1233),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1271),
.B(n_682),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1335),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1331),
.A2(n_687),
.B1(n_688),
.B2(n_683),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1336),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1271),
.A2(n_726),
.B1(n_795),
.B2(n_729),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1220),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1339),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1297),
.B(n_701),
.Y(n_1410)
);

NOR2xp33_ASAP7_75t_L g1411 ( 
.A(n_1245),
.B(n_708),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1277),
.B(n_711),
.Y(n_1412)
);

BUFx6f_ASAP7_75t_L g1413 ( 
.A(n_1337),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1267),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1287),
.Y(n_1415)
);

O2A1O1Ixp33_ASAP7_75t_L g1416 ( 
.A1(n_1229),
.A2(n_1290),
.B(n_1207),
.C(n_1252),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1256),
.Y(n_1417)
);

BUFx12f_ASAP7_75t_L g1418 ( 
.A(n_1202),
.Y(n_1418)
);

NOR2xp67_ASAP7_75t_L g1419 ( 
.A(n_1209),
.B(n_3),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1247),
.B(n_731),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1253),
.B(n_1296),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1260),
.Y(n_1422)
);

NOR2xp33_ASAP7_75t_L g1423 ( 
.A(n_1276),
.B(n_747),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1262),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1300),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1218),
.B(n_752),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1219),
.B(n_753),
.Y(n_1427)
);

OR2x6_ASAP7_75t_L g1428 ( 
.A(n_1301),
.B(n_742),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1234),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_R g1430 ( 
.A(n_1205),
.B(n_759),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1323),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1258),
.B(n_766),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1280),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1327),
.B(n_773),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1308),
.A2(n_729),
.B1(n_848),
.B2(n_795),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1342),
.A2(n_780),
.B1(n_781),
.B2(n_777),
.Y(n_1436)
);

O2A1O1Ixp5_ASAP7_75t_L g1437 ( 
.A1(n_1311),
.A2(n_794),
.B(n_809),
.C(n_787),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1305),
.B(n_783),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1231),
.B(n_1283),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1284),
.B(n_786),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1288),
.B(n_789),
.Y(n_1441)
);

AND2x2_ASAP7_75t_SL g1442 ( 
.A(n_1318),
.B(n_768),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1255),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1293),
.B(n_796),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1257),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1295),
.B(n_733),
.Y(n_1446)
);

O2A1O1Ixp5_ASAP7_75t_L g1447 ( 
.A1(n_1217),
.A2(n_794),
.B(n_809),
.C(n_787),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1285),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1215),
.A2(n_757),
.B(n_754),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1278),
.B(n_800),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1323),
.B(n_801),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1315),
.B(n_1213),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_SL g1453 ( 
.A(n_1323),
.B(n_804),
.Y(n_1453)
);

INVxp67_ASAP7_75t_SL g1454 ( 
.A(n_1208),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1303),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1312),
.A2(n_811),
.B1(n_812),
.B2(n_807),
.Y(n_1456)
);

INVx8_ASAP7_75t_L g1457 ( 
.A(n_1316),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1286),
.B(n_813),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_SL g1459 ( 
.A(n_1332),
.B(n_815),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1292),
.A2(n_848),
.B1(n_860),
.B2(n_795),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1307),
.B(n_816),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1295),
.B(n_758),
.Y(n_1462)
);

AOI22xp5_ASAP7_75t_L g1463 ( 
.A1(n_1289),
.A2(n_1299),
.B1(n_1304),
.B2(n_1223),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_R g1464 ( 
.A(n_1319),
.B(n_820),
.Y(n_1464)
);

INVxp67_ASAP7_75t_SL g1465 ( 
.A(n_1314),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1313),
.B(n_829),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1302),
.B(n_821),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1251),
.B(n_830),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1316),
.A2(n_885),
.B1(n_893),
.B2(n_860),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1236),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1348),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_SL g1472 ( 
.A(n_1251),
.B(n_845),
.Y(n_1472)
);

NOR2x1p5_ASAP7_75t_L g1473 ( 
.A(n_1230),
.B(n_970),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1321),
.B(n_859),
.Y(n_1474)
);

CKINVDCx5p33_ASAP7_75t_R g1475 ( 
.A(n_1228),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_SL g1476 ( 
.A(n_1291),
.B(n_846),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_SL g1477 ( 
.A(n_1291),
.B(n_851),
.Y(n_1477)
);

INVx3_ASAP7_75t_L g1478 ( 
.A(n_1249),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1306),
.A2(n_792),
.B1(n_797),
.B2(n_790),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1306),
.A2(n_854),
.B1(n_862),
.B2(n_858),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1259),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1261),
.B(n_867),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1294),
.B(n_869),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1310),
.B(n_1328),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1309),
.A2(n_893),
.B1(n_917),
.B2(n_885),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1241),
.B(n_879),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1237),
.B(n_1329),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1322),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1279),
.B(n_886),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_1347),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1210),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1347),
.Y(n_1492)
);

OR2x2_ASAP7_75t_L g1493 ( 
.A(n_1330),
.B(n_817),
.Y(n_1493)
);

INVx3_ASAP7_75t_L g1494 ( 
.A(n_1323),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1279),
.B(n_912),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1279),
.B(n_923),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1238),
.A2(n_917),
.B1(n_941),
.B2(n_893),
.Y(n_1497)
);

OAI22xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1331),
.A2(n_939),
.B1(n_943),
.B2(n_937),
.Y(n_1498)
);

AO22x1_ASAP7_75t_L g1499 ( 
.A1(n_1316),
.A2(n_947),
.B1(n_949),
.B2(n_946),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1240),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1330),
.B(n_948),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1238),
.A2(n_941),
.B1(n_972),
.B2(n_917),
.Y(n_1502)
);

INVx3_ASAP7_75t_L g1503 ( 
.A(n_1323),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1238),
.A2(n_941),
.B1(n_972),
.B2(n_917),
.Y(n_1504)
);

O2A1O1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1211),
.A2(n_808),
.B(n_814),
.C(n_806),
.Y(n_1505)
);

INVx8_ASAP7_75t_L g1506 ( 
.A(n_1220),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1330),
.A2(n_957),
.B1(n_965),
.B2(n_956),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1330),
.B(n_968),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1330),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1373),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_1374),
.Y(n_1511)
);

INVx4_ASAP7_75t_L g1512 ( 
.A(n_1397),
.Y(n_1512)
);

AND2x2_ASAP7_75t_SL g1513 ( 
.A(n_1361),
.B(n_941),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1402),
.A2(n_852),
.B(n_850),
.Y(n_1514)
);

INVx3_ASAP7_75t_L g1515 ( 
.A(n_1431),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1500),
.B(n_866),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1388),
.B(n_985),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1384),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1433),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1454),
.B(n_889),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_SL g1521 ( 
.A(n_1448),
.B(n_972),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1377),
.B(n_1375),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1416),
.A2(n_903),
.B(n_904),
.C(n_899),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1380),
.B(n_922),
.Y(n_1524)
);

NAND2x1p5_ASAP7_75t_L g1525 ( 
.A(n_1355),
.B(n_1491),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1471),
.A2(n_983),
.B(n_982),
.Y(n_1526)
);

INVx2_ASAP7_75t_SL g1527 ( 
.A(n_1373),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1397),
.Y(n_1528)
);

OR2x6_ASAP7_75t_SL g1529 ( 
.A(n_1415),
.B(n_5),
.Y(n_1529)
);

CKINVDCx10_ASAP7_75t_R g1530 ( 
.A(n_1390),
.Y(n_1530)
);

NOR3xp33_ASAP7_75t_L g1531 ( 
.A(n_1405),
.B(n_6),
.C(n_5),
.Y(n_1531)
);

NAND2x1p5_ASAP7_75t_L g1532 ( 
.A(n_1406),
.B(n_734),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1366),
.B(n_4),
.Y(n_1533)
);

O2A1O1Ixp5_ASAP7_75t_L g1534 ( 
.A1(n_1437),
.A2(n_874),
.B(n_959),
.C(n_750),
.Y(n_1534)
);

AOI21x1_ASAP7_75t_L g1535 ( 
.A1(n_1359),
.A2(n_874),
.B(n_750),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1364),
.B(n_4),
.Y(n_1536)
);

NOR2xp33_ASAP7_75t_SL g1537 ( 
.A(n_1418),
.B(n_750),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1381),
.A2(n_1372),
.B1(n_1498),
.B2(n_1465),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1350),
.B(n_6),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1493),
.B(n_1501),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1351),
.B(n_7),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1351),
.B(n_8),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1356),
.B(n_9),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1387),
.B(n_10),
.Y(n_1544)
);

INVx5_ASAP7_75t_L g1545 ( 
.A(n_1457),
.Y(n_1545)
);

OAI321xp33_ASAP7_75t_L g1546 ( 
.A1(n_1360),
.A2(n_1435),
.A3(n_1479),
.B1(n_1502),
.B2(n_1504),
.C(n_1497),
.Y(n_1546)
);

BUFx6f_ASAP7_75t_L g1547 ( 
.A(n_1374),
.Y(n_1547)
);

A2O1A1Ixp33_ASAP7_75t_L g1548 ( 
.A1(n_1354),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_1548)
);

AOI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1474),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1392),
.A2(n_19),
.B1(n_16),
.B2(n_18),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1390),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1425),
.B(n_19),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1365),
.B(n_20),
.Y(n_1553)
);

OAI21x1_ASAP7_75t_L g1554 ( 
.A1(n_1385),
.A2(n_465),
.B(n_464),
.Y(n_1554)
);

AO21x1_ASAP7_75t_L g1555 ( 
.A1(n_1393),
.A2(n_465),
.B(n_464),
.Y(n_1555)
);

INVx3_ASAP7_75t_L g1556 ( 
.A(n_1431),
.Y(n_1556)
);

AOI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1442),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1352),
.B(n_24),
.Y(n_1558)
);

BUFx6f_ASAP7_75t_L g1559 ( 
.A(n_1374),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_1428),
.Y(n_1560)
);

BUFx4f_ASAP7_75t_L g1561 ( 
.A(n_1506),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1353),
.B(n_1358),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1456),
.B(n_27),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1443),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1396),
.Y(n_1565)
);

OAI21xp5_ASAP7_75t_L g1566 ( 
.A1(n_1445),
.A2(n_30),
.B(n_31),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1505),
.B(n_1362),
.Y(n_1567)
);

AOI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1438),
.A2(n_34),
.B1(n_32),
.B2(n_33),
.Y(n_1568)
);

BUFx6f_ASAP7_75t_L g1569 ( 
.A(n_1490),
.Y(n_1569)
);

A2O1A1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1449),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1570)
);

BUFx6f_ASAP7_75t_L g1571 ( 
.A(n_1490),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_1475),
.Y(n_1572)
);

AOI21xp5_ASAP7_75t_L g1573 ( 
.A1(n_1368),
.A2(n_38),
.B(n_39),
.Y(n_1573)
);

A2O1A1Ixp33_ASAP7_75t_L g1574 ( 
.A1(n_1447),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1408),
.B(n_43),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1463),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_SL g1577 ( 
.A(n_1414),
.B(n_44),
.Y(n_1577)
);

OA22x2_ASAP7_75t_L g1578 ( 
.A1(n_1480),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.Y(n_1578)
);

AOI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1488),
.A2(n_50),
.B1(n_47),
.B2(n_49),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1490),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1470),
.A2(n_49),
.B(n_50),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1398),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1404),
.B(n_1409),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1417),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1363),
.B(n_51),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1422),
.B(n_52),
.Y(n_1586)
);

AOI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1434),
.A2(n_53),
.B(n_54),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1424),
.B(n_53),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1489),
.B(n_54),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1367),
.A2(n_57),
.B(n_58),
.Y(n_1590)
);

INVx1_ASAP7_75t_SL g1591 ( 
.A(n_1484),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1495),
.B(n_60),
.Y(n_1592)
);

BUFx2_ASAP7_75t_L g1593 ( 
.A(n_1430),
.Y(n_1593)
);

AND3x2_ASAP7_75t_L g1594 ( 
.A(n_1487),
.B(n_61),
.C(n_62),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_SL g1595 ( 
.A(n_1457),
.B(n_62),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1464),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1496),
.B(n_63),
.Y(n_1597)
);

INVx3_ASAP7_75t_SL g1598 ( 
.A(n_1455),
.Y(n_1598)
);

AO21x1_ASAP7_75t_L g1599 ( 
.A1(n_1383),
.A2(n_467),
.B(n_466),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1507),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1492),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1473),
.B(n_69),
.Y(n_1602)
);

AOI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1426),
.A2(n_1427),
.B(n_1482),
.Y(n_1603)
);

AO32x2_ASAP7_75t_L g1604 ( 
.A1(n_1394),
.A2(n_72),
.A3(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_1369),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1436),
.Y(n_1606)
);

INVxp67_ASAP7_75t_L g1607 ( 
.A(n_1432),
.Y(n_1607)
);

AOI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1483),
.A2(n_74),
.B(n_75),
.Y(n_1608)
);

AOI21xp5_ASAP7_75t_L g1609 ( 
.A1(n_1440),
.A2(n_76),
.B(n_77),
.Y(n_1609)
);

AOI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1499),
.A2(n_76),
.B(n_78),
.Y(n_1610)
);

AOI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1441),
.A2(n_78),
.B(n_79),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_SL g1612 ( 
.A(n_1370),
.B(n_79),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1494),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1444),
.A2(n_79),
.B(n_80),
.Y(n_1614)
);

INVx8_ASAP7_75t_L g1615 ( 
.A(n_1376),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_SL g1616 ( 
.A(n_1413),
.B(n_82),
.Y(n_1616)
);

BUFx6f_ASAP7_75t_L g1617 ( 
.A(n_1413),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_SL g1618 ( 
.A(n_1378),
.B(n_84),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1379),
.B(n_86),
.Y(n_1619)
);

OR2x6_ASAP7_75t_L g1620 ( 
.A(n_1419),
.B(n_85),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1371),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1382),
.B(n_88),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1401),
.B(n_87),
.Y(n_1623)
);

NAND2x1p5_ASAP7_75t_L g1624 ( 
.A(n_1494),
.B(n_1503),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1467),
.A2(n_90),
.B(n_91),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1420),
.B(n_90),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1399),
.B(n_92),
.Y(n_1627)
);

O2A1O1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1486),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_1628)
);

BUFx12f_ASAP7_75t_L g1629 ( 
.A(n_1446),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1395),
.B(n_94),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1412),
.B(n_96),
.Y(n_1631)
);

O2A1O1Ixp5_ASAP7_75t_L g1632 ( 
.A1(n_1468),
.A2(n_99),
.B(n_97),
.C(n_98),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1389),
.B(n_1391),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1462),
.Y(n_1634)
);

INVx3_ASAP7_75t_SL g1635 ( 
.A(n_1462),
.Y(n_1635)
);

AOI21xp5_ASAP7_75t_L g1636 ( 
.A1(n_1478),
.A2(n_101),
.B(n_102),
.Y(n_1636)
);

O2A1O1Ixp5_ASAP7_75t_L g1637 ( 
.A1(n_1472),
.A2(n_105),
.B(n_103),
.C(n_104),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1481),
.A2(n_104),
.B(n_105),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1403),
.A2(n_1452),
.B1(n_1407),
.B2(n_1458),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1466),
.B(n_106),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1376),
.Y(n_1641)
);

AOI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1450),
.A2(n_109),
.B(n_110),
.Y(n_1642)
);

AOI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1476),
.A2(n_111),
.B(n_112),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1508),
.B(n_111),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1485),
.A2(n_1423),
.B(n_1451),
.Y(n_1645)
);

AOI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1477),
.A2(n_112),
.B(n_113),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1469),
.A2(n_114),
.B1(n_112),
.B2(n_113),
.Y(n_1647)
);

AOI21x1_ASAP7_75t_L g1648 ( 
.A1(n_1453),
.A2(n_115),
.B(n_116),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1411),
.B(n_117),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1459),
.Y(n_1650)
);

NOR2xp33_ASAP7_75t_L g1651 ( 
.A(n_1461),
.B(n_117),
.Y(n_1651)
);

NAND3xp33_ASAP7_75t_L g1652 ( 
.A(n_1460),
.B(n_118),
.C(n_119),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1410),
.B(n_118),
.Y(n_1653)
);

CKINVDCx10_ASAP7_75t_R g1654 ( 
.A(n_1373),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1421),
.B(n_119),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1386),
.B(n_121),
.C(n_122),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1388),
.B(n_123),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1421),
.B(n_123),
.Y(n_1658)
);

CKINVDCx20_ASAP7_75t_R g1659 ( 
.A(n_1384),
.Y(n_1659)
);

AOI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1439),
.A2(n_124),
.B(n_125),
.Y(n_1660)
);

AND2x4_ASAP7_75t_L g1661 ( 
.A(n_1509),
.B(n_126),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1421),
.B(n_127),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1421),
.B(n_128),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1392),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1392),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.Y(n_1665)
);

INVx3_ASAP7_75t_L g1666 ( 
.A(n_1431),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1439),
.A2(n_131),
.B(n_132),
.Y(n_1667)
);

NAND2xp33_ASAP7_75t_L g1668 ( 
.A(n_1394),
.B(n_132),
.Y(n_1668)
);

CKINVDCx5p33_ASAP7_75t_R g1669 ( 
.A(n_1418),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1400),
.A2(n_469),
.B(n_468),
.Y(n_1670)
);

AO22x1_ASAP7_75t_L g1671 ( 
.A1(n_1373),
.A2(n_136),
.B1(n_137),
.B2(n_135),
.Y(n_1671)
);

NOR2xp67_ASAP7_75t_L g1672 ( 
.A(n_1509),
.B(n_134),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1397),
.Y(n_1673)
);

OAI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1392),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_1674)
);

OAI321xp33_ASAP7_75t_L g1675 ( 
.A1(n_1360),
.A2(n_141),
.A3(n_143),
.B1(n_139),
.B2(n_140),
.C(n_142),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1357),
.B(n_139),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1349),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1421),
.B(n_144),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1439),
.A2(n_145),
.B(n_146),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1421),
.B(n_145),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1421),
.B(n_146),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1349),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1392),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_1683)
);

AND2x2_ASAP7_75t_SL g1684 ( 
.A(n_1361),
.B(n_149),
.Y(n_1684)
);

NAND2x1p5_ASAP7_75t_L g1685 ( 
.A(n_1433),
.B(n_152),
.Y(n_1685)
);

AOI21xp5_ASAP7_75t_L g1686 ( 
.A1(n_1439),
.A2(n_154),
.B(n_155),
.Y(n_1686)
);

OAI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1429),
.A2(n_156),
.B(n_157),
.Y(n_1687)
);

NOR2xp67_ASAP7_75t_L g1688 ( 
.A(n_1509),
.B(n_156),
.Y(n_1688)
);

OAI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1429),
.A2(n_158),
.B(n_159),
.Y(n_1689)
);

HB1xp67_ASAP7_75t_L g1690 ( 
.A(n_1509),
.Y(n_1690)
);

CKINVDCx10_ASAP7_75t_R g1691 ( 
.A(n_1373),
.Y(n_1691)
);

INVx4_ASAP7_75t_L g1692 ( 
.A(n_1397),
.Y(n_1692)
);

AOI21xp5_ASAP7_75t_L g1693 ( 
.A1(n_1439),
.A2(n_159),
.B(n_160),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1509),
.B(n_161),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1509),
.B(n_163),
.Y(n_1695)
);

CKINVDCx10_ASAP7_75t_R g1696 ( 
.A(n_1373),
.Y(n_1696)
);

OAI321xp33_ASAP7_75t_L g1697 ( 
.A1(n_1360),
.A2(n_165),
.A3(n_168),
.B1(n_163),
.B2(n_164),
.C(n_167),
.Y(n_1697)
);

BUFx8_ASAP7_75t_SL g1698 ( 
.A(n_1418),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1439),
.A2(n_165),
.B(n_168),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1374),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1349),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_SL g1702 ( 
.A(n_1361),
.B(n_169),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1439),
.A2(n_170),
.B(n_171),
.Y(n_1703)
);

INVx3_ASAP7_75t_L g1704 ( 
.A(n_1431),
.Y(n_1704)
);

OAI21xp5_ASAP7_75t_L g1705 ( 
.A1(n_1429),
.A2(n_172),
.B(n_174),
.Y(n_1705)
);

INVx4_ASAP7_75t_L g1706 ( 
.A(n_1397),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1439),
.A2(n_175),
.B(n_176),
.Y(n_1707)
);

NOR2xp67_ASAP7_75t_L g1708 ( 
.A(n_1509),
.B(n_175),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_SL g1709 ( 
.A(n_1388),
.B(n_177),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1439),
.A2(n_176),
.B(n_177),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1349),
.Y(n_1711)
);

AOI21xp5_ASAP7_75t_L g1712 ( 
.A1(n_1439),
.A2(n_178),
.B(n_179),
.Y(n_1712)
);

AOI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1439),
.A2(n_178),
.B(n_180),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_SL g1714 ( 
.A(n_1361),
.B(n_182),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1509),
.B(n_184),
.Y(n_1715)
);

AOI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1357),
.A2(n_188),
.B1(n_185),
.B2(n_186),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1357),
.B(n_186),
.Y(n_1717)
);

NOR2xp33_ASAP7_75t_L g1718 ( 
.A(n_1357),
.B(n_189),
.Y(n_1718)
);

INVx2_ASAP7_75t_SL g1719 ( 
.A(n_1373),
.Y(n_1719)
);

AO22x1_ASAP7_75t_L g1720 ( 
.A1(n_1373),
.A2(n_192),
.B1(n_193),
.B2(n_191),
.Y(n_1720)
);

INVx2_ASAP7_75t_SL g1721 ( 
.A(n_1373),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1349),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1374),
.Y(n_1723)
);

NOR2xp33_ASAP7_75t_L g1724 ( 
.A(n_1357),
.B(n_194),
.Y(n_1724)
);

BUFx6f_ASAP7_75t_L g1725 ( 
.A(n_1374),
.Y(n_1725)
);

AND2x4_ASAP7_75t_L g1726 ( 
.A(n_1509),
.B(n_195),
.Y(n_1726)
);

INVx3_ASAP7_75t_L g1727 ( 
.A(n_1431),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1388),
.B(n_196),
.Y(n_1728)
);

BUFx6f_ASAP7_75t_L g1729 ( 
.A(n_1374),
.Y(n_1729)
);

BUFx12f_ASAP7_75t_L g1730 ( 
.A(n_1373),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1388),
.B(n_200),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1421),
.B(n_199),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_L g1733 ( 
.A(n_1394),
.B(n_202),
.Y(n_1733)
);

NAND2x1p5_ASAP7_75t_L g1734 ( 
.A(n_1433),
.B(n_201),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1349),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_1374),
.Y(n_1736)
);

NAND3xp33_ASAP7_75t_L g1737 ( 
.A(n_1386),
.B(n_203),
.C(n_204),
.Y(n_1737)
);

BUFx3_ASAP7_75t_L g1738 ( 
.A(n_1373),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1509),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.Y(n_1739)
);

O2A1O1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1357),
.A2(n_208),
.B(n_206),
.C(n_207),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1421),
.B(n_209),
.Y(n_1741)
);

NOR2xp33_ASAP7_75t_L g1742 ( 
.A(n_1357),
.B(n_210),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1357),
.B(n_211),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1388),
.B(n_212),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1429),
.A2(n_214),
.B(n_215),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1421),
.B(n_216),
.Y(n_1746)
);

NAND3xp33_ASAP7_75t_L g1747 ( 
.A(n_1386),
.B(n_218),
.C(n_219),
.Y(n_1747)
);

BUFx5_ASAP7_75t_L g1748 ( 
.A(n_1376),
.Y(n_1748)
);

BUFx6f_ASAP7_75t_L g1749 ( 
.A(n_1374),
.Y(n_1749)
);

BUFx6f_ASAP7_75t_L g1750 ( 
.A(n_1374),
.Y(n_1750)
);

AND2x4_ASAP7_75t_L g1751 ( 
.A(n_1509),
.B(n_222),
.Y(n_1751)
);

AOI21xp5_ASAP7_75t_L g1752 ( 
.A1(n_1439),
.A2(n_223),
.B(n_224),
.Y(n_1752)
);

AOI21xp5_ASAP7_75t_L g1753 ( 
.A1(n_1439),
.A2(n_223),
.B(n_224),
.Y(n_1753)
);

AOI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1439),
.A2(n_225),
.B(n_226),
.Y(n_1754)
);

AOI21xp5_ASAP7_75t_L g1755 ( 
.A1(n_1439),
.A2(n_225),
.B(n_227),
.Y(n_1755)
);

INVx3_ASAP7_75t_L g1756 ( 
.A(n_1431),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1416),
.A2(n_230),
.B(n_228),
.C(n_229),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1509),
.A2(n_230),
.B1(n_228),
.B2(n_229),
.Y(n_1758)
);

CKINVDCx10_ASAP7_75t_R g1759 ( 
.A(n_1373),
.Y(n_1759)
);

AOI21xp5_ASAP7_75t_L g1760 ( 
.A1(n_1439),
.A2(n_231),
.B(n_232),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1421),
.B(n_231),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1421),
.B(n_232),
.Y(n_1762)
);

AOI21xp5_ASAP7_75t_L g1763 ( 
.A1(n_1439),
.A2(n_233),
.B(n_234),
.Y(n_1763)
);

AOI22xp5_ASAP7_75t_L g1764 ( 
.A1(n_1509),
.A2(n_235),
.B1(n_233),
.B2(n_234),
.Y(n_1764)
);

AO21x2_ASAP7_75t_L g1765 ( 
.A1(n_1400),
.A2(n_234),
.B(n_235),
.Y(n_1765)
);

OR2x6_ASAP7_75t_L g1766 ( 
.A(n_1730),
.B(n_236),
.Y(n_1766)
);

OAI21xp5_ASAP7_75t_L g1767 ( 
.A1(n_1562),
.A2(n_236),
.B(n_237),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_SL g1768 ( 
.A1(n_1566),
.A2(n_238),
.B(n_239),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1591),
.B(n_238),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1513),
.B(n_474),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1530),
.Y(n_1771)
);

OAI22x1_ASAP7_75t_L g1772 ( 
.A1(n_1685),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_1772)
);

OAI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1567),
.A2(n_243),
.B(n_244),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1676),
.B(n_244),
.Y(n_1774)
);

OAI21x1_ASAP7_75t_L g1775 ( 
.A1(n_1535),
.A2(n_245),
.B(n_246),
.Y(n_1775)
);

OA22x2_ASAP7_75t_L g1776 ( 
.A1(n_1620),
.A2(n_1538),
.B1(n_1594),
.B2(n_1602),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1603),
.A2(n_1733),
.B(n_1668),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1698),
.B(n_247),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1512),
.B(n_1528),
.Y(n_1779)
);

OR2x6_ASAP7_75t_L g1780 ( 
.A(n_1510),
.B(n_247),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_SL g1781 ( 
.A(n_1684),
.B(n_474),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1512),
.B(n_249),
.Y(n_1782)
);

OAI22x1_ASAP7_75t_L g1783 ( 
.A1(n_1734),
.A2(n_1602),
.B1(n_1695),
.B2(n_1661),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1655),
.A2(n_252),
.B(n_253),
.Y(n_1784)
);

OAI21xp5_ASAP7_75t_L g1785 ( 
.A1(n_1523),
.A2(n_252),
.B(n_253),
.Y(n_1785)
);

BUFx6f_ASAP7_75t_L g1786 ( 
.A(n_1511),
.Y(n_1786)
);

NAND2x1_ASAP7_75t_L g1787 ( 
.A(n_1511),
.B(n_254),
.Y(n_1787)
);

AOI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1658),
.A2(n_255),
.B(n_256),
.Y(n_1788)
);

CKINVDCx5p33_ASAP7_75t_R g1789 ( 
.A(n_1654),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1511),
.A2(n_1559),
.B(n_1547),
.Y(n_1790)
);

OAI21x1_ASAP7_75t_L g1791 ( 
.A1(n_1641),
.A2(n_259),
.B(n_260),
.Y(n_1791)
);

OAI21x1_ASAP7_75t_L g1792 ( 
.A1(n_1534),
.A2(n_261),
.B(n_262),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1717),
.B(n_262),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1662),
.A2(n_263),
.B(n_264),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1718),
.B(n_263),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1724),
.B(n_265),
.Y(n_1796)
);

BUFx3_ASAP7_75t_L g1797 ( 
.A(n_1659),
.Y(n_1797)
);

NAND3xp33_ASAP7_75t_SL g1798 ( 
.A(n_1702),
.B(n_266),
.C(n_267),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1673),
.B(n_266),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1742),
.B(n_267),
.Y(n_1800)
);

OAI21x1_ASAP7_75t_L g1801 ( 
.A1(n_1554),
.A2(n_268),
.B(n_269),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1743),
.A2(n_268),
.B(n_269),
.Y(n_1802)
);

OAI21x1_ASAP7_75t_L g1803 ( 
.A1(n_1670),
.A2(n_268),
.B(n_270),
.Y(n_1803)
);

AND2x6_ASAP7_75t_L g1804 ( 
.A(n_1580),
.B(n_271),
.Y(n_1804)
);

INVxp67_ASAP7_75t_SL g1805 ( 
.A(n_1519),
.Y(n_1805)
);

NAND2x1p5_ASAP7_75t_L g1806 ( 
.A(n_1561),
.B(n_272),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1663),
.A2(n_273),
.B(n_274),
.Y(n_1807)
);

A2O1A1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1740),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_1808)
);

INVx2_ASAP7_75t_SL g1809 ( 
.A(n_1691),
.Y(n_1809)
);

NOR2xp33_ASAP7_75t_L g1810 ( 
.A(n_1606),
.B(n_276),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_SL g1811 ( 
.A(n_1714),
.B(n_475),
.Y(n_1811)
);

AND2x6_ASAP7_75t_L g1812 ( 
.A(n_1601),
.B(n_1571),
.Y(n_1812)
);

AOI21xp33_ASAP7_75t_L g1813 ( 
.A1(n_1524),
.A2(n_278),
.B(n_279),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1695),
.B(n_281),
.Y(n_1814)
);

BUFx6f_ASAP7_75t_L g1815 ( 
.A(n_1547),
.Y(n_1815)
);

HB1xp67_ASAP7_75t_L g1816 ( 
.A(n_1690),
.Y(n_1816)
);

OR2x6_ASAP7_75t_L g1817 ( 
.A(n_1738),
.B(n_282),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_L g1818 ( 
.A(n_1518),
.B(n_284),
.Y(n_1818)
);

NAND2x1p5_ASAP7_75t_L g1819 ( 
.A(n_1545),
.B(n_284),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1716),
.A2(n_287),
.B1(n_285),
.B2(n_286),
.Y(n_1820)
);

OAI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1526),
.A2(n_288),
.B(n_289),
.Y(n_1821)
);

AOI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1678),
.A2(n_1681),
.B(n_1680),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1726),
.B(n_288),
.Y(n_1823)
);

OAI21x1_ASAP7_75t_SL g1824 ( 
.A1(n_1687),
.A2(n_290),
.B(n_291),
.Y(n_1824)
);

BUFx3_ASAP7_75t_L g1825 ( 
.A(n_1598),
.Y(n_1825)
);

OA22x2_ASAP7_75t_L g1826 ( 
.A1(n_1620),
.A2(n_1557),
.B1(n_1751),
.B2(n_1549),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1677),
.Y(n_1827)
);

BUFx4_ASAP7_75t_SL g1828 ( 
.A(n_1669),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1682),
.Y(n_1829)
);

BUFx6f_ASAP7_75t_L g1830 ( 
.A(n_1547),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1560),
.B(n_294),
.Y(n_1831)
);

NAND2x1_ASAP7_75t_L g1832 ( 
.A(n_1559),
.B(n_295),
.Y(n_1832)
);

AOI21x1_ASAP7_75t_SL g1833 ( 
.A1(n_1649),
.A2(n_297),
.B(n_298),
.Y(n_1833)
);

NAND2x1p5_ASAP7_75t_L g1834 ( 
.A(n_1545),
.B(n_298),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1540),
.A2(n_301),
.B1(n_299),
.B2(n_300),
.Y(n_1835)
);

AND2x4_ASAP7_75t_L g1836 ( 
.A(n_1673),
.B(n_299),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1701),
.Y(n_1837)
);

NOR2xp33_ASAP7_75t_L g1838 ( 
.A(n_1607),
.B(n_302),
.Y(n_1838)
);

NAND2x1p5_ASAP7_75t_L g1839 ( 
.A(n_1545),
.B(n_304),
.Y(n_1839)
);

INVx4_ASAP7_75t_L g1840 ( 
.A(n_1692),
.Y(n_1840)
);

BUFx3_ASAP7_75t_L g1841 ( 
.A(n_1572),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_SL g1842 ( 
.A(n_1595),
.B(n_476),
.Y(n_1842)
);

AND2x6_ASAP7_75t_L g1843 ( 
.A(n_1559),
.B(n_308),
.Y(n_1843)
);

AOI21x1_ASAP7_75t_SL g1844 ( 
.A1(n_1640),
.A2(n_309),
.B(n_310),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1583),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_1845)
);

INVx8_ASAP7_75t_L g1846 ( 
.A(n_1629),
.Y(n_1846)
);

INVx4_ASAP7_75t_L g1847 ( 
.A(n_1706),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_SL g1848 ( 
.A1(n_1569),
.A2(n_313),
.B(n_314),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1706),
.B(n_316),
.Y(n_1849)
);

INVx4_ASAP7_75t_L g1850 ( 
.A(n_1605),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_SL g1851 ( 
.A1(n_1569),
.A2(n_318),
.B(n_319),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1696),
.Y(n_1852)
);

AOI21xp5_ASAP7_75t_SL g1853 ( 
.A1(n_1569),
.A2(n_319),
.B(n_320),
.Y(n_1853)
);

A2O1A1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1590),
.A2(n_1651),
.B(n_1573),
.C(n_1587),
.Y(n_1854)
);

O2A1O1Ixp5_ASAP7_75t_L g1855 ( 
.A1(n_1521),
.A2(n_323),
.B(n_321),
.C(n_322),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1565),
.B(n_322),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1711),
.Y(n_1857)
);

AOI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1732),
.A2(n_324),
.B(n_325),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1616),
.B(n_1537),
.Y(n_1859)
);

AOI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1741),
.A2(n_325),
.B(n_326),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1746),
.A2(n_326),
.B(n_327),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1582),
.B(n_1584),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1635),
.Y(n_1863)
);

OAI21x1_ASAP7_75t_L g1864 ( 
.A1(n_1722),
.A2(n_331),
.B(n_332),
.Y(n_1864)
);

OA21x2_ASAP7_75t_L g1865 ( 
.A1(n_1757),
.A2(n_331),
.B(n_332),
.Y(n_1865)
);

OA21x2_ASAP7_75t_L g1866 ( 
.A1(n_1689),
.A2(n_332),
.B(n_333),
.Y(n_1866)
);

AOI21xp5_ASAP7_75t_L g1867 ( 
.A1(n_1761),
.A2(n_334),
.B(n_335),
.Y(n_1867)
);

AND3x4_ASAP7_75t_L g1868 ( 
.A(n_1531),
.B(n_335),
.C(n_336),
.Y(n_1868)
);

OAI21x1_ASAP7_75t_L g1869 ( 
.A1(n_1735),
.A2(n_337),
.B(n_338),
.Y(n_1869)
);

AOI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1762),
.A2(n_339),
.B(n_340),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1639),
.A2(n_340),
.B(n_341),
.Y(n_1871)
);

AOI21xp5_ASAP7_75t_L g1872 ( 
.A1(n_1633),
.A2(n_340),
.B(n_341),
.Y(n_1872)
);

AOI21x1_ASAP7_75t_L g1873 ( 
.A1(n_1610),
.A2(n_341),
.B(n_342),
.Y(n_1873)
);

OAI22x1_ASAP7_75t_L g1874 ( 
.A1(n_1563),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1516),
.B(n_344),
.Y(n_1875)
);

AO31x2_ASAP7_75t_L g1876 ( 
.A1(n_1555),
.A2(n_347),
.A3(n_345),
.B(n_346),
.Y(n_1876)
);

BUFx4f_ASAP7_75t_L g1877 ( 
.A(n_1527),
.Y(n_1877)
);

AOI21xp5_ASAP7_75t_L g1878 ( 
.A1(n_1645),
.A2(n_1553),
.B(n_1558),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1571),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1759),
.Y(n_1880)
);

AO21x1_ASAP7_75t_L g1881 ( 
.A1(n_1576),
.A2(n_478),
.B(n_477),
.Y(n_1881)
);

NAND2xp33_ASAP7_75t_L g1882 ( 
.A(n_1615),
.B(n_349),
.Y(n_1882)
);

AND2x4_ASAP7_75t_L g1883 ( 
.A(n_1634),
.B(n_349),
.Y(n_1883)
);

NOR2xp33_ASAP7_75t_R g1884 ( 
.A(n_1551),
.B(n_350),
.Y(n_1884)
);

OAI21x1_ASAP7_75t_L g1885 ( 
.A1(n_1643),
.A2(n_350),
.B(n_351),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1586),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1694),
.B(n_351),
.Y(n_1887)
);

OAI21x1_ASAP7_75t_L g1888 ( 
.A1(n_1646),
.A2(n_353),
.B(n_354),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1715),
.B(n_354),
.Y(n_1889)
);

INVx2_ASAP7_75t_SL g1890 ( 
.A(n_1719),
.Y(n_1890)
);

AO31x2_ASAP7_75t_L g1891 ( 
.A1(n_1599),
.A2(n_358),
.A3(n_356),
.B(n_357),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_SL g1892 ( 
.A(n_1672),
.B(n_478),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1539),
.A2(n_359),
.B(n_360),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1522),
.B(n_359),
.Y(n_1894)
);

OAI22x1_ASAP7_75t_L g1895 ( 
.A1(n_1596),
.A2(n_363),
.B1(n_360),
.B2(n_362),
.Y(n_1895)
);

OAI21x1_ASAP7_75t_L g1896 ( 
.A1(n_1648),
.A2(n_362),
.B(n_363),
.Y(n_1896)
);

BUFx4_ASAP7_75t_SL g1897 ( 
.A(n_1593),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1536),
.B(n_364),
.Y(n_1898)
);

AOI21xp5_ASAP7_75t_L g1899 ( 
.A1(n_1589),
.A2(n_365),
.B(n_366),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1541),
.B(n_367),
.Y(n_1900)
);

AOI21xp33_ASAP7_75t_L g1901 ( 
.A1(n_1631),
.A2(n_370),
.B(n_371),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1542),
.B(n_371),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1543),
.B(n_372),
.Y(n_1903)
);

AOI211x1_ASAP7_75t_L g1904 ( 
.A1(n_1656),
.A2(n_1747),
.B(n_1737),
.C(n_1671),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1588),
.Y(n_1905)
);

OAI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1592),
.A2(n_375),
.B(n_376),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1533),
.B(n_376),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1525),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1765),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1597),
.A2(n_378),
.B(n_379),
.Y(n_1910)
);

INVx4_ASAP7_75t_L g1911 ( 
.A(n_1615),
.Y(n_1911)
);

OAI21x1_ASAP7_75t_L g1912 ( 
.A1(n_1515),
.A2(n_1613),
.B(n_1556),
.Y(n_1912)
);

INVx2_ASAP7_75t_SL g1913 ( 
.A(n_1721),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1575),
.B(n_380),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_SL g1915 ( 
.A1(n_1580),
.A2(n_380),
.B(n_381),
.Y(n_1915)
);

AOI21x1_ASAP7_75t_SL g1916 ( 
.A1(n_1630),
.A2(n_1627),
.B(n_1626),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1578),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1634),
.B(n_382),
.Y(n_1918)
);

INVx3_ASAP7_75t_L g1919 ( 
.A(n_1615),
.Y(n_1919)
);

AO31x2_ASAP7_75t_L g1920 ( 
.A1(n_1574),
.A2(n_386),
.A3(n_384),
.B(n_385),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1529),
.B(n_387),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1617),
.Y(n_1922)
);

AOI21x1_ASAP7_75t_L g1923 ( 
.A1(n_1623),
.A2(n_391),
.B(n_392),
.Y(n_1923)
);

INVx2_ASAP7_75t_L g1924 ( 
.A(n_1632),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1544),
.B(n_393),
.Y(n_1925)
);

AO21x2_ASAP7_75t_L g1926 ( 
.A1(n_1705),
.A2(n_395),
.B(n_396),
.Y(n_1926)
);

OAI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1568),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_1927)
);

BUFx6f_ASAP7_75t_L g1928 ( 
.A(n_1580),
.Y(n_1928)
);

OAI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1514),
.A2(n_397),
.B(n_398),
.Y(n_1929)
);

OAI21x1_ASAP7_75t_L g1930 ( 
.A1(n_1666),
.A2(n_1727),
.B(n_1704),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1644),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1585),
.B(n_403),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1666),
.B(n_403),
.Y(n_1933)
);

OAI21x1_ASAP7_75t_L g1934 ( 
.A1(n_1756),
.A2(n_406),
.B(n_407),
.Y(n_1934)
);

INVxp67_ASAP7_75t_L g1935 ( 
.A(n_1688),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1564),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1600),
.A2(n_410),
.B1(n_408),
.B2(n_409),
.Y(n_1937)
);

AO31x2_ASAP7_75t_L g1938 ( 
.A1(n_1550),
.A2(n_410),
.A3(n_408),
.B(n_409),
.Y(n_1938)
);

OAI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1756),
.A2(n_411),
.B(n_412),
.Y(n_1939)
);

NOR2xp33_ASAP7_75t_L g1940 ( 
.A(n_1520),
.B(n_411),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1621),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1577),
.B(n_415),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1708),
.B(n_415),
.Y(n_1943)
);

AOI21xp33_ASAP7_75t_L g1944 ( 
.A1(n_1546),
.A2(n_416),
.B(n_417),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1739),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1758),
.B(n_417),
.Y(n_1946)
);

BUFx2_ASAP7_75t_L g1947 ( 
.A(n_1532),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1764),
.Y(n_1948)
);

OAI21xp5_ASAP7_75t_L g1949 ( 
.A1(n_1637),
.A2(n_419),
.B(n_420),
.Y(n_1949)
);

INVx1_ASAP7_75t_SL g1950 ( 
.A(n_1624),
.Y(n_1950)
);

INVx2_ASAP7_75t_SL g1951 ( 
.A(n_1650),
.Y(n_1951)
);

BUFx8_ASAP7_75t_L g1952 ( 
.A(n_1604),
.Y(n_1952)
);

AO31x2_ASAP7_75t_L g1953 ( 
.A1(n_1664),
.A2(n_423),
.A3(n_421),
.B(n_422),
.Y(n_1953)
);

BUFx8_ASAP7_75t_L g1954 ( 
.A(n_1604),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1517),
.B(n_1653),
.Y(n_1955)
);

AOI21x1_ASAP7_75t_L g1956 ( 
.A1(n_1618),
.A2(n_1622),
.B(n_1619),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1745),
.B(n_425),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1604),
.Y(n_1958)
);

INVxp67_ASAP7_75t_L g1959 ( 
.A(n_1657),
.Y(n_1959)
);

AOI21x1_ASAP7_75t_L g1960 ( 
.A1(n_1612),
.A2(n_426),
.B(n_427),
.Y(n_1960)
);

NOR2xp33_ASAP7_75t_L g1961 ( 
.A(n_1552),
.B(n_428),
.Y(n_1961)
);

BUFx12f_ASAP7_75t_L g1962 ( 
.A(n_1617),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_SL g1963 ( 
.A1(n_1700),
.A2(n_429),
.B(n_430),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1609),
.B(n_431),
.Y(n_1964)
);

OAI22x1_ASAP7_75t_L g1965 ( 
.A1(n_1709),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1611),
.B(n_432),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1614),
.B(n_432),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1579),
.B(n_434),
.Y(n_1968)
);

NAND2x1p5_ASAP7_75t_L g1969 ( 
.A(n_1723),
.B(n_439),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1720),
.Y(n_1970)
);

BUFx6f_ASAP7_75t_L g1971 ( 
.A(n_1725),
.Y(n_1971)
);

AOI21x1_ASAP7_75t_L g1972 ( 
.A1(n_1608),
.A2(n_441),
.B(n_442),
.Y(n_1972)
);

OAI21x1_ASAP7_75t_SL g1973 ( 
.A1(n_1660),
.A2(n_444),
.B(n_445),
.Y(n_1973)
);

BUFx6f_ASAP7_75t_SL g1974 ( 
.A(n_1675),
.Y(n_1974)
);

NAND2x1p5_ASAP7_75t_L g1975 ( 
.A(n_1729),
.B(n_445),
.Y(n_1975)
);

AND3x4_ASAP7_75t_L g1976 ( 
.A(n_1697),
.B(n_446),
.C(n_447),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1777),
.A2(n_1736),
.B(n_1729),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1822),
.A2(n_1749),
.B(n_1736),
.Y(n_1978)
);

BUFx12f_ASAP7_75t_L g1979 ( 
.A(n_1771),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1816),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1828),
.Y(n_1981)
);

OR2x2_ASAP7_75t_SL g1982 ( 
.A(n_1798),
.B(n_1652),
.Y(n_1982)
);

AOI22xp33_ASAP7_75t_SL g1983 ( 
.A1(n_1776),
.A2(n_1665),
.B1(n_1683),
.B2(n_1674),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1945),
.B(n_1642),
.Y(n_1984)
);

AND2x2_ASAP7_75t_SL g1985 ( 
.A(n_1882),
.B(n_1736),
.Y(n_1985)
);

NOR2xp67_ASAP7_75t_L g1986 ( 
.A(n_1840),
.B(n_1847),
.Y(n_1986)
);

AOI22xp33_ASAP7_75t_L g1987 ( 
.A1(n_1826),
.A2(n_1731),
.B1(n_1744),
.B2(n_1728),
.Y(n_1987)
);

BUFx5_ASAP7_75t_L g1988 ( 
.A(n_1812),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1948),
.B(n_1625),
.Y(n_1989)
);

CKINVDCx20_ASAP7_75t_R g1990 ( 
.A(n_1789),
.Y(n_1990)
);

INVx3_ASAP7_75t_SL g1991 ( 
.A(n_1846),
.Y(n_1991)
);

CKINVDCx20_ASAP7_75t_R g1992 ( 
.A(n_1852),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1825),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1914),
.B(n_448),
.Y(n_1994)
);

INVx4_ASAP7_75t_L g1995 ( 
.A(n_1846),
.Y(n_1995)
);

BUFx5_ASAP7_75t_L g1996 ( 
.A(n_1812),
.Y(n_1996)
);

O2A1O1Ixp33_ASAP7_75t_L g1997 ( 
.A1(n_1854),
.A2(n_1548),
.B(n_1570),
.C(n_1628),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1878),
.A2(n_1750),
.B(n_1749),
.Y(n_1998)
);

CKINVDCx20_ASAP7_75t_R g1999 ( 
.A(n_1880),
.Y(n_1999)
);

INVx4_ASAP7_75t_SL g2000 ( 
.A(n_1804),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1849),
.A2(n_1868),
.B1(n_1810),
.B2(n_1940),
.Y(n_2001)
);

BUFx12f_ASAP7_75t_L g2002 ( 
.A(n_1809),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1797),
.B(n_1863),
.Y(n_2003)
);

INVx5_ASAP7_75t_L g2004 ( 
.A(n_1780),
.Y(n_2004)
);

NAND2x1p5_ASAP7_75t_L g2005 ( 
.A(n_1850),
.B(n_1750),
.Y(n_2005)
);

NAND2xp5_ASAP7_75t_L g2006 ( 
.A(n_1931),
.B(n_1667),
.Y(n_2006)
);

BUFx3_ASAP7_75t_L g2007 ( 
.A(n_1779),
.Y(n_2007)
);

INVx5_ASAP7_75t_L g2008 ( 
.A(n_1780),
.Y(n_2008)
);

BUFx12f_ASAP7_75t_L g2009 ( 
.A(n_1766),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1877),
.Y(n_2010)
);

OR2x6_ASAP7_75t_L g2011 ( 
.A(n_1817),
.B(n_1679),
.Y(n_2011)
);

INVx3_ASAP7_75t_L g2012 ( 
.A(n_1877),
.Y(n_2012)
);

AND2x2_ASAP7_75t_L g2013 ( 
.A(n_1769),
.B(n_448),
.Y(n_2013)
);

CKINVDCx5p33_ASAP7_75t_R g2014 ( 
.A(n_1884),
.Y(n_2014)
);

BUFx6f_ASAP7_75t_L g2015 ( 
.A(n_1962),
.Y(n_2015)
);

AND2x4_ASAP7_75t_L g2016 ( 
.A(n_1841),
.B(n_1686),
.Y(n_2016)
);

INVx2_ASAP7_75t_SL g2017 ( 
.A(n_1897),
.Y(n_2017)
);

BUFx2_ASAP7_75t_L g2018 ( 
.A(n_1908),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1814),
.B(n_449),
.Y(n_2019)
);

OR2x6_ASAP7_75t_SL g2020 ( 
.A(n_1970),
.B(n_1647),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1817),
.B(n_1693),
.Y(n_2021)
);

AOI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_1790),
.A2(n_1703),
.B(n_1699),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1823),
.B(n_449),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1783),
.B(n_1748),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1774),
.B(n_1707),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_SL g2026 ( 
.A(n_1770),
.B(n_1748),
.Y(n_2026)
);

O2A1O1Ixp33_ASAP7_75t_SL g2027 ( 
.A1(n_1859),
.A2(n_1712),
.B(n_1713),
.C(n_1710),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1827),
.Y(n_2028)
);

OA21x2_ASAP7_75t_L g2029 ( 
.A1(n_1909),
.A2(n_1753),
.B(n_1752),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1829),
.Y(n_2030)
);

OAI22xp5_ASAP7_75t_L g2031 ( 
.A1(n_1781),
.A2(n_1754),
.B1(n_1760),
.B2(n_1755),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1924),
.A2(n_1763),
.B(n_1636),
.Y(n_2032)
);

OR2x2_ASAP7_75t_L g2033 ( 
.A(n_1805),
.B(n_1581),
.Y(n_2033)
);

AND2x4_ASAP7_75t_L g2034 ( 
.A(n_1766),
.B(n_1638),
.Y(n_2034)
);

NAND3xp33_ASAP7_75t_L g2035 ( 
.A(n_1904),
.B(n_450),
.C(n_452),
.Y(n_2035)
);

INVxp67_ASAP7_75t_SL g2036 ( 
.A(n_1883),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1911),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1887),
.B(n_453),
.Y(n_2038)
);

BUFx3_ASAP7_75t_L g2039 ( 
.A(n_1890),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1913),
.B(n_454),
.Y(n_2040)
);

BUFx6f_ASAP7_75t_L g2041 ( 
.A(n_1786),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1782),
.B(n_454),
.Y(n_2042)
);

NAND4xp25_ASAP7_75t_L g2043 ( 
.A(n_1778),
.B(n_457),
.C(n_455),
.D(n_456),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1837),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1917),
.A2(n_459),
.B1(n_457),
.B2(n_458),
.Y(n_2045)
);

NAND2xp5_ASAP7_75t_L g2046 ( 
.A(n_1793),
.B(n_1795),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1857),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1974),
.A2(n_461),
.B1(n_459),
.B2(n_460),
.Y(n_2048)
);

AOI221xp5_ASAP7_75t_L g2049 ( 
.A1(n_1838),
.A2(n_462),
.B1(n_460),
.B2(n_461),
.C(n_463),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1919),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1796),
.B(n_1800),
.Y(n_2051)
);

AOI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1871),
.A2(n_1905),
.B(n_1886),
.Y(n_2052)
);

NOR2x1_ASAP7_75t_SL g2053 ( 
.A(n_1842),
.B(n_463),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1941),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1786),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_1804),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1782),
.Y(n_2057)
);

NOR2xp33_ASAP7_75t_L g2058 ( 
.A(n_1935),
.B(n_480),
.Y(n_2058)
);

AND2x2_ASAP7_75t_L g2059 ( 
.A(n_1889),
.B(n_482),
.Y(n_2059)
);

OA21x2_ASAP7_75t_L g2060 ( 
.A1(n_1958),
.A2(n_485),
.B(n_486),
.Y(n_2060)
);

OR2x6_ASAP7_75t_L g2061 ( 
.A(n_1806),
.B(n_486),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_1936),
.A2(n_487),
.B(n_488),
.Y(n_2062)
);

BUFx3_ASAP7_75t_L g2063 ( 
.A(n_1799),
.Y(n_2063)
);

AND2x4_ASAP7_75t_L g2064 ( 
.A(n_1799),
.B(n_489),
.Y(n_2064)
);

AND2x4_ASAP7_75t_L g2065 ( 
.A(n_1836),
.B(n_665),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1815),
.Y(n_2066)
);

A2O1A1Ixp33_ASAP7_75t_L g2067 ( 
.A1(n_1821),
.A2(n_492),
.B(n_490),
.C(n_491),
.Y(n_2067)
);

AND2x4_ASAP7_75t_L g2068 ( 
.A(n_1950),
.B(n_492),
.Y(n_2068)
);

AND2x4_ASAP7_75t_L g2069 ( 
.A(n_1919),
.B(n_493),
.Y(n_2069)
);

AND2x4_ASAP7_75t_L g2070 ( 
.A(n_1947),
.B(n_494),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1815),
.Y(n_2071)
);

AND2x2_ASAP7_75t_SL g2072 ( 
.A(n_1921),
.B(n_495),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1862),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1918),
.B(n_1933),
.Y(n_2074)
);

A2O1A1Ixp33_ASAP7_75t_L g2075 ( 
.A1(n_1767),
.A2(n_499),
.B(n_497),
.C(n_498),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1864),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1869),
.Y(n_2077)
);

NAND2x1_ASAP7_75t_L g2078 ( 
.A(n_1804),
.B(n_500),
.Y(n_2078)
);

CKINVDCx8_ASAP7_75t_R g2079 ( 
.A(n_1843),
.Y(n_2079)
);

OR2x2_ASAP7_75t_L g2080 ( 
.A(n_1875),
.B(n_501),
.Y(n_2080)
);

BUFx3_ASAP7_75t_L g2081 ( 
.A(n_1843),
.Y(n_2081)
);

INVx4_ASAP7_75t_SL g2082 ( 
.A(n_1843),
.Y(n_2082)
);

O2A1O1Ixp33_ASAP7_75t_L g2083 ( 
.A1(n_1808),
.A2(n_503),
.B(n_501),
.C(n_502),
.Y(n_2083)
);

OR2x6_ASAP7_75t_L g2084 ( 
.A(n_1819),
.B(n_1834),
.Y(n_2084)
);

INVx1_ASAP7_75t_SL g2085 ( 
.A(n_1839),
.Y(n_2085)
);

BUFx3_ASAP7_75t_L g2086 ( 
.A(n_1812),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_1951),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_1874),
.B(n_504),
.Y(n_2088)
);

AOI21xp5_ASAP7_75t_L g2089 ( 
.A1(n_1773),
.A2(n_505),
.B(n_506),
.Y(n_2089)
);

INVx1_ASAP7_75t_SL g2090 ( 
.A(n_1830),
.Y(n_2090)
);

CKINVDCx8_ASAP7_75t_R g2091 ( 
.A(n_1818),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1969),
.B(n_507),
.Y(n_2092)
);

INVxp67_ASAP7_75t_L g2093 ( 
.A(n_1831),
.Y(n_2093)
);

BUFx12f_ASAP7_75t_L g2094 ( 
.A(n_1975),
.Y(n_2094)
);

INVx3_ASAP7_75t_SL g2095 ( 
.A(n_1812),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_1802),
.B(n_664),
.Y(n_2096)
);

AND2x4_ASAP7_75t_L g2097 ( 
.A(n_1959),
.B(n_508),
.Y(n_2097)
);

AOI21xp5_ASAP7_75t_L g2098 ( 
.A1(n_1792),
.A2(n_509),
.B(n_510),
.Y(n_2098)
);

BUFx2_ASAP7_75t_L g2099 ( 
.A(n_1879),
.Y(n_2099)
);

NAND2xp33_ASAP7_75t_L g2100 ( 
.A(n_1772),
.B(n_511),
.Y(n_2100)
);

CKINVDCx5p33_ASAP7_75t_R g2101 ( 
.A(n_1895),
.Y(n_2101)
);

INVx3_ASAP7_75t_L g2102 ( 
.A(n_1879),
.Y(n_2102)
);

AOI21xp5_ASAP7_75t_L g2103 ( 
.A1(n_1949),
.A2(n_512),
.B(n_513),
.Y(n_2103)
);

INVx1_ASAP7_75t_SL g2104 ( 
.A(n_1928),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_1928),
.Y(n_2105)
);

AOI21xp5_ASAP7_75t_L g2106 ( 
.A1(n_1957),
.A2(n_514),
.B(n_516),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1855),
.A2(n_517),
.B(n_518),
.Y(n_2107)
);

NOR2xp33_ASAP7_75t_SL g2108 ( 
.A(n_1976),
.B(n_520),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1856),
.Y(n_2109)
);

INVx3_ASAP7_75t_L g2110 ( 
.A(n_1971),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_1943),
.B(n_522),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_1894),
.B(n_663),
.Y(n_2112)
);

AND2x4_ASAP7_75t_L g2113 ( 
.A(n_2000),
.B(n_1912),
.Y(n_2113)
);

BUFx2_ASAP7_75t_L g2114 ( 
.A(n_2000),
.Y(n_2114)
);

BUFx8_ASAP7_75t_SL g2115 ( 
.A(n_1981),
.Y(n_2115)
);

HB1xp67_ASAP7_75t_L g2116 ( 
.A(n_1980),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_1983),
.A2(n_1952),
.B1(n_1954),
.B2(n_1881),
.Y(n_2117)
);

INVx6_ASAP7_75t_L g2118 ( 
.A(n_1995),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_1991),
.Y(n_2119)
);

BUFx6f_ASAP7_75t_L g2120 ( 
.A(n_2015),
.Y(n_2120)
);

OAI21x1_ASAP7_75t_L g2121 ( 
.A1(n_1977),
.A2(n_1833),
.B(n_1844),
.Y(n_2121)
);

INVx6_ASAP7_75t_L g2122 ( 
.A(n_2015),
.Y(n_2122)
);

AOI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_2011),
.A2(n_1954),
.B1(n_1952),
.B2(n_1927),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_2082),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1979),
.Y(n_2125)
);

AO21x1_ASAP7_75t_SL g2126 ( 
.A1(n_2082),
.A2(n_1785),
.B(n_1929),
.Y(n_2126)
);

OAI21x1_ASAP7_75t_L g2127 ( 
.A1(n_1998),
.A2(n_1916),
.B(n_1775),
.Y(n_2127)
);

INVxp67_ASAP7_75t_L g2128 ( 
.A(n_2018),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_SL g2129 ( 
.A1(n_2072),
.A2(n_1824),
.B1(n_1768),
.B2(n_1866),
.Y(n_2129)
);

BUFx6f_ASAP7_75t_L g2130 ( 
.A(n_2007),
.Y(n_2130)
);

BUFx2_ASAP7_75t_SL g2131 ( 
.A(n_1986),
.Y(n_2131)
);

OR2x6_ASAP7_75t_L g2132 ( 
.A(n_2017),
.B(n_1848),
.Y(n_2132)
);

AOI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2108),
.A2(n_1955),
.B1(n_1961),
.B2(n_1820),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2028),
.Y(n_2134)
);

AND2x4_ASAP7_75t_L g2135 ( 
.A(n_2081),
.B(n_1930),
.Y(n_2135)
);

AOI22xp33_ASAP7_75t_L g2136 ( 
.A1(n_2021),
.A2(n_1937),
.B1(n_1944),
.B2(n_1968),
.Y(n_2136)
);

OAI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_2043),
.A2(n_2001),
.B1(n_2008),
.B2(n_2004),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2030),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2016),
.A2(n_1965),
.B1(n_1813),
.B2(n_1901),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_2010),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2044),
.Y(n_2141)
);

AOI21x1_ASAP7_75t_L g2142 ( 
.A1(n_2024),
.A2(n_1873),
.B(n_1923),
.Y(n_2142)
);

AOI22xp33_ASAP7_75t_SL g2143 ( 
.A1(n_1985),
.A2(n_1866),
.B1(n_1865),
.B2(n_1926),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2047),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_2056),
.Y(n_2145)
);

BUFx10_ASAP7_75t_L g2146 ( 
.A(n_1993),
.Y(n_2146)
);

BUFx4f_ASAP7_75t_SL g2147 ( 
.A(n_2002),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2038),
.B(n_525),
.Y(n_2148)
);

BUFx12f_ASAP7_75t_L g2149 ( 
.A(n_2009),
.Y(n_2149)
);

NAND2x1p5_ASAP7_75t_L g2150 ( 
.A(n_2004),
.B(n_1811),
.Y(n_2150)
);

AOI22xp33_ASAP7_75t_L g2151 ( 
.A1(n_2100),
.A2(n_1973),
.B1(n_1892),
.B2(n_1845),
.Y(n_2151)
);

OAI21x1_ASAP7_75t_L g2152 ( 
.A1(n_1978),
.A2(n_1803),
.B(n_1801),
.Y(n_2152)
);

OAI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_2089),
.A2(n_1788),
.B(n_1784),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2073),
.B(n_1938),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_2012),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_2014),
.Y(n_2156)
);

BUFx2_ASAP7_75t_R g2157 ( 
.A(n_2079),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_2019),
.B(n_526),
.Y(n_2158)
);

NAND2x1p5_ASAP7_75t_L g2159 ( 
.A(n_2037),
.B(n_1934),
.Y(n_2159)
);

OAI21x1_ASAP7_75t_L g2160 ( 
.A1(n_2076),
.A2(n_1888),
.B(n_1885),
.Y(n_2160)
);

BUFx2_ASAP7_75t_L g2161 ( 
.A(n_2036),
.Y(n_2161)
);

OAI22xp33_ASAP7_75t_L g2162 ( 
.A1(n_2061),
.A2(n_1946),
.B1(n_1906),
.B2(n_1910),
.Y(n_2162)
);

NAND2x1p5_ASAP7_75t_L g2163 ( 
.A(n_2054),
.B(n_1939),
.Y(n_2163)
);

AND2x4_ASAP7_75t_L g2164 ( 
.A(n_2074),
.B(n_1922),
.Y(n_2164)
);

INVx2_ASAP7_75t_L g2165 ( 
.A(n_2060),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_2039),
.Y(n_2166)
);

OAI21x1_ASAP7_75t_L g2167 ( 
.A1(n_2077),
.A2(n_1896),
.B(n_1791),
.Y(n_2167)
);

NAND2x1p5_ASAP7_75t_L g2168 ( 
.A(n_2078),
.B(n_1787),
.Y(n_2168)
);

CKINVDCx5p33_ASAP7_75t_R g2169 ( 
.A(n_1990),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_L g2170 ( 
.A(n_2091),
.B(n_1925),
.Y(n_2170)
);

INVx3_ASAP7_75t_L g2171 ( 
.A(n_2094),
.Y(n_2171)
);

AND2x4_ASAP7_75t_L g2172 ( 
.A(n_2086),
.B(n_1922),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2109),
.Y(n_2173)
);

NAND2x1p5_ASAP7_75t_L g2174 ( 
.A(n_2085),
.B(n_1832),
.Y(n_2174)
);

HB1xp67_ASAP7_75t_L g2175 ( 
.A(n_2057),
.Y(n_2175)
);

OAI22xp33_ASAP7_75t_L g2176 ( 
.A1(n_2084),
.A2(n_1835),
.B1(n_1942),
.B2(n_1932),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2006),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2087),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2033),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2088),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2046),
.B(n_1938),
.Y(n_2181)
);

AND2x2_ASAP7_75t_L g2182 ( 
.A(n_2023),
.B(n_527),
.Y(n_2182)
);

INVx4_ASAP7_75t_L g2183 ( 
.A(n_2095),
.Y(n_2183)
);

INVx1_ASAP7_75t_L g2184 ( 
.A(n_1984),
.Y(n_2184)
);

AOI22xp33_ASAP7_75t_L g2185 ( 
.A1(n_2034),
.A2(n_1964),
.B1(n_1967),
.B2(n_1966),
.Y(n_2185)
);

AOI22xp5_ASAP7_75t_SL g2186 ( 
.A1(n_2101),
.A2(n_1872),
.B1(n_1899),
.B2(n_1893),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1989),
.Y(n_2187)
);

AOI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_2093),
.A2(n_1900),
.B1(n_1903),
.B2(n_1902),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2041),
.Y(n_2189)
);

INVx4_ASAP7_75t_L g2190 ( 
.A(n_2063),
.Y(n_2190)
);

HB1xp67_ASAP7_75t_L g2191 ( 
.A(n_2099),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2013),
.Y(n_2192)
);

OAI21xp5_ASAP7_75t_L g2193 ( 
.A1(n_2103),
.A2(n_1807),
.B(n_1794),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1994),
.Y(n_2194)
);

HB1xp67_ASAP7_75t_L g2195 ( 
.A(n_2105),
.Y(n_2195)
);

CKINVDCx11_ASAP7_75t_R g2196 ( 
.A(n_1992),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2059),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_2055),
.Y(n_2198)
);

BUFx2_ASAP7_75t_L g2199 ( 
.A(n_1988),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_2051),
.B(n_1953),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_2055),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2069),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_2066),
.Y(n_2203)
);

INVx3_ASAP7_75t_L g2204 ( 
.A(n_2005),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2035),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2090),
.B(n_1953),
.Y(n_2206)
);

CKINVDCx5p33_ASAP7_75t_R g2207 ( 
.A(n_1999),
.Y(n_2207)
);

INVx3_ASAP7_75t_L g2208 ( 
.A(n_2070),
.Y(n_2208)
);

BUFx2_ASAP7_75t_L g2209 ( 
.A(n_2145),
.Y(n_2209)
);

HB1xp67_ASAP7_75t_L g2210 ( 
.A(n_2116),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_2180),
.B(n_2042),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2192),
.B(n_2064),
.Y(n_2212)
);

BUFx2_ASAP7_75t_L g2213 ( 
.A(n_2145),
.Y(n_2213)
);

INVx2_ASAP7_75t_SL g2214 ( 
.A(n_2118),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2173),
.B(n_2065),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2184),
.Y(n_2216)
);

OR2x2_ASAP7_75t_L g2217 ( 
.A(n_2179),
.B(n_2040),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2194),
.B(n_2111),
.Y(n_2218)
);

INVx5_ASAP7_75t_L g2219 ( 
.A(n_2118),
.Y(n_2219)
);

OA21x2_ASAP7_75t_L g2220 ( 
.A1(n_2121),
.A2(n_2127),
.B(n_2165),
.Y(n_2220)
);

INVx4_ASAP7_75t_L g2221 ( 
.A(n_2183),
.Y(n_2221)
);

BUFx2_ASAP7_75t_L g2222 ( 
.A(n_2161),
.Y(n_2222)
);

INVx3_ASAP7_75t_L g2223 ( 
.A(n_2113),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2197),
.B(n_2068),
.Y(n_2224)
);

BUFx3_ASAP7_75t_L g2225 ( 
.A(n_2120),
.Y(n_2225)
);

AOI21xp5_ASAP7_75t_L g2226 ( 
.A1(n_2162),
.A2(n_2027),
.B(n_2022),
.Y(n_2226)
);

AND2x2_ASAP7_75t_SL g2227 ( 
.A(n_2114),
.B(n_2097),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_2113),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_2134),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_2138),
.Y(n_2230)
);

OR2x6_ASAP7_75t_L g2231 ( 
.A(n_2131),
.B(n_1851),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2187),
.Y(n_2232)
);

HB1xp67_ASAP7_75t_L g2233 ( 
.A(n_2191),
.Y(n_2233)
);

INVx2_ASAP7_75t_L g2234 ( 
.A(n_2141),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_2195),
.Y(n_2235)
);

AO31x2_ASAP7_75t_L g2236 ( 
.A1(n_2181),
.A2(n_2098),
.A3(n_2031),
.B(n_2075),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2144),
.Y(n_2237)
);

AO31x2_ASAP7_75t_L g2238 ( 
.A1(n_2200),
.A2(n_2032),
.A3(n_2067),
.B(n_2052),
.Y(n_2238)
);

AOI21x1_ASAP7_75t_L g2239 ( 
.A1(n_2142),
.A2(n_2026),
.B(n_2092),
.Y(n_2239)
);

OA21x2_ASAP7_75t_L g2240 ( 
.A1(n_2152),
.A2(n_2107),
.B(n_2025),
.Y(n_2240)
);

AO21x2_ASAP7_75t_L g2241 ( 
.A1(n_2137),
.A2(n_2053),
.B(n_2062),
.Y(n_2241)
);

NAND2x1p5_ASAP7_75t_L g2242 ( 
.A(n_2119),
.B(n_2050),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_2115),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2124),
.Y(n_2244)
);

BUFx4f_ASAP7_75t_L g2245 ( 
.A(n_2149),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_2117),
.A2(n_2126),
.B1(n_2123),
.B2(n_2129),
.Y(n_2246)
);

AND2x2_ASAP7_75t_L g2247 ( 
.A(n_2148),
.B(n_2104),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2177),
.Y(n_2248)
);

AND2x6_ASAP7_75t_L g2249 ( 
.A(n_2135),
.B(n_1988),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2178),
.Y(n_2250)
);

AND2x4_ASAP7_75t_L g2251 ( 
.A(n_2206),
.B(n_2102),
.Y(n_2251)
);

BUFx6f_ASAP7_75t_L g2252 ( 
.A(n_2130),
.Y(n_2252)
);

BUFx2_ASAP7_75t_L g2253 ( 
.A(n_2199),
.Y(n_2253)
);

AO21x2_ASAP7_75t_L g2254 ( 
.A1(n_2154),
.A2(n_2096),
.B(n_2112),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2158),
.B(n_2003),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2175),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_2130),
.Y(n_2257)
);

AO21x2_ASAP7_75t_L g2258 ( 
.A1(n_2205),
.A2(n_2160),
.B(n_2167),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2182),
.B(n_2058),
.Y(n_2259)
);

INVxp67_ASAP7_75t_SL g2260 ( 
.A(n_2163),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_2128),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2202),
.Y(n_2262)
);

NOR2x1_ASAP7_75t_SL g2263 ( 
.A(n_2126),
.B(n_2071),
.Y(n_2263)
);

AND2x4_ASAP7_75t_L g2264 ( 
.A(n_2135),
.B(n_2110),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2223),
.B(n_2190),
.Y(n_2265)
);

BUFx6f_ASAP7_75t_L g2266 ( 
.A(n_2219),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2222),
.Y(n_2267)
);

AND2x2_ASAP7_75t_L g2268 ( 
.A(n_2256),
.B(n_2166),
.Y(n_2268)
);

AOI22xp33_ASAP7_75t_L g2269 ( 
.A1(n_2246),
.A2(n_2176),
.B1(n_2139),
.B2(n_2185),
.Y(n_2269)
);

AND2x2_ASAP7_75t_L g2270 ( 
.A(n_2211),
.B(n_2189),
.Y(n_2270)
);

BUFx3_ASAP7_75t_L g2271 ( 
.A(n_2219),
.Y(n_2271)
);

OR2x2_ASAP7_75t_L g2272 ( 
.A(n_2210),
.B(n_2208),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2233),
.B(n_2198),
.Y(n_2273)
);

AND2x2_ASAP7_75t_L g2274 ( 
.A(n_2235),
.B(n_2201),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2255),
.B(n_2203),
.Y(n_2275)
);

NAND2x1_ASAP7_75t_L g2276 ( 
.A(n_2221),
.B(n_2122),
.Y(n_2276)
);

OAI22xp33_ASAP7_75t_L g2277 ( 
.A1(n_2219),
.A2(n_2133),
.B1(n_2132),
.B2(n_2020),
.Y(n_2277)
);

OA21x2_ASAP7_75t_L g2278 ( 
.A1(n_2226),
.A2(n_2193),
.B(n_2153),
.Y(n_2278)
);

AND2x2_ASAP7_75t_L g2279 ( 
.A(n_2247),
.B(n_2146),
.Y(n_2279)
);

HB1xp67_ASAP7_75t_L g2280 ( 
.A(n_2209),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2261),
.B(n_2170),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2216),
.B(n_1891),
.Y(n_2282)
);

AND2x4_ASAP7_75t_L g2283 ( 
.A(n_2223),
.B(n_2132),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2250),
.B(n_2164),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_2216),
.B(n_1891),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2229),
.Y(n_2286)
);

INVx1_ASAP7_75t_SL g2287 ( 
.A(n_2213),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2228),
.B(n_2172),
.Y(n_2288)
);

AND2x2_ASAP7_75t_L g2289 ( 
.A(n_2262),
.B(n_2172),
.Y(n_2289)
);

NAND2x1p5_ASAP7_75t_L g2290 ( 
.A(n_2214),
.B(n_2227),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2232),
.B(n_1891),
.Y(n_2291)
);

AND2x2_ASAP7_75t_L g2292 ( 
.A(n_2218),
.B(n_2155),
.Y(n_2292)
);

AND2x4_ASAP7_75t_SL g2293 ( 
.A(n_2252),
.B(n_2257),
.Y(n_2293)
);

INVx2_ASAP7_75t_L g2294 ( 
.A(n_2230),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2234),
.Y(n_2295)
);

INVxp67_ASAP7_75t_SL g2296 ( 
.A(n_2237),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2224),
.B(n_2140),
.Y(n_2297)
);

OR2x2_ASAP7_75t_L g2298 ( 
.A(n_2248),
.B(n_2171),
.Y(n_2298)
);

AND2x4_ASAP7_75t_L g2299 ( 
.A(n_2228),
.B(n_2204),
.Y(n_2299)
);

AND2x2_ASAP7_75t_SL g2300 ( 
.A(n_2265),
.B(n_2245),
.Y(n_2300)
);

AOI22xp33_ASAP7_75t_L g2301 ( 
.A1(n_2269),
.A2(n_2241),
.B1(n_2254),
.B2(n_2259),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2275),
.B(n_2251),
.Y(n_2302)
);

OAI22xp5_ASAP7_75t_L g2303 ( 
.A1(n_2290),
.A2(n_2231),
.B1(n_2157),
.B2(n_2260),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2273),
.B(n_2253),
.Y(n_2304)
);

AND2x2_ASAP7_75t_L g2305 ( 
.A(n_2274),
.B(n_2264),
.Y(n_2305)
);

OAI221xp5_ASAP7_75t_SL g2306 ( 
.A1(n_2277),
.A2(n_2151),
.B1(n_2136),
.B2(n_1987),
.C(n_2217),
.Y(n_2306)
);

OAI221xp5_ASAP7_75t_L g2307 ( 
.A1(n_2276),
.A2(n_2188),
.B1(n_2215),
.B2(n_2048),
.C(n_2186),
.Y(n_2307)
);

NAND3xp33_ASAP7_75t_L g2308 ( 
.A(n_2280),
.B(n_2143),
.C(n_2212),
.Y(n_2308)
);

OAI221xp5_ASAP7_75t_L g2309 ( 
.A1(n_2272),
.A2(n_2150),
.B1(n_2242),
.B2(n_2049),
.C(n_2045),
.Y(n_2309)
);

NOR3xp33_ASAP7_75t_SL g2310 ( 
.A(n_2282),
.B(n_2243),
.C(n_2125),
.Y(n_2310)
);

OAI22xp33_ASAP7_75t_L g2311 ( 
.A1(n_2271),
.A2(n_2244),
.B1(n_2147),
.B2(n_2252),
.Y(n_2311)
);

OAI21xp5_ASAP7_75t_SL g2312 ( 
.A1(n_2266),
.A2(n_2168),
.B(n_2174),
.Y(n_2312)
);

OAI22xp5_ASAP7_75t_L g2313 ( 
.A1(n_2271),
.A2(n_2257),
.B1(n_2225),
.B2(n_2159),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2297),
.B(n_2258),
.Y(n_2314)
);

NOR2xp33_ASAP7_75t_SL g2315 ( 
.A(n_2266),
.B(n_2169),
.Y(n_2315)
);

NAND2xp5_ASAP7_75t_L g2316 ( 
.A(n_2296),
.B(n_2236),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_2296),
.B(n_2238),
.Y(n_2317)
);

OAI22xp5_ASAP7_75t_L g2318 ( 
.A1(n_2298),
.A2(n_2122),
.B1(n_2207),
.B2(n_1982),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_2270),
.B(n_2263),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2268),
.B(n_2263),
.Y(n_2320)
);

OAI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_2265),
.A2(n_1982),
.B1(n_2156),
.B2(n_2080),
.Y(n_2321)
);

NAND3xp33_ASAP7_75t_L g2322 ( 
.A(n_2278),
.B(n_2240),
.C(n_1997),
.Y(n_2322)
);

AOI22xp33_ASAP7_75t_L g2323 ( 
.A1(n_2281),
.A2(n_2283),
.B1(n_2292),
.B2(n_2284),
.Y(n_2323)
);

OAI21xp33_ASAP7_75t_L g2324 ( 
.A1(n_2287),
.A2(n_1915),
.B(n_1853),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2279),
.B(n_2249),
.Y(n_2325)
);

NAND2x1p5_ASAP7_75t_L g2326 ( 
.A(n_2300),
.B(n_2283),
.Y(n_2326)
);

AND2x2_ASAP7_75t_SL g2327 ( 
.A(n_2320),
.B(n_2288),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2305),
.B(n_2288),
.Y(n_2328)
);

OR2x6_ASAP7_75t_L g2329 ( 
.A(n_2312),
.B(n_2299),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_2304),
.B(n_2289),
.Y(n_2330)
);

INVx6_ASAP7_75t_L g2331 ( 
.A(n_2319),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2314),
.B(n_2286),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_2302),
.B(n_2267),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2316),
.Y(n_2334)
);

HB1xp67_ASAP7_75t_L g2335 ( 
.A(n_2317),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_2323),
.B(n_2325),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2310),
.B(n_2294),
.Y(n_2337)
);

AND2x2_ASAP7_75t_SL g2338 ( 
.A(n_2301),
.B(n_2293),
.Y(n_2338)
);

INVx1_ASAP7_75t_SL g2339 ( 
.A(n_2315),
.Y(n_2339)
);

OR2x2_ASAP7_75t_L g2340 ( 
.A(n_2308),
.B(n_2295),
.Y(n_2340)
);

INVx2_ASAP7_75t_SL g2341 ( 
.A(n_2313),
.Y(n_2341)
);

INVx1_ASAP7_75t_L g2342 ( 
.A(n_2318),
.Y(n_2342)
);

HB1xp67_ASAP7_75t_L g2343 ( 
.A(n_2322),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_2303),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2341),
.B(n_2285),
.Y(n_2345)
);

OR2x2_ASAP7_75t_L g2346 ( 
.A(n_2332),
.B(n_2285),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2332),
.B(n_2291),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2327),
.B(n_2321),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2331),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2343),
.B(n_2311),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2336),
.B(n_2249),
.Y(n_2351)
);

AOI21xp5_ASAP7_75t_L g2352 ( 
.A1(n_2329),
.A2(n_2306),
.B(n_2324),
.Y(n_2352)
);

HB1xp67_ASAP7_75t_L g2353 ( 
.A(n_2335),
.Y(n_2353)
);

HB1xp67_ASAP7_75t_L g2354 ( 
.A(n_2353),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_2348),
.A2(n_2338),
.B1(n_2344),
.B2(n_2342),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2351),
.B(n_2326),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2346),
.B(n_2340),
.Y(n_2357)
);

OR2x2_ASAP7_75t_L g2358 ( 
.A(n_2347),
.B(n_2334),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2345),
.B(n_2337),
.Y(n_2359)
);

INVx2_ASAP7_75t_SL g2360 ( 
.A(n_2349),
.Y(n_2360)
);

AOI22xp5_ASAP7_75t_L g2361 ( 
.A1(n_2352),
.A2(n_2339),
.B1(n_2307),
.B2(n_2329),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_2345),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2350),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2360),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2358),
.Y(n_2365)
);

AND2x4_ASAP7_75t_L g2366 ( 
.A(n_2356),
.B(n_2359),
.Y(n_2366)
);

INVx1_ASAP7_75t_SL g2367 ( 
.A(n_2362),
.Y(n_2367)
);

OAI22xp33_ASAP7_75t_L g2368 ( 
.A1(n_2361),
.A2(n_2328),
.B1(n_2330),
.B2(n_2309),
.Y(n_2368)
);

OR2x2_ASAP7_75t_L g2369 ( 
.A(n_2357),
.B(n_2333),
.Y(n_2369)
);

AND2x2_ASAP7_75t_L g2370 ( 
.A(n_2355),
.B(n_2196),
.Y(n_2370)
);

INVx1_ASAP7_75t_SL g2371 ( 
.A(n_2354),
.Y(n_2371)
);

NOR2xp67_ASAP7_75t_SL g2372 ( 
.A(n_2363),
.B(n_1963),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_L g2373 ( 
.A(n_2367),
.B(n_2371),
.Y(n_2373)
);

INVxp67_ASAP7_75t_L g2374 ( 
.A(n_2370),
.Y(n_2374)
);

OAI21xp5_ASAP7_75t_L g2375 ( 
.A1(n_2368),
.A2(n_2083),
.B(n_2106),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2364),
.Y(n_2376)
);

INVx2_ASAP7_75t_SL g2377 ( 
.A(n_2366),
.Y(n_2377)
);

OR2x2_ASAP7_75t_L g2378 ( 
.A(n_2365),
.B(n_1876),
.Y(n_2378)
);

AND2x4_ASAP7_75t_L g2379 ( 
.A(n_2377),
.B(n_2376),
.Y(n_2379)
);

INVx1_ASAP7_75t_SL g2380 ( 
.A(n_2378),
.Y(n_2380)
);

NOR2xp33_ASAP7_75t_SL g2381 ( 
.A(n_2375),
.B(n_2372),
.Y(n_2381)
);

OAI22xp5_ASAP7_75t_L g2382 ( 
.A1(n_2374),
.A2(n_2369),
.B1(n_1907),
.B2(n_1898),
.Y(n_2382)
);

INVx1_ASAP7_75t_SL g2383 ( 
.A(n_2373),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2380),
.Y(n_2384)
);

OAI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2382),
.A2(n_1860),
.B1(n_1861),
.B2(n_1858),
.Y(n_2385)
);

OAI21xp5_ASAP7_75t_SL g2386 ( 
.A1(n_2383),
.A2(n_1870),
.B(n_1867),
.Y(n_2386)
);

AOI22xp33_ASAP7_75t_L g2387 ( 
.A1(n_2379),
.A2(n_1996),
.B1(n_2220),
.B2(n_2029),
.Y(n_2387)
);

OAI221xp5_ASAP7_75t_L g2388 ( 
.A1(n_2381),
.A2(n_1972),
.B1(n_2239),
.B2(n_1956),
.C(n_1960),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2384),
.B(n_529),
.Y(n_2389)
);

NOR2x1_ASAP7_75t_L g2390 ( 
.A(n_2386),
.B(n_530),
.Y(n_2390)
);

NOR4xp75_ASAP7_75t_L g2391 ( 
.A(n_2388),
.B(n_535),
.C(n_533),
.D(n_534),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_2387),
.B(n_533),
.Y(n_2392)
);

AOI211xp5_ASAP7_75t_L g2393 ( 
.A1(n_2385),
.A2(n_538),
.B(n_536),
.C(n_537),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2389),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2392),
.Y(n_2395)
);

OAI211xp5_ASAP7_75t_SL g2396 ( 
.A1(n_2390),
.A2(n_542),
.B(n_540),
.C(n_541),
.Y(n_2396)
);

NAND3xp33_ASAP7_75t_SL g2397 ( 
.A(n_2391),
.B(n_545),
.C(n_546),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_2394),
.Y(n_2398)
);

NOR2x1_ASAP7_75t_L g2399 ( 
.A(n_2395),
.B(n_2393),
.Y(n_2399)
);

NOR3xp33_ASAP7_75t_L g2400 ( 
.A(n_2396),
.B(n_546),
.C(n_547),
.Y(n_2400)
);

AOI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2397),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_2401)
);

OAI221xp5_ASAP7_75t_L g2402 ( 
.A1(n_2401),
.A2(n_554),
.B1(n_552),
.B2(n_553),
.C(n_555),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2400),
.B(n_552),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_2398),
.Y(n_2404)
);

XNOR2x1_ASAP7_75t_L g2405 ( 
.A(n_2399),
.B(n_556),
.Y(n_2405)
);

INVx2_ASAP7_75t_L g2406 ( 
.A(n_2404),
.Y(n_2406)
);

INVx2_ASAP7_75t_SL g2407 ( 
.A(n_2405),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2403),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2402),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_2406),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2409),
.Y(n_2411)
);

NOR3xp33_ASAP7_75t_L g2412 ( 
.A(n_2410),
.B(n_2408),
.C(n_2407),
.Y(n_2412)
);

OR3x1_ASAP7_75t_L g2413 ( 
.A(n_2411),
.B(n_560),
.C(n_562),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2412),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.Y(n_2414)
);

XOR2xp5_ASAP7_75t_L g2415 ( 
.A(n_2414),
.B(n_2413),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2415),
.Y(n_2416)
);

OR2x2_ASAP7_75t_L g2417 ( 
.A(n_2416),
.B(n_569),
.Y(n_2417)
);

OAI22xp5_ASAP7_75t_L g2418 ( 
.A1(n_2417),
.A2(n_1920),
.B1(n_573),
.B2(n_571),
.Y(n_2418)
);

AOI221xp5_ASAP7_75t_L g2419 ( 
.A1(n_2418),
.A2(n_575),
.B1(n_572),
.B2(n_574),
.C(n_576),
.Y(n_2419)
);

AOI211xp5_ASAP7_75t_L g2420 ( 
.A1(n_2419),
.A2(n_579),
.B(n_577),
.C(n_578),
.Y(n_2420)
);


endmodule