module real_aes_8810_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_182;
wire n_93;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_166;
wire n_103;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
A2O1A1Ixp33_ASAP7_75t_SL g252 ( .A1(n_0), .A2(n_253), .B(n_256), .C(n_260), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_1), .B(n_244), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_2), .B(n_254), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_3), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_4), .A2(n_213), .B(n_309), .Y(n_308) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_5), .A2(n_246), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g199 ( .A(n_6), .Y(n_199) );
AND2x6_ASAP7_75t_L g218 ( .A(n_6), .B(n_197), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_6), .B(n_531), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_L g334 ( .A1(n_7), .A2(n_218), .B(n_220), .C(n_335), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_8), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_9), .Y(n_100) );
AO22x2_ASAP7_75t_L g89 ( .A1(n_10), .A2(n_26), .B1(n_90), .B2(n_91), .Y(n_89) );
INVx1_ASAP7_75t_L g238 ( .A(n_11), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_12), .B(n_254), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_13), .A2(n_42), .B1(n_154), .B2(n_157), .Y(n_153) );
AO22x2_ASAP7_75t_L g93 ( .A1(n_14), .A2(n_28), .B1(n_90), .B2(n_94), .Y(n_93) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_15), .A2(n_68), .B1(n_171), .B2(n_173), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_16), .A2(n_220), .B(n_223), .C(n_231), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_17), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_18), .Y(n_132) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_19), .A2(n_220), .B(n_231), .C(n_321), .Y(n_320) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_20), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_21), .A2(n_80), .B1(n_81), .B2(n_177), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_21), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_22), .A2(n_213), .B(n_249), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g144 ( .A1(n_23), .A2(n_24), .B1(n_145), .B2(n_149), .Y(n_144) );
INVx2_ASAP7_75t_L g216 ( .A(n_25), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g269 ( .A1(n_27), .A2(n_270), .B(n_271), .C(n_275), .Y(n_269) );
OAI221xp5_ASAP7_75t_L g190 ( .A1(n_28), .A2(n_44), .B1(n_54), .B2(n_191), .C(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g193 ( .A(n_28), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_29), .Y(n_107) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_30), .A2(n_70), .B1(n_163), .B2(n_166), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g183 ( .A1(n_31), .A2(n_37), .B1(n_184), .B2(n_185), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_31), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_31), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_32), .B(n_212), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g339 ( .A(n_33), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_34), .B(n_254), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_35), .B(n_213), .Y(n_319) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_36), .A2(n_270), .B(n_275), .C(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g185 ( .A(n_37), .Y(n_185) );
INVx1_ASAP7_75t_L g257 ( .A(n_38), .Y(n_257) );
INVx1_ASAP7_75t_L g301 ( .A(n_39), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_39), .A2(n_80), .B1(n_81), .B2(n_301), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_40), .B(n_213), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_41), .A2(n_80), .B1(n_81), .B2(n_537), .Y(n_536) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_41), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_43), .Y(n_240) );
AO22x2_ASAP7_75t_L g97 ( .A1(n_44), .A2(n_61), .B1(n_90), .B2(n_94), .Y(n_97) );
INVxp67_ASAP7_75t_L g194 ( .A(n_44), .Y(n_194) );
INVx1_ASAP7_75t_L g197 ( .A(n_45), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_46), .B(n_213), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_47), .B(n_244), .Y(n_314) );
A2O1A1Ixp33_ASAP7_75t_L g311 ( .A1(n_48), .A2(n_230), .B(n_286), .C(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g237 ( .A(n_49), .Y(n_237) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_50), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_51), .B(n_254), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_52), .B(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_53), .B(n_255), .Y(n_336) );
AO22x2_ASAP7_75t_L g99 ( .A1(n_54), .A2(n_67), .B1(n_90), .B2(n_91), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_55), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_56), .B(n_225), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_57), .A2(n_220), .B(n_275), .C(n_284), .Y(n_283) );
CKINVDCx16_ASAP7_75t_R g310 ( .A(n_58), .Y(n_310) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_59), .B(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g277 ( .A(n_60), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_62), .A2(n_76), .B1(n_181), .B2(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_62), .Y(n_182) );
INVx2_ASAP7_75t_L g235 ( .A(n_63), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_64), .Y(n_293) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_65), .B(n_259), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_66), .B(n_213), .Y(n_268) );
INVx1_ASAP7_75t_L g272 ( .A(n_69), .Y(n_272) );
INVxp67_ASAP7_75t_L g313 ( .A(n_71), .Y(n_313) );
INVx1_ASAP7_75t_L g90 ( .A(n_72), .Y(n_90) );
INVx1_ASAP7_75t_L g92 ( .A(n_72), .Y(n_92) );
INVx1_ASAP7_75t_L g285 ( .A(n_73), .Y(n_285) );
INVx1_ASAP7_75t_L g332 ( .A(n_74), .Y(n_332) );
AND2x2_ASAP7_75t_L g303 ( .A(n_75), .B(n_234), .Y(n_303) );
INVx1_ASAP7_75t_L g181 ( .A(n_76), .Y(n_181) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_187), .B1(n_200), .B2(n_522), .C(n_526), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_178), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
HB1xp67_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g82 ( .A(n_83), .B(n_142), .Y(n_82) );
NOR3xp33_ASAP7_75t_L g83 ( .A(n_84), .B(n_115), .C(n_131), .Y(n_83) );
OAI221xp5_ASAP7_75t_L g84 ( .A1(n_85), .A2(n_100), .B1(n_101), .B2(n_107), .C(n_108), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_87), .Y(n_86) );
AND2x6_ASAP7_75t_L g87 ( .A(n_88), .B(n_95), .Y(n_87) );
AND2x4_ASAP7_75t_L g112 ( .A(n_88), .B(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g88 ( .A(n_89), .B(n_93), .Y(n_88) );
AND2x2_ASAP7_75t_L g106 ( .A(n_89), .B(n_97), .Y(n_106) );
INVx2_ASAP7_75t_L g122 ( .A(n_89), .Y(n_122) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g94 ( .A(n_92), .Y(n_94) );
OR2x2_ASAP7_75t_L g121 ( .A(n_93), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g130 ( .A(n_93), .B(n_122), .Y(n_130) );
INVx2_ASAP7_75t_L g137 ( .A(n_93), .Y(n_137) );
INVx1_ASAP7_75t_L g176 ( .A(n_93), .Y(n_176) );
AND2x6_ASAP7_75t_L g147 ( .A(n_95), .B(n_148), .Y(n_147) );
AND2x2_ASAP7_75t_L g156 ( .A(n_95), .B(n_152), .Y(n_156) );
AND2x4_ASAP7_75t_L g165 ( .A(n_95), .B(n_130), .Y(n_165) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_98), .Y(n_95) );
AND2x2_ASAP7_75t_L g124 ( .A(n_96), .B(n_99), .Y(n_124) );
INVx2_ASAP7_75t_L g96 ( .A(n_97), .Y(n_96) );
AND2x2_ASAP7_75t_L g151 ( .A(n_97), .B(n_114), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_97), .B(n_99), .Y(n_160) );
INVx1_ASAP7_75t_L g98 ( .A(n_99), .Y(n_98) );
INVx1_ASAP7_75t_L g105 ( .A(n_99), .Y(n_105) );
INVx1_ASAP7_75t_L g114 ( .A(n_99), .Y(n_114) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
BUFx6f_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AND2x2_ASAP7_75t_L g136 ( .A(n_105), .B(n_137), .Y(n_136) );
AND2x4_ASAP7_75t_L g135 ( .A(n_106), .B(n_136), .Y(n_135) );
NAND2x1p5_ASAP7_75t_L g140 ( .A(n_106), .B(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
INVx1_ASAP7_75t_SL g110 ( .A(n_111), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B1(n_125), .B2(n_126), .Y(n_115) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_123), .Y(n_120) );
INVx2_ASAP7_75t_L g148 ( .A(n_121), .Y(n_148) );
AND2x2_ASAP7_75t_L g152 ( .A(n_122), .B(n_137), .Y(n_152) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g129 ( .A(n_124), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g172 ( .A(n_124), .B(n_152), .Y(n_172) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g169 ( .A(n_130), .B(n_151), .Y(n_169) );
OAI22xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_133), .B1(n_138), .B2(n_139), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g141 ( .A(n_137), .Y(n_141) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g142 ( .A(n_143), .B(n_161), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_153), .Y(n_143) );
INVx2_ASAP7_75t_SL g145 ( .A(n_146), .Y(n_145) );
INVx11_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_152), .Y(n_150) );
AND2x4_ASAP7_75t_L g158 ( .A(n_152), .B(n_159), .Y(n_158) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx2_ASAP7_75t_SL g157 ( .A(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
OR2x6_ASAP7_75t_L g175 ( .A(n_160), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_170), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx6_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx5_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx8_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
BUFx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx6_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
OAI22xp5_ASAP7_75t_SL g178 ( .A1(n_179), .A2(n_180), .B1(n_183), .B2(n_186), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_183), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g187 ( .A(n_188), .Y(n_187) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_189), .Y(n_188) );
AND3x1_ASAP7_75t_SL g189 ( .A(n_190), .B(n_195), .C(n_198), .Y(n_189) );
INVxp67_ASAP7_75t_L g531 ( .A(n_190), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_193), .B(n_194), .Y(n_192) );
INVx1_ASAP7_75t_L g532 ( .A(n_195), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_195), .A2(n_524), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_196), .B(n_199), .Y(n_535) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_SL g540 ( .A(n_198), .B(n_532), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_SL g201 ( .A(n_202), .B(n_477), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_203), .B(n_412), .Y(n_202) );
NAND4xp25_ASAP7_75t_SL g203 ( .A(n_204), .B(n_357), .C(n_381), .D(n_404), .Y(n_203) );
AOI221xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_294), .B1(n_328), .B2(n_341), .C(n_344), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_264), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_207), .A2(n_242), .B1(n_295), .B2(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_207), .B(n_265), .Y(n_415) );
AND2x2_ASAP7_75t_L g434 ( .A(n_207), .B(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_207), .B(n_418), .Y(n_504) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_242), .Y(n_207) );
AND2x2_ASAP7_75t_L g372 ( .A(n_208), .B(n_265), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_208), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g395 ( .A(n_208), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g400 ( .A(n_208), .B(n_243), .Y(n_400) );
INVx2_ASAP7_75t_L g432 ( .A(n_208), .Y(n_432) );
HB1xp67_ASAP7_75t_L g476 ( .A(n_208), .Y(n_476) );
AND2x2_ASAP7_75t_L g493 ( .A(n_208), .B(n_370), .Y(n_493) );
INVx5_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g411 ( .A(n_209), .B(n_370), .Y(n_411) );
AND2x4_ASAP7_75t_L g425 ( .A(n_209), .B(n_242), .Y(n_425) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_209), .Y(n_429) );
AND2x2_ASAP7_75t_L g449 ( .A(n_209), .B(n_364), .Y(n_449) );
AND2x2_ASAP7_75t_L g499 ( .A(n_209), .B(n_266), .Y(n_499) );
AND2x2_ASAP7_75t_L g509 ( .A(n_209), .B(n_243), .Y(n_509) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_239), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_219), .B(n_232), .Y(n_210) );
BUFx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
AND2x4_ASAP7_75t_L g213 ( .A(n_214), .B(n_218), .Y(n_213) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_214), .B(n_218), .Y(n_333) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
INVx1_ASAP7_75t_L g230 ( .A(n_215), .Y(n_230) );
INVx1_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g221 ( .A(n_216), .Y(n_221) );
INVx1_ASAP7_75t_L g327 ( .A(n_216), .Y(n_327) );
INVx1_ASAP7_75t_L g222 ( .A(n_217), .Y(n_222) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_217), .Y(n_226) );
INVx3_ASAP7_75t_L g255 ( .A(n_217), .Y(n_255) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_217), .Y(n_259) );
INVx1_ASAP7_75t_L g323 ( .A(n_217), .Y(n_323) );
BUFx3_ASAP7_75t_L g231 ( .A(n_218), .Y(n_231) );
INVx4_ASAP7_75t_SL g262 ( .A(n_218), .Y(n_262) );
INVx5_ASAP7_75t_L g251 ( .A(n_220), .Y(n_251) );
AND2x6_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
BUFx3_ASAP7_75t_L g261 ( .A(n_221), .Y(n_261) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_227), .B(n_229), .Y(n_223) );
INVx2_ASAP7_75t_L g228 ( .A(n_225), .Y(n_228) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx4_ASAP7_75t_L g287 ( .A(n_226), .Y(n_287) );
O2A1O1Ixp33_ASAP7_75t_L g271 ( .A1(n_228), .A2(n_272), .B(n_273), .C(n_274), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g300 ( .A1(n_228), .A2(n_274), .B(n_301), .C(n_302), .Y(n_300) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_228), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_229), .B(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_231), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g241 ( .A(n_234), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_234), .A2(n_268), .B(n_269), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_234), .A2(n_298), .B(n_299), .Y(n_297) );
AND2x2_ASAP7_75t_SL g234 ( .A(n_235), .B(n_236), .Y(n_234) );
AND2x2_ASAP7_75t_L g247 ( .A(n_235), .B(n_236), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_L g365 ( .A(n_242), .B(n_265), .Y(n_365) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_242), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_242), .B(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g455 ( .A(n_242), .Y(n_455) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g343 ( .A(n_243), .B(n_280), .Y(n_343) );
AND2x2_ASAP7_75t_L g370 ( .A(n_243), .B(n_281), .Y(n_370) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_244), .A2(n_248), .B(n_263), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g276 ( .A(n_245), .B(n_277), .Y(n_276) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_245), .A2(n_282), .B(n_292), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_245), .B(n_293), .Y(n_292) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_245), .A2(n_331), .B(n_338), .Y(n_330) );
INVx4_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_246), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_246), .A2(n_319), .B(n_320), .Y(n_318) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g340 ( .A(n_247), .Y(n_340) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_251), .B(n_252), .C(n_262), .Y(n_249) );
INVx2_ASAP7_75t_L g270 ( .A(n_251), .Y(n_270) );
O2A1O1Ixp33_ASAP7_75t_L g309 ( .A1(n_251), .A2(n_262), .B(n_310), .C(n_311), .Y(n_309) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_254), .B(n_313), .Y(n_312) );
INVx5_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx4_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_261), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_262), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_264), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_278), .Y(n_264) );
OR2x2_ASAP7_75t_L g396 ( .A(n_265), .B(n_279), .Y(n_396) );
AND2x2_ASAP7_75t_L g433 ( .A(n_265), .B(n_343), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_265), .B(n_364), .Y(n_444) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_265), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_265), .B(n_400), .Y(n_517) );
INVx5_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
BUFx2_ASAP7_75t_L g342 ( .A(n_266), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_266), .B(n_279), .Y(n_351) );
AND2x2_ASAP7_75t_L g467 ( .A(n_266), .B(n_362), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_266), .B(n_400), .Y(n_489) );
OR2x6_ASAP7_75t_L g266 ( .A(n_267), .B(n_276), .Y(n_266) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_279), .Y(n_435) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_280), .Y(n_387) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx2_ASAP7_75t_L g364 ( .A(n_281), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_291), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_286), .B(n_288), .C(n_289), .Y(n_284) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_295), .B(n_304), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_295), .B(n_377), .Y(n_496) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NOR2xp33_ASAP7_75t_L g328 ( .A(n_296), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g348 ( .A(n_296), .B(n_349), .Y(n_348) );
INVx5_ASAP7_75t_SL g356 ( .A(n_296), .Y(n_356) );
OR2x2_ASAP7_75t_L g379 ( .A(n_296), .B(n_349), .Y(n_379) );
OR2x2_ASAP7_75t_L g389 ( .A(n_296), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g452 ( .A(n_296), .B(n_306), .Y(n_452) );
AND2x2_ASAP7_75t_SL g490 ( .A(n_296), .B(n_305), .Y(n_490) );
NOR4xp25_ASAP7_75t_L g511 ( .A(n_296), .B(n_432), .C(n_512), .D(n_513), .Y(n_511) );
AND2x2_ASAP7_75t_L g521 ( .A(n_296), .B(n_353), .Y(n_521) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_303), .Y(n_296) );
OAI322xp33_ASAP7_75t_L g526 ( .A1(n_301), .A2(n_527), .A3(n_528), .B1(n_532), .B2(n_533), .C1(n_536), .C2(n_538), .Y(n_526) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g346 ( .A(n_305), .B(n_342), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_305), .B(n_348), .Y(n_515) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_315), .Y(n_305) );
OR2x2_ASAP7_75t_L g355 ( .A(n_306), .B(n_356), .Y(n_355) );
INVx3_ASAP7_75t_L g362 ( .A(n_306), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_306), .B(n_330), .Y(n_374) );
INVxp67_ASAP7_75t_L g377 ( .A(n_306), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_306), .B(n_349), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_306), .B(n_316), .Y(n_443) );
AND2x2_ASAP7_75t_L g458 ( .A(n_306), .B(n_353), .Y(n_458) );
OR2x2_ASAP7_75t_L g487 ( .A(n_306), .B(n_316), .Y(n_487) );
OA21x2_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B(n_314), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_315), .B(n_392), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_315), .B(n_356), .Y(n_495) );
OR2x2_ASAP7_75t_L g516 ( .A(n_315), .B(n_393), .Y(n_516) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g329 ( .A(n_316), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_349), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g368 ( .A(n_316), .B(n_330), .Y(n_368) );
AND2x2_ASAP7_75t_L g438 ( .A(n_316), .B(n_362), .Y(n_438) );
AND2x2_ASAP7_75t_L g472 ( .A(n_316), .B(n_356), .Y(n_472) );
INVx2_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_317), .B(n_356), .Y(n_375) );
AND2x2_ASAP7_75t_L g403 ( .A(n_317), .B(n_330), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B(n_325), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_325), .A2(n_336), .B(n_337), .Y(n_335) );
INVx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_328), .B(n_411), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_329), .A2(n_418), .B1(n_454), .B2(n_471), .C(n_473), .Y(n_470) );
INVx5_ASAP7_75t_SL g349 ( .A(n_330), .Y(n_349) );
OAI21xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_333), .B(n_334), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
OAI33xp33_ASAP7_75t_L g369 ( .A1(n_342), .A2(n_370), .A3(n_371), .B1(n_373), .B2(n_376), .B3(n_380), .Y(n_369) );
OR2x2_ASAP7_75t_L g385 ( .A(n_342), .B(n_386), .Y(n_385) );
AOI322xp5_ASAP7_75t_L g494 ( .A1(n_342), .A2(n_411), .A3(n_418), .B1(n_495), .B2(n_496), .C1(n_497), .C2(n_500), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_342), .B(n_370), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_SL g518 ( .A1(n_342), .A2(n_370), .B(n_519), .C(n_521), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g357 ( .A1(n_343), .A2(n_358), .B1(n_363), .B2(n_366), .C(n_369), .Y(n_357) );
INVx1_ASAP7_75t_L g450 ( .A(n_343), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_343), .B(n_499), .Y(n_498) );
OAI22xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B1(n_350), .B2(n_352), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g427 ( .A(n_348), .B(n_362), .Y(n_427) );
AND2x2_ASAP7_75t_L g485 ( .A(n_348), .B(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g393 ( .A(n_349), .B(n_356), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_349), .B(n_362), .Y(n_421) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_351), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_351), .B(n_429), .Y(n_483) );
OAI321xp33_ASAP7_75t_L g502 ( .A1(n_351), .A2(n_424), .A3(n_503), .B1(n_504), .B2(n_505), .C(n_506), .Y(n_502) );
INVx1_ASAP7_75t_L g469 ( .A(n_352), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_353), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g408 ( .A(n_353), .B(n_356), .Y(n_408) );
AOI321xp33_ASAP7_75t_L g466 ( .A1(n_353), .A2(n_370), .A3(n_467), .B1(n_468), .B2(n_469), .C(n_470), .Y(n_466) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g383 ( .A(n_355), .B(n_368), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_356), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_356), .B(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_356), .B(n_442), .Y(n_479) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x4_ASAP7_75t_L g402 ( .A(n_360), .B(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g367 ( .A(n_361), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g475 ( .A(n_362), .Y(n_475) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_365), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g398 ( .A(n_370), .Y(n_398) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_372), .B(n_407), .Y(n_456) );
OR2x2_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
OR2x2_ASAP7_75t_L g420 ( .A(n_375), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_SL g465 ( .A(n_375), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_376), .A2(n_423), .B1(n_426), .B2(n_428), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
OR2x2_ASAP7_75t_L g520 ( .A(n_379), .B(n_443), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_384), .B1(n_388), .B2(n_394), .C(n_397), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx2_ASAP7_75t_L g418 ( .A(n_387), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_391), .Y(n_388) );
INVx1_ASAP7_75t_SL g464 ( .A(n_390), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_392), .B(n_442), .Y(n_441) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_392), .A2(n_460), .B(n_462), .Y(n_459) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x2_ASAP7_75t_L g505 ( .A(n_393), .B(n_487), .Y(n_505) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_SL g407 ( .A(n_396), .Y(n_407) );
AOI21xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g451 ( .A(n_403), .B(n_452), .Y(n_451) );
INVxp67_ASAP7_75t_L g513 ( .A(n_403), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_408), .B(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_407), .B(n_425), .Y(n_461) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g482 ( .A(n_411), .Y(n_482) );
NAND5xp2_ASAP7_75t_L g412 ( .A(n_413), .B(n_430), .C(n_439), .D(n_459), .E(n_466), .Y(n_412) );
O2A1O1Ixp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B(n_419), .C(n_422), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_426), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g468 ( .A(n_428), .Y(n_468) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_431), .A2(n_434), .B(n_436), .Y(n_430) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_431), .A2(n_485), .B1(n_488), .B2(n_490), .C(n_491), .Y(n_484) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
AOI321xp33_ASAP7_75t_L g439 ( .A1(n_432), .A2(n_440), .A3(n_444), .B1(n_445), .B2(n_451), .C(n_453), .Y(n_439) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g510 ( .A(n_444), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g445 ( .A(n_446), .B(n_450), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g462 ( .A(n_447), .B(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
NOR2xp67_ASAP7_75t_SL g474 ( .A(n_448), .B(n_455), .Y(n_474) );
AOI321xp33_ASAP7_75t_SL g506 ( .A1(n_451), .A2(n_507), .A3(n_508), .B1(n_509), .B2(n_510), .C(n_511), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_456), .C(n_457), .Y(n_453) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_464), .B(n_472), .Y(n_501) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .C(n_476), .Y(n_473) );
NOR3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_502), .C(n_514), .Y(n_477) );
OAI211xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .B(n_484), .C(n_494), .Y(n_478) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_482), .B(n_483), .Y(n_481) );
OAI221xp5_ASAP7_75t_L g514 ( .A1(n_483), .A2(n_515), .B1(n_516), .B2(n_517), .C(n_518), .Y(n_514) );
INVx1_ASAP7_75t_L g503 ( .A(n_485), .Y(n_503) );
INVx1_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_SL g507 ( .A(n_505), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
CKINVDCx14_ASAP7_75t_R g519 ( .A(n_520), .Y(n_519) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_523), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_540), .Y(n_539) );
endmodule