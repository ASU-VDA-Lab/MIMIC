module fake_jpeg_3557_n_552 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_552);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_552;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_55),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_42),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_58),
.B(n_76),
.Y(n_119)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_59),
.Y(n_137)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_60),
.Y(n_158)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_63),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_27),
.B(n_17),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_85),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

INVx6_ASAP7_75t_SL g75 ( 
.A(n_22),
.Y(n_75)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_20),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_77),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_22),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_78),
.B(n_86),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_27),
.B(n_17),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_20),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_103),
.Y(n_139)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_54),
.Y(n_97)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_99),
.B(n_101),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_100),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_30),
.B(n_16),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_21),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_32),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_22),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_105),
.B(n_107),
.Y(n_152)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_24),
.Y(n_106)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_24),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_48),
.C(n_32),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_111),
.B(n_31),
.C(n_49),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_89),
.A2(n_45),
.B1(n_37),
.B2(n_36),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_113),
.A2(n_159),
.B1(n_34),
.B2(n_23),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_130),
.Y(n_180)
);

BUFx12_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_121),
.B(n_165),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx12_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_131),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_104),
.B(n_48),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_65),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_91),
.A2(n_45),
.B1(n_48),
.B2(n_50),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_154),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_56),
.A2(n_50),
.B1(n_37),
.B2(n_47),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_62),
.A2(n_45),
.B1(n_40),
.B2(n_49),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_67),
.A2(n_50),
.B1(n_53),
.B2(n_21),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_64),
.A2(n_53),
.B1(n_26),
.B2(n_47),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_57),
.B(n_29),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_84),
.B(n_36),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_168),
.B(n_23),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

INVx3_ASAP7_75t_SL g239 ( 
.A(n_169),
.Y(n_239)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_170),
.Y(n_234)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_173),
.Y(n_255)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_174),
.Y(n_240)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_82),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g270 ( 
.A1(n_178),
.A2(n_183),
.B(n_214),
.Y(n_270)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_119),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_181),
.B(n_223),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_139),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_182),
.B(n_187),
.Y(n_228)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_184),
.Y(n_243)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_185),
.Y(n_271)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_127),
.Y(n_186)
);

BUFx2_ASAP7_75t_SL g254 ( 
.A(n_186),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_133),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_79),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_188),
.B(n_189),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_73),
.Y(n_189)
);

CKINVDCx12_ASAP7_75t_R g190 ( 
.A(n_110),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_190),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_209),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_26),
.B1(n_29),
.B2(n_39),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_219),
.B1(n_220),
.B2(n_109),
.Y(n_227)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_194),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_81),
.B1(n_69),
.B2(n_93),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_195),
.A2(n_215),
.B1(n_132),
.B2(n_160),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_152),
.A2(n_28),
.B1(n_49),
.B2(n_40),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_196),
.A2(n_199),
.B1(n_141),
.B2(n_123),
.Y(n_260)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_197),
.Y(n_268)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_198),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_125),
.A2(n_28),
.B1(n_40),
.B2(n_34),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_143),
.B(n_107),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_203),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g202 ( 
.A1(n_162),
.A2(n_106),
.B1(n_105),
.B2(n_101),
.Y(n_202)
);

AO21x2_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_221),
.B(n_117),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_143),
.B(n_39),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_163),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_206),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_110),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_207),
.B(n_208),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_167),
.Y(n_208)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_135),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_150),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_210),
.B(n_217),
.Y(n_261)
);

NAND3xp33_ASAP7_75t_SL g211 ( 
.A(n_118),
.B(n_31),
.C(n_19),
.Y(n_211)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_218),
.Y(n_231)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_212),
.B(n_141),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_112),
.B(n_34),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_141),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_128),
.B(n_99),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_109),
.A2(n_96),
.B1(n_92),
.B2(n_88),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_100),
.C(n_83),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_202),
.C(n_150),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_113),
.A2(n_31),
.B1(n_23),
.B2(n_28),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_125),
.A2(n_19),
.B1(n_22),
.B2(n_90),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_158),
.A2(n_19),
.B1(n_51),
.B2(n_41),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_128),
.B(n_16),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_225),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_126),
.B(n_15),
.Y(n_223)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_138),
.B(n_14),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_262),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_229),
.B(n_241),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_224),
.A2(n_158),
.B1(n_145),
.B2(n_120),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_250),
.B1(n_237),
.B2(n_247),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_237),
.A2(n_238),
.B1(n_247),
.B2(n_257),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_219),
.A2(n_132),
.B1(n_160),
.B2(n_153),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_245),
.B(n_214),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_195),
.A2(n_120),
.B1(n_166),
.B2(n_153),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_213),
.B(n_123),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_267),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_253),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_182),
.B(n_14),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_256),
.Y(n_306)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_218),
.A2(n_134),
.B1(n_114),
.B2(n_136),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_191),
.A2(n_134),
.B1(n_114),
.B2(n_136),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_258),
.A2(n_215),
.B1(n_209),
.B2(n_198),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_260),
.A2(n_265),
.B(n_192),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_178),
.B(n_123),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_175),
.B(n_14),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_186),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_210),
.A2(n_164),
.B1(n_117),
.B2(n_131),
.Y(n_265)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_221),
.A2(n_178),
.B1(n_202),
.B2(n_173),
.Y(n_266)
);

NOR2x1_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_237),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_172),
.B(n_1),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_274),
.Y(n_322)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_254),
.Y(n_275)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_241),
.B(n_180),
.C(n_216),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_276),
.B(n_294),
.C(n_314),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_277),
.A2(n_52),
.B1(n_51),
.B2(n_41),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_225),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_278),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_223),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_279),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_262),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_208),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_285),
.Y(n_317)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_244),
.Y(n_283)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_243),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_295),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_179),
.Y(n_285)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_286),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g349 ( 
.A(n_287),
.B(n_297),
.Y(n_349)
);

A2O1A1Ixp33_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_171),
.B(n_214),
.C(n_202),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_288),
.B(n_290),
.Y(n_319)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_289),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_241),
.B(n_236),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_304),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_228),
.B(n_174),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_293),
.B(n_298),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_229),
.B(n_170),
.C(n_194),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_273),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_246),
.B(n_212),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_300),
.Y(n_343)
);

NOR2x1p5_ASAP7_75t_L g297 ( 
.A(n_231),
.B(n_169),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_267),
.B(n_176),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_259),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_242),
.B(n_264),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_301),
.B(n_311),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_237),
.A2(n_177),
.B1(n_206),
.B2(n_205),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_302),
.A2(n_308),
.B1(n_309),
.B2(n_315),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_259),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_248),
.Y(n_307)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_237),
.A2(n_197),
.B1(n_184),
.B2(n_185),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_253),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_310),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_231),
.B(n_204),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_253),
.B(n_249),
.Y(n_323)
);

INVx13_ASAP7_75t_L g313 ( 
.A(n_239),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_313),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_258),
.B(n_201),
.C(n_192),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_266),
.A2(n_201),
.B1(n_131),
.B2(n_52),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_255),
.B(n_1),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_316),
.B(n_248),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_323),
.A2(n_333),
.B(n_345),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_281),
.B(n_294),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_337),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_282),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_332),
.B(n_298),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_297),
.A2(n_262),
.B(n_266),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_336),
.B(n_341),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_337),
.B(n_351),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_233),
.B(n_255),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_338),
.A2(n_340),
.B(n_349),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_299),
.A2(n_249),
.B1(n_235),
.B2(n_268),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_339),
.A2(n_277),
.B1(n_302),
.B2(n_329),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_287),
.A2(n_233),
.B(n_232),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_280),
.B(n_271),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_271),
.B(n_240),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g347 ( 
.A1(n_285),
.A2(n_252),
.A3(n_234),
.B1(n_240),
.B2(n_235),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_347),
.B(n_309),
.Y(n_356)
);

AOI32xp33_ASAP7_75t_L g348 ( 
.A1(n_292),
.A2(n_268),
.A3(n_272),
.B1(n_252),
.B2(n_234),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_350),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_276),
.B(n_232),
.C(n_272),
.Y(n_351)
);

NOR2xp67_ASAP7_75t_L g352 ( 
.A(n_280),
.B(n_239),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_303),
.A2(n_239),
.B1(n_52),
.B2(n_51),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_312),
.B(n_308),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_355),
.A2(n_299),
.B1(n_291),
.B2(n_310),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_356),
.B(n_364),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_333),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_358),
.B(n_359),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_360),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_361),
.A2(n_371),
.B1(n_353),
.B2(n_319),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_284),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g399 ( 
.A(n_363),
.B(n_368),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_322),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_377),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_300),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_374),
.C(n_351),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_287),
.Y(n_370)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_332),
.A2(n_318),
.B1(n_320),
.B2(n_315),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_372),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_345),
.Y(n_373)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_373),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_290),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_318),
.B(n_304),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_346),
.Y(n_378)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_378),
.Y(n_410)
);

AOI21xp33_ASAP7_75t_SL g380 ( 
.A1(n_320),
.A2(n_314),
.B(n_303),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_380),
.A2(n_388),
.B(n_389),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_317),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_385),
.Y(n_398)
);

AOI32xp33_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_296),
.A3(n_295),
.B1(n_288),
.B2(n_303),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_382),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_317),
.B(n_341),
.Y(n_383)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_383),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_316),
.Y(n_384)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_384),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_338),
.Y(n_385)
);

INVx13_ASAP7_75t_L g386 ( 
.A(n_328),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_386),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_275),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_387),
.B(n_330),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_344),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_330),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_369),
.B(n_342),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_393),
.B(n_404),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_356),
.A2(n_339),
.B1(n_319),
.B2(n_329),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_395),
.A2(n_412),
.B1(n_416),
.B2(n_423),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_306),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_400),
.B(n_406),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_388),
.A2(n_323),
.B(n_340),
.Y(n_401)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_401),
.Y(n_440)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_403),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_366),
.B(n_342),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_367),
.B(n_326),
.Y(n_406)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_409),
.B(n_366),
.C(n_358),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_SL g431 ( 
.A1(n_411),
.A2(n_383),
.B1(n_384),
.B2(n_379),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_362),
.A2(n_352),
.B1(n_349),
.B2(n_350),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_377),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_413),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_346),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_379),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_375),
.A2(n_348),
.B1(n_321),
.B2(n_347),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_368),
.Y(n_418)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_418),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_361),
.A2(n_381),
.B1(n_360),
.B2(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_419),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_373),
.A2(n_321),
.B1(n_328),
.B2(n_307),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_402),
.A2(n_380),
.B(n_363),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_427),
.B(n_421),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_433),
.Y(n_462)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_365),
.C(n_385),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_432),
.B(n_436),
.C(n_442),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g434 ( 
.A(n_415),
.B(n_365),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_439),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_382),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_435),
.B(n_450),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_370),
.C(n_378),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_395),
.A2(n_370),
.B1(n_389),
.B2(n_364),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_438),
.A2(n_414),
.B1(n_398),
.B2(n_416),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_411),
.B(n_376),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_441),
.Y(n_459)
);

XOR2x1_ASAP7_75t_SL g442 ( 
.A(n_414),
.B(n_386),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_443),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_392),
.Y(n_444)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_444),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_405),
.B(n_372),
.C(n_357),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_445),
.B(n_448),
.C(n_417),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_423),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_446),
.B(n_451),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_357),
.C(n_359),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_392),
.B(n_331),
.Y(n_450)
);

NOR2xp67_ASAP7_75t_L g451 ( 
.A(n_391),
.B(n_386),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_452),
.A2(n_455),
.B1(n_470),
.B2(n_440),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_437),
.A2(n_414),
.B1(n_391),
.B2(n_398),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_449),
.B(n_421),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_456),
.B(n_439),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_447),
.B(n_399),
.Y(n_457)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_457),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_444),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_469),
.Y(n_493)
);

AOI221xp5_ASAP7_75t_L g487 ( 
.A1(n_464),
.A2(n_445),
.B1(n_434),
.B2(n_396),
.C(n_435),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_465),
.B(n_433),
.Y(n_489)
);

BUFx24_ASAP7_75t_SL g466 ( 
.A(n_424),
.Y(n_466)
);

BUFx24_ASAP7_75t_SL g483 ( 
.A(n_466),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_402),
.C(n_417),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_473),
.C(n_436),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_429),
.A2(n_412),
.B1(n_420),
.B2(n_422),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_426),
.A2(n_438),
.B1(n_450),
.B2(n_420),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_430),
.Y(n_471)
);

INVx6_ASAP7_75t_L g488 ( 
.A(n_471),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_428),
.B(n_401),
.C(n_422),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_425),
.A2(n_396),
.B1(n_408),
.B2(n_397),
.Y(n_474)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_474),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_476),
.B(n_479),
.Y(n_494)
);

INVx8_ASAP7_75t_L g477 ( 
.A(n_472),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_477),
.B(n_481),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_491),
.B1(n_454),
.B2(n_461),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_465),
.B(n_432),
.C(n_448),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_453),
.A2(n_426),
.B1(n_440),
.B2(n_442),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_480),
.A2(n_410),
.B1(n_408),
.B2(n_397),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_455),
.Y(n_481)
);

INVx13_ASAP7_75t_L g484 ( 
.A(n_471),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_484),
.Y(n_504)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_463),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_489),
.Y(n_503)
);

BUFx12_ASAP7_75t_L g486 ( 
.A(n_467),
.Y(n_486)
);

CKINVDCx16_ASAP7_75t_R g498 ( 
.A(n_486),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_487),
.A2(n_492),
.B1(n_2),
.B2(n_3),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_490),
.B(n_354),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_470),
.A2(n_452),
.B1(n_460),
.B2(n_459),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_473),
.A2(n_461),
.B(n_454),
.Y(n_492)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_496),
.Y(n_516)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_497),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_462),
.C(n_468),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_499),
.B(n_500),
.Y(n_521)
);

FAx1_ASAP7_75t_SL g500 ( 
.A(n_478),
.B(n_456),
.CI(n_468),
.CON(n_500),
.SN(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_489),
.B(n_462),
.C(n_331),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_501),
.B(n_502),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_476),
.B(n_354),
.C(n_410),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_509),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_482),
.A2(n_305),
.B1(n_283),
.B2(n_313),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_506),
.B(n_508),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_488),
.B(n_286),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_507),
.B(n_484),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_41),
.C(n_25),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_493),
.B(n_2),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g513 ( 
.A(n_510),
.B(n_491),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_495),
.A2(n_477),
.B1(n_475),
.B2(n_480),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_512),
.B(n_513),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_514),
.B(n_515),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g515 ( 
.A(n_494),
.B(n_483),
.Y(n_515)
);

AO21x1_ASAP7_75t_L g518 ( 
.A1(n_496),
.A2(n_490),
.B(n_486),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_518),
.B(n_499),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g520 ( 
.A1(n_498),
.A2(n_488),
.B1(n_486),
.B2(n_6),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g533 ( 
.A(n_520),
.B(n_523),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_502),
.B(n_3),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_522),
.B(n_504),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_509),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_SL g524 ( 
.A1(n_503),
.A2(n_4),
.B(n_6),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_524),
.A2(n_497),
.B(n_508),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_526),
.B(n_527),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_501),
.C(n_506),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_530),
.B(n_531),
.Y(n_540)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_517),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_516),
.B(n_504),
.Y(n_532)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_532),
.A2(n_534),
.B(n_535),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_519),
.C(n_525),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_531),
.A2(n_518),
.B(n_500),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_536),
.A2(n_541),
.B(n_4),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_527),
.B(n_511),
.C(n_505),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_537),
.B(n_25),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g541 ( 
.A1(n_529),
.A2(n_500),
.B(n_524),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_539),
.B(n_528),
.Y(n_542)
);

AOI322xp5_ASAP7_75t_L g546 ( 
.A1(n_542),
.A2(n_543),
.A3(n_544),
.B1(n_545),
.B2(n_540),
.C1(n_25),
.C2(n_8),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_538),
.A2(n_511),
.B(n_533),
.Y(n_543)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_546),
.B(n_547),
.Y(n_548)
);

AOI322xp5_ASAP7_75t_L g547 ( 
.A1(n_542),
.A2(n_25),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_6),
.C2(n_11),
.Y(n_547)
);

AOI221xp5_ASAP7_75t_L g549 ( 
.A1(n_548),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_549)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_549),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_550),
.B(n_11),
.C(n_12),
.Y(n_551)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_12),
.B(n_13),
.Y(n_552)
);


endmodule