module fake_jpeg_31360_n_542 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_542);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_480;
wire n_267;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx8_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_0),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_55),
.Y(n_134)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_56),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_61),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_62),
.Y(n_158)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_64),
.Y(n_169)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_67),
.Y(n_151)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_68),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_83),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_0),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_76),
.B(n_82),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_77),
.Y(n_156)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_78),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_34),
.Y(n_79)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_18),
.B(n_0),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_87),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_19),
.Y(n_88)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_19),
.Y(n_91)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_2),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_103),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_2),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_106),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_22),
.Y(n_101)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_102),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_105),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_49),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_107),
.B(n_25),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_30),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_72),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

AO22x1_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_36),
.B1(n_25),
.B2(n_31),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_115),
.A2(n_166),
.B(n_50),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_100),
.A2(n_54),
.B1(n_52),
.B2(n_40),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_162),
.B1(n_42),
.B2(n_32),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_54),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_132),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_83),
.B(n_52),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_136),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_73),
.A2(n_24),
.B1(n_20),
.B2(n_46),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_140),
.A2(n_142),
.B1(n_157),
.B2(n_36),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_75),
.A2(n_24),
.B1(n_20),
.B2(n_46),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_90),
.B(n_23),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_155),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_60),
.B(n_40),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_93),
.A2(n_41),
.B1(n_38),
.B2(n_44),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_25),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_108),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_172),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_74),
.A2(n_48),
.B1(n_32),
.B2(n_42),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_99),
.B(n_38),
.C(n_35),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_165),
.B(n_29),
.C(n_50),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_L g166 ( 
.A1(n_109),
.A2(n_31),
.B(n_35),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_55),
.B(n_48),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_175),
.B(n_191),
.Y(n_231)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_176),
.Y(n_267)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

INVx13_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_133),
.A2(n_44),
.B(n_41),
.Y(n_180)
);

OR2x2_ASAP7_75t_SL g253 ( 
.A(n_180),
.B(n_171),
.Y(n_253)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_181),
.Y(n_264)
);

INVx8_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx11_ASAP7_75t_L g273 ( 
.A(n_182),
.Y(n_273)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx8_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_171),
.Y(n_185)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_185),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_123),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_186),
.B(n_192),
.Y(n_246)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

CKINVDCx6p67_ASAP7_75t_R g271 ( 
.A(n_188),
.Y(n_271)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

OA22x2_ASAP7_75t_SL g190 ( 
.A1(n_115),
.A2(n_36),
.B1(n_110),
.B2(n_96),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g242 ( 
.A(n_190),
.B(n_197),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_126),
.B(n_50),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_201),
.B1(n_221),
.B2(n_225),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_166),
.A2(n_65),
.B(n_68),
.C(n_102),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_29),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_198),
.B(n_203),
.Y(n_247)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_164),
.Y(n_199)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_156),
.A2(n_101),
.B1(n_84),
.B2(n_94),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_128),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_204),
.B(n_205),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_137),
.B(n_29),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_207),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_144),
.B(n_118),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_163),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_208),
.B(n_210),
.Y(n_254)
);

BUFx2_ASAP7_75t_SL g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_209),
.Y(n_268)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_170),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_212),
.Y(n_275)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_140),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_214),
.Y(n_235)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

CKINVDCx6p67_ASAP7_75t_R g215 ( 
.A(n_145),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_215),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_216),
.B(n_219),
.Y(n_259)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_146),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_220),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_148),
.B(n_29),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_223),
.Y(n_236)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_149),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_152),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_167),
.B(n_29),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_142),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_224),
.B(n_226),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_156),
.A2(n_87),
.B1(n_86),
.B2(n_79),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_136),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_169),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_125),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_244)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_134),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_121),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_238),
.B(n_185),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_161),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_239),
.B(n_256),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_241),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_174),
.B(n_121),
.C(n_122),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_245),
.B(n_257),
.C(n_188),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_253),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_177),
.B(n_124),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_222),
.B(n_122),
.C(n_151),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_197),
.B(n_124),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_57),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_219),
.B(n_157),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_17),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_222),
.A2(n_150),
.B1(n_134),
.B2(n_169),
.Y(n_265)
);

BUFx2_ASAP7_75t_SL g292 ( 
.A(n_265),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_196),
.A2(n_139),
.B1(n_151),
.B2(n_170),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_266),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_190),
.A2(n_129),
.B1(n_143),
.B2(n_158),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_270),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_190),
.A2(n_129),
.B1(n_143),
.B2(n_158),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_274),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_176),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_276),
.B(n_288),
.Y(n_320)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_277),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_231),
.A2(n_97),
.B1(n_225),
.B2(n_201),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_278),
.A2(n_306),
.B1(n_237),
.B2(n_242),
.Y(n_323)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_279),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_261),
.A2(n_62),
.B1(n_58),
.B2(n_69),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_280),
.A2(n_295),
.B1(n_269),
.B2(n_251),
.Y(n_317)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_281),
.Y(n_324)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_262),
.Y(n_282)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_282),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_262),
.Y(n_286)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_260),
.A2(n_215),
.B(n_195),
.C(n_206),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_289),
.A2(n_296),
.B(n_308),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_183),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_290),
.B(n_293),
.Y(n_327)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_184),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_250),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_294),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_261),
.A2(n_210),
.B1(n_208),
.B2(n_200),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_238),
.A2(n_215),
.B(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_297),
.B(n_309),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_259),
.B(n_182),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_246),
.B(n_3),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_300),
.B(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_193),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_303),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_246),
.B(n_3),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_247),
.B(n_50),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_305),
.B(n_254),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_231),
.A2(n_227),
.B1(n_4),
.B2(n_5),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_307),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_241),
.A2(n_50),
.B(n_179),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_234),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_317),
.A2(n_326),
.B1(n_338),
.B2(n_306),
.Y(n_367)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_259),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_319),
.B(n_285),
.C(n_312),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_284),
.B(n_247),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_339),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_323),
.A2(n_332),
.B1(n_333),
.B2(n_335),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_283),
.A2(n_259),
.B1(n_235),
.B2(n_231),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_292),
.A2(n_269),
.B1(n_268),
.B2(n_243),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_328),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_290),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_343),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_283),
.A2(n_242),
.B1(n_257),
.B2(n_245),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_311),
.A2(n_242),
.B1(n_253),
.B2(n_256),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_311),
.A2(n_239),
.B1(n_244),
.B2(n_252),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_295),
.A2(n_252),
.B1(n_254),
.B2(n_233),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_272),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_341),
.B(n_286),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_301),
.B(n_268),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_282),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_276),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_284),
.Y(n_347)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_348),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_317),
.A2(n_278),
.B1(n_298),
.B2(n_288),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_349),
.A2(n_357),
.B1(n_364),
.B2(n_367),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_303),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_368),
.C(n_315),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_329),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_351),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_316),
.A2(n_310),
.B(n_326),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_352),
.A2(n_362),
.B(n_373),
.Y(n_409)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_332),
.B(n_293),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_353),
.B(n_319),
.Y(n_385)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_318),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_354),
.Y(n_406)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_329),
.Y(n_356)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_356),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_317),
.A2(n_326),
.B1(n_342),
.B2(n_338),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

OAI32xp33_ASAP7_75t_L g361 ( 
.A1(n_327),
.A2(n_302),
.A3(n_305),
.B1(n_277),
.B2(n_279),
.Y(n_361)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_361),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_345),
.A2(n_299),
.B(n_308),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_343),
.A2(n_310),
.B1(n_302),
.B2(n_287),
.Y(n_364)
);

OAI32xp33_ASAP7_75t_L g365 ( 
.A1(n_327),
.A2(n_289),
.A3(n_280),
.B1(n_304),
.B2(n_300),
.Y(n_365)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_320),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_366),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_369),
.Y(n_399)
);

AO21x1_ASAP7_75t_L g370 ( 
.A1(n_345),
.A2(n_285),
.B(n_296),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_370),
.B(n_371),
.Y(n_408)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_340),
.Y(n_372)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_372),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_344),
.A2(n_281),
.B(n_297),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_330),
.B(n_309),
.Y(n_374)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_374),
.Y(n_396)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_318),
.Y(n_375)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_375),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_322),
.B(n_249),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_376),
.B(n_377),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_322),
.B(n_249),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_357),
.A2(n_323),
.B1(n_335),
.B2(n_333),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_379),
.A2(n_392),
.B1(n_393),
.B2(n_356),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_359),
.A2(n_334),
.B1(n_321),
.B2(n_315),
.Y(n_382)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_382),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_387),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_319),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_391),
.C(n_398),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_314),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_389),
.B(n_394),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_359),
.A2(n_314),
.B1(n_320),
.B2(n_328),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_349),
.A2(n_313),
.B1(n_316),
.B2(n_336),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_339),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_353),
.B(n_337),
.Y(n_398)
);

AOI21x1_ASAP7_75t_SL g401 ( 
.A1(n_370),
.A2(n_271),
.B(n_336),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_401),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_331),
.C(n_337),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_403),
.C(n_373),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_346),
.B(n_362),
.C(n_367),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_369),
.B(n_324),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_404),
.B(n_405),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_351),
.B(n_331),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_408),
.A2(n_352),
.B(n_355),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_410),
.A2(n_427),
.B(n_421),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_412),
.B(n_436),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_413),
.A2(n_388),
.B1(n_384),
.B2(n_382),
.Y(n_441)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_389),
.Y(n_414)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_414),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_389),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_418),
.Y(n_454)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_394),
.Y(n_417)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_386),
.B(n_346),
.Y(n_418)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_407),
.B(n_366),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_419),
.A2(n_421),
.B1(n_426),
.B2(n_430),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_399),
.B(n_365),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_420),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g421 ( 
.A(n_380),
.B(n_370),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_394),
.B(n_374),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_422),
.B(n_423),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_380),
.B(n_371),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_396),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_425),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

INVx13_ASAP7_75t_L g426 ( 
.A(n_406),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_SL g427 ( 
.A(n_409),
.B(n_361),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_388),
.A2(n_355),
.B1(n_364),
.B2(n_372),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_429),
.A2(n_416),
.B1(n_425),
.B2(n_414),
.Y(n_445)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_396),
.Y(n_430)
);

BUFx12_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_431),
.B(n_432),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_395),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_381),
.B(n_360),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_434),
.A2(n_438),
.B1(n_383),
.B2(n_291),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_391),
.B(n_294),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_437),
.B(n_428),
.C(n_402),
.Y(n_439)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_383),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_439),
.B(n_433),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_441),
.A2(n_443),
.B1(n_452),
.B2(n_459),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_442),
.A2(n_458),
.B(n_427),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_411),
.A2(n_384),
.B1(n_378),
.B2(n_398),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_445),
.B(n_271),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_403),
.C(n_385),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_451),
.C(n_453),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_428),
.B(n_378),
.C(n_393),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_379),
.B1(n_408),
.B2(n_390),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_436),
.B(n_400),
.C(n_390),
.Y(n_453)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_455),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_416),
.A2(n_419),
.B1(n_429),
.B2(n_410),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_456),
.A2(n_433),
.B1(n_430),
.B2(n_424),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_412),
.B(n_397),
.C(n_354),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_457),
.B(n_460),
.C(n_243),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_417),
.A2(n_397),
.B1(n_375),
.B2(n_358),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_358),
.C(n_325),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_SL g462 ( 
.A(n_461),
.B(n_435),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_462),
.B(n_463),
.Y(n_483)
);

CKINVDCx14_ASAP7_75t_R g463 ( 
.A(n_454),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_446),
.B(n_422),
.Y(n_464)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_464),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_456),
.B(n_426),
.Y(n_468)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_468),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_474),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_470),
.A2(n_443),
.B1(n_460),
.B2(n_441),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_471),
.B(n_472),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_448),
.B(n_423),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_448),
.A2(n_438),
.B1(n_431),
.B2(n_325),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_473),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_452),
.A2(n_431),
.B1(n_233),
.B2(n_251),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_449),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_478),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_477),
.C(n_479),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_234),
.C(n_232),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_232),
.C(n_240),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_240),
.C(n_258),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_480),
.B(n_450),
.C(n_459),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_485),
.Y(n_505)
);

BUFx24_ASAP7_75t_SL g485 ( 
.A(n_471),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_440),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_488),
.B(n_490),
.Y(n_501)
);

BUFx24_ASAP7_75t_SL g489 ( 
.A(n_469),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_267),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_465),
.A2(n_451),
.B1(n_447),
.B2(n_444),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_464),
.A2(n_442),
.B(n_440),
.Y(n_491)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_491),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_493),
.B(n_264),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_466),
.B(n_476),
.C(n_479),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_494),
.B(n_478),
.C(n_467),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_480),
.B(n_477),
.Y(n_496)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_496),
.Y(n_509)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_470),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_498),
.A2(n_499),
.B(n_506),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_481),
.A2(n_445),
.B(n_474),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_500),
.B(n_502),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g502 ( 
.A1(n_492),
.A2(n_467),
.B(n_271),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_495),
.A2(n_271),
.B1(n_273),
.B2(n_243),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_497),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_271),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_504),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_482),
.A2(n_240),
.B(n_273),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_255),
.C(n_258),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_487),
.C(n_486),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_487),
.A2(n_255),
.B1(n_264),
.B2(n_267),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_510),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_3),
.Y(n_519)
);

XNOR2x1_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_4),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_515),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_508),
.A2(n_497),
.B1(n_264),
.B2(n_267),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_516),
.B(n_519),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_509),
.A2(n_3),
.B(n_4),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_518),
.A2(n_502),
.B(n_8),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_506),
.C(n_510),
.Y(n_528)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_501),
.A2(n_5),
.B(n_6),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_522),
.A2(n_7),
.B(n_10),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_523),
.B(n_503),
.Y(n_525)
);

XNOR2x1_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_500),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_524),
.B(n_525),
.Y(n_531)
);

NAND4xp25_ASAP7_75t_SL g534 ( 
.A(n_528),
.B(n_530),
.C(n_520),
.D(n_507),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_529),
.A2(n_519),
.B(n_499),
.Y(n_533)
);

AOI211xp5_ASAP7_75t_L g532 ( 
.A1(n_527),
.A2(n_513),
.B(n_520),
.C(n_505),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_532),
.A2(n_526),
.B(n_504),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_534),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_536),
.A2(n_531),
.B1(n_10),
.B2(n_11),
.Y(n_537)
);

AOI322xp5_ASAP7_75t_L g538 ( 
.A1(n_537),
.A2(n_535),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C1(n_15),
.C2(n_16),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g539 ( 
.A1(n_538),
.A2(n_7),
.B(n_12),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_539),
.A2(n_7),
.B(n_13),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_540),
.A2(n_13),
.B(n_15),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_16),
.Y(n_542)
);


endmodule