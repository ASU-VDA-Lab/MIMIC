module fake_jpeg_31121_n_16 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_16);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_16;

wire n_13;
wire n_11;
wire n_14;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_15;
wire n_7;

OAI22xp5_ASAP7_75t_L g7 ( 
.A1(n_3),
.A2(n_6),
.B1(n_1),
.B2(n_4),
.Y(n_7)
);

AO22x1_ASAP7_75t_SL g8 ( 
.A1(n_4),
.A2(n_5),
.B1(n_0),
.B2(n_6),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_9),
.B(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

FAx1_ASAP7_75t_SL g11 ( 
.A(n_7),
.B(n_0),
.CI(n_2),
.CON(n_11),
.SN(n_11)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_11),
.A2(n_12),
.B1(n_8),
.B2(n_5),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_8),
.A2(n_0),
.B(n_2),
.Y(n_12)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_14),
.B(n_12),
.Y(n_15)
);

A2O1A1Ixp33_ASAP7_75t_L g16 ( 
.A1(n_15),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_16)
);


endmodule