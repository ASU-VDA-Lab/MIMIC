module real_aes_6681_n_271 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_271);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_271;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_528;
wire n_372;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_755;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_527;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_288;
wire n_756;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_649;
wire n_275;
wire n_385;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g731 ( .A(n_0), .Y(n_731) );
AOI22xp5_ASAP7_75t_SL g402 ( .A1(n_1), .A2(n_225), .B1(n_403), .B2(n_404), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g787 ( .A1(n_2), .A2(n_16), .B1(n_416), .B2(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g429 ( .A(n_3), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_4), .A2(n_110), .B1(n_336), .B2(n_785), .Y(n_784) );
AOI22xp5_ASAP7_75t_L g841 ( .A1(n_5), .A2(n_52), .B1(n_417), .B2(n_612), .Y(n_841) );
CKINVDCx20_ASAP7_75t_R g481 ( .A(n_6), .Y(n_481) );
INVx1_ASAP7_75t_L g718 ( .A(n_7), .Y(n_718) );
INVx1_ASAP7_75t_L g494 ( .A(n_8), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_9), .Y(n_486) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_10), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g293 ( .A(n_11), .Y(n_293) );
AOI22xp33_ASAP7_75t_SL g774 ( .A1(n_12), .A2(n_134), .B1(n_440), .B2(n_775), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_13), .A2(n_126), .B1(n_589), .B2(n_682), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_14), .A2(n_141), .B1(n_620), .B2(n_678), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_15), .A2(n_211), .B1(n_770), .B2(n_772), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g506 ( .A1(n_17), .A2(n_107), .B1(n_507), .B2(n_508), .C(n_509), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_18), .Y(n_410) );
CKINVDCx20_ASAP7_75t_R g478 ( .A(n_19), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g679 ( .A1(n_20), .A2(n_158), .B1(n_585), .B2(n_622), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_21), .B(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_22), .A2(n_102), .B1(n_503), .B2(n_556), .Y(n_657) );
INVx1_ASAP7_75t_L g725 ( .A(n_23), .Y(n_725) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_24), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_25), .Y(n_458) );
AO22x2_ASAP7_75t_L g299 ( .A1(n_26), .A2(n_83), .B1(n_300), .B2(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g830 ( .A(n_26), .Y(n_830) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_27), .B(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_28), .A2(n_268), .B1(n_404), .B2(n_440), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_29), .A2(n_200), .B1(n_327), .B2(n_416), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g582 ( .A1(n_30), .A2(n_151), .B1(n_400), .B2(n_406), .Y(n_582) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_31), .A2(n_269), .B1(n_360), .B2(n_678), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g847 ( .A1(n_32), .A2(n_246), .B1(n_397), .B2(n_805), .Y(n_847) );
INVx1_ASAP7_75t_L g724 ( .A(n_33), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g613 ( .A(n_34), .Y(n_613) );
INVx1_ASAP7_75t_L g843 ( .A(n_35), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g674 ( .A1(n_36), .A2(n_167), .B1(n_417), .B2(n_675), .Y(n_674) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_37), .A2(n_86), .B1(n_300), .B2(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g831 ( .A(n_37), .Y(n_831) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_38), .A2(n_129), .B1(n_337), .B2(n_413), .Y(n_467) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_39), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_40), .A2(n_154), .B1(n_403), .B2(n_440), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_41), .A2(n_255), .B1(n_420), .B2(n_518), .Y(n_789) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_42), .A2(n_153), .B1(n_406), .B2(n_407), .Y(n_405) );
CKINVDCx20_ASAP7_75t_R g344 ( .A(n_43), .Y(n_344) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_44), .A2(n_106), .B1(n_514), .B2(n_553), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g668 ( .A(n_45), .Y(n_668) );
AOI22xp33_ASAP7_75t_SL g549 ( .A1(n_46), .A2(n_65), .B1(n_370), .B2(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_47), .B(n_526), .Y(n_646) );
AOI22xp33_ASAP7_75t_SL g544 ( .A1(n_48), .A2(n_150), .B1(n_545), .B2(n_546), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_49), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_50), .A2(n_112), .B1(n_514), .B2(n_659), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g813 ( .A1(n_51), .A2(n_181), .B1(n_250), .B2(n_327), .C1(n_575), .C2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_53), .A2(n_55), .B1(n_380), .B2(n_559), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_54), .A2(n_70), .B1(n_440), .B2(n_711), .Y(n_710) );
AOI22xp5_ASAP7_75t_SL g398 ( .A1(n_56), .A2(n_147), .B1(n_399), .B2(n_400), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_57), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_57), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_58), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_59), .A2(n_498), .B1(n_499), .B2(n_528), .Y(n_497) );
INVx1_ASAP7_75t_L g528 ( .A(n_59), .Y(n_528) );
AOI221xp5_ASAP7_75t_L g516 ( .A1(n_60), .A2(n_94), .B1(n_517), .B2(n_518), .C(n_519), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_61), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_62), .A2(n_262), .B1(n_434), .B2(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_63), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_64), .A2(n_184), .B1(n_622), .B2(n_623), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g811 ( .A1(n_66), .A2(n_179), .B1(n_407), .B2(n_678), .Y(n_811) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_67), .B(n_420), .Y(n_543) );
AOI22xp33_ASAP7_75t_SL g677 ( .A1(n_68), .A2(n_189), .B1(n_587), .B2(n_678), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_69), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_71), .A2(n_157), .B1(n_365), .B2(n_655), .Y(n_778) );
AOI22xp5_ASAP7_75t_SL g394 ( .A1(n_72), .A2(n_136), .B1(n_395), .B2(n_397), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_73), .A2(n_213), .B1(n_420), .B2(n_423), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_74), .Y(n_570) );
AO22x2_ASAP7_75t_L g562 ( .A1(n_75), .A2(n_563), .B1(n_590), .B2(n_591), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g591 ( .A(n_75), .Y(n_591) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_76), .A2(n_224), .B1(n_584), .B2(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g644 ( .A(n_77), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g605 ( .A(n_78), .Y(n_605) );
AOI211xp5_ASAP7_75t_L g603 ( .A1(n_79), .A2(n_572), .B(n_604), .C(n_609), .Y(n_603) );
AOI22xp5_ASAP7_75t_SL g432 ( .A1(n_80), .A2(n_140), .B1(n_397), .B2(n_406), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_81), .A2(n_142), .B1(n_360), .B2(n_682), .Y(n_792) );
INVx1_ASAP7_75t_L g859 ( .A(n_82), .Y(n_859) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_84), .Y(n_474) );
AOI222xp33_ASAP7_75t_L g524 ( .A1(n_85), .A2(n_109), .B1(n_132), .B2(n_325), .C1(n_525), .C2(n_526), .Y(n_524) );
INVx1_ASAP7_75t_L g640 ( .A(n_87), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_88), .A2(n_194), .B1(n_381), .B2(n_515), .Y(n_796) );
AOI211xp5_ASAP7_75t_L g271 ( .A1(n_89), .A2(n_272), .B(n_280), .C(n_832), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_90), .Y(n_815) );
INVx1_ASAP7_75t_L g279 ( .A(n_91), .Y(n_279) );
INVx1_ASAP7_75t_L g712 ( .A(n_92), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_93), .A2(n_144), .B1(n_354), .B2(n_360), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_95), .A2(n_192), .B1(n_678), .B2(n_777), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_96), .B(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_SL g437 ( .A1(n_97), .A2(n_228), .B1(n_360), .B2(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g452 ( .A1(n_98), .A2(n_177), .B1(n_453), .B2(n_454), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_99), .A2(n_195), .B1(n_618), .B2(n_620), .Y(n_617) );
INVx1_ASAP7_75t_L g275 ( .A(n_100), .Y(n_275) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_101), .A2(n_135), .B1(n_354), .B2(n_559), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g669 ( .A1(n_103), .A2(n_139), .B1(n_327), .B2(n_337), .Y(n_669) );
AOI22xp33_ASAP7_75t_SL g795 ( .A1(n_104), .A2(n_159), .B1(n_384), .B2(n_655), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g840 ( .A(n_105), .B(n_518), .Y(n_840) );
INVx1_ASAP7_75t_L g469 ( .A(n_108), .Y(n_469) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_111), .A2(n_155), .B1(n_675), .B2(n_809), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g424 ( .A(n_113), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_114), .A2(n_210), .B1(n_327), .B2(n_416), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_115), .A2(n_163), .B1(n_371), .B2(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_116), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g733 ( .A(n_117), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_118), .A2(n_169), .B1(n_376), .B2(n_682), .Y(n_706) );
INVx1_ASAP7_75t_L g742 ( .A(n_119), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_120), .A2(n_199), .B1(n_374), .B2(n_380), .Y(n_373) );
XNOR2xp5_ASAP7_75t_L g532 ( .A(n_121), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_122), .B(n_541), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_123), .A2(n_715), .B1(n_743), .B2(n_744), .Y(n_714) );
CKINVDCx16_ASAP7_75t_R g743 ( .A(n_123), .Y(n_743) );
INVx1_ASAP7_75t_L g512 ( .A(n_124), .Y(n_512) );
INVx1_ASAP7_75t_L g702 ( .A(n_125), .Y(n_702) );
INVx1_ASAP7_75t_L g495 ( .A(n_127), .Y(n_495) );
AOI22xp5_ASAP7_75t_SL g635 ( .A1(n_128), .A2(n_636), .B1(n_660), .B2(n_661), .Y(n_635) );
INVx1_ASAP7_75t_L g661 ( .A(n_128), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_130), .A2(n_172), .B1(n_336), .B2(n_413), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g501 ( .A1(n_131), .A2(n_188), .B1(n_365), .B2(n_395), .C(n_502), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_133), .A2(n_204), .B1(n_545), .B2(n_546), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_137), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g278 ( .A(n_138), .B(n_279), .Y(n_278) );
AOI22xp33_ASAP7_75t_SL g538 ( .A1(n_143), .A2(n_212), .B1(n_325), .B2(n_453), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g610 ( .A(n_145), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_146), .A2(n_234), .B1(n_623), .B2(n_727), .Y(n_726) );
AND2x6_ASAP7_75t_L g274 ( .A(n_148), .B(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_148), .Y(n_824) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_149), .A2(n_221), .B1(n_300), .B2(n_304), .Y(n_309) );
CKINVDCx16_ASAP7_75t_R g601 ( .A(n_152), .Y(n_601) );
INVx1_ASAP7_75t_L g639 ( .A(n_156), .Y(n_639) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_160), .A2(n_193), .B1(n_395), .B2(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_161), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_162), .Y(n_483) );
CKINVDCx20_ASAP7_75t_R g451 ( .A(n_164), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g849 ( .A1(n_165), .A2(n_251), .B1(n_406), .B2(n_777), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_166), .B(n_335), .Y(n_334) );
CKINVDCx20_ASAP7_75t_R g456 ( .A(n_168), .Y(n_456) );
AOI22xp33_ASAP7_75t_SL g709 ( .A1(n_170), .A2(n_191), .B1(n_370), .B2(n_384), .Y(n_709) );
CKINVDCx20_ASAP7_75t_R g797 ( .A(n_171), .Y(n_797) );
INVx1_ASAP7_75t_L g649 ( .A(n_173), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_174), .A2(n_197), .B1(n_654), .B2(n_655), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_175), .A2(n_247), .B1(n_376), .B2(n_589), .Y(n_588) );
AO22x1_ASAP7_75t_L g502 ( .A1(n_176), .A2(n_215), .B1(n_503), .B2(n_504), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g681 ( .A1(n_178), .A2(n_241), .B1(n_360), .B2(n_682), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g684 ( .A(n_180), .Y(n_684) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_182), .A2(n_237), .B1(n_300), .B2(n_301), .Y(n_307) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_183), .A2(n_257), .B1(n_336), .B2(n_675), .Y(n_703) );
INVx1_ASAP7_75t_L g645 ( .A(n_185), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_186), .A2(n_242), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g631 ( .A(n_187), .Y(n_631) );
INVx1_ASAP7_75t_L g466 ( .A(n_190), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_196), .A2(n_263), .B1(n_527), .B2(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g491 ( .A(n_198), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_201), .B(n_699), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_202), .A2(n_243), .B1(n_395), .B2(n_400), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_203), .A2(n_220), .B1(n_556), .B2(n_557), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_205), .Y(n_333) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_206), .B(n_404), .Y(n_479) );
INVx1_ASAP7_75t_L g763 ( .A(n_207), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_208), .A2(n_240), .B1(n_515), .B2(n_584), .Y(n_812) );
INVx1_ASAP7_75t_L g737 ( .A(n_209), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g580 ( .A(n_214), .Y(n_580) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_216), .Y(n_627) );
AOI22xp33_ASAP7_75t_SL g848 ( .A1(n_217), .A2(n_226), .B1(n_380), .B2(n_711), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g340 ( .A(n_218), .Y(n_340) );
INVx1_ASAP7_75t_L g759 ( .A(n_219), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_221), .B(n_829), .Y(n_828) );
XOR2xp5_ASAP7_75t_L g833 ( .A(n_222), .B(n_834), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g671 ( .A(n_223), .B(n_518), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_227), .A2(n_266), .B1(n_365), .B2(n_368), .Y(n_364) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_229), .Y(n_488) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_230), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_231), .A2(n_245), .B1(n_518), .B2(n_607), .Y(n_807) );
INVx1_ASAP7_75t_L g648 ( .A(n_232), .Y(n_648) );
INVx1_ASAP7_75t_L g741 ( .A(n_233), .Y(n_741) );
INVx1_ASAP7_75t_L g510 ( .A(n_235), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_236), .A2(n_249), .B1(n_383), .B2(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g827 ( .A(n_237), .Y(n_827) );
AOI22xp33_ASAP7_75t_SL g766 ( .A1(n_238), .A2(n_239), .B1(n_767), .B2(n_768), .Y(n_766) );
INVx1_ASAP7_75t_L g721 ( .A(n_244), .Y(n_721) );
OA22x2_ASAP7_75t_L g288 ( .A1(n_248), .A2(n_289), .B1(n_290), .B2(n_390), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_248), .Y(n_289) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_252), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_253), .Y(n_521) );
INVx1_ASAP7_75t_L g300 ( .A(n_254), .Y(n_300) );
INVx1_ASAP7_75t_L g302 ( .A(n_254), .Y(n_302) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_256), .Y(n_537) );
INVx1_ASAP7_75t_L g756 ( .A(n_258), .Y(n_756) );
INVx1_ASAP7_75t_L g735 ( .A(n_259), .Y(n_735) );
INVx1_ASAP7_75t_L g755 ( .A(n_260), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_261), .A2(n_270), .B1(n_327), .B2(n_453), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_264), .Y(n_783) );
INVx1_ASAP7_75t_L g762 ( .A(n_265), .Y(n_762) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_267), .Y(n_310) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_275), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g857 ( .A1(n_276), .A2(n_822), .B(n_858), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g276 ( .A(n_277), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI221xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_595), .B1(n_817), .B2(n_818), .C(n_819), .Y(n_280) );
INVx1_ASAP7_75t_L g817 ( .A(n_281), .Y(n_817) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_283), .B1(n_459), .B2(n_594), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI22xp5_ASAP7_75t_SL g283 ( .A1(n_284), .A2(n_285), .B1(n_426), .B2(n_427), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
HB1xp67_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_391), .B1(n_392), .B2(n_425), .Y(n_287) );
INVx1_ASAP7_75t_L g425 ( .A(n_288), .Y(n_425) );
INVx1_ASAP7_75t_L g390 ( .A(n_290), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_351), .Y(n_290) );
NOR3xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_316), .C(n_339), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_294), .B1(n_310), .B2(n_311), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_294), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_754) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g567 ( .A(n_295), .Y(n_567) );
INVx1_ASAP7_75t_SL g732 ( .A(n_295), .Y(n_732) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_296), .Y(n_450) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_296), .A2(n_466), .B(n_467), .Y(n_465) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_305), .Y(n_296) );
INVx2_ASAP7_75t_L g379 ( .A(n_297), .Y(n_379) );
OR2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_303), .Y(n_297) );
AND2x2_ASAP7_75t_L g315 ( .A(n_298), .B(n_303), .Y(n_315) );
AND2x2_ASAP7_75t_L g359 ( .A(n_298), .B(n_331), .Y(n_359) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g320 ( .A(n_299), .B(n_303), .Y(n_320) );
AND2x2_ASAP7_75t_L g332 ( .A(n_299), .B(n_309), .Y(n_332) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g304 ( .A(n_302), .Y(n_304) );
INVx2_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
INVx1_ASAP7_75t_L g389 ( .A(n_303), .Y(n_389) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2x1p5_ASAP7_75t_L g314 ( .A(n_306), .B(n_315), .Y(n_314) );
AND2x4_ASAP7_75t_L g381 ( .A(n_306), .B(n_359), .Y(n_381) );
AND2x4_ASAP7_75t_L g422 ( .A(n_306), .B(n_379), .Y(n_422) );
AND2x6_ASAP7_75t_L g423 ( .A(n_306), .B(n_315), .Y(n_423) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
INVx1_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
INVx1_ASAP7_75t_L g350 ( .A(n_307), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_307), .B(n_309), .Y(n_363) );
AND2x2_ASAP7_75t_L g321 ( .A(n_308), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g358 ( .A(n_309), .B(n_350), .Y(n_358) );
OAI211xp5_ASAP7_75t_L g604 ( .A1(n_311), .A2(n_605), .B(n_606), .C(n_608), .Y(n_604) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_313), .A2(n_342), .B1(n_469), .B2(n_470), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_313), .A2(n_731), .B1(n_732), .B2(n_733), .Y(n_730) );
BUFx3_ASAP7_75t_L g757 ( .A(n_313), .Y(n_757) );
BUFx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g444 ( .A(n_314), .Y(n_444) );
AND2x4_ASAP7_75t_L g371 ( .A(n_315), .B(n_321), .Y(n_371) );
AND2x2_ASAP7_75t_L g386 ( .A(n_315), .B(n_358), .Y(n_386) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_315), .B(n_358), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_323), .B1(n_324), .B2(n_333), .C(n_334), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI22xp5_ASAP7_75t_SL g455 ( .A1(n_318), .A2(n_456), .B1(n_457), .B2(n_458), .Y(n_455) );
INVx4_ASAP7_75t_L g814 ( .A(n_318), .Y(n_814) );
INVx4_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g411 ( .A(n_319), .Y(n_411) );
INVx2_ASAP7_75t_SL g473 ( .A(n_319), .Y(n_473) );
BUFx6f_ASAP7_75t_L g525 ( .A(n_319), .Y(n_525) );
BUFx3_ASAP7_75t_L g572 ( .A(n_319), .Y(n_572) );
INVx2_ASAP7_75t_L g667 ( .A(n_319), .Y(n_667) );
AND2x6_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g347 ( .A(n_320), .Y(n_347) );
AND2x4_ASAP7_75t_L g413 ( .A(n_320), .B(n_349), .Y(n_413) );
AND2x2_ASAP7_75t_L g367 ( .A(n_321), .B(n_359), .Y(n_367) );
AND2x6_ASAP7_75t_L g378 ( .A(n_321), .B(n_379), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_324), .A2(n_643), .B1(n_644), .B2(n_645), .C(n_646), .Y(n_642) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI22xp5_ASAP7_75t_L g471 ( .A1(n_326), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_471) );
INVx4_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx2_ASAP7_75t_L g457 ( .A(n_327), .Y(n_457) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx2_ASAP7_75t_L g574 ( .A(n_328), .Y(n_574) );
BUFx6f_ASAP7_75t_L g612 ( .A(n_328), .Y(n_612) );
BUFx4f_ASAP7_75t_SL g788 ( .A(n_328), .Y(n_788) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_332), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g338 ( .A(n_330), .Y(n_338) );
INVx1_ASAP7_75t_L g343 ( .A(n_331), .Y(n_343) );
AND2x4_ASAP7_75t_L g337 ( .A(n_332), .B(n_338), .Y(n_337) );
NAND2x1p5_ASAP7_75t_L g342 ( .A(n_332), .B(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g417 ( .A(n_332), .B(n_418), .Y(n_417) );
BUFx4f_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g576 ( .A(n_336), .Y(n_576) );
BUFx12f_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_337), .Y(n_453) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_337), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B1(n_344), .B2(n_345), .Y(n_339) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx4_ASAP7_75t_L g447 ( .A(n_342), .Y(n_447) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_342), .A2(n_520), .B1(n_521), .B2(n_522), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_342), .A2(n_345), .B1(n_762), .B2(n_763), .Y(n_761) );
AND2x2_ASAP7_75t_L g404 ( .A(n_343), .B(n_362), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_345), .A2(n_446), .B1(n_648), .B2(n_649), .Y(n_647) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_346), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g577 ( .A1(n_346), .A2(n_578), .B1(n_579), .B2(n_580), .Y(n_577) );
OR2x6_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NOR2xp67_ASAP7_75t_L g351 ( .A(n_352), .B(n_372), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_364), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx4f_ASAP7_75t_SL g767 ( .A(n_356), .Y(n_767) );
BUFx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g406 ( .A(n_357), .Y(n_406) );
BUFx3_ASAP7_75t_L g682 ( .A(n_357), .Y(n_682) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_358), .B(n_359), .Y(n_492) );
AND2x4_ASAP7_75t_L g361 ( .A(n_359), .B(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx3_ASAP7_75t_L g403 ( .A(n_361), .Y(n_403) );
INVx1_ASAP7_75t_L g487 ( .A(n_361), .Y(n_487) );
BUFx3_ASAP7_75t_L g505 ( .A(n_361), .Y(n_505) );
BUFx3_ASAP7_75t_L g589 ( .A(n_361), .Y(n_589) );
BUFx2_ASAP7_75t_L g620 ( .A(n_361), .Y(n_620) );
BUFx2_ASAP7_75t_SL g768 ( .A(n_361), .Y(n_768) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
OR2x6_ASAP7_75t_L g388 ( .A(n_363), .B(n_389), .Y(n_388) );
INVx1_ASAP7_75t_SL g630 ( .A(n_365), .Y(n_630) );
BUFx6f_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx3_ASAP7_75t_L g556 ( .A(n_366), .Y(n_556) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_SL g399 ( .A(n_367), .Y(n_399) );
INVx2_ASAP7_75t_L g435 ( .A(n_367), .Y(n_435) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx3_ASAP7_75t_L g400 ( .A(n_371), .Y(n_400) );
INVx6_ASAP7_75t_L g482 ( .A(n_371), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_382), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_377), .B(n_494), .Y(n_493) );
INVx4_ASAP7_75t_L g557 ( .A(n_377), .Y(n_557) );
INVx2_ASAP7_75t_L g654 ( .A(n_377), .Y(n_654) );
INVx5_ASAP7_75t_SL g777 ( .A(n_377), .Y(n_777) );
INVx11_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx11_ASAP7_75t_L g396 ( .A(n_378), .Y(n_396) );
BUFx2_ASAP7_75t_L g503 ( .A(n_380), .Y(n_503) );
BUFx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx3_ASAP7_75t_L g407 ( .A(n_381), .Y(n_407) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_381), .Y(n_440) );
INVx2_ASAP7_75t_L g477 ( .A(n_381), .Y(n_477) );
BUFx3_ASAP7_75t_L g587 ( .A(n_381), .Y(n_587) );
BUFx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_384), .Y(n_659) );
INVx5_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g397 ( .A(n_385), .Y(n_397) );
INVx4_ASAP7_75t_L g554 ( .A(n_385), .Y(n_554) );
INVx2_ASAP7_75t_L g584 ( .A(n_385), .Y(n_584) );
INVx1_ASAP7_75t_L g622 ( .A(n_385), .Y(n_622) );
BUFx3_ASAP7_75t_L g728 ( .A(n_385), .Y(n_728) );
INVx8_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx6_ASAP7_75t_SL g515 ( .A(n_388), .Y(n_515) );
INVx1_ASAP7_75t_SL g623 ( .A(n_388), .Y(n_623) );
INVx1_ASAP7_75t_SL g711 ( .A(n_388), .Y(n_711) );
INVx1_ASAP7_75t_L g418 ( .A(n_389), .Y(n_418) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
XOR2x2_ASAP7_75t_L g392 ( .A(n_393), .B(n_424), .Y(n_392) );
NAND4xp75_ASAP7_75t_SL g393 ( .A(n_394), .B(n_398), .C(n_401), .D(n_408), .Y(n_393) );
INVx1_ASAP7_75t_L g626 ( .A(n_395), .Y(n_626) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx4_ASAP7_75t_L g438 ( .A(n_396), .Y(n_438) );
INVx2_ASAP7_75t_SL g720 ( .A(n_396), .Y(n_720) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_405), .Y(n_401) );
BUFx2_ASAP7_75t_L g508 ( .A(n_406), .Y(n_508) );
INVx1_ASAP7_75t_L g551 ( .A(n_406), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g408 ( .A(n_409), .B(n_414), .Y(n_408) );
OAI21xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B(n_412), .Y(n_409) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_413), .Y(n_454) );
BUFx3_ASAP7_75t_L g675 ( .A(n_413), .Y(n_675) );
BUFx2_ASAP7_75t_SL g785 ( .A(n_413), .Y(n_785) );
BUFx2_ASAP7_75t_SL g845 ( .A(n_413), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_419), .Y(n_414) );
BUFx3_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx2_ASAP7_75t_L g545 ( .A(n_417), .Y(n_545) );
BUFx2_ASAP7_75t_L g809 ( .A(n_417), .Y(n_809) );
BUFx6f_ASAP7_75t_L g517 ( .A(n_420), .Y(n_517) );
INVx5_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g607 ( .A(n_421), .Y(n_607) );
INVx2_ASAP7_75t_L g673 ( .A(n_421), .Y(n_673) );
INVx2_ASAP7_75t_L g699 ( .A(n_421), .Y(n_699) );
INVx4_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
BUFx4f_ASAP7_75t_L g518 ( .A(n_423), .Y(n_518) );
BUFx2_ASAP7_75t_L g697 ( .A(n_423), .Y(n_697) );
INVx1_ASAP7_75t_SL g426 ( .A(n_427), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
XNOR2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
NAND3x1_ASAP7_75t_SL g430 ( .A(n_431), .B(n_436), .C(n_441), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx3_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI22xp5_ASAP7_75t_SL g480 ( .A1(n_435), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_480) );
INVx3_ASAP7_75t_L g678 ( .A(n_435), .Y(n_678) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_439), .Y(n_436) );
INVx4_ASAP7_75t_L g619 ( .A(n_440), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_449), .C(n_455), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_445), .B1(n_446), .B2(n_448), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_443), .A2(n_566), .B1(n_567), .B2(n_568), .Y(n_565) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_SL g641 ( .A(n_444), .Y(n_641) );
INVx3_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g579 ( .A(n_447), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_450), .A2(n_451), .B(n_452), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g638 ( .A1(n_450), .A2(n_639), .B1(n_640), .B2(n_641), .Y(n_638) );
BUFx4f_ASAP7_75t_L g739 ( .A(n_453), .Y(n_739) );
INVx1_ASAP7_75t_SL g547 ( .A(n_454), .Y(n_547) );
INVx1_ASAP7_75t_L g594 ( .A(n_459), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_461), .B1(n_496), .B2(n_593), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
XNOR2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_495), .Y(n_462) );
AND3x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .C(n_484), .Y(n_463) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_468), .C(n_471), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
OAI21xp5_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_478), .B(n_479), .Y(n_476) );
INVx2_ASAP7_75t_L g507 ( .A(n_482), .Y(n_507) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_482), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
INVx3_ASAP7_75t_L g655 ( .A(n_482), .Y(n_655) );
OAI221xp5_ASAP7_75t_SL g723 ( .A1(n_482), .A2(n_632), .B1(n_724), .B2(n_725), .C(n_726), .Y(n_723) );
INVx2_ASAP7_75t_L g805 ( .A(n_482), .Y(n_805) );
NOR3xp33_ASAP7_75t_L g484 ( .A(n_485), .B(n_490), .C(n_493), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B1(n_488), .B2(n_489), .Y(n_485) );
BUFx2_ASAP7_75t_R g511 ( .A(n_489), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx1_ASAP7_75t_L g633 ( .A(n_492), .Y(n_633) );
INVx1_ASAP7_75t_L g593 ( .A(n_496), .Y(n_593) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_497), .A2(n_529), .B1(n_530), .B2(n_592), .Y(n_496) );
INVx1_ASAP7_75t_L g592 ( .A(n_497), .Y(n_592) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND4x1_ASAP7_75t_L g500 ( .A(n_501), .B(n_506), .C(n_516), .D(n_524), .Y(n_500) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_L g560 ( .A(n_505), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_512), .B2(n_513), .Y(n_509) );
CKINVDCx20_ASAP7_75t_R g513 ( .A(n_514), .Y(n_513) );
BUFx4f_ASAP7_75t_SL g514 ( .A(n_515), .Y(n_514) );
BUFx2_ASAP7_75t_L g585 ( .A(n_515), .Y(n_585) );
BUFx2_ASAP7_75t_L g772 ( .A(n_515), .Y(n_772) );
INVx1_ASAP7_75t_L g542 ( .A(n_518), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_522), .A2(n_579), .B1(n_741), .B2(n_742), .Y(n_740) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g536 ( .A(n_525), .Y(n_536) );
INVx2_ASAP7_75t_SL g643 ( .A(n_525), .Y(n_643) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
AO22x1_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_532), .B1(n_561), .B2(n_562), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
NAND4xp75_ASAP7_75t_SL g533 ( .A(n_534), .B(n_548), .C(n_555), .D(n_558), .Y(n_533) );
NOR2xp67_ASAP7_75t_L g534 ( .A(n_535), .B(n_539), .Y(n_534) );
OAI21xp5_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_537), .B(n_538), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .C(n_544), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g771 ( .A(n_554), .Y(n_771) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g590 ( .A(n_563), .Y(n_590) );
AND2x2_ASAP7_75t_SL g563 ( .A(n_564), .B(n_581), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_569), .C(n_577), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g569 ( .A1(n_570), .A2(n_571), .B(n_573), .Y(n_569) );
INVx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g736 ( .A(n_574), .Y(n_736) );
INVx1_ASAP7_75t_L g614 ( .A(n_575), .Y(n_614) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND4x1_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .C(n_586), .D(n_588), .Y(n_581) );
INVx1_ASAP7_75t_L g818 ( .A(n_595), .Y(n_818) );
XNOR2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_687), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B1(n_634), .B2(n_686), .Y(n_596) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
XNOR2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_615), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B1(n_613), .B2(n_614), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NOR3xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_624), .C(n_628), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_621), .Y(n_616) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_628) );
OAI221xp5_ASAP7_75t_SL g717 ( .A1(n_630), .A2(n_718), .B1(n_719), .B2(n_721), .C(n_722), .Y(n_717) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_SL g686 ( .A(n_634), .Y(n_686) );
OA22x2_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_662), .B1(n_663), .B2(n_685), .Y(n_634) );
INVx1_ASAP7_75t_L g685 ( .A(n_635), .Y(n_685) );
INVx2_ASAP7_75t_SL g660 ( .A(n_636), .Y(n_660) );
AND2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_650), .Y(n_636) );
NOR3xp33_ASAP7_75t_L g637 ( .A(n_638), .B(n_642), .C(n_647), .Y(n_637) );
OAI221xp5_ASAP7_75t_SL g734 ( .A1(n_643), .A2(n_735), .B1(n_736), .B2(n_737), .C(n_738), .Y(n_734) );
OAI21xp33_ASAP7_75t_SL g758 ( .A1(n_643), .A2(n_759), .B(n_760), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_651), .B(n_656), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx4_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
XOR2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_684), .Y(n_663) );
NAND3x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .C(n_680), .Y(n_664) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_670), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_668), .B(n_669), .Y(n_666) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_667), .A2(n_702), .B(n_703), .Y(n_701) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_667), .A2(n_783), .B(n_784), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g842 ( .A1(n_667), .A2(n_843), .B(n_844), .Y(n_842) );
NAND3xp33_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .C(n_674), .Y(n_670) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_681), .B(n_683), .Y(n_680) );
AOI22xp5_ASAP7_75t_SL g687 ( .A1(n_688), .A2(n_799), .B1(n_800), .B2(n_816), .Y(n_687) );
INVx1_ASAP7_75t_L g816 ( .A(n_688), .Y(n_816) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_745), .B2(n_746), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
XOR2x2_ASAP7_75t_L g690 ( .A(n_691), .B(n_713), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
XOR2x2_ASAP7_75t_SL g692 ( .A(n_693), .B(n_712), .Y(n_692) );
NAND2x1p5_ASAP7_75t_L g693 ( .A(n_694), .B(n_704), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_701), .Y(n_694) );
NAND3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_698), .C(n_700), .Y(n_695) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_705), .B(n_708), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_707), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g744 ( .A(n_715), .Y(n_744) );
AND2x2_ASAP7_75t_SL g715 ( .A(n_716), .B(n_729), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_723), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
NOR3xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_734), .C(n_740), .Y(n_729) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AO22x1_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B1(n_779), .B2(n_798), .Y(n_747) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g751 ( .A(n_752), .Y(n_751) );
AND2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_764), .Y(n_752) );
NOR3xp33_ASAP7_75t_L g753 ( .A(n_754), .B(n_758), .C(n_761), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_773), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_769), .Y(n_765) );
INVx3_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_774), .B(n_778), .Y(n_773) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx3_ASAP7_75t_SL g798 ( .A(n_779), .Y(n_798) );
XOR2x2_ASAP7_75t_L g779 ( .A(n_780), .B(n_797), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g780 ( .A(n_781), .B(n_790), .Y(n_780) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_782), .B(n_786), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_789), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx2_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
XOR2x2_ASAP7_75t_L g800 ( .A(n_801), .B(n_815), .Y(n_800) );
NAND4xp75_ASAP7_75t_L g801 ( .A(n_802), .B(n_806), .C(n_810), .D(n_813), .Y(n_801) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AND2x2_ASAP7_75t_SL g806 ( .A(n_807), .B(n_808), .Y(n_806) );
AND2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
INVx1_ASAP7_75t_SL g819 ( .A(n_820), .Y(n_819) );
NOR2x1_ASAP7_75t_L g820 ( .A(n_821), .B(n_825), .Y(n_820) );
OR2x2_ASAP7_75t_SL g863 ( .A(n_821), .B(n_826), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_823), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_823), .B(n_855), .Y(n_858) );
CKINVDCx16_ASAP7_75t_R g855 ( .A(n_824), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_826), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_827), .B(n_828), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_831), .Y(n_829) );
OAI322xp33_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_851), .A3(n_852), .B1(n_856), .B2(n_859), .C1(n_860), .C2(n_861), .Y(n_832) );
CKINVDCx20_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
HB1xp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
XOR2x2_ASAP7_75t_L g860 ( .A(n_836), .B(n_859), .Y(n_860) );
NAND4xp75_ASAP7_75t_SL g836 ( .A(n_837), .B(n_846), .C(n_849), .D(n_850), .Y(n_836) );
NOR2xp67_ASAP7_75t_SL g837 ( .A(n_838), .B(n_842), .Y(n_837) );
NAND3xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_840), .C(n_841), .Y(n_838) );
AND2x2_ASAP7_75t_L g846 ( .A(n_847), .B(n_848), .Y(n_846) );
HB1xp67_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
HB1xp67_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
CKINVDCx20_ASAP7_75t_R g856 ( .A(n_857), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_863), .Y(n_862) );
endmodule