module fake_jpeg_6188_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_1),
.B(n_0),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_2),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.C(n_1),
.Y(n_18)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_8),
.B(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_1),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_24),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_29),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_14),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_30),
.Y(n_35)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_12),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_11),
.C(n_16),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_23),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_30),
.A2(n_22),
.B1(n_9),
.B2(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_10),
.B1(n_15),
.B2(n_8),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_29),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_38),
.A2(n_33),
.B(n_35),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_22),
.B1(n_9),
.B2(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_41),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_22),
.B1(n_9),
.B2(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_21),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_36),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_7),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_39),
.C(n_42),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_2),
.C(n_3),
.Y(n_54)
);

OAI21x1_ASAP7_75t_SL g52 ( 
.A1(n_49),
.A2(n_45),
.B(n_48),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_54),
.Y(n_55)
);

OAI221xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_40),
.B1(n_17),
.B2(n_13),
.C(n_21),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_53),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_56),
.B(n_3),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_4),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_55),
.B(n_5),
.Y(n_59)
);

AOI322xp5_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_5),
.A3(n_6),
.B1(n_55),
.B2(n_57),
.C1(n_46),
.C2(n_47),
.Y(n_60)
);


endmodule