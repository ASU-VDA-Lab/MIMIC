module fake_jpeg_5041_n_44 (n_3, n_2, n_1, n_0, n_4, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_4),
.Y(n_7)
);

INVx2_ASAP7_75t_SL g8 ( 
.A(n_5),
.Y(n_8)
);

INVx5_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx2_ASAP7_75t_SL g11 ( 
.A(n_4),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_0),
.B(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_13),
.B(n_2),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_15),
.B(n_16),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_10),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_6),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_20),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_6),
.A2(n_1),
.B1(n_5),
.B2(n_10),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_6),
.A2(n_12),
.B1(n_9),
.B2(n_8),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_7),
.C(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_12),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_20),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_14),
.B(n_17),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_21),
.C(n_26),
.Y(n_34)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_7),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_28),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_SL g35 ( 
.A(n_32),
.B(n_8),
.C(n_11),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_34),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_16),
.B(n_19),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_39),
.B(n_22),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_26),
.B(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.C(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_33),
.Y(n_41)
);

OAI321xp33_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_8),
.A3(n_11),
.B1(n_18),
.B2(n_40),
.C(n_39),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_8),
.Y(n_44)
);


endmodule