module fake_jpeg_21791_n_49 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_49);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_49;

wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_40;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_32;

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_24),
.A2(n_13),
.B1(n_21),
.B2(n_20),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_30),
.B1(n_27),
.B2(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_26),
.A2(n_9),
.B1(n_19),
.B2(n_18),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_30),
.B(n_22),
.Y(n_32)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_1),
.Y(n_34)
);

XNOR2x1_ASAP7_75t_SL g39 ( 
.A(n_34),
.B(n_35),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_25),
.B(n_27),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_31),
.A2(n_8),
.B1(n_16),
.B2(n_3),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_42),
.B(n_43),
.C(n_35),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_42),
.A2(n_41),
.B1(n_38),
.B2(n_33),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_45),
.C(n_37),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_2),
.C(n_5),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_6),
.C(n_10),
.Y(n_49)
);


endmodule