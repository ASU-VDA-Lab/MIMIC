module fake_jpeg_955_n_200 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_200);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_200;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx10_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_6),
.A2(n_13),
.B(n_46),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_4),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_16),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_14),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_73),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_71),
.B(n_50),
.Y(n_80)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_48),
.B(n_45),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_52),
.Y(n_78)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_86),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_69),
.A2(n_56),
.B1(n_55),
.B2(n_63),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_80),
.B(n_85),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_50),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g93 ( 
.A1(n_81),
.A2(n_88),
.B(n_73),
.C(n_56),
.Y(n_93)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_71),
.B(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_53),
.Y(n_88)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_89),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_88),
.C(n_57),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_68),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_100),
.Y(n_113)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_108),
.C(n_77),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_57),
.B(n_55),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_67),
.C(n_54),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_30),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_105),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_69),
.B1(n_68),
.B2(n_75),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_84),
.B1(n_89),
.B2(n_47),
.Y(n_122)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_53),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_107),
.B(n_91),
.Y(n_111)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_110),
.B(n_111),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_112),
.A2(n_47),
.B(n_62),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_63),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_49),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_118),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_97),
.B(n_49),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_96),
.B(n_94),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_119),
.A2(n_102),
.B(n_108),
.Y(n_133)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_95),
.B(n_75),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_125),
.C(n_96),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_60),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_126),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_6),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_101),
.B(n_59),
.C(n_60),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_65),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_136),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_131),
.B(n_8),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_102),
.B1(n_61),
.B2(n_47),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_138),
.B1(n_9),
.B2(n_10),
.Y(n_160)
);

INVxp33_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_98),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_109),
.C(n_122),
.Y(n_151)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_47),
.B1(n_1),
.B2(n_2),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_119),
.A2(n_0),
.B(n_2),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_142),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_165)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_26),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_148),
.B(n_12),
.C(n_13),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_125),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_150),
.B(n_161),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_155),
.C(n_156),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_7),
.C(n_8),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_153),
.B(n_141),
.Y(n_170)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_23),
.B(n_43),
.C(n_42),
.D(n_39),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_20),
.C(n_38),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_44),
.C(n_37),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_163),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_160),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_12),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_141),
.B(n_144),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_169),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_170),
.B(n_172),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_164),
.A2(n_140),
.B1(n_147),
.B2(n_134),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_148),
.C(n_140),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_155),
.C(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_178),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_172),
.A2(n_157),
.B(n_151),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_182),
.A2(n_187),
.B(n_184),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_186),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_150),
.Y(n_186)
);

AOI322xp5_ASAP7_75t_L g187 ( 
.A1(n_174),
.A2(n_153),
.A3(n_167),
.B1(n_156),
.B2(n_35),
.C1(n_25),
.C2(n_33),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_180),
.A2(n_171),
.B1(n_173),
.B2(n_168),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_188),
.B(n_189),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_171),
.B1(n_168),
.B2(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_190),
.B(n_191),
.C(n_182),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_193),
.B(n_36),
.C(n_195),
.Y(n_197)
);

NOR3xp33_ASAP7_75t_SL g194 ( 
.A(n_189),
.B(n_186),
.C(n_185),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_192),
.B(n_28),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_196),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_198),
.B(n_197),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g200 ( 
.A(n_199),
.Y(n_200)
);


endmodule