module fake_jpeg_14939_n_82 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_82);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_82;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_6),
.B(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_11),
.B(n_3),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_21),
.B(n_29),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_25),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_23),
.A2(n_24),
.B1(n_26),
.B2(n_19),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_1),
.B1(n_5),
.B2(n_4),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_20),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_14),
.C(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_13),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_35),
.Y(n_45)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_27),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_17),
.B(n_14),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_14),
.C(n_19),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_34),
.B(n_30),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_57),
.C(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_41),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_56),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_31),
.B(n_33),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_SL g62 ( 
.A(n_52),
.B(n_45),
.C(n_49),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_62),
.A2(n_10),
.B(n_47),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_64),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_33),
.B1(n_41),
.B2(n_48),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_47),
.C(n_39),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_63),
.C(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_74),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_65),
.C(n_64),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_67),
.B1(n_44),
.B2(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_73),
.A2(n_68),
.B(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_68),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_76),
.B(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_78),
.Y(n_82)
);


endmodule