module real_jpeg_25021_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_150;
wire n_74;
wire n_32;
wire n_20;
wire n_80;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_4),
.B(n_46),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_4),
.B(n_49),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_54),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_4),
.B(n_64),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_4),
.B(n_28),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_4),
.B(n_17),
.Y(n_208)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_5),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_5),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_5),
.B(n_64),
.Y(n_94)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_6),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_7),
.B(n_64),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_7),
.B(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_7),
.B(n_54),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_7),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_7),
.B(n_28),
.Y(n_180)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_8),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_9),
.B(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_9),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_9),
.B(n_64),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_9),
.B(n_49),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_9),
.B(n_54),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_28),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_9),
.B(n_82),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_9),
.B(n_41),
.Y(n_235)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_11),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_41),
.Y(n_69)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_11),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_11),
.B(n_34),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_11),
.B(n_64),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_11),
.B(n_28),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_54),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_11),
.B(n_194),
.Y(n_193)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_13),
.B(n_28),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_13),
.B(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_13),
.B(n_49),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_13),
.B(n_17),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_54),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_14),
.B(n_41),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_14),
.B(n_28),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_14),
.B(n_174),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_15),
.B(n_28),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_15),
.B(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_16),
.B(n_49),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_41),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_16),
.B(n_64),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_16),
.B(n_28),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_16),
.B(n_46),
.Y(n_233)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_17),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_151),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_128),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_70),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_51),
.C(n_57),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_22),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.C(n_44),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_23),
.B(n_265),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_24),
.B(n_53),
.C(n_56),
.Y(n_117)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_30),
.CI(n_33),
.CON(n_24),
.SN(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_79),
.Y(n_78)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_36),
.A2(n_37),
.B(n_40),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_36),
.B(n_44),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_39),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.C(n_50),
.Y(n_44)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_45),
.B(n_48),
.CI(n_50),
.CON(n_132),
.SN(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_51),
.B(n_57),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_54),
.Y(n_214)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_66),
.C(n_68),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_58),
.B(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_62),
.C(n_63),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_59),
.B(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_60),
.B(n_214),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_62),
.B(n_63),
.Y(n_254)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_96),
.B2(n_127),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_86),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_77),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_76),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B1(n_84),
.B2(n_85),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_79),
.B(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_84),
.B1(n_88),
.B2(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_88),
.C(n_89),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_90),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_92),
.Y(n_276)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.CI(n_95),
.CON(n_92),
.SN(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_96),
.Y(n_273)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_117),
.CI(n_118),
.CON(n_96),
.SN(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_107),
.C(n_113),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_98),
.B(n_148),
.Y(n_147)
);

BUFx24_ASAP7_75t_SL g271 ( 
.A(n_98),
.Y(n_271)
);

FAx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_102),
.CI(n_105),
.CON(n_98),
.SN(n_98)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_102),
.C(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_113),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_111),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_126),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_122),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_147),
.C(n_149),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_129),
.A2(n_130),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_143),
.C(n_145),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_131),
.B(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.C(n_139),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_132),
.B(n_247),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g272 ( 
.A(n_132),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_133),
.A2(n_134),
.B1(n_139),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_135),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_139),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.C(n_142),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_140),
.B(n_141),
.CI(n_142),
.CON(n_228),
.SN(n_228)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_143),
.B(n_145),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_147),
.B(n_149),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_267),
.C(n_268),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_257),
.C(n_258),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_240),
.C(n_241),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_222),
.C(n_223),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_184),
.C(n_197),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_170),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_165),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_158),
.B(n_165),
.C(n_170),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.C(n_163),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_160),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_161),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_168),
.C(n_169),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_171),
.B(n_178),
.C(n_179),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_196)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_180),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_181),
.B(n_183),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.C(n_196),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_189),
.B1(n_196),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_218),
.C(n_219),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_206),
.C(n_211),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_204),
.C(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.C(n_215),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_230),
.C(n_239),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g274 ( 
.A(n_228),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_239),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_237),
.B2(n_238),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_236),
.C(n_238),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_237),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_249),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_244),
.B(n_245),
.C(n_249),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_253),
.C(n_255),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_252),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_266),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_263),
.C(n_264),
.Y(n_267)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_269),
.Y(n_270)
);


endmodule