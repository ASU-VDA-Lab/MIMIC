module fake_jpeg_15364_n_36 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_36);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_9),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_18),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_12),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_16),
.B(n_1),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_17),
.A2(n_16),
.B1(n_14),
.B2(n_4),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_21),
.A2(n_25),
.B1(n_3),
.B2(n_4),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_14),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_2),
.Y(n_28)
);

CKINVDCx10_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_26),
.A2(n_2),
.B(n_5),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_13),
.B1(n_3),
.B2(n_5),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_29),
.B(n_23),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_32),
.B(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_6),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_34),
.B(n_11),
.Y(n_36)
);


endmodule