module fake_jpeg_242_n_179 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_179);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_16),
.B(n_44),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_6),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_24),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_11),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_66),
.Y(n_73)
);

AOI21xp33_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_19),
.B(n_40),
.Y(n_67)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_67),
.A2(n_0),
.B(n_2),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_57),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_62),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_74),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_70),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_53),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_80),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_77),
.B(n_81),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_57),
.B1(n_53),
.B2(n_49),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_65),
.B1(n_66),
.B2(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_84),
.B(n_93),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_81),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_87),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_79),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_58),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_90),
.A2(n_63),
.B1(n_50),
.B2(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_50),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_94),
.Y(n_103)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_97),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_76),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_73),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_22),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_73),
.B1(n_58),
.B2(n_56),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_100),
.A2(n_106),
.B1(n_115),
.B2(n_10),
.Y(n_135)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

CKINVDCx6p67_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_56),
.B1(n_51),
.B2(n_65),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_63),
.B(n_59),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_5),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_108),
.A2(n_113),
.B1(n_116),
.B2(n_112),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_88),
.A2(n_61),
.B(n_47),
.C(n_63),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_114),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_45),
.B(n_2),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_9),
.B(n_10),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_88),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_96),
.B1(n_92),
.B2(n_94),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_91),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_101),
.C(n_109),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_119),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_86),
.C(n_25),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_129),
.B(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_104),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_6),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_124),
.B(n_125),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_111),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_126),
.A2(n_135),
.B1(n_12),
.B2(n_13),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_26),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_11),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_23),
.C(n_38),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_131),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_113),
.A2(n_110),
.B(n_100),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_7),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_7),
.Y(n_131)
);

CKINVDCx12_ASAP7_75t_R g134 ( 
.A(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_103),
.B(n_30),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_145),
.A2(n_149),
.B1(n_147),
.B2(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g146 ( 
.A(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_32),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_153),
.Y(n_155)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g153 ( 
.A1(n_137),
.A2(n_31),
.B(n_36),
.C(n_35),
.D(n_34),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_142),
.B(n_127),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_154),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_135),
.B1(n_120),
.B2(n_133),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_144),
.B1(n_150),
.B2(n_146),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_159),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_128),
.C(n_29),
.Y(n_160)
);

AO221x1_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_161),
.B1(n_153),
.B2(n_14),
.C(n_15),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_43),
.C(n_33),
.Y(n_161)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_163),
.A2(n_167),
.B1(n_157),
.B2(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_155),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_150),
.B1(n_138),
.B2(n_152),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_154),
.C(n_139),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_171),
.A2(n_170),
.B1(n_165),
.B2(n_168),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_148),
.C(n_166),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_172),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_172),
.B(n_14),
.C(n_15),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_13),
.C(n_17),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_177),
.A2(n_17),
.B(n_18),
.Y(n_178)
);

FAx1_ASAP7_75t_SL g179 ( 
.A(n_178),
.B(n_18),
.CI(n_177),
.CON(n_179),
.SN(n_179)
);


endmodule