module fake_jpeg_19995_n_236 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_236);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_236;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_2),
.B(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g88 ( 
.A(n_38),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx12f_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_60),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_24),
.Y(n_79)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_23),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_13),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_52),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_25),
.B(n_0),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_37),
.B1(n_21),
.B2(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_61),
.A2(n_82),
.B1(n_5),
.B2(n_7),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_63),
.B(n_72),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_37),
.B1(n_21),
.B2(n_30),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_68),
.Y(n_116)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_77),
.Y(n_107)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_26),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_80),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_17),
.Y(n_103)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_84),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_37),
.B1(n_19),
.B2(n_28),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_28),
.B1(n_20),
.B2(n_31),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_111)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_94),
.B(n_95),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_31),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_100),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_59),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_97),
.B(n_106),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_90),
.B(n_53),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_98),
.B(n_103),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_86),
.A2(n_19),
.B1(n_17),
.B2(n_22),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_104),
.B1(n_105),
.B2(n_88),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_66),
.Y(n_100)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_102),
.A2(n_111),
.B1(n_116),
.B2(n_91),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_34),
.B1(n_22),
.B2(n_3),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_34),
.B1(n_1),
.B2(n_3),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_0),
.Y(n_106)
);

OAI22x1_ASAP7_75t_L g135 ( 
.A1(n_108),
.A2(n_88),
.B1(n_76),
.B2(n_11),
.Y(n_135)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_117),
.Y(n_129)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_62),
.A2(n_68),
.B(n_82),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_114),
.B(n_118),
.C(n_9),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_74),
.B(n_13),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_8),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_65),
.B(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_124),
.Y(n_132)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

INVx3_ASAP7_75t_SL g123 ( 
.A(n_66),
.Y(n_123)
);

INVx5_ASAP7_75t_SL g139 ( 
.A(n_123),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_65),
.B(n_9),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_111),
.B1(n_114),
.B2(n_91),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_131),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_127),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_138),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_89),
.B1(n_70),
.B2(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_75),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_140),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_98),
.B(n_105),
.Y(n_161)
);

NAND2x1_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_118),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_109),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_15),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_142),
.B(n_103),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_145),
.Y(n_156)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_144),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_146),
.B(n_98),
.Y(n_159)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_149),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_102),
.B(n_121),
.C(n_100),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_165),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_132),
.C(n_125),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_167),
.Y(n_186)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_148),
.Y(n_154)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_159),
.B(n_160),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_161),
.A2(n_135),
.B1(n_127),
.B2(n_131),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_126),
.B1(n_67),
.B2(n_139),
.C(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_148),
.Y(n_163)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_124),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_106),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_168),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_118),
.C(n_83),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_102),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_170),
.B(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_172),
.A2(n_178),
.B(n_179),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_157),
.B(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_156),
.Y(n_200)
);

BUFx24_ASAP7_75t_SL g175 ( 
.A(n_160),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_153),
.Y(n_189)
);

OAI32xp33_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_130),
.A3(n_137),
.B1(n_149),
.B2(n_136),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_178),
.B(n_174),
.Y(n_192)
);

A2O1A1O1Ixp25_ASAP7_75t_L g178 ( 
.A1(n_162),
.A2(n_145),
.B(n_139),
.C(n_136),
.D(n_126),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_96),
.B1(n_139),
.B2(n_84),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_180),
.A2(n_184),
.B1(n_188),
.B2(n_151),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_141),
.B1(n_144),
.B2(n_83),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_158),
.A2(n_141),
.B1(n_123),
.B2(n_11),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_190),
.A2(n_193),
.B(n_195),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_174),
.A2(n_161),
.B1(n_155),
.B2(n_168),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_198),
.B1(n_199),
.B2(n_202),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_185),
.B(n_156),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_165),
.C(n_166),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_194),
.B(n_196),
.C(n_200),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_182),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_171),
.C(n_169),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_187),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_167),
.C(n_159),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_181),
.C(n_162),
.Y(n_208)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_197),
.A2(n_176),
.B(n_183),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_210),
.B(n_199),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_211),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_184),
.C(n_170),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_209),
.B(n_195),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_197),
.A2(n_192),
.B(n_202),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_172),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_188),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_198),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_204),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_214),
.B(n_216),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_218),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_190),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_213),
.Y(n_224)
);

A2O1A1Ixp33_ASAP7_75t_SL g219 ( 
.A1(n_207),
.A2(n_151),
.B(n_180),
.C(n_152),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_219),
.A2(n_152),
.B1(n_163),
.B2(n_154),
.Y(n_220)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_219),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_222),
.A2(n_150),
.B1(n_123),
.B2(n_85),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_224),
.B(n_225),
.C(n_150),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_213),
.B(n_210),
.C(n_203),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_223),
.A2(n_217),
.B(n_219),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_226),
.A2(n_225),
.B(n_221),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_227),
.B(n_229),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_228),
.A2(n_224),
.B(n_229),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_231),
.A2(n_9),
.B(n_85),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_233),
.B(n_232),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_235),
.B(n_234),
.Y(n_236)
);


endmodule