module fake_jpeg_3137_n_218 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_218);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_218;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_20),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_14),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_0),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_4),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_13),
.Y(n_76)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

CKINVDCx9p33_ASAP7_75t_R g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_51),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_60),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_76),
.B1(n_73),
.B2(n_66),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_81),
.B1(n_65),
.B2(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_55),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_95),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_67),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_97),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_66),
.Y(n_97)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_92),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_76),
.B1(n_73),
.B2(n_82),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_106),
.B1(n_79),
.B2(n_77),
.Y(n_119)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_98),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_108),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_86),
.A2(n_81),
.B1(n_60),
.B2(n_62),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_115),
.B(n_100),
.C(n_103),
.Y(n_126)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_94),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_116),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_64),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_114),
.B(n_72),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_91),
.A2(n_81),
.B1(n_69),
.B2(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_61),
.B1(n_57),
.B2(n_3),
.Y(n_135)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_1),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_120),
.B1(n_129),
.B2(n_135),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_62),
.B1(n_70),
.B2(n_79),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_59),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_124),
.B(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_54),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_128),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_112),
.B(n_75),
.C(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_111),
.B(n_56),
.Y(n_128)
);

AOI22x1_ASAP7_75t_SL g129 ( 
.A1(n_109),
.A2(n_71),
.B1(n_61),
.B2(n_57),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_58),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_0),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_SL g132 ( 
.A(n_108),
.B(n_61),
.C(n_57),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_132),
.B(n_48),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_124),
.B(n_1),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_142),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_123),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

BUFx24_ASAP7_75t_SL g144 ( 
.A(n_128),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_145),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_2),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_147),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_2),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_153),
.B1(n_154),
.B2(n_29),
.Y(n_162)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_3),
.B(n_4),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_6),
.B(n_7),
.Y(n_161)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_43),
.B1(n_42),
.B2(n_36),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_133),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_129),
.A2(n_132),
.B(n_137),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_155),
.A2(n_160),
.B(n_154),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_5),
.Y(n_159)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_5),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_169),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_165)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_165),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_28),
.C(n_27),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_175),
.C(n_178),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_150),
.B1(n_156),
.B2(n_148),
.Y(n_168)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_152),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_180),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_141),
.A2(n_25),
.B(n_23),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_158),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_11),
.C(n_12),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_153),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_168),
.A2(n_138),
.B(n_145),
.C(n_17),
.D(n_18),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_164),
.B(n_170),
.Y(n_200)
);

XOR2x2_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_15),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_172),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_15),
.C(n_16),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_16),
.C(n_18),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_19),
.C(n_178),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_173),
.Y(n_194)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_195),
.B(n_196),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_187),
.A2(n_165),
.B1(n_162),
.B2(n_180),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_174),
.B1(n_170),
.B2(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_184),
.B(n_19),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_199),
.A2(n_200),
.B(n_181),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_164),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_182),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_201),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_204),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_210),
.C(n_207),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_206),
.A2(n_182),
.B1(n_195),
.B2(n_186),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_211),
.A2(n_212),
.B(n_188),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_203),
.B(n_205),
.Y(n_212)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_213),
.B(n_214),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_215),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_209),
.C(n_202),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_202),
.Y(n_218)
);


endmodule