module fake_jpeg_8600_n_92 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_92);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx6_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_17),
.B(n_13),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

AND2x6_ASAP7_75t_SL g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp67_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_0),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_5),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

OAI21xp33_ASAP7_75t_SL g49 ( 
.A1(n_28),
.A2(n_1),
.B(n_2),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_68)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_51),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_1),
.B1(n_6),
.B2(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g55 ( 
.A(n_45),
.Y(n_55)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_9),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_12),
.B1(n_36),
.B2(n_43),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_40),
.A2(n_47),
.B1(n_35),
.B2(n_36),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_62),
.C(n_63),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_43),
.A2(n_34),
.B1(n_25),
.B2(n_32),
.Y(n_61)
);

AND2x6_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_64),
.Y(n_73)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_27),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_26),
.B(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_56),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_79),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_70),
.B(n_64),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_52),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_78),
.A2(n_67),
.B1(n_71),
.B2(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_75),
.A2(n_73),
.B1(n_49),
.B2(n_68),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_71),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_73),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_84),
.B1(n_80),
.B2(n_81),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_86),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_84),
.A2(n_72),
.B1(n_65),
.B2(n_74),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_76),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_87),
.B(n_61),
.Y(n_89)
);

OAI21x1_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_90),
.B(n_87),
.Y(n_91)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_74),
.A3(n_63),
.B1(n_46),
.B2(n_66),
.C1(n_37),
.C2(n_31),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_66),
.Y(n_92)
);


endmodule