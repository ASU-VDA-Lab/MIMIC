module fake_jpeg_4216_n_166 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_23),
.Y(n_35)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_24),
.B(n_27),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_33),
.A2(n_29),
.B(n_13),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_27),
.B(n_22),
.C(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_43),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

OR2x4_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_27),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_19),
.A3(n_40),
.B1(n_18),
.B2(n_13),
.Y(n_63)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_45),
.B(n_50),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_29),
.B1(n_23),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_47),
.A2(n_40),
.B1(n_23),
.B2(n_32),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_51),
.C(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_21),
.B(n_12),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_28),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_65),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_51),
.B(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_67),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_39),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_23),
.B1(n_14),
.B2(n_19),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_53),
.C(n_38),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_80),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_18),
.B(n_12),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_74),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_17),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_61),
.A2(n_32),
.B1(n_14),
.B2(n_21),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_25),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_81),
.A2(n_90),
.B(n_73),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_78),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_84),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_79),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_32),
.B1(n_61),
.B2(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_56),
.B1(n_13),
.B2(n_18),
.Y(n_105)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_64),
.Y(n_103)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_89),
.Y(n_96)
);

XNOR2x1_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_60),
.Y(n_91)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_69),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_102),
.C(n_87),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_71),
.B1(n_68),
.B2(n_70),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_101),
.B1(n_17),
.B2(n_16),
.Y(n_113)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_76),
.C(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_30),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_106),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_85),
.B(n_30),
.Y(n_106)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_88),
.B1(n_92),
.B2(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_107),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_94),
.B(n_97),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.C(n_113),
.Y(n_124)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_88),
.C(n_92),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_112),
.C(n_119),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_15),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_26),
.C(n_21),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_55),
.B1(n_34),
.B2(n_26),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_96),
.B1(n_34),
.B2(n_26),
.Y(n_121)
);

XNOR2x1_ASAP7_75t_L g119 ( 
.A(n_106),
.B(n_17),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_123),
.B1(n_34),
.B2(n_11),
.Y(n_140)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_119),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_125),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_128),
.C(n_129),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVxp67_ASAP7_75t_SL g131 ( 
.A(n_127),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_110),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_17),
.C(n_16),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_114),
.B(n_17),
.C(n_15),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_114),
.C(n_115),
.Y(n_134)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_136),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_137),
.C(n_138),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_116),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_109),
.C(n_17),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_15),
.C(n_20),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_20),
.C(n_11),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_1),
.C(n_2),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_140),
.B(n_11),
.Y(n_144)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_9),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_135),
.B(n_120),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_143),
.B(n_6),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g143 ( 
.A(n_131),
.B(n_10),
.C(n_1),
.Y(n_143)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_0),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_145),
.A2(n_3),
.B(n_5),
.Y(n_150)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_146),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_143),
.C(n_8),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_152),
.A2(n_153),
.B(n_7),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_147),
.A2(n_5),
.B(n_6),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_156),
.B(n_158),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_141),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_7),
.B(n_8),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_152),
.B(n_9),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_157),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

NAND2x1_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_162),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_164),
.Y(n_166)
);


endmodule