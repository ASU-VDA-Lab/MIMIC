module fake_jpeg_25577_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_14),
.B(n_12),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_45),
.B(n_30),
.Y(n_55)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_36),
.B1(n_23),
.B2(n_18),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_54),
.Y(n_77)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_59),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_65),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_32),
.B1(n_37),
.B2(n_40),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_57),
.A2(n_37),
.B1(n_48),
.B2(n_42),
.Y(n_86)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_64),
.B(n_27),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_36),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_89),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_38),
.C(n_44),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_105),
.Y(n_141)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_30),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_88),
.Y(n_128)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_84),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_86),
.A2(n_28),
.B1(n_19),
.B2(n_17),
.Y(n_122)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_30),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_60),
.B(n_23),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_37),
.B1(n_42),
.B2(n_32),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_111),
.B1(n_114),
.B2(n_39),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_60),
.B(n_20),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_92),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_66),
.B(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_63),
.B(n_33),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_94),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_97),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_99),
.B(n_103),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_72),
.Y(n_103)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_48),
.B(n_44),
.C(n_41),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_30),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_44),
.Y(n_135)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_108),
.Y(n_124)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_50),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_42),
.B1(n_47),
.B2(n_41),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_75),
.A2(n_42),
.B1(n_58),
.B2(n_43),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_74),
.B1(n_57),
.B2(n_68),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_116),
.A2(n_95),
.B1(n_84),
.B2(n_96),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_117),
.B(n_101),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_47),
.B1(n_27),
.B2(n_41),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_118),
.A2(n_120),
.B1(n_125),
.B2(n_129),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_88),
.A2(n_34),
.B1(n_26),
.B2(n_47),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_122),
.B1(n_109),
.B2(n_108),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_80),
.A2(n_47),
.B1(n_27),
.B2(n_41),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_79),
.A2(n_77),
.B1(n_90),
.B2(n_83),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_47),
.B1(n_44),
.B2(n_26),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_132),
.A2(n_143),
.B1(n_39),
.B2(n_24),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_82),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_44),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_105),
.A2(n_26),
.B1(n_34),
.B2(n_35),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_76),
.B(n_34),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_107),
.Y(n_168)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_145),
.B(n_146),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_138),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_147),
.B(n_151),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_118),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_152),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_141),
.A2(n_114),
.B(n_102),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_149),
.A2(n_155),
.B(n_159),
.Y(n_192)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_136),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_134),
.B(n_85),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_85),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_157),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_81),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_158),
.B(n_162),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_160),
.B(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_161),
.A2(n_165),
.B1(n_166),
.B2(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_130),
.B(n_104),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_163),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_115),
.B(n_28),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_135),
.A2(n_95),
.B1(n_97),
.B2(n_96),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_29),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_167),
.B(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_116),
.A2(n_94),
.B1(n_34),
.B2(n_26),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_29),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_35),
.B1(n_19),
.B2(n_17),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_171),
.A2(n_173),
.B1(n_131),
.B2(n_117),
.Y(n_193)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_172),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_115),
.B(n_24),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_22),
.B(n_24),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_22),
.B(n_107),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_121),
.B(n_0),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_179),
.Y(n_211)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_180),
.B(n_184),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_182),
.Y(n_229)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_147),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_132),
.C(n_143),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_186),
.C(n_207),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_126),
.C(n_140),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_122),
.C(n_133),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_202),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_193),
.A2(n_206),
.B1(n_155),
.B2(n_169),
.Y(n_213)
);

AOI21x1_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_125),
.B(n_140),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_101),
.B(n_98),
.Y(n_221)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_1),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_165),
.B(n_127),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_1),
.B(n_3),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_150),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_201),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_167),
.B(n_22),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_156),
.A2(n_139),
.B1(n_127),
.B2(n_138),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_153),
.B(n_139),
.C(n_131),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_189),
.B(n_177),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_209),
.B(n_218),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_153),
.Y(n_210)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_178),
.A2(n_156),
.B1(n_148),
.B2(n_173),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_223),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_155),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_214),
.B(n_219),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_159),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_227),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_204),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_159),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_178),
.A2(n_145),
.B1(n_151),
.B2(n_123),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_198),
.B1(n_184),
.B2(n_180),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_225),
.B(n_230),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_182),
.Y(n_224)
);

NOR4xp25_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_233),
.C(n_195),
.D(n_188),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_0),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_208),
.B(n_192),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_199),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_232),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_3),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_191),
.B(n_4),
.Y(n_231)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_231),
.Y(n_235)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_237),
.B(n_239),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_221),
.A2(n_192),
.B(n_200),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_213),
.A2(n_185),
.B1(n_200),
.B2(n_183),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_247),
.B1(n_255),
.B2(n_225),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_183),
.B(n_208),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_241),
.B(n_214),
.Y(n_266)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_211),
.B(n_226),
.Y(n_247)
);

AO22x1_ASAP7_75t_L g248 ( 
.A1(n_220),
.A2(n_190),
.B1(n_202),
.B2(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_186),
.C(n_6),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_222),
.C(n_234),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_211),
.A2(n_230),
.B1(n_232),
.B2(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_251),
.B(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_4),
.Y(n_252)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_252),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_SL g255 ( 
.A(n_215),
.B(n_4),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_256),
.A2(n_266),
.B(n_247),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_257),
.B(n_258),
.Y(n_278)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_272),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_219),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_268),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_222),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_271),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_245),
.B(n_217),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_229),
.C(n_8),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_273),
.C(n_252),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_253),
.B(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_270),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_7),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_7),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_7),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_259),
.A2(n_242),
.B1(n_254),
.B2(n_243),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_275),
.A2(n_276),
.B1(n_248),
.B2(n_10),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_261),
.A2(n_242),
.B1(n_243),
.B2(n_236),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_9),
.C(n_10),
.Y(n_297)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_269),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_256),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_285),
.Y(n_293)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_286),
.A2(n_260),
.B1(n_246),
.B2(n_251),
.Y(n_288)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_262),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_238),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_291),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_274),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_289),
.B(n_292),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_278),
.B(n_257),
.C(n_268),
.Y(n_291)
);

A2O1A1O1Ixp25_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_237),
.B(n_248),
.C(n_264),
.D(n_239),
.Y(n_294)
);

NOR2x1_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_297),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_238),
.B(n_235),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_9),
.B(n_10),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_298),
.B(n_11),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_276),
.C(n_279),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_300),
.B(n_304),
.Y(n_308)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_301),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_275),
.B1(n_286),
.B2(n_277),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_274),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_306),
.A2(n_11),
.B(n_12),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_302),
.A2(n_297),
.B1(n_279),
.B2(n_14),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_311),
.B1(n_312),
.B2(n_15),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_309),
.B(n_310),
.Y(n_313)
);

AND2x2_ASAP7_75t_SL g310 ( 
.A(n_300),
.B(n_12),
.Y(n_310)
);

AO21x1_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_299),
.B(n_303),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_308),
.A2(n_304),
.B1(n_15),
.B2(n_16),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_315),
.A2(n_14),
.B(n_16),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_313),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_314),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_316),
.Y(n_321)
);


endmodule