module real_jpeg_32240_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_0),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22x1_ASAP7_75t_L g158 ( 
.A1(n_0),
.A2(n_51),
.B1(n_159),
.B2(n_163),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_0),
.A2(n_51),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_0),
.B(n_83),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g295 ( 
.A1(n_0),
.A2(n_296),
.A3(n_301),
.B1(n_304),
.B2(n_312),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_0),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_0),
.B(n_156),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_1),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_1),
.Y(n_120)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_1),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_2),
.A2(n_15),
.B(n_414),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_2),
.B(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_5),
.Y(n_106)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_5),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_5),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_6),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_107)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_6),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_6),
.A2(n_111),
.B1(n_172),
.B2(n_174),
.Y(n_171)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_7),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_7),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_8),
.Y(n_89)
);

OAI22x1_ASAP7_75t_SL g53 ( 
.A1(n_9),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_9),
.A2(n_56),
.B1(n_65),
.B2(n_68),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_9),
.A2(n_56),
.B1(n_149),
.B2(n_152),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_9),
.A2(n_56),
.B1(n_251),
.B2(n_252),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_10),
.A2(n_123),
.B1(n_124),
.B2(n_126),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_10),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_123),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_11),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_13),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_233),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_231),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_200),
.B(n_201),
.Y(n_17)
);

NOR3xp33_ASAP7_75t_L g232 ( 
.A(n_18),
.B(n_200),
.C(n_201),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_167),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_19),
.B(n_167),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_61),
.C(n_96),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_20),
.A2(n_62),
.B1(n_63),
.B2(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_20),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_20),
.A2(n_204),
.B1(n_328),
.B2(n_333),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_20),
.A2(n_204),
.B1(n_207),
.B2(n_360),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_20),
.B(n_328),
.C(n_393),
.Y(n_392)
);

AOI22x1_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_47),
.B1(n_53),
.B2(n_60),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_21),
.Y(n_189)
);

AND2x4_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_37),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_32),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_32),
.Y(n_300)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_36),
.Y(n_311)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_37),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_37),
.A2(n_189),
.B(n_190),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_37),
.B(n_51),
.Y(n_355)
);

OA22x2_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B1(n_42),
.B2(n_45),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_40),
.Y(n_166)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_40),
.Y(n_317)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_44),
.Y(n_135)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_44),
.Y(n_155)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_47),
.Y(n_190)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_50),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_50),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_51),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_51),
.B(n_341),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_L g347 ( 
.A1(n_51),
.A2(n_136),
.B(n_348),
.Y(n_347)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_53),
.Y(n_188)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_61),
.Y(n_276)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_63),
.B(n_198),
.Y(n_397)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_71),
.B1(n_90),
.B2(n_95),
.Y(n_63)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_64),
.A2(n_95),
.B(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_67),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2x1p5_ASAP7_75t_L g184 ( 
.A(n_71),
.B(n_95),
.Y(n_184)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_72),
.B(n_91),
.Y(n_226)
);

NOR2x1_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_83),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_76),
.B1(n_79),
.B2(n_82),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g270 ( 
.A(n_82),
.Y(n_270)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_88),
.Y(n_83)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_88),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_91),
.B(n_184),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_93),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_97),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_129),
.Y(n_97)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_98),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_107),
.B1(n_117),
.B2(n_121),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_99),
.B(n_101),
.Y(n_181)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_100),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_100),
.A2(n_212),
.B1(n_217),
.B2(n_250),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_104),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_105),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_106),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_107),
.A2(n_211),
.B(n_216),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_116),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_122),
.B(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_128),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_129),
.B(n_243),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_129),
.B(n_285),
.C(n_293),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_129),
.A2(n_130),
.B1(n_354),
.B2(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_129),
.B(n_248),
.C(n_355),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_129),
.A2(n_293),
.B1(n_294),
.B2(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_130),
.Y(n_383)
);

AOI22x1_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_147),
.B1(n_156),
.B2(n_157),
.Y(n_130)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_131),
.A2(n_156),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_131),
.A2(n_156),
.B1(n_157),
.B2(n_209),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_136),
.B(n_141),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_132),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_134),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_135),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_136),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_139),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_138),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_141),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_171),
.B1(n_178),
.B2(n_179),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_141),
.B(n_330),
.C(n_331),
.Y(n_329)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_142),
.Y(n_253)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_155),
.Y(n_177)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_162),
.Y(n_303)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_185),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_182),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_170),
.A2(n_180),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_179),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_180),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_181),
.B(n_217),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

NAND2xp33_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_187),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_187),
.A2(n_198),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_195),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_198),
.B(n_246),
.C(n_276),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_198),
.B(n_288),
.C(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.C(n_227),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_202),
.A2(n_227),
.B1(n_228),
.B2(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_202),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_204),
.B(n_207),
.C(n_376),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_205),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_221),
.C(n_223),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_239),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_207),
.B(n_339),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_207),
.A2(n_339),
.B1(n_359),
.B2(n_360),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_207),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_207),
.A2(n_210),
.B1(n_360),
.B2(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g395 ( 
.A(n_210),
.Y(n_395)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_214),
.Y(n_290)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_216),
.A2(n_290),
.B(n_291),
.Y(n_289)
);

OAI211xp5_ASAP7_75t_L g292 ( 
.A1(n_216),
.A2(n_288),
.B(n_290),
.C(n_291),
.Y(n_292)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_225),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_223),
.B(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_225),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_280),
.B(n_412),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_277),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_236),
.B(n_277),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_242),
.C(n_244),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_238),
.B(n_242),
.Y(n_405)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_240),
.Y(n_393)
);

INVxp33_ASAP7_75t_SL g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_245),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_247),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_254),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_248),
.B(n_255),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_248),
.B(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_249),
.B(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_249),
.B(n_369),
.Y(n_370)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_250),
.Y(n_291)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21x1_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_259),
.B(n_268),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_386),
.B(n_406),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

OAI21x1_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_334),
.B(n_385),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_319),
.Y(n_283)
);

OR2x2_ASAP7_75t_L g385 ( 
.A(n_284),
.B(n_319),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_285),
.B(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_289),
.B(n_292),
.Y(n_287)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_289),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_289),
.B(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_318),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_295),
.B(n_318),
.Y(n_376)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

BUFx4f_ASAP7_75t_SL g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_308),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_326),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_324),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_321),
.B(n_326),
.C(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_324),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g357 ( 
.A(n_325),
.B(n_358),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_325),
.B(n_358),
.Y(n_371)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_328),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

AOI21x1_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_379),
.B(n_384),
.Y(n_334)
);

OAI21x1_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_373),
.B(n_378),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_356),
.B(n_372),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_352),
.Y(n_337)
);

NOR2xp67_ASAP7_75t_SL g372 ( 
.A(n_338),
.B(n_352),
.Y(n_372)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_339),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_343),
.B(n_347),
.Y(n_339)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

OAI21x1_ASAP7_75t_SL g356 ( 
.A1(n_357),
.A2(n_361),
.B(n_371),
.Y(n_356)
);

AOI21x1_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_368),
.B(n_370),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_367),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_374),
.B(n_375),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_377),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g384 ( 
.A(n_380),
.B(n_381),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_398),
.Y(n_386)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_390),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_396),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_402),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_402),
.Y(n_403)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_396),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_404),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g410 ( 
.A(n_399),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g399 ( 
.A1(n_400),
.A2(n_401),
.B(n_403),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_404),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_R g406 ( 
.A(n_407),
.B(n_409),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_411),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);


endmodule