module fake_ariane_502_n_798 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_798);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_798;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_754;
wire n_731;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_664;
wire n_629;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_61),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_118),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_36),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_138),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_56),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_35),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_16),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_23),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_4),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_16),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_47),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_102),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_27),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_103),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_82),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_112),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_10),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_104),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_97),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_19),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_73),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_57),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_88),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_58),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_45),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_51),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_142),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_30),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_133),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_90),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_78),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_21),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_48),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_69),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_28),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_53),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_17),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_110),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_33),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_98),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_5),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_147),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_86),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_15),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_152),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_100),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

AND2x4_ASAP7_75t_L g215 ( 
.A(n_167),
.B(n_0),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_0),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_200),
.Y(n_218)
);

OAI22x1_ASAP7_75t_R g219 ( 
.A1(n_169),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_197),
.Y(n_222)
);

AOI22x1_ASAP7_75t_SL g223 ( 
.A1(n_200),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_207),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

AND2x2_ASAP7_75t_R g226 ( 
.A(n_205),
.B(n_210),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_159),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

OAI22x1_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_6),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_165),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_163),
.Y(n_235)
);

AND2x4_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_7),
.Y(n_236)
);

BUFx8_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

OAI22x1_ASAP7_75t_SL g239 ( 
.A1(n_163),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_8),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

CKINVDCx11_ASAP7_75t_R g242 ( 
.A(n_161),
.Y(n_242)
);

AND2x4_ASAP7_75t_L g243 ( 
.A(n_179),
.B(n_9),
.Y(n_243)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_160),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_191),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_180),
.A2(n_11),
.B(n_12),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_11),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_192),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_191),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_166),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_211),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_171),
.B(n_172),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_218),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_220),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_222),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_242),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_218),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_176),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_242),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_216),
.A2(n_212),
.B1(n_209),
.B2(n_206),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_217),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_235),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_229),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_234),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_238),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_244),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_244),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_174),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_222),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_225),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_225),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_248),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_256),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_257),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_237),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_225),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_253),
.B(n_257),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_217),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_226),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_230),
.B(n_177),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_254),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_254),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_R g295 ( 
.A(n_233),
.B(n_181),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_254),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_225),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_251),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_227),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_254),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_237),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_251),
.Y(n_303)
);

NAND2xp33_ASAP7_75t_R g304 ( 
.A(n_246),
.B(n_182),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_251),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_251),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_243),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_280),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_282),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_282),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_261),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_243),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_278),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_265),
.B(n_232),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_285),
.B(n_232),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_273),
.B(n_274),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_282),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_268),
.Y(n_320)
);

NAND2xp33_ASAP7_75t_L g321 ( 
.A(n_275),
.B(n_293),
.Y(n_321)
);

AND2x6_ASAP7_75t_SL g322 ( 
.A(n_290),
.B(n_247),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_265),
.B(n_236),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_292),
.B(n_236),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_272),
.Y(n_326)
);

NAND2xp33_ASAP7_75t_L g327 ( 
.A(n_294),
.B(n_240),
.Y(n_327)
);

NAND2xp33_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_240),
.Y(n_328)
);

NOR3xp33_ASAP7_75t_L g329 ( 
.A(n_267),
.B(n_247),
.C(n_241),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_260),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_270),
.B(n_241),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_263),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_276),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_292),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_269),
.B(n_221),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_277),
.Y(n_337)
);

NAND2x1p5_ASAP7_75t_L g338 ( 
.A(n_262),
.B(n_215),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_303),
.B(n_250),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_271),
.B(n_221),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_283),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_228),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_295),
.B(n_215),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_249),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_302),
.B(n_231),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_279),
.B(n_227),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_282),
.B(n_288),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_297),
.B(n_227),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_258),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_299),
.B(n_227),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_288),
.B(n_301),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_288),
.B(n_185),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_186),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_298),
.B(n_187),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_298),
.B(n_188),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_264),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_300),
.Y(n_360)
);

INVxp33_ASAP7_75t_L g361 ( 
.A(n_266),
.Y(n_361)
);

NAND3xp33_ASAP7_75t_L g362 ( 
.A(n_304),
.B(n_246),
.C(n_199),
.Y(n_362)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_291),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_287),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_286),
.B(n_189),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_261),
.Y(n_367)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_286),
.B(n_190),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_286),
.B(n_193),
.Y(n_370)
);

AO221x1_ASAP7_75t_L g371 ( 
.A1(n_267),
.A2(n_219),
.B1(n_239),
.B2(n_223),
.C(n_15),
.Y(n_371)
);

NOR3xp33_ASAP7_75t_SL g372 ( 
.A(n_366),
.B(n_204),
.C(n_201),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_334),
.B(n_314),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_310),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_329),
.A2(n_198),
.B(n_196),
.C(n_195),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_12),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_313),
.B(n_13),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_329),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_379)
);

NOR2xp67_ASAP7_75t_L g380 ( 
.A(n_326),
.B(n_18),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_341),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_354),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_359),
.Y(n_384)
);

NAND3xp33_ASAP7_75t_SL g385 ( 
.A(n_307),
.B(n_14),
.C(n_20),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_342),
.B(n_158),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_349),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_324),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_370),
.B(n_26),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_309),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_29),
.Y(n_391)
);

OR2x6_ASAP7_75t_L g392 ( 
.A(n_332),
.B(n_31),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_322),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_319),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_324),
.A2(n_32),
.B1(n_34),
.B2(n_37),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_342),
.B(n_157),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_336),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_315),
.B(n_38),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_344),
.B(n_343),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_156),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g404 ( 
.A1(n_362),
.A2(n_39),
.B(n_40),
.Y(n_404)
);

OR2x6_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_41),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_343),
.B(n_155),
.Y(n_406)
);

AND2x6_ASAP7_75t_SL g407 ( 
.A(n_335),
.B(n_42),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_320),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_339),
.B(n_151),
.Y(n_409)
);

OR2x6_ASAP7_75t_L g410 ( 
.A(n_323),
.B(n_331),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_323),
.B(n_43),
.Y(n_411)
);

INVx4_ASAP7_75t_L g412 ( 
.A(n_319),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_325),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_318),
.B(n_44),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_319),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_318),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_338),
.B(n_46),
.Y(n_420)
);

AND2x4_ASAP7_75t_SL g421 ( 
.A(n_363),
.B(n_49),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_346),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_369),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_310),
.Y(n_424)
);

CKINVDCx8_ASAP7_75t_R g425 ( 
.A(n_361),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_360),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_338),
.B(n_50),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_369),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

NAND2x1p5_ASAP7_75t_L g430 ( 
.A(n_317),
.B(n_52),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_317),
.B(n_54),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_355),
.B(n_55),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_311),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_337),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_350),
.B(n_59),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_345),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_358),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_327),
.B(n_64),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_328),
.B(n_150),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_308),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_308),
.Y(n_441)
);

O2A1O1Ixp33_ASAP7_75t_L g442 ( 
.A1(n_376),
.A2(n_321),
.B(n_358),
.C(n_353),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_402),
.B(n_355),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_381),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_410),
.B(n_352),
.Y(n_445)
);

A2O1A1Ixp33_ASAP7_75t_L g446 ( 
.A1(n_403),
.A2(n_353),
.B(n_352),
.C(n_356),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_375),
.B(n_371),
.Y(n_447)
);

OA22x2_ASAP7_75t_L g448 ( 
.A1(n_394),
.A2(n_347),
.B1(n_357),
.B2(n_356),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_413),
.B(n_308),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_378),
.B(n_308),
.Y(n_450)
);

AOI21xp33_ASAP7_75t_L g451 ( 
.A1(n_411),
.A2(n_347),
.B(n_311),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_308),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_425),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_383),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_417),
.B(n_308),
.Y(n_455)
);

BUFx8_ASAP7_75t_L g456 ( 
.A(n_384),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_428),
.B(n_65),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_149),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_400),
.B(n_66),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_434),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_418),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_379),
.A2(n_67),
.B1(n_68),
.B2(n_70),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_426),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_439),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_377),
.B(n_75),
.Y(n_466)
);

O2A1O1Ixp33_ASAP7_75t_L g467 ( 
.A1(n_373),
.A2(n_76),
.B(n_77),
.C(n_79),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_395),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_434),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_387),
.B(n_81),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_386),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_398),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_372),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_422),
.B(n_87),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_410),
.B(n_89),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_436),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_382),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_429),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_416),
.B(n_95),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_405),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

BUFx3_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_393),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_397),
.B(n_96),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_399),
.A2(n_99),
.B1(n_101),
.B2(n_105),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_408),
.Y(n_489)
);

OA22x2_ASAP7_75t_L g490 ( 
.A1(n_392),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_441),
.A2(n_109),
.B(n_111),
.Y(n_491)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_421),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_113),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_392),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_R g495 ( 
.A(n_395),
.B(n_114),
.Y(n_495)
);

O2A1O1Ixp33_ASAP7_75t_L g496 ( 
.A1(n_385),
.A2(n_115),
.B(n_116),
.C(n_119),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_382),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_440),
.A2(n_121),
.B(n_122),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_380),
.B(n_123),
.Y(n_499)
);

INVx6_ASAP7_75t_SL g500 ( 
.A(n_407),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_445),
.B(n_395),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_461),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g503 ( 
.A1(n_446),
.A2(n_404),
.B(n_409),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_456),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_479),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_459),
.A2(n_420),
.B(n_427),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_453),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_445),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_470),
.A2(n_406),
.B(n_438),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_479),
.Y(n_513)
);

AO21x2_ASAP7_75t_L g514 ( 
.A1(n_450),
.A2(n_401),
.B(n_432),
.Y(n_514)
);

BUFx4_ASAP7_75t_SL g515 ( 
.A(n_484),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_482),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_464),
.Y(n_517)
);

OAI21xp33_ASAP7_75t_SL g518 ( 
.A1(n_493),
.A2(n_414),
.B(n_431),
.Y(n_518)
);

AND2x4_ASAP7_75t_L g519 ( 
.A(n_468),
.B(n_412),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_490),
.A2(n_391),
.B1(n_430),
.B2(n_388),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_485),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_460),
.Y(n_522)
);

INVx1_ASAP7_75t_SL g523 ( 
.A(n_447),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_469),
.Y(n_524)
);

NAND2x1p5_ASAP7_75t_L g525 ( 
.A(n_468),
.B(n_412),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_476),
.A2(n_389),
.B(n_374),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_494),
.B(n_374),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_472),
.B(n_433),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_485),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_474),
.Y(n_530)
);

BUFx2_ASAP7_75t_R g531 ( 
.A(n_466),
.Y(n_531)
);

OAI21x1_ASAP7_75t_L g532 ( 
.A1(n_499),
.A2(n_396),
.B(n_437),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_449),
.A2(n_491),
.B(n_498),
.Y(n_533)
);

AO21x2_ASAP7_75t_L g534 ( 
.A1(n_451),
.A2(n_391),
.B(n_415),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_443),
.A2(n_391),
.B(n_424),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g536 ( 
.A(n_477),
.Y(n_536)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_485),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_500),
.Y(n_538)
);

AOI22x1_ASAP7_75t_L g539 ( 
.A1(n_473),
.A2(n_475),
.B1(n_424),
.B2(n_433),
.Y(n_539)
);

NAND2x1p5_ASAP7_75t_L g540 ( 
.A(n_497),
.B(n_433),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_480),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_448),
.A2(n_391),
.B(n_415),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_497),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_455),
.B(n_424),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_442),
.A2(n_415),
.B(n_125),
.Y(n_545)
);

BUFx2_ASAP7_75t_SL g546 ( 
.A(n_492),
.Y(n_546)
);

AND2x4_ASAP7_75t_L g547 ( 
.A(n_497),
.B(n_124),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_458),
.Y(n_548)
);

AOI22x1_ASAP7_75t_L g549 ( 
.A1(n_487),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_508),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_SL g551 ( 
.A1(n_548),
.A2(n_457),
.B1(n_463),
.B2(n_452),
.Y(n_551)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_506),
.Y(n_552)
);

INVx6_ASAP7_75t_L g553 ( 
.A(n_529),
.Y(n_553)
);

INVx2_ASAP7_75t_SL g554 ( 
.A(n_515),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_548),
.A2(n_481),
.B1(n_478),
.B2(n_465),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_502),
.B(n_489),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_523),
.A2(n_489),
.B1(n_483),
.B2(n_486),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_510),
.B(n_454),
.Y(n_558)
);

INVx4_ASAP7_75t_L g559 ( 
.A(n_508),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_520),
.A2(n_500),
.B1(n_444),
.B2(n_488),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_522),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_517),
.Y(n_562)
);

AO21x1_ASAP7_75t_SL g563 ( 
.A1(n_520),
.A2(n_496),
.B(n_495),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_536),
.A2(n_471),
.B1(n_467),
.B2(n_134),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_502),
.A2(n_131),
.B1(n_132),
.B2(n_135),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_544),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_544),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_511),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_519),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_524),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_538),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_541),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_509),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_536),
.A2(n_136),
.B1(n_137),
.B2(n_139),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_SL g576 ( 
.A1(n_549),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_576)
);

BUFx8_ASAP7_75t_SL g577 ( 
.A(n_538),
.Y(n_577)
);

OAI21x1_ASAP7_75t_L g578 ( 
.A1(n_533),
.A2(n_144),
.B(n_146),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_501),
.B(n_148),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_513),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_501),
.A2(n_503),
.B1(n_518),
.B2(n_546),
.Y(n_581)
);

INVx5_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_501),
.A2(n_503),
.B1(n_530),
.B2(n_516),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_513),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_519),
.B(n_509),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_547),
.Y(n_586)
);

OAI21x1_ASAP7_75t_L g587 ( 
.A1(n_545),
.A2(n_507),
.B(n_512),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_515),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_547),
.Y(n_589)
);

AND2x4_ASAP7_75t_L g590 ( 
.A(n_519),
.B(n_537),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_547),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_534),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_526),
.A2(n_532),
.B(n_535),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_551),
.A2(n_516),
.B1(n_530),
.B2(n_542),
.Y(n_595)
);

AND2x4_ASAP7_75t_L g596 ( 
.A(n_585),
.B(n_537),
.Y(n_596)
);

AND2x4_ASAP7_75t_L g597 ( 
.A(n_585),
.B(n_543),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_562),
.B(n_568),
.Y(n_598)
);

BUFx4f_ASAP7_75t_SL g599 ( 
.A(n_588),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_583),
.B(n_543),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_577),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_592),
.Y(n_602)
);

NOR2x1p5_ASAP7_75t_L g603 ( 
.A(n_571),
.B(n_504),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_572),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_583),
.B(n_543),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_577),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_556),
.B(n_534),
.Y(n_607)
);

INVx3_ASAP7_75t_L g608 ( 
.A(n_552),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_592),
.Y(n_609)
);

BUFx2_ASAP7_75t_L g610 ( 
.A(n_566),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_555),
.A2(n_504),
.B1(n_505),
.B2(n_539),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_575),
.B(n_543),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_580),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_575),
.B(n_506),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_560),
.A2(n_505),
.B1(n_514),
.B2(n_531),
.Y(n_615)
);

OR2x2_ASAP7_75t_L g616 ( 
.A(n_566),
.B(n_506),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_561),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_R g618 ( 
.A(n_579),
.B(n_529),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_R g619 ( 
.A(n_554),
.B(n_521),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_584),
.B(n_521),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_561),
.Y(n_621)
);

NAND2xp33_ASAP7_75t_R g622 ( 
.A(n_579),
.B(n_540),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_560),
.A2(n_525),
.B1(n_540),
.B2(n_521),
.Y(n_623)
);

HB1xp67_ASAP7_75t_L g624 ( 
.A(n_573),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_570),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_573),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_581),
.B(n_521),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_593),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_581),
.B(n_525),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_586),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_567),
.B(n_514),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_567),
.B(n_594),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_550),
.Y(n_634)
);

NOR3xp33_ASAP7_75t_SL g635 ( 
.A(n_571),
.B(n_565),
.C(n_559),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_594),
.B(n_591),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_585),
.B(n_590),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_587),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_590),
.B(n_558),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_SL g640 ( 
.A(n_559),
.B(n_590),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_578),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_553),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_552),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_625),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_617),
.Y(n_645)
);

OA21x2_ASAP7_75t_L g646 ( 
.A1(n_638),
.A2(n_564),
.B(n_574),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_632),
.B(n_552),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_625),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_632),
.B(n_552),
.Y(n_649)
);

INVxp67_ASAP7_75t_SL g650 ( 
.A(n_607),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_604),
.B(n_569),
.Y(n_651)
);

BUFx3_ASAP7_75t_L g652 ( 
.A(n_642),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_598),
.B(n_569),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_627),
.B(n_582),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_621),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_613),
.B(n_633),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_610),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_621),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_610),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_607),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_630),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_630),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_620),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_640),
.A2(n_564),
.B(n_576),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_612),
.B(n_579),
.Y(n_665)
);

OAI221xp5_ASAP7_75t_L g666 ( 
.A1(n_611),
.A2(n_574),
.B1(n_557),
.B2(n_563),
.C(n_553),
.Y(n_666)
);

OAI221xp5_ASAP7_75t_L g667 ( 
.A1(n_615),
.A2(n_553),
.B1(n_582),
.B2(n_595),
.C(n_635),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_643),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_631),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_636),
.B(n_582),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_597),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_639),
.B(n_582),
.Y(n_672)
);

HB1xp67_ASAP7_75t_L g673 ( 
.A(n_620),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_631),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_602),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_609),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_624),
.B(n_626),
.Y(n_677)
);

AND2x4_ASAP7_75t_SL g678 ( 
.A(n_597),
.B(n_596),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_643),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_612),
.B(n_614),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_659),
.B(n_656),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_644),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_656),
.B(n_614),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_657),
.Y(n_684)
);

NAND3xp33_ASAP7_75t_L g685 ( 
.A(n_677),
.B(n_616),
.C(n_634),
.Y(n_685)
);

OAI22xp5_ASAP7_75t_L g686 ( 
.A1(n_664),
.A2(n_634),
.B1(n_642),
.B2(n_603),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_654),
.B(n_627),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_653),
.B(n_616),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_652),
.B(n_599),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_659),
.B(n_628),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_663),
.B(n_605),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_644),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_648),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_673),
.B(n_651),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_647),
.B(n_628),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_647),
.B(n_629),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_646),
.B(n_629),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_651),
.B(n_600),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_649),
.B(n_638),
.Y(n_699)
);

AOI22xp33_ASAP7_75t_L g700 ( 
.A1(n_666),
.A2(n_600),
.B1(n_605),
.B2(n_636),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_680),
.B(n_608),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_648),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_650),
.B(n_637),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_645),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_645),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_649),
.B(n_608),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_672),
.B(n_608),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_668),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_652),
.B(n_619),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_668),
.B(n_679),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_660),
.B(n_597),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_675),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_710),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_681),
.B(n_660),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_681),
.B(n_665),
.Y(n_715)
);

NOR3xp33_ASAP7_75t_L g716 ( 
.A(n_686),
.B(n_667),
.C(n_668),
.Y(n_716)
);

INVx3_ASAP7_75t_L g717 ( 
.A(n_710),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_682),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_692),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_692),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_702),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_689),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_687),
.B(n_654),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_684),
.B(n_679),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_684),
.B(n_679),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_702),
.Y(n_726)
);

AND2x4_ASAP7_75t_L g727 ( 
.A(n_687),
.B(n_654),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_706),
.B(n_665),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_704),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_682),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_704),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_688),
.B(n_670),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_716),
.A2(n_700),
.B1(n_622),
.B2(n_618),
.Y(n_733)
);

NAND2x1_ASAP7_75t_L g734 ( 
.A(n_713),
.B(n_706),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_732),
.B(n_683),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_718),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_729),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_730),
.Y(n_738)
);

OAI22xp5_ASAP7_75t_L g739 ( 
.A1(n_722),
.A2(n_685),
.B1(n_709),
.B2(n_697),
.Y(n_739)
);

INVx1_ASAP7_75t_SL g740 ( 
.A(n_723),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_719),
.Y(n_741)
);

OAI32xp33_ASAP7_75t_L g742 ( 
.A1(n_724),
.A2(n_697),
.A3(n_694),
.B1(n_691),
.B2(n_698),
.Y(n_742)
);

AOI22xp5_ASAP7_75t_L g743 ( 
.A1(n_723),
.A2(n_697),
.B1(n_687),
.B2(n_696),
.Y(n_743)
);

OAI21xp5_ASAP7_75t_L g744 ( 
.A1(n_733),
.A2(n_724),
.B(n_725),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_736),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_734),
.Y(n_746)
);

OAI22xp5_ASAP7_75t_L g747 ( 
.A1(n_733),
.A2(n_713),
.B1(n_717),
.B2(n_715),
.Y(n_747)
);

INVxp67_ASAP7_75t_L g748 ( 
.A(n_739),
.Y(n_748)
);

OAI21xp5_ASAP7_75t_L g749 ( 
.A1(n_742),
.A2(n_725),
.B(n_715),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_738),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_749),
.B(n_748),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_750),
.B(n_735),
.Y(n_752)
);

OAI311xp33_ASAP7_75t_L g753 ( 
.A1(n_744),
.A2(n_743),
.A3(n_707),
.B1(n_701),
.C1(n_711),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_747),
.A2(n_741),
.B1(n_646),
.B2(n_737),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_745),
.A2(n_695),
.B1(n_696),
.B2(n_699),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_746),
.A2(n_695),
.B1(n_699),
.B2(n_740),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_751),
.A2(n_601),
.B(n_606),
.Y(n_757)
);

AOI221xp5_ASAP7_75t_L g758 ( 
.A1(n_753),
.A2(n_726),
.B1(n_721),
.B2(n_720),
.C(n_719),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_752),
.A2(n_754),
.B(n_601),
.Y(n_759)
);

OAI21xp33_ASAP7_75t_SL g760 ( 
.A1(n_756),
.A2(n_714),
.B(n_713),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_755),
.B(n_714),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_757),
.B(n_728),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_761),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_759),
.B(n_728),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_763),
.A2(n_760),
.B1(n_758),
.B2(n_646),
.Y(n_765)
);

O2A1O1Ixp33_ASAP7_75t_L g766 ( 
.A1(n_764),
.A2(n_646),
.B(n_623),
.C(n_717),
.Y(n_766)
);

AOI221xp5_ASAP7_75t_L g767 ( 
.A1(n_762),
.A2(n_693),
.B1(n_712),
.B2(n_726),
.C(n_721),
.Y(n_767)
);

INVxp67_ASAP7_75t_SL g768 ( 
.A(n_766),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_765),
.A2(n_606),
.B1(n_727),
.B2(n_723),
.Y(n_769)
);

NOR4xp25_ASAP7_75t_L g770 ( 
.A(n_767),
.B(n_712),
.C(n_717),
.D(n_720),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_767),
.B(n_727),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_767),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_768),
.B(n_690),
.Y(n_773)
);

AOI221xp5_ASAP7_75t_L g774 ( 
.A1(n_772),
.A2(n_729),
.B1(n_731),
.B2(n_641),
.C(n_690),
.Y(n_774)
);

OA21x2_ASAP7_75t_L g775 ( 
.A1(n_769),
.A2(n_771),
.B(n_770),
.Y(n_775)
);

AOI221xp5_ASAP7_75t_L g776 ( 
.A1(n_768),
.A2(n_731),
.B1(n_641),
.B2(n_708),
.C(n_662),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_768),
.Y(n_777)
);

NAND3x2_ASAP7_75t_L g778 ( 
.A(n_772),
.B(n_727),
.C(n_703),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_777),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_773),
.Y(n_780)
);

BUFx2_ASAP7_75t_L g781 ( 
.A(n_775),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_778),
.Y(n_782)
);

NOR2xp67_ASAP7_75t_L g783 ( 
.A(n_776),
.B(n_774),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_781),
.A2(n_703),
.B1(n_670),
.B2(n_671),
.Y(n_784)
);

XNOR2xp5_ASAP7_75t_L g785 ( 
.A(n_779),
.B(n_596),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_780),
.Y(n_786)
);

AO22x2_ASAP7_75t_L g787 ( 
.A1(n_782),
.A2(n_596),
.B1(n_676),
.B2(n_675),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_782),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_788),
.Y(n_789)
);

AOI31xp33_ASAP7_75t_L g790 ( 
.A1(n_786),
.A2(n_783),
.A3(n_669),
.B(n_674),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_784),
.A2(n_674),
.B1(n_662),
.B2(n_661),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_789),
.A2(n_785),
.B1(n_787),
.B2(n_678),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_791),
.A2(n_661),
.B1(n_669),
.B2(n_671),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_792),
.A2(n_790),
.B1(n_678),
.B2(n_671),
.Y(n_794)
);

OAI21xp5_ASAP7_75t_L g795 ( 
.A1(n_794),
.A2(n_793),
.B(n_676),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_795),
.A2(n_705),
.B1(n_671),
.B2(n_658),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_796),
.B(n_671),
.Y(n_797)
);

AOI211xp5_ASAP7_75t_L g798 ( 
.A1(n_797),
.A2(n_655),
.B(n_658),
.C(n_705),
.Y(n_798)
);


endmodule