module fake_jpeg_10693_n_202 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_202);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_139;
wire n_45;
wire n_61;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_3),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_12),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_41),
.B1(n_18),
.B2(n_28),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_24),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx2_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_4),
.B1(n_8),
.B2(n_9),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_35),
.B1(n_28),
.B2(n_26),
.Y(n_54)
);

NAND2x1_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_31),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_46),
.C(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_47),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_60),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2x1_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_66),
.Y(n_74)
);

BUFx12_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_53),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_26),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_64),
.B(n_28),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_37),
.B(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_38),
.B(n_20),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_62),
.B(n_63),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_36),
.B(n_17),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_29),
.B(n_23),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_36),
.B(n_20),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_19),
.B1(n_25),
.B2(n_21),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_68),
.A2(n_18),
.B(n_35),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_26),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_70),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_41),
.B(n_35),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_77),
.CON(n_102),
.SN(n_102)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_84),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_50),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_80),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_46),
.B1(n_39),
.B2(n_42),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_83),
.B1(n_86),
.B2(n_90),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_43),
.C(n_42),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_54),
.A2(n_39),
.B1(n_43),
.B2(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AO21x2_ASAP7_75t_SL g85 ( 
.A1(n_53),
.A2(n_43),
.B(n_22),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_85),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_30),
.B1(n_27),
.B2(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_89),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_58),
.A2(n_30),
.B1(n_34),
.B2(n_24),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_91),
.B(n_64),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_55),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_21),
.B(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_95),
.B(n_60),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_110),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_52),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_117),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_69),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_114),
.A2(n_85),
.B1(n_88),
.B2(n_53),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_115),
.A2(n_116),
.B(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_17),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_76),
.B(n_91),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_33),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_94),
.B(n_68),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_126),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_105),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_101),
.B(n_94),
.C(n_77),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_135),
.C(n_139),
.Y(n_140)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_133),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_97),
.A2(n_85),
.B1(n_56),
.B2(n_83),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_85),
.B1(n_97),
.B2(n_65),
.Y(n_154)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_115),
.A2(n_88),
.B(n_80),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_85),
.B(n_79),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_138),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_119),
.A2(n_72),
.B(n_80),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_98),
.B(n_106),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_110),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_103),
.C(n_117),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_142),
.C(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_110),
.C(n_112),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_111),
.B(n_113),
.C(n_102),
.D(n_118),
.Y(n_144)
);

OAI322xp33_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_145),
.A3(n_153),
.B1(n_157),
.B2(n_151),
.C1(n_156),
.C2(n_147),
.Y(n_164)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_123),
.A2(n_109),
.B(n_108),
.C(n_107),
.D(n_116),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_149),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_96),
.C(n_114),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_155),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_SL g153 ( 
.A1(n_125),
.A2(n_98),
.A3(n_16),
.B1(n_90),
.B2(n_86),
.C1(n_114),
.C2(n_97),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_154),
.A2(n_133),
.B1(n_120),
.B2(n_131),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_128),
.A2(n_89),
.B1(n_65),
.B2(n_25),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_152),
.B(n_137),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_16),
.C(n_8),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_159),
.A2(n_155),
.B1(n_143),
.B2(n_61),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_142),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_162),
.A2(n_170),
.B(n_32),
.C(n_22),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_154),
.A2(n_138),
.B1(n_136),
.B2(n_126),
.Y(n_163)
);

AOI321xp33_ASAP7_75t_L g182 ( 
.A1(n_164),
.A2(n_9),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_124),
.C(n_135),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_127),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_169),
.C(n_171),
.Y(n_175)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_168),
.B(n_4),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_132),
.Y(n_169)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_149),
.B(n_120),
.CON(n_170),
.SN(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_122),
.C(n_130),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g172 ( 
.A1(n_145),
.A2(n_59),
.A3(n_84),
.B1(n_65),
.B2(n_87),
.C1(n_93),
.C2(n_30),
.Y(n_172)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_172),
.A2(n_59),
.A3(n_61),
.B1(n_57),
.B2(n_32),
.C1(n_22),
.C2(n_24),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_159),
.Y(n_186)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_174),
.A2(n_61),
.A3(n_170),
.B1(n_32),
.B2(n_166),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_57),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_161),
.B(n_32),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_171),
.Y(n_178)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_178),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_166),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_179),
.B(n_180),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_59),
.B(n_32),
.Y(n_181)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_182),
.B(n_169),
.Y(n_184)
);

NAND4xp25_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_190),
.C(n_177),
.D(n_160),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_185),
.A2(n_186),
.B1(n_188),
.B2(n_181),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_165),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_193),
.Y(n_196)
);

A2O1A1Ixp33_ASAP7_75t_SL g192 ( 
.A1(n_186),
.A2(n_177),
.B(n_176),
.C(n_175),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_189),
.B(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

AOI322xp5_ASAP7_75t_L g197 ( 
.A1(n_192),
.A2(n_187),
.A3(n_183),
.B1(n_190),
.B2(n_14),
.C1(n_11),
.C2(n_13),
.Y(n_197)
);

AOI322xp5_ASAP7_75t_L g198 ( 
.A1(n_192),
.A2(n_12),
.A3(n_13),
.B1(n_14),
.B2(n_15),
.C1(n_163),
.C2(n_191),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

AO21x2_ASAP7_75t_L g201 ( 
.A1(n_200),
.A2(n_195),
.B(n_197),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_199),
.Y(n_202)
);


endmodule