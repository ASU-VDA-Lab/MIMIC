module real_jpeg_12628_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_126;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx2_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx4f_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_3),
.A2(n_42),
.B1(n_45),
.B2(n_48),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_42),
.B1(n_59),
.B2(n_65),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_4),
.A2(n_59),
.B1(n_65),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_4),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_5),
.A2(n_26),
.B(n_32),
.C(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_71),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_5),
.B(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_5),
.B(n_27),
.Y(n_139)
);

AOI21xp33_ASAP7_75t_SL g154 ( 
.A1(n_5),
.A2(n_27),
.B(n_139),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_5),
.B(n_59),
.C(n_76),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_5),
.A2(n_45),
.B1(n_48),
.B2(n_71),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_5),
.A2(n_58),
.B1(n_61),
.B2(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_5),
.B(n_54),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_9),
.A2(n_37),
.B1(n_45),
.B2(n_48),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_9),
.A2(n_37),
.B1(n_59),
.B2(n_65),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_10),
.A2(n_59),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_10),
.A2(n_45),
.B1(n_48),
.B2(n_64),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_11),
.A2(n_45),
.B1(n_48),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_11),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_11),
.A2(n_59),
.B1(n_65),
.B2(n_82),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_13),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_13),
.A2(n_39),
.B1(n_45),
.B2(n_48),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_13),
.A2(n_39),
.B1(n_59),
.B2(n_65),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_14),
.A2(n_45),
.B1(n_48),
.B2(n_53),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_14),
.A2(n_53),
.B1(n_59),
.B2(n_65),
.Y(n_143)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_122),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_120),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_106),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_38),
.Y(n_23)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_31),
.Y(n_24)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_26),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_26),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_27),
.A2(n_28),
.B1(n_46),
.B2(n_47),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_30),
.B(n_71),
.Y(n_70)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND3xp33_ASAP7_75t_SL g140 ( 
.A(n_28),
.B(n_46),
.C(n_48),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_36),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_43),
.B(n_50),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_41),
.A2(n_43),
.B1(n_44),
.B2(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_43),
.A2(n_44),
.B1(n_100),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_43),
.A2(n_44),
.B1(n_119),
.B2(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_45),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_48),
.B1(n_76),
.B2(n_77),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g137 ( 
.A1(n_45),
.A2(n_47),
.B(n_138),
.C(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_45),
.B(n_163),
.Y(n_162)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_54),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_68),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_56),
.A2(n_68),
.B1(n_69),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_57),
.A2(n_88),
.B(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_57),
.A2(n_62),
.B1(n_168),
.B2(n_170),
.Y(n_167)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_58),
.B(n_89),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_58),
.A2(n_61),
.B1(n_169),
.B2(n_177),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_58),
.A2(n_171),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.Y(n_58)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_59),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_65),
.B1(n_76),
.B2(n_77),
.Y(n_75)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_61),
.B(n_71),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_62),
.A2(n_63),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_62),
.B(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_65),
.B(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_71),
.B(n_75),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_90),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_85),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_79),
.B(n_80),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_SL g76 ( 
.A(n_77),
.Y(n_76)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_83),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_83),
.A2(n_97),
.B1(n_133),
.B2(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_83),
.A2(n_97),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_83),
.A2(n_97),
.B1(n_156),
.B2(n_166),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_98),
.C(n_101),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_91),
.A2(n_92),
.B1(n_98),
.B2(n_99),
.Y(n_108)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_93),
.A2(n_94),
.B(n_96),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_93),
.A2(n_132),
.B(n_134),
.Y(n_131)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_95),
.B(n_97),
.Y(n_134)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_101),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_109),
.C(n_112),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_126),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_116),
.C(n_118),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_130)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_130),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_201),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_144),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_128),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_131),
.C(n_135),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_131),
.A2(n_135),
.B1(n_136),
.B2(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_141),
.B1(n_142),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_157),
.B(n_200),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_149),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_152),
.C(n_155),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_152),
.A2(n_153),
.B1(n_155),
.B2(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_194),
.B(n_199),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_183),
.B(n_193),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_172),
.B(n_182),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_167),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_167),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_164),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_178),
.B(n_181),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_184),
.B(n_185),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_186),
.B(n_189),
.C(n_192),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_198),
.Y(n_199)
);


endmodule