module fake_jpeg_13224_n_448 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_448);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_448;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_8),
.Y(n_32)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_4),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_58),
.B(n_61),
.Y(n_132)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_17),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_62),
.B(n_99),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_25),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_63),
.B(n_64),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_65),
.B(n_75),
.Y(n_160)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_69),
.Y(n_139)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_70),
.Y(n_173)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_73),
.Y(n_123)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_79),
.B(n_83),
.Y(n_164)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_81),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_82),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_33),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_38),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_84),
.B(n_87),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_85),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_86),
.Y(n_187)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_88),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_90),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_91),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_17),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_94),
.B(n_108),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_95),
.Y(n_161)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_26),
.Y(n_96)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_97),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_29),
.B(n_15),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_26),
.Y(n_100)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_100),
.Y(n_176)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_SL g181 ( 
.A(n_101),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_38),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_102),
.B(n_107),
.Y(n_184)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_103),
.Y(n_177)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_105),
.Y(n_155)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_106),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_29),
.B(n_15),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_109),
.B(n_110),
.Y(n_179)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_38),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_111),
.A2(n_113),
.B(n_116),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_47),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_112),
.B(n_0),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g113 ( 
.A(n_52),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_114),
.A2(n_32),
.B1(n_46),
.B2(n_51),
.Y(n_118)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g185 ( 
.A1(n_115),
.A2(n_105),
.B1(n_101),
.B2(n_97),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_52),
.B(n_12),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_57),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_66),
.A2(n_32),
.B1(n_43),
.B2(n_36),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_120),
.A2(n_125),
.B1(n_134),
.B2(n_141),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_43),
.B1(n_36),
.B2(n_54),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_121),
.A2(n_131),
.B1(n_159),
.B2(n_185),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_81),
.A2(n_18),
.B1(n_46),
.B2(n_57),
.Y(n_125)
);

INVxp33_ASAP7_75t_L g229 ( 
.A(n_127),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_108),
.A2(n_18),
.B1(n_54),
.B2(n_49),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_129),
.A2(n_144),
.B1(n_165),
.B2(n_182),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_56),
.B1(n_49),
.B2(n_42),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_59),
.A2(n_53),
.B1(n_56),
.B2(n_42),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_74),
.B(n_53),
.C(n_35),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_136),
.B(n_169),
.C(n_32),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_110),
.A2(n_35),
.B1(n_30),
.B2(n_27),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_143),
.B(n_157),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_112),
.A2(n_30),
.B1(n_27),
.B2(n_12),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_76),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_168),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_93),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_82),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_73),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_156),
.A2(n_114),
.B1(n_117),
.B2(n_157),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_77),
.B(n_6),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_157),
.B(n_183),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_78),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_85),
.A2(n_11),
.B1(n_95),
.B2(n_91),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_82),
.A2(n_11),
.B1(n_86),
.B2(n_70),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_100),
.B(n_115),
.C(n_106),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_86),
.A2(n_109),
.B1(n_71),
.B2(n_69),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_171),
.A2(n_188),
.B1(n_32),
.B2(n_82),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_89),
.A2(n_113),
.B1(n_88),
.B2(n_90),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_67),
.B(n_92),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_180),
.B1(n_173),
.B2(n_181),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_98),
.A2(n_32),
.B1(n_33),
.B2(n_23),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_172),
.B(n_133),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_189),
.B(n_191),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_184),
.B(n_117),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_192),
.A2(n_215),
.B1(n_221),
.B2(n_227),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_128),
.B(n_136),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_193),
.B(n_196),
.Y(n_253)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_127),
.A2(n_169),
.B(n_183),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_195),
.A2(n_223),
.B(n_244),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_166),
.B(n_164),
.Y(n_196)
);

FAx1_ASAP7_75t_SL g197 ( 
.A(n_143),
.B(n_179),
.CI(n_160),
.CON(n_197),
.SN(n_197)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_197),
.B(n_199),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_132),
.B(n_146),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_200),
.B(n_209),
.Y(n_269)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_158),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_201),
.Y(n_281)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_202),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_163),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_203),
.Y(n_251)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_205),
.A2(n_222),
.B(n_223),
.Y(n_286)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_156),
.A2(n_161),
.B1(n_177),
.B2(n_137),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_206),
.A2(n_213),
.B(n_219),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_129),
.A2(n_161),
.B1(n_122),
.B2(n_177),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g272 ( 
.A1(n_207),
.A2(n_211),
.B1(n_212),
.B2(n_222),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_126),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_137),
.B(n_148),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_122),
.A2(n_119),
.B1(n_123),
.B2(n_124),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_119),
.A2(n_123),
.B1(n_124),
.B2(n_154),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_130),
.A2(n_154),
.B1(n_170),
.B2(n_167),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_130),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_170),
.A2(n_167),
.B1(n_151),
.B2(n_176),
.Y(n_215)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_147),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_238),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_176),
.A2(n_138),
.B1(n_135),
.B2(n_142),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_142),
.A2(n_135),
.B1(n_152),
.B2(n_174),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_180),
.A2(n_187),
.B(n_152),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_138),
.A2(n_173),
.B1(n_174),
.B2(n_140),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_224),
.A2(n_225),
.B1(n_240),
.B2(n_228),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_140),
.A2(n_162),
.B1(n_139),
.B2(n_187),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_162),
.A2(n_133),
.B1(n_157),
.B2(n_121),
.Y(n_227)
);

INVx3_ASAP7_75t_SL g228 ( 
.A(n_139),
.Y(n_228)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_228),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_126),
.B(n_113),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_232),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_146),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_233),
.B(n_239),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_126),
.Y(n_234)
);

BUFx5_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_241),
.Y(n_268)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_181),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_184),
.B(n_166),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_157),
.B(n_143),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_157),
.A2(n_143),
.B1(n_133),
.B2(n_156),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_151),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_172),
.B(n_133),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_242),
.B(n_243),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_119),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_127),
.A2(n_128),
.B(n_134),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_166),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_217),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_166),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_247),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_184),
.B(n_166),
.Y(n_247)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_226),
.Y(n_261)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_195),
.A2(n_220),
.B1(n_193),
.B2(n_244),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_250),
.A2(n_255),
.B1(n_275),
.B2(n_282),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_200),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_252),
.B(n_260),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_229),
.A2(n_220),
.B1(n_190),
.B2(n_197),
.Y(n_255)
);

OR2x4_ASAP7_75t_L g257 ( 
.A(n_229),
.B(n_197),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_257),
.A2(n_233),
.B(n_231),
.Y(n_291)
);

AND2x6_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_198),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_261),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_196),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_262),
.B(n_264),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_191),
.B(n_230),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_224),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_266),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_209),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_276),
.Y(n_293)
);

INVx13_ASAP7_75t_L g271 ( 
.A(n_228),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_272),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_239),
.B(n_233),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_198),
.A2(n_240),
.B1(n_231),
.B2(n_227),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_210),
.B(n_202),
.Y(n_285)
);

NAND3xp33_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_287),
.C(n_205),
.Y(n_288)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_288),
.B(n_310),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_291),
.A2(n_258),
.B(n_265),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_192),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_296),
.Y(n_323)
);

A2O1A1Ixp33_ASAP7_75t_SL g295 ( 
.A1(n_279),
.A2(n_205),
.B(n_206),
.C(n_219),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_295),
.A2(n_304),
.B(n_286),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_206),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g297 ( 
.A1(n_270),
.A2(n_206),
.B1(n_225),
.B2(n_249),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_315),
.B1(n_284),
.B2(n_261),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_241),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_298),
.B(n_305),
.Y(n_330)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_256),
.Y(n_299)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_299),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_215),
.C(n_201),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_300),
.B(n_302),
.C(n_306),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_213),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_270),
.A2(n_214),
.B1(n_243),
.B2(n_216),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_303),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_279),
.A2(n_208),
.B(n_234),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_284),
.A2(n_204),
.B1(n_194),
.B2(n_237),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_235),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_260),
.B(n_250),
.C(n_282),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_312),
.C(n_317),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_267),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_308),
.B(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_273),
.Y(n_309)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_283),
.B(n_257),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_269),
.B(n_253),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_284),
.A2(n_269),
.B1(n_261),
.B2(n_266),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_277),
.Y(n_316)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_316),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_253),
.B(n_258),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_318),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_278),
.B(n_287),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_280),
.Y(n_321)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_321),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_324),
.B(n_295),
.C(n_321),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_308),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_293),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_278),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_339),
.C(n_344),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_331),
.A2(n_313),
.B(n_263),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_314),
.B(n_291),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_333),
.A2(n_346),
.B(n_280),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_317),
.B(n_283),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_334),
.B(n_341),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_315),
.Y(n_354)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_306),
.B(n_275),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_290),
.B(n_251),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_342),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_289),
.B(n_251),
.C(n_265),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_319),
.B(n_254),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_345),
.B(n_347),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_311),
.A2(n_314),
.B(n_313),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_312),
.B(n_259),
.Y(n_347)
);

BUFx4f_ASAP7_75t_SL g349 ( 
.A(n_322),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_364),
.Y(n_384)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

AOI321xp33_ASAP7_75t_L g353 ( 
.A1(n_347),
.A2(n_293),
.A3(n_310),
.B1(n_298),
.B2(n_294),
.C(n_296),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_353),
.A2(n_368),
.B(n_343),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_354),
.A2(n_360),
.B1(n_365),
.B2(n_333),
.Y(n_371)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_329),
.Y(n_355)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_355),
.Y(n_385)
);

OAI21xp33_ASAP7_75t_L g356 ( 
.A1(n_325),
.A2(n_304),
.B(n_320),
.Y(n_356)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_356),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_336),
.B(n_302),
.Y(n_357)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_358),
.A2(n_343),
.B(n_335),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_323),
.A2(n_301),
.B1(n_295),
.B2(n_297),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_361),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_326),
.A2(n_301),
.B1(n_305),
.B2(n_295),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_345),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_329),
.Y(n_362)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_362),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_331),
.A2(n_263),
.B(n_300),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_363),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_323),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_281),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_338),
.C(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_342),
.Y(n_367)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_367),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_334),
.B(n_292),
.Y(n_370)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_370),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_371),
.A2(n_359),
.B1(n_330),
.B2(n_363),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_340),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_379),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_338),
.C(n_328),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_381),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_339),
.C(n_346),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_386),
.B(n_388),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_339),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_358),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_374),
.A2(n_361),
.B1(n_341),
.B2(n_344),
.Y(n_391)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_378),
.A2(n_354),
.B1(n_364),
.B2(n_352),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_392),
.A2(n_395),
.B1(n_372),
.B2(n_387),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_378),
.A2(n_368),
.B1(n_330),
.B2(n_326),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_384),
.Y(n_396)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_396),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_388),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_389),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_398),
.B(n_324),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_399),
.A2(n_400),
.B1(n_404),
.B2(n_386),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_382),
.A2(n_348),
.B1(n_353),
.B2(n_369),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_382),
.A2(n_348),
.B1(n_369),
.B2(n_355),
.Y(n_401)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_401),
.Y(n_415)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_376),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_375),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_372),
.A2(n_367),
.B1(n_350),
.B2(n_362),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_405),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_408),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_375),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_404),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_395),
.A2(n_373),
.B1(n_383),
.B2(n_376),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_393),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_379),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_412),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_411),
.A2(n_381),
.B(n_397),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_380),
.C(n_377),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_416),
.A2(n_400),
.B(n_399),
.Y(n_422)
);

OAI221xp5_ASAP7_75t_L g417 ( 
.A1(n_414),
.A2(n_393),
.B1(n_396),
.B2(n_373),
.C(n_390),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_417),
.A2(n_415),
.B1(n_413),
.B2(n_405),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_411),
.Y(n_433)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_420),
.Y(n_432)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_421),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_422),
.B(n_406),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_412),
.B(n_394),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_424),
.B(n_410),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_426),
.Y(n_439)
);

AO21x1_ASAP7_75t_L g427 ( 
.A1(n_419),
.A2(n_407),
.B(n_409),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_427),
.A2(n_428),
.B(n_430),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_425),
.B(n_408),
.Y(n_430)
);

NOR2xp67_ASAP7_75t_SL g438 ( 
.A(n_431),
.B(n_433),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_432),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_434),
.B(n_435),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_432),
.B(n_425),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_433),
.A2(n_423),
.B(n_419),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_437),
.A2(n_390),
.B(n_418),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_439),
.A2(n_427),
.B1(n_385),
.B2(n_350),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_441),
.A2(n_337),
.B1(n_332),
.B2(n_327),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_438),
.B(n_402),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_442),
.A2(n_443),
.B(n_436),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_444),
.A2(n_445),
.B(n_440),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_446),
.A2(n_322),
.B(n_403),
.Y(n_447)
);

BUFx24_ASAP7_75t_SL g448 ( 
.A(n_447),
.Y(n_448)
);


endmodule