module fake_jpeg_21947_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_3),
.Y(n_7)
);

INVx6_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_4),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_L g11 ( 
.A1(n_2),
.A2(n_5),
.B1(n_3),
.B2(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_14),
.Y(n_15)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_12),
.B(n_5),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_14),
.B(n_13),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_8),
.A2(n_12),
.B1(n_7),
.B2(n_13),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_20),
.B(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_26),
.B(n_18),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_22),
.A2(n_17),
.B1(n_16),
.B2(n_8),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_22),
.B1(n_23),
.B2(n_8),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_29),
.B1(n_11),
.B2(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_35),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_24),
.C(n_15),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_31),
.B(n_15),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_39),
.C(n_35),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_6),
.B(n_1),
.Y(n_39)
);

AO221x1_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.C(n_3),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B(n_6),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_42),
.A2(n_6),
.B(n_1),
.Y(n_43)
);


endmodule