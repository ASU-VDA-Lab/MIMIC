module fake_jpeg_23728_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx5p33_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_40),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_20),
.B(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_44),
.B(n_25),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_58),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_41),
.A2(n_18),
.B1(n_22),
.B2(n_25),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_31),
.B1(n_20),
.B2(n_22),
.Y(n_70)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_61),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_64),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_69),
.Y(n_84)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_24),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_45),
.B(n_27),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_70),
.A2(n_80),
.B1(n_20),
.B2(n_21),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_31),
.B1(n_19),
.B2(n_29),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_96),
.B1(n_49),
.B2(n_47),
.Y(n_99)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_51),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_88),
.Y(n_123)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_77),
.B(n_66),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_53),
.A2(n_31),
.B1(n_29),
.B2(n_40),
.Y(n_80)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_91),
.Y(n_106)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_89),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_28),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_94),
.Y(n_107)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_95),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_68),
.B1(n_29),
.B2(n_47),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_74),
.A2(n_77),
.B(n_80),
.C(n_70),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_109),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_66),
.B(n_45),
.C(n_29),
.Y(n_98)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx11_ASAP7_75t_L g136 ( 
.A(n_101),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_30),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_84),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_81),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_79),
.A2(n_30),
.B1(n_21),
.B2(n_29),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_43),
.A3(n_30),
.B1(n_21),
.B2(n_32),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_17),
.Y(n_131)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_115),
.Y(n_146)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_116),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_89),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_122),
.B1(n_92),
.B2(n_82),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g119 ( 
.A(n_79),
.B(n_65),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_121),
.C(n_81),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_62),
.C(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_125),
.B(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_106),
.B(n_23),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_129),
.B(n_76),
.C(n_100),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_121),
.A2(n_82),
.B(n_55),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_133),
.B(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_132),
.Y(n_156)
);

AOI22x1_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_118),
.B1(n_104),
.B2(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_76),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_138),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_145),
.B1(n_101),
.B2(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_27),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_139),
.B(n_142),
.Y(n_159)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_98),
.B(n_52),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_85),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_148),
.Y(n_161)
);

AOI22x1_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_17),
.B1(n_32),
.B2(n_52),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_58),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_111),
.A2(n_52),
.B(n_36),
.C(n_37),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_120),
.Y(n_150)
);

OAI22x1_ASAP7_75t_L g151 ( 
.A1(n_134),
.A2(n_141),
.B1(n_145),
.B2(n_149),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_151),
.A2(n_144),
.B1(n_17),
.B2(n_32),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_134),
.A2(n_126),
.B1(n_131),
.B2(n_142),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_154),
.A2(n_164),
.B1(n_174),
.B2(n_173),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_155),
.A2(n_158),
.B1(n_169),
.B2(n_170),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_136),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_104),
.B1(n_110),
.B2(n_100),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_103),
.Y(n_162)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_162),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_95),
.B1(n_115),
.B2(n_75),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_146),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_171),
.B(n_172),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_130),
.A2(n_114),
.B1(n_60),
.B2(n_55),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_133),
.A2(n_56),
.B(n_61),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_0),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_124),
.A2(n_88),
.B1(n_86),
.B2(n_114),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_175),
.B(n_176),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_125),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_174),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_177),
.B(n_192),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_163),
.A2(n_139),
.B(n_124),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_178),
.A2(n_182),
.B(n_184),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_161),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_183),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_140),
.B(n_132),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_140),
.B(n_127),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_147),
.A3(n_150),
.B1(n_148),
.B2(n_138),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_186),
.Y(n_222)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_128),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_196),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_160),
.Y(n_189)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_152),
.B(n_23),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_191),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_152),
.B(n_33),
.Y(n_192)
);

OAI21xp33_ASAP7_75t_SL g225 ( 
.A1(n_193),
.A2(n_194),
.B(n_199),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_167),
.B(n_38),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_201),
.Y(n_208)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_144),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_164),
.A2(n_107),
.B1(n_116),
.B2(n_33),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_199),
.A2(n_32),
.B1(n_17),
.B2(n_26),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_166),
.Y(n_200)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_163),
.A2(n_33),
.B(n_28),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_202),
.B(n_0),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_198),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_213),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_203),
.A2(n_173),
.B1(n_151),
.B2(n_168),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_206),
.B1(n_207),
.B2(n_215),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_169),
.B1(n_170),
.B2(n_165),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_203),
.A2(n_159),
.B1(n_175),
.B2(n_167),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_159),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_219),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_172),
.C(n_52),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_212),
.C(n_221),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_39),
.C(n_107),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_217),
.A2(n_225),
.B(n_177),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_39),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_28),
.C(n_26),
.Y(n_221)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_227),
.Y(n_230)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_28),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_228),
.B(n_180),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_190),
.C(n_189),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_234),
.C(n_242),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_190),
.C(n_182),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_181),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_235),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_218),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_243),
.B(n_244),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_200),
.Y(n_239)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_240),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_179),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_184),
.C(n_178),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_218),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_224),
.B(n_179),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_246),
.B(n_247),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_188),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g271 ( 
.A(n_248),
.B(n_235),
.CI(n_241),
.CON(n_271),
.SN(n_271)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_229),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_249),
.A2(n_250),
.B1(n_209),
.B2(n_215),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_188),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_207),
.A2(n_205),
.B1(n_222),
.B2(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_216),
.B1(n_222),
.B2(n_220),
.Y(n_252)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_252),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_251),
.B(n_208),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_259),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_230),
.C(n_234),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_257),
.C(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_220),
.C(n_223),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_219),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_214),
.C(n_221),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_250),
.Y(n_263)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_263),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_201),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_232),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_236),
.B(n_232),
.C(n_238),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_270),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_194),
.B1(n_187),
.B2(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_268),
.Y(n_287)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_245),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_254),
.B(n_244),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_15),
.C(n_14),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_276),
.B(n_0),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_282),
.B(n_286),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_248),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_279),
.B(n_28),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_257),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_258),
.B1(n_262),
.B2(n_255),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_283),
.A2(n_284),
.B1(n_15),
.B2(n_14),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_271),
.B1(n_261),
.B2(n_243),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_237),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_288),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_269),
.B(n_267),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_194),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_253),
.B(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

FAx1_ASAP7_75t_L g290 ( 
.A(n_288),
.B(n_265),
.CI(n_253),
.CON(n_290),
.SN(n_290)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_290),
.A2(n_302),
.B1(n_11),
.B2(n_3),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_192),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_299),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_191),
.Y(n_294)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_294),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_276),
.B(n_26),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_300),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_301),
.C(n_12),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_14),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_13),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_272),
.B(n_287),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_277),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_280),
.C(n_2),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_281),
.B1(n_279),
.B2(n_275),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_305),
.A2(n_310),
.B1(n_314),
.B2(n_5),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_313),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_280),
.B1(n_12),
.B2(n_11),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_292),
.C(n_290),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_311),
.A2(n_2),
.B(n_3),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_5),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_293),
.B(n_1),
.Y(n_313)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_316),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_315),
.B(n_2),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_318),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_4),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_4),
.B(n_5),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_319),
.B(n_321),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_4),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_324),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_4),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_307),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_323),
.B(n_311),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_327),
.A2(n_328),
.B(n_320),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_304),
.B(n_307),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_5),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_333),
.C(n_334),
.Y(n_335)
);

AOI211x1_ASAP7_75t_L g333 ( 
.A1(n_325),
.A2(n_329),
.B(n_326),
.C(n_331),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_330),
.B(n_7),
.C(n_8),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_6),
.C(n_7),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

O2A1O1Ixp33_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_6),
.B(n_7),
.C(n_9),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_10),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_SL g341 ( 
.A1(n_340),
.A2(n_10),
.B(n_322),
.C(n_338),
.Y(n_341)
);


endmodule