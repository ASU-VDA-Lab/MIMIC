module real_jpeg_5276_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_0),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_0),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_0),
.Y(n_152)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_0),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_0),
.Y(n_228)
);

INVx6_ASAP7_75t_L g463 ( 
.A(n_0),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_1),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_1),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_1),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_1),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_1),
.B(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_1),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_1),
.B(n_460),
.Y(n_459)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_3),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_3),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_3),
.B(n_242),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_3),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_3),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_3),
.B(n_240),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_3),
.B(n_384),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_4),
.A2(n_232),
.B(n_234),
.Y(n_231)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_4),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_4),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_4),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_4),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_4),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_4),
.B(n_393),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_5),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_6),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_6),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_6),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_6),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_6),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_6),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_6),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_6),
.B(n_407),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_7),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_7),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_7),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_7),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_7),
.B(n_255),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_7),
.B(n_240),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_7),
.B(n_389),
.Y(n_388)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_9),
.Y(n_147)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_9),
.Y(n_238)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_9),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_10),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_10),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_10),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_10),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_10),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_10),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_10),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_10),
.B(n_462),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_11),
.B(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_11),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_11),
.B(n_106),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_11),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_11),
.B(n_144),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_11),
.B(n_178),
.Y(n_177)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_12),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_12),
.Y(n_233)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_14),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_39),
.Y(n_38)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_14),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_14),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_14),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_14),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_14),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_15),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_15),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_15),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_442),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_198),
.B(n_440),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_165),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_20),
.B(n_165),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_93),
.C(n_123),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_21),
.B(n_93),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_58),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_23),
.B(n_40),
.C(n_58),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.C(n_38),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_24),
.B(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_27),
.C(n_31),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_25),
.B(n_50),
.C(n_54),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_25),
.A2(n_54),
.B1(n_89),
.B2(n_90),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_25),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_25),
.A2(n_31),
.B1(n_89),
.B2(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_25),
.A2(n_89),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_25),
.B(n_367),
.Y(n_409)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_26),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_27),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_27),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_27),
.A2(n_126),
.B1(n_193),
.B2(n_197),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_30),
.Y(n_150)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_30),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_31),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_31),
.B(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_31),
.A2(n_129),
.B1(n_262),
.B2(n_263),
.Y(n_331)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_32),
.Y(n_358)
);

INVx8_ASAP7_75t_L g382 ( 
.A(n_32),
.Y(n_382)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g391 ( 
.A(n_33),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_34),
.A2(n_38),
.B1(n_48),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_34),
.Y(n_164)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_38),
.A2(n_42),
.B1(n_43),
.B2(n_48),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

OA22x2_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_40)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_43),
.B(n_48),
.C(n_57),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_47),
.Y(n_134)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_47),
.Y(n_322)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_50),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_50),
.B(n_221),
.C(n_225),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_50),
.A2(n_91),
.B1(n_221),
.B2(n_292),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_54),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_77),
.C(n_87),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_59),
.B(n_77),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_68),
.C(n_72),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_60),
.A2(n_61),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_60),
.B(n_116),
.C(n_122),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_60),
.A2(n_61),
.B1(n_142),
.B2(n_143),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_61),
.B(n_143),
.Y(n_299)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_62),
.Y(n_137)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_68),
.B1(n_72),
.B2(n_76),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_71),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_71),
.Y(n_348)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_72),
.A2(n_76),
.B1(n_454),
.B2(n_455),
.Y(n_453)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.C(n_85),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_85),
.Y(n_139)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g373 ( 
.A(n_84),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_87),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_113),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_95),
.B(n_96),
.C(n_113),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_110),
.B2(n_111),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_105),
.B1(n_108),
.B2(n_109),
.Y(n_98)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_103),
.Y(n_224)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_104),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_108),
.C(n_111),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_105),
.B(n_132),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_131),
.C(n_135),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_112),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_122),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_119),
.A2(n_122),
.B1(n_177),
.B2(n_180),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_119),
.B(n_254),
.C(n_258),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_119),
.A2(n_122),
.B1(n_258),
.B2(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_122),
.B(n_173),
.C(n_177),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_123),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_140),
.C(n_162),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_124),
.B(n_278),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_138),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_125),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_126),
.B(n_188),
.C(n_193),
.Y(n_452)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_130),
.B(n_138),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_135),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_140),
.B(n_162),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_153),
.C(n_157),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_141),
.B(n_244),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.C(n_151),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_142),
.A2(n_143),
.B1(n_151),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_147),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_147),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_148),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_148),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_148),
.A2(n_172),
.B1(n_173),
.B2(n_267),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_151),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_153),
.A2(n_157),
.B1(n_158),
.B2(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_153),
.Y(n_245)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_156),
.Y(n_325)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_161),
.Y(n_191)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_161),
.Y(n_242)
);

BUFx24_ASAP7_75t_SL g468 ( 
.A(n_165),
.Y(n_468)
);

FAx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_167),
.CI(n_181),
.CON(n_165),
.SN(n_165)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_166),
.B(n_167),
.C(n_181),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_209),
.C(n_214),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_172),
.A2(n_173),
.B1(n_209),
.B2(n_210),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_177),
.Y(n_180)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_182),
.B(n_184),
.C(n_187),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_192),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_190),
.Y(n_460)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_193),
.Y(n_197)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI221xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_337),
.B1(n_433),
.B2(n_438),
.C(n_439),
.Y(n_199)
);

NOR3xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_280),
.C(n_284),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_201),
.A2(n_434),
.B(n_437),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_273),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_202),
.B(n_273),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_246),
.C(n_249),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_203),
.B(n_246),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_229),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_204),
.B(n_230),
.C(n_243),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.C(n_219),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_206),
.B(n_220),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_208),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_214),
.B(n_252),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_218),
.Y(n_366)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_225),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_243),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_239),
.C(n_241),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_231),
.B(n_272),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_231),
.A2(n_234),
.B(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx5_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_241),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_266),
.C(n_271),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_288),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.C(n_260),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_251),
.B(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_253),
.A2(n_260),
.B1(n_261),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_253),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_254),
.B(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

INVx6_ASAP7_75t_L g329 ( 
.A(n_259),
.Y(n_329)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_266),
.B(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_279),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_281)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_280),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_281),
.B(n_282),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_310),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_285),
.A2(n_435),
.B(n_436),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_308),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_286),
.B(n_308),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_289),
.C(n_306),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_306),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.C(n_297),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_293),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_295),
.B(n_371),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_297),
.B(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.C(n_303),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_298),
.A2(n_299),
.B1(n_421),
.B2(n_422),
.Y(n_420)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_300),
.A2(n_301),
.B1(n_303),
.B2(n_304),
.Y(n_421)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_335),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_311),
.B(n_335),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_314),
.C(n_332),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_312),
.B(n_431),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_314),
.B(n_332),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.C(n_330),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g423 ( 
.A(n_315),
.B(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_318),
.A2(n_330),
.B1(n_331),
.B2(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_318),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_323),
.C(n_326),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_319),
.A2(n_320),
.B1(n_326),
.B2(n_327),
.Y(n_413)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_323),
.B(n_413),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_428),
.B(n_432),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_415),
.B(n_427),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_402),
.B(n_414),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_376),
.B(n_401),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_368),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_342),
.B(n_368),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_354),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_343),
.B(n_355),
.C(n_364),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_349),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_344),
.B(n_350),
.C(n_351),
.Y(n_411)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_364),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_359),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_356),
.B(n_359),
.Y(n_369)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_365),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_370),
.C(n_374),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_369),
.B(n_398),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_370),
.A2(n_374),
.B1(n_375),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_395),
.B(n_400),
.Y(n_376)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_378),
.A2(n_387),
.B(n_394),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_379),
.B(n_386),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_386),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_383),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_383),
.Y(n_396)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_SL g384 ( 
.A(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_392),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_396),
.B(n_397),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_404),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_410),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_405),
.A2(n_418),
.B1(n_419),
.B2(n_420),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_405),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_405),
.B(n_411),
.C(n_412),
.Y(n_426)
);

FAx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.B(n_408),
.CI(n_409),
.CON(n_405),
.SN(n_405)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_416),
.B(n_426),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_416),
.B(n_426),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_423),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_418),
.B(n_420),
.C(n_423),
.Y(n_429)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_421),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_430),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_429),
.B(n_430),
.Y(n_432)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_466),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_445),
.B(n_446),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_456),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_459),
.A2(n_461),
.B1(n_464),
.B2(n_465),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_459),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_461),
.Y(n_465)
);

INVx8_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);


endmodule