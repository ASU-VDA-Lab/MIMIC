module fake_jpeg_15272_n_368 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_368);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_368;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx3_ASAP7_75t_SL g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx11_ASAP7_75t_SL g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_60),
.Y(n_72)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_21),
.B(n_10),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_57),
.B(n_58),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_11),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_28),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_11),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_42),
.B1(n_24),
.B2(n_44),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_70),
.A2(n_93),
.B1(n_35),
.B2(n_37),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_42),
.B1(n_41),
.B2(n_30),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_30),
.B1(n_53),
.B2(n_28),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_85),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_25),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_80),
.B(n_81),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_60),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_42),
.B1(n_44),
.B2(n_29),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_105)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx2_ASAP7_75t_SL g100 ( 
.A(n_91),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_61),
.A2(n_28),
.B1(n_29),
.B2(n_44),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_22),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_46),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_99),
.A2(n_118),
.B1(n_123),
.B2(n_127),
.Y(n_153)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

BUFx4f_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_104),
.B(n_32),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_105),
.A2(n_130),
.B1(n_30),
.B2(n_31),
.Y(n_134)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_109),
.Y(n_131)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_46),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_114),
.B(n_31),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_69),
.B(n_43),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_117),
.Y(n_145)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_76),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_122),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_88),
.A2(n_30),
.B1(n_62),
.B2(n_63),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_124),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_98),
.B(n_30),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_65),
.C(n_52),
.Y(n_156)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_126),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_88),
.A2(n_30),
.B1(n_55),
.B2(n_51),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

BUFx10_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_75),
.A2(n_38),
.B1(n_22),
.B2(n_43),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_134),
.A2(n_128),
.B1(n_101),
.B2(n_103),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_102),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_120),
.A2(n_75),
.B1(n_86),
.B2(n_38),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_136),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_120),
.A2(n_86),
.B1(n_39),
.B2(n_89),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_141),
.B(n_143),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_39),
.B1(n_92),
.B2(n_89),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_144),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_91),
.B1(n_82),
.B2(n_35),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_0),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_104),
.A2(n_92),
.B1(n_82),
.B2(n_45),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_37),
.A3(n_45),
.B1(n_48),
.B2(n_40),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_147),
.B(n_99),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_97),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_148),
.B(n_157),
.Y(n_179)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_36),
.CON(n_149),
.SN(n_149)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_149),
.A2(n_151),
.B(n_0),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_94),
.C(n_129),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_71),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_100),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_110),
.A2(n_85),
.B1(n_32),
.B2(n_36),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_109),
.B(n_117),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_164),
.Y(n_196)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_140),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_163),
.Y(n_198)
);

INVxp33_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_185),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_143),
.A2(n_127),
.B1(n_111),
.B2(n_112),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_168),
.A2(n_178),
.B1(n_139),
.B2(n_144),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_119),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_169),
.B(n_182),
.Y(n_192)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_170),
.Y(n_193)
);

O2A1O1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_143),
.A2(n_116),
.B(n_107),
.C(n_122),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_171),
.A2(n_177),
.B(n_174),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_SL g197 ( 
.A(n_174),
.B(n_175),
.C(n_176),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g175 ( 
.A(n_143),
.B(n_124),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_137),
.A2(n_103),
.B(n_119),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_16),
.B1(n_20),
.B2(n_19),
.Y(n_178)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_180),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_181),
.B(n_146),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_160),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_157),
.B(n_32),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_173),
.A2(n_153),
.B1(n_156),
.B2(n_147),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_200),
.B1(n_172),
.B2(n_168),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_188),
.A2(n_171),
.B1(n_185),
.B2(n_175),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_170),
.Y(n_190)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_204),
.B(n_207),
.Y(n_219)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_177),
.Y(n_195)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_195),
.Y(n_224)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_177),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_173),
.A2(n_152),
.B1(n_145),
.B2(n_146),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_150),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_203),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_172),
.A2(n_150),
.B(n_145),
.Y(n_204)
);

AND2x4_ASAP7_75t_L g205 ( 
.A(n_171),
.B(n_161),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_205),
.A2(n_142),
.B(n_131),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_152),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_233),
.B1(n_197),
.B2(n_208),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_214),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_195),
.A2(n_183),
.B1(n_173),
.B2(n_164),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_211),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_169),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_222),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_190),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_199),
.A2(n_182),
.B1(n_178),
.B2(n_166),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_205),
.A2(n_186),
.B1(n_194),
.B2(n_203),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_205),
.A2(n_162),
.B1(n_181),
.B2(n_161),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_220),
.B1(n_223),
.B2(n_227),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_161),
.B1(n_140),
.B2(n_133),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_192),
.B(n_74),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_155),
.B1(n_132),
.B2(n_133),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_206),
.B(n_131),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_225),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_191),
.A2(n_155),
.B1(n_154),
.B2(n_159),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_194),
.B(n_131),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_231),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_236),
.B(n_193),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_204),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_186),
.B(n_159),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_155),
.B1(n_159),
.B2(n_142),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_196),
.B(n_32),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_234),
.B(n_36),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_202),
.B(n_32),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_244),
.B1(n_248),
.B2(n_215),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_224),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_249),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_197),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_256),
.B(n_260),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_242),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_189),
.B(n_207),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_209),
.A2(n_189),
.B1(n_188),
.B2(n_193),
.Y(n_244)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_94),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_250),
.C(n_257),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_210),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_198),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_198),
.Y(n_250)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_214),
.Y(n_251)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_251),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_129),
.Y(n_254)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_254),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_1),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_129),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_246),
.C(n_247),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_231),
.A2(n_13),
.B(n_20),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_221),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_221),
.Y(n_266)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_264),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_250),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_237),
.A2(n_229),
.B1(n_224),
.B2(n_211),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_271),
.A2(n_239),
.B1(n_248),
.B2(n_256),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_261),
.B(n_226),
.Y(n_272)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_226),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_273),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_240),
.A2(n_229),
.B1(n_233),
.B2(n_227),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_282),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_240),
.A2(n_236),
.B1(n_220),
.B2(n_213),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_234),
.B1(n_2),
.B2(n_3),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_246),
.B(n_124),
.C(n_36),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_241),
.C(n_245),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_260),
.B(n_15),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_1),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.Y(n_285)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_292),
.C(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_289),
.B(n_290),
.C(n_294),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_268),
.B(n_258),
.C(n_239),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_271),
.B(n_255),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_291),
.B(n_302),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_257),
.C(n_242),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_256),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_297),
.B(n_300),
.Y(n_314)
);

NOR2xp67_ASAP7_75t_SL g298 ( 
.A(n_263),
.B(n_15),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_269),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_124),
.C(n_36),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_284),
.C(n_275),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_269),
.A2(n_281),
.B1(n_273),
.B2(n_266),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_303),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_33),
.Y(n_303)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_308),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_274),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_279),
.C(n_277),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_285),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_311),
.A2(n_270),
.B1(n_296),
.B2(n_286),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_276),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_318),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_279),
.C(n_281),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_313),
.B(n_316),
.Y(n_331)
);

AND2x2_ASAP7_75t_SL g315 ( 
.A(n_295),
.B(n_275),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_317),
.C(n_299),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_267),
.C(n_283),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_267),
.C(n_270),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_321),
.A2(n_322),
.B1(n_5),
.B2(n_12),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_303),
.C(n_301),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_325),
.C(n_327),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_272),
.C(n_278),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_312),
.B(n_300),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_282),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_318),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_33),
.C(n_5),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_5),
.C(n_9),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_319),
.A2(n_13),
.B1(n_6),
.B2(n_7),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_330),
.B(n_16),
.Y(n_342)
);

AOI21x1_ASAP7_75t_L g332 ( 
.A1(n_311),
.A2(n_16),
.B(n_7),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_17),
.B(n_9),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_331),
.A2(n_315),
.B(n_314),
.Y(n_333)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_333),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_334),
.B(n_336),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_324),
.B(n_310),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_343),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_325),
.A2(n_315),
.B1(n_9),
.B2(n_12),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_320),
.B(n_17),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_338),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_340),
.B(n_341),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_342),
.A2(n_18),
.B(n_19),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_327),
.A2(n_18),
.B1(n_19),
.B2(n_33),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_339),
.B(n_326),
.C(n_321),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_349),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_348),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_323),
.C(n_324),
.Y(n_349)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_341),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_352),
.B(n_343),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_347),
.B(n_340),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_353),
.B(n_351),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_350),
.A2(n_335),
.B(n_329),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_358),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_334),
.C(n_328),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_357),
.A2(n_345),
.B(n_354),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_361),
.Y(n_362)
);

NOR3xp33_ASAP7_75t_L g363 ( 
.A(n_362),
.B(n_360),
.C(n_355),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_363),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_364),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_351),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g367 ( 
.A(n_366),
.B(n_345),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_367),
.A2(n_33),
.B(n_361),
.Y(n_368)
);


endmodule