module fake_jpeg_14026_n_198 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_198);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_11),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_33),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_14),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_32),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_18),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_0),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_66),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_86),
.Y(n_92)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_66),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_73),
.B(n_23),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_58),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_57),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_85),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_93),
.B(n_105),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_64),
.B(n_53),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_59),
.B(n_63),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_86),
.B(n_70),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_88),
.A2(n_77),
.B1(n_65),
.B2(n_62),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_106),
.A2(n_67),
.B1(n_69),
.B2(n_78),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_76),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_107),
.B(n_71),
.Y(n_115)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_106),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_110),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_1),
.Y(n_144)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_115),
.B(n_120),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_89),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_81),
.Y(n_136)
);

OR2x4_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_61),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_119),
.B(n_56),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_99),
.A2(n_69),
.B1(n_83),
.B2(n_78),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_119),
.A2(n_127),
.B1(n_58),
.B2(n_56),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_72),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_75),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_123),
.Y(n_135)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_54),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_93),
.A2(n_67),
.B1(n_84),
.B2(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_128),
.Y(n_141)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_109),
.B(n_118),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g170 ( 
.A1(n_134),
.A2(n_146),
.B(n_11),
.C(n_12),
.D(n_15),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_68),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_138),
.B(n_149),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_112),
.B(n_79),
.C(n_60),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_7),
.C(n_8),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_142),
.A2(n_144),
.B1(n_7),
.B2(n_8),
.Y(n_164)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_145),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_1),
.B(n_2),
.C(n_3),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_6),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_2),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_28),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_128),
.B(n_3),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_26),
.B(n_47),
.C(n_46),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g166 ( 
.A(n_151),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_153),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_155),
.A2(n_164),
.B1(n_169),
.B2(n_151),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_156),
.B(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_4),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_167),
.Y(n_180)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_170),
.C(n_16),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_139),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_10),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_134),
.B1(n_147),
.B2(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_175),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_158),
.B(n_135),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_176),
.B(n_178),
.Y(n_183)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_181),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_140),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_166),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_184),
.B(n_173),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_177),
.A2(n_170),
.B1(n_152),
.B2(n_131),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_186),
.B1(n_183),
.B2(n_187),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_152),
.B1(n_131),
.B2(n_154),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

XNOR2x1_ASAP7_75t_SL g192 ( 
.A(n_191),
.B(n_183),
.Y(n_192)
);

OAI221xp5_ASAP7_75t_L g193 ( 
.A1(n_192),
.A2(n_178),
.B1(n_180),
.B2(n_165),
.C(n_30),
.Y(n_193)
);

A2O1A1O1Ixp25_ASAP7_75t_L g194 ( 
.A1(n_193),
.A2(n_20),
.B(n_22),
.C(n_25),
.D(n_31),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_195),
.A2(n_172),
.B(n_39),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_165),
.B1(n_41),
.B2(n_42),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_38),
.Y(n_198)
);


endmodule