module fake_aes_11658_n_29 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_5), .B(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_9), .Y(n_16) );
INVx6_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
BUFx6f_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_15), .B(n_0), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
AO21x2_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_19), .B(n_13), .Y(n_21) );
AND2x2_ASAP7_75t_SL g22 ( .A(n_21), .B(n_16), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
BUFx6f_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
OAI322xp33_ASAP7_75t_L g25 ( .A1(n_23), .A2(n_14), .A3(n_12), .B1(n_0), .B2(n_17), .C1(n_6), .C2(n_11), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_24), .Y(n_26) );
INVxp67_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
NOR2x1p5_ASAP7_75t_L g28 ( .A(n_26), .B(n_25), .Y(n_28) );
AOI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_27), .B1(n_4), .B2(n_10), .Y(n_29) );
endmodule