module real_jpeg_9199_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_2),
.A2(n_58),
.B(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_2),
.B(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_2),
.B(n_92),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_30),
.B1(n_33),
.B2(n_37),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_5),
.B(n_46),
.C(n_110),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g129 ( 
.A1(n_2),
.A2(n_4),
.B(n_30),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_2),
.B(n_40),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_37),
.B1(n_44),
.B2(n_46),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

O2A1O1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_4),
.A2(n_24),
.B(n_28),
.C(n_29),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_4),
.B(n_24),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_4),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_41),
.B(n_46),
.C(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_5),
.B(n_46),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_7),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_7),
.A2(n_11),
.B1(n_45),
.B2(n_58),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_7),
.A2(n_30),
.B1(n_33),
.B2(n_45),
.Y(n_125)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_9),
.A2(n_30),
.B1(n_33),
.B2(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_9),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_10),
.A2(n_44),
.B1(n_46),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_10),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_10),
.A2(n_30),
.B1(n_33),
.B2(n_53),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_53),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_11),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_117),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_116),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_102),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_16),
.B(n_102),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_67),
.B2(n_101),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_55),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_38),
.B2(n_54),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_34),
.B(n_35),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_23),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_23),
.B(n_36),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_23),
.B(n_154),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_24),
.A2(n_37),
.B(n_42),
.Y(n_110)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_25),
.A2(n_32),
.B(n_37),
.C(n_129),
.Y(n_128)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_29),
.B(n_36),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_29),
.B(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_29),
.B(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_30),
.B(n_71),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_33),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_34),
.B(n_37),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_37),
.B(n_71),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_47),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_39),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_43),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_41),
.B(n_52),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_46),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_44),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_61),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_48),
.B(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_49),
.B(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_58),
.A2(n_59),
.B(n_60),
.C(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_60),
.Y(n_64)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_64),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_67),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B1(n_86),
.B2(n_100),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_80),
.B1(n_81),
.B2(n_85),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_73),
.B(n_75),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_79),
.B(n_97),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_72),
.B(n_78),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_72),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_72),
.B(n_96),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_76),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVxp33_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_86),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_91),
.C(n_93),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_91),
.A2(n_93),
.B1(n_94),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_91),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_95),
.B(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_98),
.B(n_125),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_107),
.C(n_112),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_103),
.A2(n_104),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_107),
.A2(n_108),
.B1(n_112),
.B2(n_180),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_109),
.A2(n_111),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_112),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_114),
.B(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_175),
.B(n_181),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_158),
.B(n_174),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_145),
.B(n_157),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_134),
.B(n_144),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_126),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_126),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_130),
.B2(n_131),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_128),
.B(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_139),
.B(n_143),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_147),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_149),
.B(n_152),
.C(n_155),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_160),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_164),
.B1(n_165),
.B2(n_173),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_161),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_168),
.B1(n_169),
.B2(n_172),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_172),
.C(n_173),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_177),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);


endmodule