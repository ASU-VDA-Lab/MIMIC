module real_jpeg_29443_n_18 (n_17, n_8, n_0, n_2, n_10, n_338, n_9, n_12, n_6, n_337, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_338;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_0),
.B(n_50),
.Y(n_89)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_0),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_171),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_1),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_SL g176 ( 
.A1(n_1),
.A2(n_28),
.B(n_32),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_1),
.B(n_30),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_1),
.A2(n_56),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_1),
.B(n_56),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_1),
.B(n_70),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_1),
.A2(n_88),
.B1(n_92),
.B2(n_254),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_1),
.A2(n_31),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_2),
.A2(n_36),
.B1(n_56),
.B2(n_57),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_36),
.B1(n_50),
.B2(n_51),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_4),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_100),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g168 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_100),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_100),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_5),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_131),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_131),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_131),
.Y(n_274)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_45),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_8),
.A2(n_45),
.B1(n_56),
.B2(n_57),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_45),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_8),
.A2(n_45),
.B1(n_50),
.B2(n_51),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_9),
.A2(n_24),
.B1(n_25),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_43),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_9),
.A2(n_43),
.B1(n_56),
.B2(n_57),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_9),
.A2(n_43),
.B1(n_50),
.B2(n_51),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_10),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_173),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_10),
.A2(n_56),
.B1(n_57),
.B2(n_173),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_173),
.Y(n_254)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_11),
.A2(n_51),
.A3(n_56),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_31),
.B1(n_32),
.B2(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_12),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_12),
.A2(n_24),
.B1(n_25),
.B2(n_162),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_162),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_162),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_13),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_13),
.A2(n_56),
.B1(n_57),
.B2(n_98),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_98),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_98),
.Y(n_243)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_15),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_16),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_16),
.A2(n_26),
.B1(n_56),
.B2(n_57),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_16),
.A2(n_26),
.B1(n_50),
.B2(n_51),
.Y(n_123)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_17),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_78),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_37),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_37),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_23),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_28),
.Y(n_29)
);

A2O1A1Ixp33_ASAP7_75t_L g175 ( 
.A1(n_25),
.A2(n_34),
.B(n_171),
.C(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_30),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_27),
.A2(n_30),
.B1(n_97),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_27),
.A2(n_30),
.B1(n_170),
.B2(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_27),
.A2(n_30),
.B1(n_130),
.B2(n_202),
.Y(n_216)
);

AO22x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_30)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_30),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_31),
.A2(n_64),
.B(n_66),
.C(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_64),
.Y(n_66)
);

OAI32xp33_ASAP7_75t_L g278 ( 
.A1(n_31),
.A2(n_57),
.A3(n_64),
.B1(n_271),
.B2(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_32),
.B(n_171),
.Y(n_271)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_71),
.C(n_73),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_38),
.A2(n_39),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.C(n_60),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_40),
.B(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_42),
.A2(n_75),
.B1(n_77),
.B2(n_99),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_44),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_46),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_46),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_46),
.A2(n_60),
.B1(n_140),
.B2(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_54),
.B(n_59),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_47),
.A2(n_54),
.B1(n_59),
.B2(n_109),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_47),
.A2(n_54),
.B1(n_106),
.B2(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_47),
.A2(n_54),
.B1(n_126),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_47),
.A2(n_54),
.B1(n_227),
.B2(n_229),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_47),
.A2(n_54),
.B1(n_229),
.B2(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_47),
.B(n_171),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_47),
.A2(n_54),
.B1(n_167),
.B2(n_296),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_49),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_49),
.B(n_50),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_50),
.B(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_56),
.B(n_280),
.Y(n_279)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_60),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_61),
.A2(n_62),
.B1(n_70),
.B2(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_70),
.B1(n_115),
.B2(n_128),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_62),
.A2(n_70),
.B1(n_161),
.B2(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_62),
.A2(n_70),
.B1(n_128),
.B2(n_205),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_67),
.B(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_63),
.A2(n_67),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_63),
.A2(n_67),
.B1(n_160),
.B2(n_163),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_63),
.A2(n_67),
.B1(n_163),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_63),
.A2(n_67),
.B1(n_185),
.B2(n_269),
.Y(n_268)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_64),
.Y(n_280)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_69),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_71),
.A2(n_73),
.B1(n_74),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_71),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_75),
.A2(n_77),
.B1(n_96),
.B2(n_99),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_75),
.A2(n_77),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_327),
.B(n_333),
.Y(n_80)
);

OAI321xp33_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_143),
.A3(n_152),
.B1(n_325),
.B2(n_326),
.C(n_337),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_132),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_83),
.B(n_132),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_112),
.C(n_119),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_84),
.B(n_112),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_101),
.B1(n_102),
.B2(n_111),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_94),
.B2(n_95),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_86),
.A2(n_95),
.B(n_101),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_86),
.A2(n_87),
.B1(n_103),
.B2(n_104),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_87),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B(n_93),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_93),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_88),
.A2(n_123),
.B1(n_124),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_88),
.A2(n_90),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_88),
.A2(n_90),
.B1(n_248),
.B2(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_88),
.A2(n_124),
.B1(n_243),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_89),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_89),
.A2(n_91),
.B1(n_178),
.B2(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_89),
.A2(n_91),
.B1(n_247),
.B2(n_249),
.Y(n_246)
);

INVx5_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_107),
.B1(n_108),
.B2(n_110),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_107),
.A2(n_110),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_107),
.A2(n_110),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_117),
.B(n_118),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_117),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

FAx1_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_133),
.CI(n_142),
.CON(n_132),
.SN(n_132)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_133),
.C(n_142),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_119),
.A2(n_120),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_127),
.C(n_129),
.Y(n_120)
);

FAx1_ASAP7_75t_SL g308 ( 
.A(n_121),
.B(n_127),
.CI(n_129),
.CON(n_308),
.SN(n_308)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_125),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_122),
.B(n_125),
.Y(n_212)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_132),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_141),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_135),
.B1(n_147),
.B2(n_150),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_135),
.B(n_137),
.C(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_135),
.B(n_150),
.C(n_151),
.Y(n_328)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_137),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_144),
.B(n_145),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_151),
.Y(n_145)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

AOI321xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_306),
.A3(n_314),
.B1(n_319),
.B2(n_324),
.C(n_338),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_207),
.C(n_219),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_189),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_155),
.B(n_189),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_174),
.C(n_181),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_156),
.B(n_303),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_169),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_164),
.B2(n_165),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_165),
.C(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_171),
.B(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_172),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_174),
.A2(n_181),
.B1(n_182),
.B2(n_304),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_174),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_175),
.B(n_177),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_180),
.Y(n_195)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_188),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_183),
.B(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_186),
.B(n_188),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_187),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_197),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_191),
.B(n_196),
.C(n_197),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_192),
.B(n_194),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_206),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_203),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_203),
.C(n_206),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g320 ( 
.A1(n_208),
.A2(n_321),
.B(n_322),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_209),
.B(n_210),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_218),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_212),
.B(n_213),
.C(n_218),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_214),
.B(n_216),
.C(n_217),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_300),
.B(n_305),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_286),
.B(n_299),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_264),
.B(n_285),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_244),
.B(n_263),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_234),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_224),
.B(n_234),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_225),
.A2(n_226),
.B1(n_230),
.B2(n_231),
.Y(n_250)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_228),
.Y(n_232)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_241),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_240),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_242),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_251),
.B(n_262),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_250),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_256),
.B(n_261),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_253),
.B(n_255),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_265),
.B(n_266),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_277),
.B1(n_283),
.B2(n_284),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_272),
.B1(n_275),
.B2(n_276),
.Y(n_267)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_268),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_276),
.C(n_284),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_274),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_277),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_281),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_288),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_295),
.C(n_297),
.Y(n_301)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_297),
.B2(n_298),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_295),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_311),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_311),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.C(n_310),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_308),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_315),
.A2(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_316),
.B(n_317),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_329),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);


endmodule