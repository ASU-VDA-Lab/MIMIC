module fake_jpeg_22746_n_321 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_4),
.B(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_0),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_46),
.Y(n_80)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_2),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_45),
.A2(n_25),
.B1(n_28),
.B2(n_22),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_50),
.A2(n_51),
.B1(n_76),
.B2(n_85),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_45),
.A2(n_25),
.B1(n_22),
.B2(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_25),
.B1(n_36),
.B2(n_29),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_53),
.A2(n_54),
.B1(n_59),
.B2(n_66),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_29),
.B1(n_36),
.B2(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_57),
.B(n_17),
.Y(n_114)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_65),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_19),
.B1(n_37),
.B2(n_34),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_62),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_4),
.Y(n_62)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_41),
.A2(n_40),
.B1(n_26),
.B2(n_24),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_67),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g68 ( 
.A(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_69),
.Y(n_100)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_73),
.Y(n_109)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_41),
.A2(n_37),
.B1(n_34),
.B2(n_21),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_39),
.A2(n_33),
.B1(n_32),
.B2(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_79),
.A2(n_82),
.B1(n_23),
.B2(n_35),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_40),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_82)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g119 ( 
.A(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_42),
.B(n_18),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_31),
.B1(n_30),
.B2(n_33),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_86),
.A2(n_20),
.B1(n_23),
.B2(n_10),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_71),
.B(n_4),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_87),
.B(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_38),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_102),
.Y(n_136)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_80),
.Y(n_90)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_91),
.B(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_83),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_38),
.C(n_35),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_38),
.C(n_35),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_60),
.B(n_5),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_94),
.B(n_114),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_101),
.Y(n_131)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_61),
.B(n_38),
.Y(n_102)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_106),
.B(n_108),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_64),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_54),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_116),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_64),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_62),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_118),
.Y(n_144)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

BUFx10_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_120),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_53),
.B(n_5),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_121),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_110),
.A2(n_63),
.B1(n_62),
.B2(n_81),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_122),
.A2(n_126),
.B1(n_102),
.B2(n_106),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_127),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_81),
.B1(n_78),
.B2(n_56),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_145),
.B1(n_147),
.B2(n_91),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_74),
.B1(n_68),
.B2(n_75),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_80),
.C(n_73),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_128),
.B(n_130),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_107),
.Y(n_130)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_105),
.B(n_90),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_132),
.A2(n_144),
.B(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_150),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_152),
.C(n_99),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_17),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_148),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_96),
.A2(n_72),
.B1(n_55),
.B2(n_35),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_6),
.Y(n_146)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_146),
.A2(n_104),
.A3(n_114),
.B1(n_97),
.B2(n_11),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_89),
.A2(n_20),
.B1(n_23),
.B2(n_10),
.Y(n_147)
);

BUFx8_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_111),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_151),
.Y(n_177)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_7),
.C(n_8),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_153),
.B(n_103),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_155),
.A2(n_169),
.B1(n_168),
.B2(n_133),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_156),
.A2(n_88),
.B1(n_137),
.B2(n_112),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_158),
.B(n_161),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_94),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_164),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_121),
.B(n_95),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_170),
.B(n_179),
.Y(n_203)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_131),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_107),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_103),
.C(n_92),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_183),
.C(n_152),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_118),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_175),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_148),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_145),
.A2(n_88),
.B1(n_119),
.B2(n_101),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_119),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_172),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_112),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_139),
.B(n_7),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_176),
.B(n_186),
.Y(n_211)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_123),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_184),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_119),
.Y(n_182)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_126),
.B(n_8),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_154),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_187),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_138),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_134),
.A2(n_98),
.B(n_10),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_8),
.B(n_11),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_128),
.B(n_146),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_191),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_204),
.C(n_183),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g195 ( 
.A(n_164),
.B(n_140),
.CI(n_153),
.CON(n_195),
.SN(n_195)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_197),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_196),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_169),
.B1(n_158),
.B2(n_157),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_199),
.A2(n_206),
.B1(n_217),
.B2(n_163),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_137),
.C(n_120),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_209),
.Y(n_220)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_174),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_210),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_120),
.Y(n_212)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_173),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_214),
.Y(n_226)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_12),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_156),
.A2(n_143),
.B1(n_151),
.B2(n_14),
.Y(n_217)
);

AOI21x1_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_12),
.B(n_13),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_218),
.B(n_188),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_224),
.C(n_239),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_SL g249 ( 
.A1(n_221),
.A2(n_218),
.B(n_216),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_211),
.B(n_176),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_223),
.B(n_235),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_198),
.B(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_231),
.Y(n_251)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_189),
.B(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_232),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_178),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_236),
.A2(n_199),
.B1(n_214),
.B2(n_201),
.Y(n_245)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_237),
.A2(n_238),
.B(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_190),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_204),
.B(n_181),
.C(n_186),
.Y(n_239)
);

INVxp33_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_210),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_193),
.B(n_181),
.C(n_184),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_242),
.C(n_219),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_160),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_253),
.B1(n_257),
.B2(n_230),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_250),
.C(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_189),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_248),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_229),
.B(n_203),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_258),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_239),
.B(n_191),
.C(n_212),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_252),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_234),
.A2(n_208),
.B1(n_202),
.B2(n_213),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_202),
.C(n_192),
.Y(n_254)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_256),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_209),
.B(n_207),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_206),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_220),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_261),
.Y(n_266)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_226),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_247),
.B(n_232),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_269),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_228),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_228),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_271),
.A2(n_200),
.B(n_185),
.Y(n_290)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

INVxp67_ASAP7_75t_SL g280 ( 
.A(n_272),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_226),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.C(n_275),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_244),
.B(n_227),
.C(n_231),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_227),
.C(n_225),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_245),
.A2(n_222),
.B1(n_220),
.B2(n_225),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_205),
.B1(n_195),
.B2(n_181),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_248),
.A2(n_238),
.B(n_237),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_215),
.B(n_195),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_272),
.A2(n_250),
.B1(n_251),
.B2(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_263),
.B(n_254),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_285),
.C(n_291),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_290),
.B(n_277),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_263),
.B(n_246),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_236),
.C(n_205),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_267),
.C(n_274),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_289),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_268),
.B(n_200),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_197),
.B(n_221),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_291),
.B(n_266),
.C(n_278),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_287),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_279),
.C(n_267),
.Y(n_307)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_295),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_265),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_297),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_167),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_273),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_279),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_306),
.C(n_307),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_296),
.B(n_280),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_308),
.B(n_282),
.C(n_262),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_303),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_310),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_298),
.Y(n_311)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_311),
.A2(n_304),
.A3(n_292),
.B1(n_302),
.B2(n_262),
.C1(n_13),
.C2(n_15),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_307),
.C(n_285),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_314),
.B(n_309),
.C(n_12),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_315),
.B(n_312),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_318),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_319),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_316),
.Y(n_321)
);


endmodule