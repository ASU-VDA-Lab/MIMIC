module fake_netlist_6_3110_n_891 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_891);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_891;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_872;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_707;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_361;
wire n_508;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_26),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_38),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_88),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_107),
.Y(n_175)
);

BUFx5_ASAP7_75t_L g176 ( 
.A(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_52),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_32),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_27),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_168),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_83),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_15),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_95),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_106),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_39),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_152),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_92),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_127),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_99),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_67),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_1),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_55),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_34),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_149),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_129),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_17),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_1),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_57),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_166),
.Y(n_209)
);

BUFx5_ASAP7_75t_L g210 ( 
.A(n_151),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_102),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_121),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_0),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_161),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_159),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_96),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_165),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_85),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_71),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_132),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_21),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_160),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_23),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_163),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_70),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_150),
.B(n_25),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_77),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_53),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_20),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_47),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_141),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_148),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_153),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_28),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_157),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_14),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_137),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_64),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_146),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_118),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_11),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_15),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_42),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_147),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_60),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_87),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_36),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_155),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_169),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_142),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_3),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_50),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_109),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_4),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_91),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_44),
.Y(n_260)
);

INVx5_ASAP7_75t_L g261 ( 
.A(n_217),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_176),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_176),
.Y(n_263)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_217),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_176),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_213),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_197),
.B(n_0),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_220),
.B(n_2),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_172),
.B(n_19),
.Y(n_269)
);

OA21x2_ASAP7_75t_L g270 ( 
.A1(n_244),
.A2(n_177),
.B(n_173),
.Y(n_270)
);

BUFx8_ASAP7_75t_SL g271 ( 
.A(n_187),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_189),
.B(n_2),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_213),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_179),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_180),
.Y(n_275)
);

OAI22x1_ASAP7_75t_R g276 ( 
.A1(n_185),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_191),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_224),
.B(n_22),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_216),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_280)
);

CKINVDCx6p67_ASAP7_75t_R g281 ( 
.A(n_195),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_176),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_203),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_205),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_181),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_176),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_226),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_190),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_198),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_186),
.B(n_6),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_199),
.A2(n_8),
.B(n_9),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_202),
.B(n_24),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_254),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_190),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_208),
.Y(n_300)
);

INVx5_ASAP7_75t_L g301 ( 
.A(n_190),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_190),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_209),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_190),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_249),
.Y(n_306)
);

BUFx8_ASAP7_75t_SL g307 ( 
.A(n_215),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_210),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_252),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_210),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_210),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_253),
.B(n_30),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_228),
.B(n_31),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_255),
.Y(n_315)
);

CKINVDCx6p67_ASAP7_75t_R g316 ( 
.A(n_240),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_219),
.B(n_10),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

OA21x2_ASAP7_75t_L g319 ( 
.A1(n_260),
.A2(n_10),
.B(n_11),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_171),
.Y(n_320)
);

BUFx8_ASAP7_75t_SL g321 ( 
.A(n_242),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_175),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_R g325 ( 
.A(n_284),
.B(n_12),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_287),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_271),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_271),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_279),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_307),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_R g333 ( 
.A(n_293),
.B(n_251),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_285),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_307),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_321),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_321),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_316),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_285),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_285),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_281),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_281),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_320),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_320),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_261),
.Y(n_349)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_292),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_298),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_298),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_261),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_275),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_261),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_277),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_273),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_300),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_261),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_293),
.B(n_178),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_288),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_303),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_264),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_264),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_305),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_264),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_283),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_264),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

NOR2xp67_ASAP7_75t_L g374 ( 
.A(n_301),
.B(n_182),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_283),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_266),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_290),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_323),
.B(n_269),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_354),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_269),
.Y(n_380)
);

NAND2xp33_ASAP7_75t_L g381 ( 
.A(n_347),
.B(n_314),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_269),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_332),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_278),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_332),
.B(n_322),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_341),
.B(n_278),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_290),
.Y(n_387)
);

NAND3xp33_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_317),
.C(n_268),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_278),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_365),
.B(n_377),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_324),
.B(n_295),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_336),
.B(n_295),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_329),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_359),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_375),
.B(n_295),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_361),
.B(n_313),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_313),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_374),
.B(n_313),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_362),
.A2(n_268),
.B(n_310),
.C(n_315),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_352),
.Y(n_401)
);

NAND2xp33_ASAP7_75t_L g402 ( 
.A(n_333),
.B(n_314),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_369),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_SL g406 ( 
.A(n_360),
.B(n_267),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_376),
.B(n_280),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_329),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_351),
.B(n_270),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_270),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_349),
.B(n_355),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_331),
.B(n_306),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_358),
.B(n_306),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_331),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_329),
.B(n_270),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_360),
.Y(n_417)
);

AND2x6_ASAP7_75t_L g418 ( 
.A(n_334),
.B(n_262),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_363),
.B(n_183),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_325),
.Y(n_420)
);

NAND3xp33_ASAP7_75t_L g421 ( 
.A(n_325),
.B(n_291),
.C(n_300),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_334),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_334),
.B(n_314),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_367),
.B(n_368),
.Y(n_425)
);

NOR3xp33_ASAP7_75t_L g426 ( 
.A(n_340),
.B(n_188),
.C(n_184),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_334),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_L g428 ( 
.A(n_370),
.B(n_314),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_344),
.B(n_192),
.Y(n_429)
);

NAND2xp33_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_314),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_350),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_350),
.Y(n_432)
);

INVxp33_ASAP7_75t_L g433 ( 
.A(n_326),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_327),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_335),
.B(n_193),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_345),
.B(n_194),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_342),
.B(n_301),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_328),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_337),
.B(n_301),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_339),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_330),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_338),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_332),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_323),
.B(n_301),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_354),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_378),
.B(n_294),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_404),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_379),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_392),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g451 ( 
.A1(n_420),
.A2(n_319),
.B1(n_294),
.B2(n_243),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_380),
.B(n_294),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_396),
.B(n_196),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_420),
.A2(n_319),
.B1(n_241),
.B2(n_238),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_384),
.B(n_319),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_L g456 ( 
.A1(n_410),
.A2(n_299),
.B1(n_312),
.B2(n_311),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_382),
.B(n_200),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

BUFx4f_ASAP7_75t_L g459 ( 
.A(n_439),
.Y(n_459)
);

OR2x2_ASAP7_75t_SL g460 ( 
.A(n_388),
.B(n_276),
.Y(n_460)
);

INVx5_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_SL g462 ( 
.A(n_407),
.B(n_204),
.C(n_201),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_411),
.A2(n_299),
.B1(n_312),
.B2(n_311),
.Y(n_463)
);

AND3x1_ASAP7_75t_L g464 ( 
.A(n_413),
.B(n_289),
.C(n_263),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_387),
.B(n_207),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_395),
.B(n_211),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_212),
.Y(n_467)
);

INVx5_ASAP7_75t_L g468 ( 
.A(n_418),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_421),
.B(n_214),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_405),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_383),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_444),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_446),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_390),
.B(n_218),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_400),
.B(n_221),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_397),
.B(n_222),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_391),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_417),
.B(n_223),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_393),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_437),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_415),
.Y(n_482)
);

AND3x1_ASAP7_75t_SL g483 ( 
.A(n_431),
.B(n_13),
.C(n_16),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_422),
.A2(n_250),
.B1(n_227),
.B2(n_229),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_432),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_225),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_414),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_394),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_394),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_R g493 ( 
.A(n_434),
.B(n_230),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_385),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_416),
.B(n_262),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_422),
.A2(n_257),
.B1(n_232),
.B2(n_233),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_389),
.B(n_231),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_413),
.B(n_234),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_399),
.B(n_235),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_423),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_408),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_408),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_426),
.B(n_236),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_427),
.B(n_246),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_L g506 ( 
.A1(n_381),
.A2(n_282),
.B1(n_309),
.B2(n_263),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_445),
.B(n_247),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_424),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_402),
.B(n_248),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_440),
.B(n_256),
.Y(n_511)
);

BUFx2_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_418),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_430),
.B(n_265),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_406),
.B(n_16),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_428),
.B(n_438),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_495),
.A2(n_419),
.B(n_412),
.Y(n_518)
);

NOR3xp33_ASAP7_75t_SL g519 ( 
.A(n_462),
.B(n_436),
.C(n_429),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

AO22x1_ASAP7_75t_L g521 ( 
.A1(n_498),
.A2(n_433),
.B1(n_435),
.B2(n_441),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_489),
.B(n_418),
.Y(n_522)
);

O2A1O1Ixp33_ASAP7_75t_L g523 ( 
.A1(n_486),
.A2(n_425),
.B(n_289),
.C(n_309),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_482),
.B(n_259),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_477),
.B(n_265),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_450),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_479),
.B(n_282),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_488),
.B(n_442),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_481),
.B(n_286),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_514),
.A2(n_304),
.B(n_286),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_459),
.B(n_304),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_492),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_480),
.B(n_17),
.Y(n_533)
);

O2A1O1Ixp5_ASAP7_75t_L g534 ( 
.A1(n_452),
.A2(n_318),
.B(n_308),
.C(n_302),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_454),
.A2(n_318),
.B1(n_308),
.B2(n_302),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_501),
.Y(n_536)
);

A2O1A1Ixp33_ASAP7_75t_L g537 ( 
.A1(n_508),
.A2(n_453),
.B(n_494),
.C(n_452),
.Y(n_537)
);

NOR3xp33_ASAP7_75t_SL g538 ( 
.A(n_496),
.B(n_18),
.C(n_33),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_512),
.B(n_18),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_470),
.Y(n_540)
);

O2A1O1Ixp33_ASAP7_75t_L g541 ( 
.A1(n_469),
.A2(n_318),
.B(n_308),
.C(n_302),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_447),
.A2(n_318),
.B1(n_308),
.B2(n_302),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_516),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_543)
);

A2O1A1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_455),
.A2(n_473),
.B(n_454),
.C(n_514),
.Y(n_544)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_455),
.A2(n_43),
.B(n_45),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_502),
.B(n_505),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_464),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_515),
.B(n_51),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_465),
.B(n_54),
.Y(n_549)
);

AOI21xp33_ASAP7_75t_L g550 ( 
.A1(n_485),
.A2(n_497),
.B(n_499),
.Y(n_550)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_485),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_476),
.B(n_61),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_458),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_496),
.B(n_62),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_492),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_478),
.B(n_63),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_510),
.A2(n_65),
.B(n_66),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_474),
.B(n_68),
.Y(n_558)
);

O2A1O1Ixp5_ASAP7_75t_L g559 ( 
.A1(n_507),
.A2(n_69),
.B(n_72),
.C(n_73),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_475),
.Y(n_560)
);

A2O1A1Ixp33_ASAP7_75t_L g561 ( 
.A1(n_475),
.A2(n_74),
.B(n_75),
.C(n_78),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_464),
.B(n_80),
.Y(n_562)
);

O2A1O1Ixp33_ASAP7_75t_SL g563 ( 
.A1(n_451),
.A2(n_81),
.B(n_82),
.C(n_84),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_500),
.Y(n_564)
);

BUFx4f_ASAP7_75t_L g565 ( 
.A(n_487),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_492),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_448),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_504),
.B(n_86),
.Y(n_568)
);

BUFx12f_ASAP7_75t_L g569 ( 
.A(n_460),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_471),
.B(n_89),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_461),
.A2(n_468),
.B(n_506),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_448),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_484),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_459),
.B(n_90),
.Y(n_575)
);

BUFx3_ASAP7_75t_L g576 ( 
.A(n_553),
.Y(n_576)
);

CKINVDCx8_ASAP7_75t_R g577 ( 
.A(n_532),
.Y(n_577)
);

AO21x2_ASAP7_75t_L g578 ( 
.A1(n_544),
.A2(n_451),
.B(n_457),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_560),
.B(n_487),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_520),
.B(n_503),
.Y(n_580)
);

INVx6_ASAP7_75t_L g581 ( 
.A(n_532),
.Y(n_581)
);

OAI21x1_ASAP7_75t_L g582 ( 
.A1(n_517),
.A2(n_513),
.B(n_509),
.Y(n_582)
);

CKINVDCx11_ASAP7_75t_R g583 ( 
.A(n_569),
.Y(n_583)
);

AO21x2_ASAP7_75t_L g584 ( 
.A1(n_550),
.A2(n_466),
.B(n_467),
.Y(n_584)
);

OAI21x1_ASAP7_75t_L g585 ( 
.A1(n_534),
.A2(n_491),
.B(n_490),
.Y(n_585)
);

NOR2xp67_ASAP7_75t_R g586 ( 
.A(n_566),
.B(n_468),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_528),
.B(n_503),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_565),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_536),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_526),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_456),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_564),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_546),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_575),
.B(n_573),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_532),
.Y(n_596)
);

INVxp33_ASAP7_75t_L g597 ( 
.A(n_533),
.Y(n_597)
);

NOR2xp67_ASAP7_75t_SL g598 ( 
.A(n_555),
.B(n_461),
.Y(n_598)
);

BUFx6f_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_574),
.Y(n_600)
);

INVx8_ASAP7_75t_L g601 ( 
.A(n_555),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_567),
.Y(n_602)
);

AND2x4_ASAP7_75t_L g603 ( 
.A(n_519),
.B(n_572),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_565),
.Y(n_604)
);

BUFx2_ASAP7_75t_R g605 ( 
.A(n_562),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_566),
.Y(n_606)
);

AO21x2_ASAP7_75t_L g607 ( 
.A1(n_537),
.A2(n_511),
.B(n_493),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_538),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_525),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_524),
.Y(n_610)
);

AO21x1_ASAP7_75t_L g611 ( 
.A1(n_554),
.A2(n_558),
.B(n_556),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_527),
.Y(n_612)
);

NAND2x1_ASAP7_75t_L g613 ( 
.A(n_522),
.B(n_491),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_568),
.A2(n_463),
.B(n_468),
.Y(n_614)
);

AO21x2_ASAP7_75t_L g615 ( 
.A1(n_518),
.A2(n_483),
.B(n_461),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_529),
.B(n_170),
.Y(n_616)
);

BUFx4_ASAP7_75t_SL g617 ( 
.A(n_521),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_570),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_548),
.B(n_93),
.Y(n_619)
);

BUFx3_ASAP7_75t_L g620 ( 
.A(n_549),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_543),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_559),
.Y(n_622)
);

AO21x2_ASAP7_75t_L g623 ( 
.A1(n_552),
.A2(n_94),
.B(n_97),
.Y(n_623)
);

INVx3_ASAP7_75t_SL g624 ( 
.A(n_531),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_589),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_590),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_593),
.B(n_523),
.Y(n_627)
);

BUFx2_ASAP7_75t_R g628 ( 
.A(n_576),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_592),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_593),
.B(n_547),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_576),
.Y(n_631)
);

NAND2x1p5_ASAP7_75t_L g632 ( 
.A(n_621),
.B(n_613),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_577),
.Y(n_633)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_594),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_577),
.Y(n_635)
);

OAI22xp33_ASAP7_75t_L g636 ( 
.A1(n_597),
.A2(n_621),
.B1(n_608),
.B2(n_580),
.Y(n_636)
);

OAI22xp5_ASAP7_75t_L g637 ( 
.A1(n_621),
.A2(n_571),
.B1(n_551),
.B2(n_535),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g638 ( 
.A(n_595),
.Y(n_638)
);

OAI21x1_ASAP7_75t_SL g639 ( 
.A1(n_611),
.A2(n_545),
.B(n_557),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_589),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_606),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_609),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_582),
.Y(n_643)
);

OA21x2_ASAP7_75t_L g644 ( 
.A1(n_614),
.A2(n_530),
.B(n_561),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_600),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_587),
.A2(n_535),
.B1(n_542),
.B2(n_563),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_582),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_602),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_585),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_612),
.B(n_98),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_585),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_591),
.B(n_100),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_591),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_578),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_578),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_606),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_616),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_616),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_622),
.A2(n_541),
.B(n_103),
.Y(n_659)
);

AOI21x1_ASAP7_75t_L g660 ( 
.A1(n_622),
.A2(n_101),
.B(n_104),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_615),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_614),
.A2(n_619),
.B(n_579),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_603),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_615),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_599),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_619),
.A2(n_108),
.B(n_110),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_601),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_595),
.Y(n_668)
);

OAI21xp5_ASAP7_75t_SL g669 ( 
.A1(n_636),
.A2(n_587),
.B(n_597),
.Y(n_669)
);

NOR3xp33_ASAP7_75t_SL g670 ( 
.A(n_663),
.B(n_617),
.C(n_608),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_642),
.B(n_595),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_579),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_626),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_634),
.Y(n_674)
);

INVx3_ASAP7_75t_L g675 ( 
.A(n_667),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_629),
.Y(n_676)
);

BUFx6f_ASAP7_75t_L g677 ( 
.A(n_633),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_657),
.A2(n_603),
.B1(n_610),
.B2(n_604),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_638),
.B(n_588),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_628),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_645),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_631),
.B(n_588),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_634),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_631),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_657),
.A2(n_603),
.B1(n_624),
.B2(n_620),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_668),
.B(n_605),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_652),
.B(n_624),
.Y(n_687)
);

CKINVDCx16_ASAP7_75t_R g688 ( 
.A(n_633),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_652),
.B(n_581),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_R g690 ( 
.A(n_650),
.B(n_583),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_642),
.B(n_620),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_635),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_635),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_640),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_650),
.B(n_653),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_625),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_625),
.Y(n_697)
);

AO31x2_ASAP7_75t_L g698 ( 
.A1(n_643),
.A2(n_596),
.A3(n_607),
.B(n_584),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_653),
.B(n_658),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_SL g700 ( 
.A(n_658),
.B(n_646),
.C(n_630),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_640),
.Y(n_701)
);

AOI21xp33_ASAP7_75t_L g702 ( 
.A1(n_637),
.A2(n_584),
.B(n_607),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_639),
.A2(n_607),
.B1(n_584),
.B2(n_618),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_648),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_667),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_667),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_641),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_641),
.B(n_581),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_632),
.A2(n_618),
.B1(n_581),
.B2(n_606),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_SL g710 ( 
.A1(n_639),
.A2(n_623),
.B1(n_601),
.B2(n_606),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_641),
.B(n_599),
.Y(n_711)
);

AO31x2_ASAP7_75t_L g712 ( 
.A1(n_643),
.A2(n_596),
.A3(n_623),
.B(n_586),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_SL g713 ( 
.A(n_632),
.B(n_596),
.C(n_583),
.Y(n_713)
);

OR2x6_ASAP7_75t_L g714 ( 
.A(n_656),
.B(n_601),
.Y(n_714)
);

AOI211xp5_ASAP7_75t_L g715 ( 
.A1(n_627),
.A2(n_662),
.B(n_664),
.C(n_661),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_665),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_665),
.Y(n_717)
);

NAND2x1p5_ASAP7_75t_L g718 ( 
.A(n_685),
.B(n_662),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_694),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_695),
.B(n_664),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_701),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_683),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_676),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_681),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_672),
.B(n_661),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_699),
.B(n_654),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_698),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_704),
.B(n_654),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_702),
.A2(n_715),
.B(n_700),
.Y(n_730)
);

OR2x2_ASAP7_75t_L g731 ( 
.A(n_698),
.B(n_655),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_698),
.B(n_655),
.Y(n_732)
);

NAND3xp33_ASAP7_75t_L g733 ( 
.A(n_669),
.B(n_644),
.C(n_656),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_696),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_697),
.Y(n_735)
);

OAI211xp5_ASAP7_75t_L g736 ( 
.A1(n_678),
.A2(n_666),
.B(n_660),
.C(n_644),
.Y(n_736)
);

HB1xp67_ASAP7_75t_L g737 ( 
.A(n_674),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_703),
.B(n_647),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_712),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_691),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_671),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_717),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_707),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_685),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_687),
.B(n_656),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_678),
.B(n_665),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_711),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_689),
.B(n_647),
.Y(n_748)
);

NOR4xp25_ASAP7_75t_SL g749 ( 
.A(n_690),
.B(n_666),
.C(n_660),
.D(n_632),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_679),
.B(n_665),
.Y(n_750)
);

AO21x2_ASAP7_75t_L g751 ( 
.A1(n_713),
.A2(n_651),
.B(n_649),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_679),
.B(n_665),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_712),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_708),
.B(n_651),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_712),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_719),
.Y(n_756)
);

HB1xp67_ASAP7_75t_L g757 ( 
.A(n_728),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_728),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_740),
.B(n_688),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_719),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_722),
.B(n_686),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_720),
.B(n_649),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_720),
.B(n_710),
.Y(n_763)
);

HB1xp67_ASAP7_75t_L g764 ( 
.A(n_729),
.Y(n_764)
);

AOI221xp5_ASAP7_75t_L g765 ( 
.A1(n_730),
.A2(n_670),
.B1(n_709),
.B2(n_677),
.C(n_692),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_747),
.B(n_677),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_721),
.B(n_682),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_723),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_741),
.B(n_677),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_722),
.B(n_693),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_724),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_721),
.B(n_682),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_726),
.B(n_748),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_725),
.B(n_675),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_738),
.B(n_644),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_726),
.B(n_684),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_738),
.B(n_644),
.Y(n_777)
);

NOR2x1_ASAP7_75t_L g778 ( 
.A(n_733),
.B(n_706),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_748),
.B(n_716),
.Y(n_779)
);

OAI22xp5_ASAP7_75t_L g780 ( 
.A1(n_744),
.A2(n_680),
.B1(n_705),
.B2(n_714),
.Y(n_780)
);

NAND3xp33_ASAP7_75t_L g781 ( 
.A(n_765),
.B(n_746),
.C(n_745),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_756),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_760),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_764),
.B(n_718),
.Y(n_784)
);

OR2x2_ASAP7_75t_L g785 ( 
.A(n_764),
.B(n_731),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_773),
.B(n_763),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_763),
.B(n_718),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_768),
.Y(n_788)
);

BUFx2_ASAP7_75t_L g789 ( 
.A(n_767),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_771),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_775),
.B(n_718),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_775),
.B(n_729),
.Y(n_792)
);

INVxp67_ASAP7_75t_L g793 ( 
.A(n_759),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_777),
.B(n_739),
.Y(n_794)
);

INVxp67_ASAP7_75t_L g795 ( 
.A(n_770),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_777),
.B(n_739),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_767),
.B(n_737),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_767),
.Y(n_798)
);

OAI33xp33_ASAP7_75t_L g799 ( 
.A1(n_788),
.A2(n_769),
.A3(n_761),
.B1(n_780),
.B2(n_742),
.B3(n_743),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_789),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_782),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_792),
.B(n_762),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_790),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_783),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_798),
.Y(n_805)
);

NOR4xp25_ASAP7_75t_L g806 ( 
.A(n_781),
.B(n_736),
.C(n_776),
.D(n_734),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_785),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_785),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_804),
.Y(n_809)
);

XNOR2xp5_ASAP7_75t_L g810 ( 
.A(n_806),
.B(n_766),
.Y(n_810)
);

OAI21xp5_ASAP7_75t_L g811 ( 
.A1(n_806),
.A2(n_778),
.B(n_793),
.Y(n_811)
);

AO21x1_ASAP7_75t_L g812 ( 
.A1(n_801),
.A2(n_808),
.B(n_807),
.Y(n_812)
);

OAI221xp5_ASAP7_75t_SL g813 ( 
.A1(n_800),
.A2(n_795),
.B1(n_791),
.B2(n_787),
.C(n_797),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_803),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_810),
.B(n_786),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_812),
.Y(n_816)
);

NOR3xp33_ASAP7_75t_L g817 ( 
.A(n_811),
.B(n_799),
.C(n_752),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_809),
.B(n_805),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_814),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_813),
.A2(n_787),
.B1(n_802),
.B2(n_784),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_809),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_819),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_815),
.B(n_811),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_816),
.B(n_774),
.C(n_772),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_817),
.B(n_786),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_818),
.B(n_784),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_823),
.B(n_817),
.C(n_820),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_825),
.B(n_821),
.Y(n_828)
);

NOR4xp25_ASAP7_75t_L g829 ( 
.A(n_822),
.B(n_824),
.C(n_802),
.D(n_826),
.Y(n_829)
);

NAND4xp25_ASAP7_75t_SL g830 ( 
.A(n_827),
.B(n_792),
.C(n_794),
.D(n_796),
.Y(n_830)
);

NAND4xp25_ASAP7_75t_L g831 ( 
.A(n_828),
.B(n_750),
.C(n_772),
.D(n_774),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_829),
.A2(n_772),
.B1(n_774),
.B2(n_779),
.Y(n_832)
);

NOR2xp33_ASAP7_75t_SL g833 ( 
.A(n_827),
.B(n_754),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_833),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_831),
.Y(n_835)
);

OR2x2_ASAP7_75t_L g836 ( 
.A(n_830),
.B(n_832),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_830),
.B(n_714),
.Y(n_837)
);

AND2x4_ASAP7_75t_L g838 ( 
.A(n_832),
.B(n_796),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_832),
.B(n_794),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_832),
.A2(n_749),
.B1(n_758),
.B2(n_757),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_834),
.A2(n_754),
.B1(n_762),
.B2(n_757),
.Y(n_841)
);

NOR3xp33_ASAP7_75t_L g842 ( 
.A(n_835),
.B(n_675),
.C(n_659),
.Y(n_842)
);

OAI211xp5_ASAP7_75t_SL g843 ( 
.A1(n_836),
.A2(n_735),
.B(n_755),
.C(n_753),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_838),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_839),
.B(n_727),
.Y(n_845)
);

NOR2xp33_ASAP7_75t_L g846 ( 
.A(n_837),
.B(n_111),
.Y(n_846)
);

NAND3xp33_ASAP7_75t_SL g847 ( 
.A(n_840),
.B(n_735),
.C(n_727),
.Y(n_847)
);

NAND4xp75_ASAP7_75t_L g848 ( 
.A(n_837),
.B(n_601),
.C(n_598),
.D(n_115),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_835),
.B(n_113),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_844),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_849),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_R g852 ( 
.A(n_846),
.B(n_114),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_847),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_841),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_848),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_845),
.Y(n_856)
);

CKINVDCx20_ASAP7_75t_R g857 ( 
.A(n_843),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_850),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_857),
.A2(n_842),
.B1(n_758),
.B2(n_716),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_856),
.Y(n_860)
);

XNOR2xp5_ASAP7_75t_L g861 ( 
.A(n_851),
.B(n_117),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_856),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_852),
.A2(n_855),
.B(n_853),
.Y(n_863)
);

AO22x2_ASAP7_75t_L g864 ( 
.A1(n_854),
.A2(n_755),
.B1(n_753),
.B2(n_732),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_853),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_857),
.A2(n_716),
.B1(n_755),
.B2(n_753),
.Y(n_866)
);

OR3x1_ASAP7_75t_L g867 ( 
.A(n_850),
.B(n_119),
.C(n_120),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_867),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_865),
.A2(n_599),
.B1(n_732),
.B2(n_731),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_863),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_858),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_860),
.B(n_751),
.Y(n_872)
);

OAI22xp5_ASAP7_75t_SL g873 ( 
.A1(n_862),
.A2(n_599),
.B1(n_123),
.B2(n_125),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_861),
.A2(n_859),
.B1(n_866),
.B2(n_864),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_864),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_860),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_860),
.B(n_751),
.Y(n_877)
);

XOR2xp5_ASAP7_75t_L g878 ( 
.A(n_868),
.B(n_122),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_871),
.A2(n_659),
.B(n_128),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_876),
.Y(n_880)
);

CKINVDCx20_ASAP7_75t_R g881 ( 
.A(n_870),
.Y(n_881)
);

OAI22xp5_ASAP7_75t_L g882 ( 
.A1(n_874),
.A2(n_751),
.B1(n_130),
.B2(n_134),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_872),
.A2(n_877),
.B(n_875),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_880),
.Y(n_884)
);

AND3x4_ASAP7_75t_L g885 ( 
.A(n_881),
.B(n_873),
.C(n_869),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_878),
.Y(n_886)
);

NAND3xp33_ASAP7_75t_L g887 ( 
.A(n_884),
.B(n_883),
.C(n_886),
.Y(n_887)
);

NAND3xp33_ASAP7_75t_L g888 ( 
.A(n_885),
.B(n_882),
.C(n_879),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_887),
.A2(n_126),
.B1(n_135),
.B2(n_136),
.Y(n_889)
);

AOI221xp5_ASAP7_75t_L g890 ( 
.A1(n_889),
.A2(n_888),
.B1(n_139),
.B2(n_140),
.C(n_143),
.Y(n_890)
);

AOI22xp33_ASAP7_75t_L g891 ( 
.A1(n_890),
.A2(n_138),
.B1(n_144),
.B2(n_145),
.Y(n_891)
);


endmodule