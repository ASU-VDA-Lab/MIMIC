module fake_jpeg_16804_n_301 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx11_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_13),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_41),
.B(n_47),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_26),
.B(n_11),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_11),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_51),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_25),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_70),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_57),
.Y(n_79)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_24),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_65),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_62),
.Y(n_75)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_24),
.B(n_9),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_64),
.B(n_8),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_28),
.B(n_30),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_67),
.Y(n_110)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_69),
.B(n_20),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_0),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_50),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_39),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_67),
.A2(n_29),
.B1(n_14),
.B2(n_16),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_88),
.A2(n_95),
.B(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_31),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_102),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_40),
.B(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_90),
.B(n_113),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_29),
.B1(n_32),
.B2(n_38),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_92),
.A2(n_84),
.B1(n_96),
.B2(n_103),
.Y(n_155)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_58),
.A2(n_33),
.B1(n_38),
.B2(n_27),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_100),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_59),
.A2(n_33),
.B1(n_27),
.B2(n_19),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_34),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_45),
.A2(n_19),
.B1(n_17),
.B2(n_34),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_107),
.B1(n_112),
.B2(n_57),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_55),
.A2(n_31),
.B1(n_28),
.B2(n_35),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_69),
.A2(n_39),
.B1(n_23),
.B2(n_2),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_56),
.B(n_8),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_48),
.Y(n_115)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g174 ( 
.A1(n_119),
.A2(n_120),
.B(n_147),
.C(n_133),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_43),
.B(n_39),
.C(n_2),
.Y(n_120)
);

O2A1O1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_144),
.B(n_152),
.C(n_156),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_121),
.B(n_127),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_73),
.B(n_8),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_123),
.B(n_64),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_0),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_125),
.A2(n_157),
.B(n_159),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_81),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_132),
.B1(n_133),
.B2(n_139),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_113),
.B(n_1),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_125),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_110),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_86),
.A2(n_5),
.B1(n_111),
.B2(n_80),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_98),
.B(n_5),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_137),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_71),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_88),
.A2(n_112),
.B1(n_101),
.B2(n_95),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_141),
.B(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_82),
.B(n_100),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_143),
.B(n_145),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_92),
.A2(n_72),
.B1(n_74),
.B2(n_80),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_85),
.B(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_154),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_72),
.A2(n_104),
.B1(n_93),
.B2(n_87),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_150),
.B(n_132),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_74),
.A2(n_106),
.B1(n_75),
.B2(n_97),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_85),
.B(n_97),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_158),
.Y(n_185)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_84),
.B(n_96),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_75),
.B(n_116),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_115),
.B(n_73),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_160),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_163),
.A2(n_161),
.B(n_174),
.Y(n_208)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

NOR3xp33_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_129),
.C(n_123),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_165),
.B(n_173),
.Y(n_195)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_166),
.Y(n_197)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_125),
.B(n_159),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_168),
.A2(n_174),
.B(n_161),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_180),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_159),
.C(n_128),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_193),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_138),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_181),
.B(n_186),
.Y(n_206)
);

AOI211xp5_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_155),
.B(n_117),
.C(n_157),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_183),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_135),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_187),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_118),
.B(n_134),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_131),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_131),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_175),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_122),
.B(n_149),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

INVxp67_ASAP7_75t_SL g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_190),
.Y(n_201)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_156),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_183),
.B1(n_174),
.B2(n_180),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_196),
.A2(n_205),
.B1(n_215),
.B2(n_193),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_202),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_176),
.A2(n_174),
.B1(n_163),
.B2(n_160),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_208),
.A2(n_170),
.B(n_167),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_173),
.B(n_186),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_219),
.Y(n_231)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_212),
.A2(n_213),
.B(n_198),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_168),
.A2(n_162),
.B(n_185),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_181),
.B(n_162),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_214),
.B(n_195),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_174),
.A2(n_179),
.B1(n_188),
.B2(n_177),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_165),
.B(n_172),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_170),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_218),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_225),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_222),
.A2(n_224),
.B(n_230),
.Y(n_248)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_171),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_220),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_191),
.B1(n_164),
.B2(n_182),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_227),
.B1(n_212),
.B2(n_205),
.Y(n_246)
);

NOR4xp25_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_192),
.C(n_219),
.D(n_194),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_208),
.C(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_199),
.C(n_209),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_237),
.Y(n_249)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_216),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_238),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_199),
.C(n_215),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_196),
.B(n_216),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_241),
.B(n_242),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_196),
.B(n_194),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_255),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_246),
.B(n_259),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_242),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_250),
.Y(n_264)
);

AO221x1_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_204),
.B1(n_200),
.B2(n_197),
.C(n_217),
.Y(n_251)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_241),
.A2(n_202),
.B1(n_201),
.B2(n_200),
.Y(n_252)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_252),
.Y(n_269)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_238),
.A2(n_242),
.B(n_240),
.C(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_233),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_225),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_272),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_254),
.B1(n_247),
.B2(n_258),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_248),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_237),
.C(n_234),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_265),
.C(n_268),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_237),
.C(n_234),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_253),
.B(n_227),
.C(n_229),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_229),
.C(n_231),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_252),
.C(n_231),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g279 ( 
.A1(n_271),
.A2(n_230),
.B(n_232),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_224),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_273),
.B(n_274),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_269),
.A2(n_222),
.B1(n_259),
.B2(n_243),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_277),
.C(n_278),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_248),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_282),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_245),
.B1(n_255),
.B2(n_250),
.Y(n_280)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

AOI31xp67_ASAP7_75t_L g282 ( 
.A1(n_268),
.A2(n_226),
.A3(n_244),
.B(n_239),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_203),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_285),
.Y(n_291)
);

OAI21x1_ASAP7_75t_L g285 ( 
.A1(n_279),
.A2(n_270),
.B(n_262),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_267),
.B1(n_265),
.B2(n_226),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_288),
.A2(n_274),
.B1(n_266),
.B2(n_210),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_290),
.B(n_292),
.C(n_293),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_275),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_275),
.C(n_277),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_294),
.B(n_286),
.C(n_288),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_296),
.B(n_297),
.Y(n_298)
);

AOI31xp67_ASAP7_75t_SL g297 ( 
.A1(n_291),
.A2(n_294),
.A3(n_289),
.B(n_293),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_292),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_210),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_298),
.Y(n_301)
);


endmodule