module fake_jpeg_1039_n_9 (n_0, n_1, n_9);

input n_0;
input n_1;

output n_9;

wire n_3;
wire n_2;
wire n_4;
wire n_8;
wire n_6;
wire n_5;
wire n_7;

INVx6_ASAP7_75t_SL g2 ( 
.A(n_0),
.Y(n_2)
);

BUFx2_ASAP7_75t_L g3 ( 
.A(n_1),
.Y(n_3)
);

MAJIxp5_ASAP7_75t_L g4 ( 
.A(n_3),
.B(n_0),
.C(n_1),
.Y(n_4)
);

INVx1_ASAP7_75t_L g5 ( 
.A(n_4),
.Y(n_5)
);

INVx11_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_6),
.B(n_3),
.Y(n_7)
);

NAND2xp5_ASAP7_75t_L g8 ( 
.A(n_7),
.B(n_2),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_8),
.B(n_6),
.Y(n_9)
);


endmodule