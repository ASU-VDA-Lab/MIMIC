module real_aes_7820_n_398 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_398);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_398;
wire n_480;
wire n_1177;
wire n_1073;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_1066;
wire n_1178;
wire n_1096;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_1170;
wire n_1175;
wire n_1205;
wire n_778;
wire n_522;
wire n_800;
wire n_838;
wire n_933;
wire n_1092;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_503;
wire n_635;
wire n_673;
wire n_792;
wire n_1192;
wire n_518;
wire n_905;
wire n_878;
wire n_1067;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1197;
wire n_657;
wire n_1106;
wire n_900;
wire n_718;
wire n_841;
wire n_1129;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1218;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_852;
wire n_766;
wire n_1113;
wire n_974;
wire n_857;
wire n_919;
wire n_1089;
wire n_1122;
wire n_1217;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_1123;
wire n_923;
wire n_1034;
wire n_1219;
wire n_952;
wire n_429;
wire n_976;
wire n_1166;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_1110;
wire n_593;
wire n_1137;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_666;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_1094;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_1146;
wire n_983;
wire n_1220;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_1147;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_1093;
wire n_1109;
wire n_870;
wire n_961;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_564;
wire n_519;
wire n_638;
wire n_1116;
wire n_573;
wire n_510;
wire n_1140;
wire n_1099;
wire n_709;
wire n_786;
wire n_512;
wire n_743;
wire n_816;
wire n_626;
wire n_400;
wire n_539;
wire n_795;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_550;
wire n_1108;
wire n_966;
wire n_1160;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_994;
wire n_1078;
wire n_1072;
wire n_744;
wire n_938;
wire n_1128;
wire n_935;
wire n_1098;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_1199;
wire n_992;
wire n_774;
wire n_813;
wire n_1213;
wire n_981;
wire n_791;
wire n_1049;
wire n_466;
wire n_1182;
wire n_872;
wire n_636;
wire n_559;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_1086;
wire n_726;
wire n_1189;
wire n_1070;
wire n_1180;
wire n_517;
wire n_931;
wire n_780;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_904;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_1117;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_1210;
wire n_1082;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_1168;
wire n_1025;
wire n_755;
wire n_1148;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_523;
wire n_996;
wire n_909;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_1152;
wire n_801;
wire n_1126;
wire n_529;
wire n_1115;
wire n_455;
wire n_973;
wire n_504;
wire n_725;
wire n_671;
wire n_1084;
wire n_960;
wire n_1081;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_925;
wire n_608;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1121;
wire n_1207;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_1196;
wire n_1013;
wire n_737;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_1215;
wire n_620;
wire n_582;
wire n_641;
wire n_1063;
wire n_1135;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_1100;
wire n_1193;
wire n_1167;
wire n_1174;
wire n_688;
wire n_425;
wire n_609;
wire n_1042;
wire n_879;
wire n_417;
wire n_754;
wire n_607;
wire n_449;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_1198;
wire n_499;
wire n_508;
wire n_1142;
wire n_1141;
wire n_706;
wire n_901;
wire n_561;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_1112;
wire n_428;
wire n_405;
wire n_1149;
wire n_621;
wire n_783;
wire n_1107;
wire n_1012;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_1212;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_1134;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_1083;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1103;
wire n_1031;
wire n_1037;
wire n_1131;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_1095;
wire n_1060;
wire n_859;
wire n_695;
wire n_1181;
wire n_685;
wire n_881;
wire n_1154;
wire n_1080;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_1145;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_1222;
wire n_1077;
wire n_501;
wire n_488;
wire n_1041;
wire n_1111;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_1125;
wire n_957;
wire n_995;
wire n_1124;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_1202;
wire n_464;
wire n_1163;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_562;
wire n_1022;
wire n_756;
wire n_404;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_1201;
wire n_1179;
wire n_569;
wire n_997;
wire n_785;
wire n_563;
wire n_1171;
wire n_1203;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_1105;
wire n_1158;
wire n_1157;
wire n_1132;
wire n_853;
wire n_810;
wire n_843;
wire n_1079;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1028;
wire n_1187;
wire n_1000;
wire n_1003;
wire n_727;
wire n_1014;
wire n_1056;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_1155;
wire n_934;
wire n_1165;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1169;
wire n_1058;
wire n_1139;
wire n_927;
wire n_1038;
wire n_965;
wire n_1216;
wire n_723;
wire n_662;
wire n_1085;
wire n_845;
wire n_850;
wire n_1043;
wire n_1136;
wire n_720;
wire n_972;
wire n_968;
wire n_435;
wire n_1127;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_747;
wire n_1204;
wire n_486;
wire n_930;
wire n_1209;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_1005;
wire n_939;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_928;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1087;
wire n_1051;
wire n_1194;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_942;
wire n_1048;
wire n_472;
wire n_1120;
wire n_971;
wire n_866;
wire n_452;
wire n_1071;
wire n_1052;
wire n_787;
wire n_630;
wire n_1214;
wire n_806;
wire n_689;
wire n_820;
wire n_1097;
wire n_959;
wire n_715;
wire n_1208;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_1130;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_717;
wire n_456;
wire n_1090;
wire n_1133;
wire n_1164;
wire n_712;
wire n_1183;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_1162;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1195;
wire n_762;
wire n_575;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1186;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_1172;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_674;
wire n_644;
wire n_888;
wire n_836;
wire n_793;
wire n_1150;
wire n_1184;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_1161;
wire n_929;
wire n_1143;
wire n_686;
wire n_1190;
wire n_776;
wire n_1138;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_1114;
wire n_837;
wire n_967;
wire n_871;
wire n_1045;
wire n_1156;
wire n_474;
wire n_1159;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_1088;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1176;
wire n_1151;
wire n_1036;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_1211;
wire n_710;
wire n_650;
wire n_823;
wire n_652;
wire n_703;
wire n_1040;
wire n_500;
wire n_1101;
wire n_601;
wire n_661;
wire n_463;
wire n_1185;
wire n_804;
wire n_1076;
wire n_447;
wire n_1102;
wire n_1173;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_1119;
wire n_802;
wire n_868;
wire n_877;
wire n_1039;
wire n_574;
wire n_1069;
wire n_1024;
wire n_1104;
wire n_842;
wire n_1144;
wire n_849;
wire n_1061;
wire n_475;
wire n_554;
wire n_897;
wire n_1153;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g626 ( .A1(n_0), .A2(n_63), .B1(n_627), .B2(n_631), .Y(n_626) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_1), .A2(n_305), .B1(n_541), .B2(n_543), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_2), .Y(n_491) );
CKINVDCx20_ASAP7_75t_R g913 ( .A(n_3), .Y(n_913) );
CKINVDCx20_ASAP7_75t_R g849 ( .A(n_4), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_5), .Y(n_517) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_6), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g1123 ( .A1(n_7), .A2(n_57), .B1(n_634), .B2(n_1124), .Y(n_1123) );
AOI221xp5_ASAP7_75t_L g1097 ( .A1(n_8), .A2(n_16), .B1(n_959), .B2(n_1098), .C(n_1099), .Y(n_1097) );
AOI221xp5_ASAP7_75t_L g1083 ( .A1(n_9), .A2(n_293), .B1(n_695), .B2(n_992), .C(n_1084), .Y(n_1083) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_10), .A2(n_349), .B1(n_754), .B2(n_794), .C(n_1211), .Y(n_1210) );
AOI22x1_ASAP7_75t_L g1000 ( .A1(n_11), .A2(n_1001), .B1(n_1029), .B2(n_1030), .Y(n_1000) );
INVx1_ASAP7_75t_L g1029 ( .A(n_11), .Y(n_1029) );
CKINVDCx20_ASAP7_75t_R g920 ( .A(n_12), .Y(n_920) );
AO22x2_ASAP7_75t_L g433 ( .A1(n_13), .A2(n_241), .B1(n_425), .B2(n_430), .Y(n_433) );
INVx1_ASAP7_75t_L g1164 ( .A(n_13), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_14), .A2(n_170), .B1(n_419), .B2(n_436), .Y(n_418) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_15), .Y(n_1027) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_17), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_18), .A2(n_309), .B1(n_545), .B2(n_546), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_19), .A2(n_100), .B1(n_436), .B2(n_756), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g597 ( .A(n_20), .Y(n_597) );
AOI222xp33_ASAP7_75t_L g632 ( .A1(n_21), .A2(n_58), .B1(n_156), .B2(n_482), .C1(n_633), .C2(n_634), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_22), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_23), .A2(n_165), .B1(n_648), .B2(n_830), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_24), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_25), .Y(n_574) );
CKINVDCx20_ASAP7_75t_R g1116 ( .A(n_26), .Y(n_1116) );
AOI221xp5_ASAP7_75t_L g1215 ( .A1(n_27), .A2(n_38), .B1(n_688), .B2(n_959), .C(n_1216), .Y(n_1215) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_28), .A2(n_378), .B1(n_688), .B2(n_689), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_29), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_30), .Y(n_812) );
AOI222xp33_ASAP7_75t_L g1048 ( .A1(n_31), .A2(n_62), .B1(n_364), .B2(n_480), .C1(n_631), .C2(n_1049), .Y(n_1048) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_32), .A2(n_129), .B1(n_534), .B2(n_665), .Y(n_935) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_33), .Y(n_653) );
AO22x2_ASAP7_75t_L g435 ( .A1(n_34), .A2(n_112), .B1(n_425), .B2(n_426), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g1081 ( .A1(n_35), .A2(n_1082), .B1(n_1103), .B2(n_1104), .Y(n_1081) );
INVx1_ASAP7_75t_L g1103 ( .A(n_35), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_36), .A2(n_391), .B1(n_461), .B2(n_794), .Y(n_939) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_37), .A2(n_226), .B1(n_698), .B2(n_700), .Y(n_697) );
AOI22xp5_ASAP7_75t_L g784 ( .A1(n_39), .A2(n_785), .B1(n_815), .B2(n_816), .Y(n_784) );
CKINVDCx20_ASAP7_75t_R g815 ( .A(n_39), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_40), .A2(n_266), .B1(n_534), .B2(n_594), .Y(n_1046) );
INVx1_ASAP7_75t_L g1063 ( .A(n_41), .Y(n_1063) );
AOI22xp33_ASAP7_75t_L g704 ( .A1(n_42), .A2(n_59), .B1(n_453), .B2(n_455), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_43), .A2(n_116), .B1(n_420), .B2(n_612), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g1111 ( .A1(n_44), .A2(n_172), .B1(n_615), .B2(n_735), .Y(n_1111) );
CKINVDCx20_ASAP7_75t_R g1187 ( .A(n_45), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_46), .B(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g1213 ( .A(n_47), .Y(n_1213) );
AOI22xp5_ASAP7_75t_SL g710 ( .A1(n_48), .A2(n_711), .B1(n_712), .B2(n_740), .Y(n_710) );
INVx1_ASAP7_75t_L g740 ( .A(n_48), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_49), .A2(n_204), .B1(n_419), .B2(n_594), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_50), .A2(n_315), .B1(n_523), .B2(n_572), .Y(n_571) );
AOI222xp33_ASAP7_75t_L g1219 ( .A1(n_51), .A2(n_132), .B1(n_141), .B2(n_493), .C1(n_680), .C2(n_1124), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_52), .A2(n_359), .B1(n_607), .B2(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_53), .A2(n_263), .B1(n_734), .B2(n_735), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_54), .B(n_881), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g1023 ( .A(n_55), .Y(n_1023) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_56), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_60), .Y(n_773) );
AOI22xp33_ASAP7_75t_SL g886 ( .A1(n_61), .A2(n_396), .B1(n_887), .B2(n_888), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_64), .A2(n_260), .B1(n_452), .B2(n_455), .Y(n_451) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_65), .A2(n_750), .B1(n_781), .B2(n_782), .Y(n_749) );
INVx1_ASAP7_75t_L g781 ( .A(n_65), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_66), .A2(n_137), .B1(n_465), .B2(n_1016), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g982 ( .A(n_67), .B(n_493), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_68), .A2(n_343), .B1(n_619), .B2(n_762), .Y(n_1112) );
AOI22xp33_ASAP7_75t_SL g834 ( .A1(n_69), .A2(n_294), .B1(n_661), .B2(n_835), .Y(n_834) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_70), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_71), .A2(n_322), .B1(n_666), .B2(n_1009), .Y(n_1073) );
CKINVDCx20_ASAP7_75t_R g1056 ( .A(n_72), .Y(n_1056) );
AOI22xp33_ASAP7_75t_SL g890 ( .A1(n_73), .A2(n_200), .B1(n_760), .B2(n_891), .Y(n_890) );
CKINVDCx20_ASAP7_75t_R g798 ( .A(n_74), .Y(n_798) );
CKINVDCx20_ASAP7_75t_R g1185 ( .A(n_75), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_76), .A2(n_106), .B1(n_534), .B2(n_680), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g1171 ( .A(n_77), .Y(n_1171) );
INVx1_ASAP7_75t_L g621 ( .A(n_78), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_79), .A2(n_101), .B1(n_659), .B2(n_662), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_80), .A2(n_269), .B1(n_686), .B2(n_719), .Y(n_1174) );
AOI22xp5_ASAP7_75t_L g901 ( .A1(n_81), .A2(n_279), .B1(n_523), .B2(n_572), .Y(n_901) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_82), .A2(n_314), .B1(n_446), .B2(n_536), .Y(n_1047) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_83), .A2(n_337), .B1(n_494), .B2(n_633), .Y(n_877) );
AOI22xp5_ASAP7_75t_L g954 ( .A1(n_84), .A2(n_231), .B1(n_494), .B2(n_631), .Y(n_954) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_85), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g1085 ( .A(n_86), .Y(n_1085) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_87), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_88), .A2(n_140), .B1(n_726), .B2(n_727), .Y(n_1129) );
AO22x2_ASAP7_75t_L g429 ( .A1(n_89), .A2(n_270), .B1(n_425), .B2(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g1161 ( .A(n_89), .Y(n_1161) );
CKINVDCx20_ASAP7_75t_R g1135 ( .A(n_90), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_91), .A2(n_92), .B1(n_446), .B2(n_545), .Y(n_860) );
CKINVDCx20_ASAP7_75t_R g586 ( .A(n_93), .Y(n_586) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_94), .A2(n_246), .B1(n_495), .B2(n_523), .Y(n_522) );
OA22x2_ASAP7_75t_L g555 ( .A1(n_95), .A2(n_556), .B1(n_557), .B2(n_558), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_95), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_96), .A2(n_157), .B1(n_659), .B2(n_700), .Y(n_1183) );
AOI222xp33_ASAP7_75t_L g1102 ( .A1(n_97), .A2(n_109), .B1(n_144), .B2(n_480), .C1(n_528), .C2(n_1049), .Y(n_1102) );
CKINVDCx20_ASAP7_75t_R g928 ( .A(n_98), .Y(n_928) );
CKINVDCx20_ASAP7_75t_R g780 ( .A(n_99), .Y(n_780) );
INVx1_ASAP7_75t_L g502 ( .A(n_102), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_103), .A2(n_150), .B1(n_717), .B2(n_719), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_104), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_105), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_107), .A2(n_196), .B1(n_576), .B2(n_830), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_108), .A2(n_233), .B1(n_452), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_SL g730 ( .A1(n_110), .A2(n_377), .B1(n_731), .B2(n_732), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_111), .A2(n_159), .B1(n_438), .B2(n_835), .Y(n_912) );
INVx1_ASAP7_75t_L g1165 ( .A(n_112), .Y(n_1165) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_113), .A2(n_177), .B1(n_576), .B2(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g1122 ( .A(n_114), .Y(n_1122) );
CKINVDCx20_ASAP7_75t_R g930 ( .A(n_115), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_117), .A2(n_238), .B1(n_461), .B2(n_835), .Y(n_995) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_118), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_119), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g823 ( .A(n_120), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g1013 ( .A(n_121), .Y(n_1013) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_122), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g909 ( .A1(n_123), .A2(n_308), .B1(n_536), .B2(n_757), .Y(n_909) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_124), .A2(n_292), .B1(n_731), .B2(n_760), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g1020 ( .A(n_125), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1181 ( .A1(n_126), .A2(n_333), .B1(n_695), .B2(n_1182), .Y(n_1181) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_127), .A2(n_243), .B1(n_465), .B2(n_762), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_128), .A2(n_142), .B1(n_441), .B2(n_992), .Y(n_991) );
AOI22xp33_ASAP7_75t_SL g880 ( .A1(n_130), .A2(n_251), .B1(n_689), .B2(n_881), .Y(n_880) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_131), .A2(n_329), .B1(n_443), .B2(n_534), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g922 ( .A(n_133), .Y(n_922) );
AOI22xp33_ASAP7_75t_SL g1141 ( .A1(n_134), .A2(n_190), .B1(n_648), .B2(n_724), .Y(n_1141) );
NAND2xp5_ASAP7_75t_L g1173 ( .A(n_135), .B(n_1098), .Y(n_1173) );
AOI22xp33_ASAP7_75t_SL g1144 ( .A1(n_136), .A2(n_324), .B1(n_545), .B2(n_942), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_138), .A2(n_186), .B1(n_615), .B2(n_616), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_139), .A2(n_358), .B1(n_495), .B2(n_724), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g829 ( .A1(n_143), .A2(n_352), .B1(n_523), .B2(n_830), .Y(n_829) );
AOI22xp33_ASAP7_75t_SL g685 ( .A1(n_145), .A2(n_209), .B1(n_631), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g1039 ( .A1(n_146), .A2(n_356), .B1(n_698), .B2(n_738), .Y(n_1039) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_147), .A2(n_332), .B1(n_964), .B2(n_1009), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g892 ( .A1(n_148), .A2(n_334), .B1(n_452), .B2(n_455), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_149), .A2(n_222), .B1(n_436), .B2(n_970), .Y(n_969) );
CKINVDCx20_ASAP7_75t_R g1101 ( .A(n_151), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_152), .B(n_827), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_153), .A2(n_257), .B1(n_609), .B2(n_612), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_154), .A2(n_220), .B1(n_591), .B2(n_937), .Y(n_936) );
AND2x6_ASAP7_75t_L g401 ( .A(n_155), .B(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g1158 ( .A(n_155), .Y(n_1158) );
AOI22xp33_ASAP7_75t_SL g883 ( .A1(n_158), .A2(n_180), .B1(n_446), .B2(n_884), .Y(n_883) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_160), .A2(n_254), .B1(n_760), .B2(n_990), .Y(n_989) );
AOI22xp33_ASAP7_75t_SL g1127 ( .A1(n_161), .A2(n_299), .B1(n_719), .B2(n_1128), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g859 ( .A1(n_162), .A2(n_188), .B1(n_462), .B2(n_536), .Y(n_859) );
INVx1_ASAP7_75t_L g985 ( .A(n_163), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_164), .A2(n_283), .B1(n_486), .B2(n_668), .Y(n_857) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_166), .Y(n_640) );
AO22x1_ASAP7_75t_L g1209 ( .A1(n_167), .A2(n_176), .B1(n_990), .B2(n_1009), .Y(n_1209) );
CKINVDCx20_ASAP7_75t_R g1100 ( .A(n_168), .Y(n_1100) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_169), .A2(n_280), .B1(n_453), .B2(n_582), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_171), .A2(n_198), .B1(n_964), .B2(n_965), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g1208 ( .A1(n_173), .A2(n_357), .B1(n_615), .B2(n_731), .C(n_1209), .Y(n_1208) );
AOI22xp33_ASAP7_75t_SL g824 ( .A1(n_174), .A2(n_301), .B1(n_572), .B2(n_633), .Y(n_824) );
NAND2xp5_ASAP7_75t_SL g1140 ( .A(n_175), .B(n_688), .Y(n_1140) );
AO22x2_ASAP7_75t_L g424 ( .A1(n_178), .A2(n_258), .B1(n_425), .B2(n_426), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g1162 ( .A(n_178), .B(n_1163), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_179), .B(n_775), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g1025 ( .A(n_181), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_182), .A2(n_212), .B1(n_438), .B2(n_703), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_183), .A2(n_194), .B1(n_465), .B2(n_698), .Y(n_1068) );
AOI22xp33_ASAP7_75t_SL g1147 ( .A1(n_184), .A2(n_278), .B1(n_588), .B2(n_735), .Y(n_1147) );
CKINVDCx20_ASAP7_75t_R g1190 ( .A(n_185), .Y(n_1190) );
AOI211xp5_ASAP7_75t_L g1169 ( .A1(n_187), .A2(n_570), .B(n_1170), .C(n_1175), .Y(n_1169) );
AOI22xp33_ASAP7_75t_SL g1136 ( .A1(n_189), .A2(n_289), .B1(n_494), .B2(n_523), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_191), .A2(n_199), .B1(n_606), .B2(n_607), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g900 ( .A(n_192), .Y(n_900) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_193), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_195), .Y(n_644) );
CKINVDCx20_ASAP7_75t_R g1177 ( .A(n_197), .Y(n_1177) );
CKINVDCx20_ASAP7_75t_R g515 ( .A(n_201), .Y(n_515) );
AOI22xp33_ASAP7_75t_SL g908 ( .A1(n_202), .A2(n_242), .B1(n_456), .B2(n_703), .Y(n_908) );
AOI22xp33_ASAP7_75t_SL g1146 ( .A1(n_203), .A2(n_218), .B1(n_441), .B2(n_456), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_205), .A2(n_244), .B1(n_726), .B2(n_727), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_206), .A2(n_1052), .B1(n_1074), .B2(n_1075), .Y(n_1051) );
INVx1_ASAP7_75t_L g1074 ( .A(n_206), .Y(n_1074) );
AOI22xp33_ASAP7_75t_SL g737 ( .A1(n_207), .A2(n_379), .B1(n_582), .B2(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g715 ( .A(n_208), .Y(n_715) );
CKINVDCx20_ASAP7_75t_R g1096 ( .A(n_210), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_211), .A2(n_340), .B1(n_461), .B2(n_465), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_213), .B(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g932 ( .A(n_214), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g1050 ( .A(n_215), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_216), .A2(n_384), .B1(n_545), .B2(n_546), .Y(n_1040) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_217), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_219), .A2(n_313), .B1(n_546), .B2(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_221), .A2(n_323), .B1(n_453), .B2(n_661), .Y(n_911) );
AOI22xp33_ASAP7_75t_SL g1143 ( .A1(n_223), .A2(n_374), .B1(n_698), .B2(n_794), .Y(n_1143) );
CKINVDCx20_ASAP7_75t_R g1042 ( .A(n_224), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_225), .B(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_227), .A2(n_275), .B1(n_534), .B2(n_536), .Y(n_833) );
CKINVDCx20_ASAP7_75t_R g925 ( .A(n_228), .Y(n_925) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_229), .Y(n_475) );
CKINVDCx20_ASAP7_75t_R g1007 ( .A(n_230), .Y(n_1007) );
CKINVDCx20_ASAP7_75t_R g978 ( .A(n_232), .Y(n_978) );
AOI211xp5_ASAP7_75t_L g398 ( .A1(n_234), .A2(n_399), .B(n_407), .C(n_1166), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_235), .A2(n_240), .B1(n_494), .B2(n_647), .Y(n_646) );
XNOR2x2_ASAP7_75t_L g602 ( .A(n_236), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g1201 ( .A(n_237), .Y(n_1201) );
AOI22xp5_ASAP7_75t_L g1204 ( .A1(n_237), .A2(n_1201), .B1(n_1205), .B2(n_1206), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_239), .A2(n_273), .B1(n_441), .B2(n_446), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_245), .A2(n_350), .B1(n_545), .B2(n_546), .Y(n_739) );
OA22x2_ASAP7_75t_L g841 ( .A1(n_247), .A2(n_842), .B1(n_843), .B2(n_861), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_247), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_248), .A2(n_390), .B1(n_618), .B2(n_619), .Y(n_617) );
CKINVDCx20_ASAP7_75t_R g813 ( .A(n_249), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g1138 ( .A(n_250), .B(n_1139), .Y(n_1138) );
XNOR2x2_ASAP7_75t_L g1107 ( .A(n_252), .B(n_1108), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_253), .A2(n_382), .B1(n_538), .B2(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g405 ( .A(n_255), .B(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_256), .A2(n_415), .B1(n_509), .B2(n_510), .Y(n_414) );
INVx1_ASAP7_75t_L g509 ( .A(n_256), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_259), .A2(n_272), .B1(n_665), .B2(n_666), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g904 ( .A(n_261), .B(n_727), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_262), .Y(n_771) );
AOI22xp33_ASAP7_75t_SL g879 ( .A1(n_264), .A2(n_295), .B1(n_524), .B2(n_686), .Y(n_879) );
AOI22xp33_ASAP7_75t_SL g839 ( .A1(n_265), .A2(n_393), .B1(n_438), .B2(n_538), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g1114 ( .A(n_267), .Y(n_1114) );
AOI22xp33_ASAP7_75t_SL g837 ( .A1(n_268), .A2(n_388), .B1(n_607), .B2(n_838), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_271), .A2(n_368), .B1(n_629), .B2(n_633), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_274), .A2(n_1168), .B1(n_1192), .B2(n_1193), .Y(n_1167) );
CKINVDCx20_ASAP7_75t_R g1192 ( .A(n_274), .Y(n_1192) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_276), .Y(n_795) );
CKINVDCx20_ASAP7_75t_R g1088 ( .A(n_277), .Y(n_1088) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_281), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g984 ( .A(n_282), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_284), .A2(n_327), .B1(n_453), .B2(n_455), .Y(n_994) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_285), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_286), .A2(n_389), .B1(n_588), .B2(n_591), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_287), .B(n_957), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_288), .A2(n_371), .B1(n_619), .B2(n_790), .Y(n_789) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_290), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g846 ( .A(n_291), .Y(n_846) );
OA22x2_ASAP7_75t_L g870 ( .A1(n_296), .A2(n_871), .B1(n_872), .B2(n_893), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_296), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_297), .B(n_623), .Y(n_622) );
OA22x2_ASAP7_75t_L g672 ( .A1(n_298), .A2(n_673), .B1(n_674), .B2(n_705), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_298), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_300), .A2(n_326), .B1(n_941), .B2(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g425 ( .A(n_302), .Y(n_425) );
INVx1_ASAP7_75t_L g427 ( .A(n_302), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_303), .A2(n_387), .B1(n_534), .B2(n_668), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_304), .Y(n_577) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_306), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g1028 ( .A(n_307), .Y(n_1028) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_310), .Y(n_767) );
CKINVDCx20_ASAP7_75t_R g1217 ( .A(n_311), .Y(n_1217) );
CKINVDCx20_ASAP7_75t_R g1189 ( .A(n_312), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1090 ( .A1(n_316), .A2(n_336), .B1(n_666), .B2(n_1091), .C(n_1094), .Y(n_1090) );
CKINVDCx20_ASAP7_75t_R g977 ( .A(n_317), .Y(n_977) );
CKINVDCx20_ASAP7_75t_R g943 ( .A(n_318), .Y(n_943) );
CKINVDCx20_ASAP7_75t_R g1022 ( .A(n_319), .Y(n_1022) );
CKINVDCx20_ASAP7_75t_R g678 ( .A(n_320), .Y(n_678) );
INVx1_ASAP7_75t_L g471 ( .A(n_321), .Y(n_471) );
INVx1_ASAP7_75t_L g765 ( .A(n_325), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g1043 ( .A(n_328), .B(n_957), .Y(n_1043) );
CKINVDCx20_ASAP7_75t_R g563 ( .A(n_330), .Y(n_563) );
AOI22xp33_ASAP7_75t_SL g968 ( .A1(n_331), .A2(n_381), .B1(n_541), .B2(n_543), .Y(n_968) );
AOI22xp33_ASAP7_75t_L g1067 ( .A1(n_335), .A2(n_355), .B1(n_419), .B2(n_443), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_338), .A2(n_373), .B1(n_536), .B2(n_538), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g1060 ( .A(n_339), .Y(n_1060) );
INVx1_ASAP7_75t_L g406 ( .A(n_341), .Y(n_406) );
INVx1_ASAP7_75t_L g1064 ( .A(n_342), .Y(n_1064) );
CKINVDCx20_ASAP7_75t_R g980 ( .A(n_344), .Y(n_980) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_345), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g1148 ( .A(n_346), .Y(n_1148) );
INVx1_ASAP7_75t_L g402 ( .A(n_347), .Y(n_402) );
CKINVDCx20_ASAP7_75t_R g1118 ( .A(n_348), .Y(n_1118) );
CKINVDCx20_ASAP7_75t_R g1095 ( .A(n_351), .Y(n_1095) );
OA22x2_ASAP7_75t_L g818 ( .A1(n_353), .A2(n_819), .B1(n_820), .B2(n_840), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_353), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_354), .B(n_623), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g800 ( .A(n_360), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g1119 ( .A(n_361), .Y(n_1119) );
CKINVDCx20_ASAP7_75t_R g1004 ( .A(n_362), .Y(n_1004) );
CKINVDCx20_ASAP7_75t_R g1176 ( .A(n_363), .Y(n_1176) );
CKINVDCx20_ASAP7_75t_R g953 ( .A(n_365), .Y(n_953) );
CKINVDCx20_ASAP7_75t_R g981 ( .A(n_366), .Y(n_981) );
INVx1_ASAP7_75t_L g669 ( .A(n_367), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_369), .B(n_719), .Y(n_923) );
CKINVDCx20_ASAP7_75t_R g778 ( .A(n_370), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_372), .Y(n_650) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_375), .Y(n_568) );
CKINVDCx20_ASAP7_75t_R g1014 ( .A(n_376), .Y(n_1014) );
INVx1_ASAP7_75t_L g547 ( .A(n_380), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g971 ( .A(n_383), .Y(n_971) );
INVx1_ASAP7_75t_L g1212 ( .A(n_385), .Y(n_1212) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_386), .B(n_494), .Y(n_1061) );
OA22x2_ASAP7_75t_SL g972 ( .A1(n_392), .A2(n_973), .B1(n_974), .B2(n_996), .Y(n_972) );
INVx1_ASAP7_75t_L g996 ( .A(n_392), .Y(n_996) );
CKINVDCx20_ASAP7_75t_R g1218 ( .A(n_394), .Y(n_1218) );
CKINVDCx20_ASAP7_75t_R g1055 ( .A(n_395), .Y(n_1055) );
CKINVDCx20_ASAP7_75t_R g1059 ( .A(n_397), .Y(n_1059) );
INVx1_ASAP7_75t_SL g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
HB1xp67_ASAP7_75t_L g1157 ( .A(n_402), .Y(n_1157) );
OAI21xp5_ASAP7_75t_L g1199 ( .A1(n_403), .A2(n_1156), .B(n_1200), .Y(n_1199) );
CKINVDCx20_ASAP7_75t_R g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_998), .B1(n_1151), .B2(n_1152), .C(n_1153), .Y(n_407) );
INVx1_ASAP7_75t_L g1151 ( .A(n_408), .Y(n_1151) );
XNOR2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_746), .Y(n_408) );
AOI22xp5_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_549), .B2(n_745), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_511), .B2(n_548), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g510 ( .A(n_415), .Y(n_510) );
AND2x2_ASAP7_75t_SL g415 ( .A(n_416), .B(n_469), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_450), .Y(n_416) );
NAND2xp33_ASAP7_75t_SL g417 ( .A(n_418), .B(n_440), .Y(n_417) );
BUFx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_420), .Y(n_615) );
INVx3_ASAP7_75t_L g696 ( .A(n_420), .Y(n_696) );
BUFx3_ASAP7_75t_L g760 ( .A(n_420), .Y(n_760) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx2_ASAP7_75t_L g537 ( .A(n_421), .Y(n_537) );
BUFx2_ASAP7_75t_SL g588 ( .A(n_421), .Y(n_588) );
BUFx2_ASAP7_75t_SL g734 ( .A(n_421), .Y(n_734) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_431), .Y(n_421) );
AND2x6_ASAP7_75t_L g443 ( .A(n_422), .B(n_444), .Y(n_443) );
AND2x4_ASAP7_75t_L g453 ( .A(n_422), .B(n_454), .Y(n_453) );
AND2x6_ASAP7_75t_L g482 ( .A(n_422), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_428), .Y(n_422) );
AND2x2_ASAP7_75t_L g439 ( .A(n_423), .B(n_429), .Y(n_439) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_424), .B(n_429), .Y(n_449) );
AND2x2_ASAP7_75t_L g458 ( .A(n_424), .B(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g490 ( .A(n_424), .B(n_433), .Y(n_490) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g430 ( .A(n_427), .Y(n_430) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g459 ( .A(n_429), .Y(n_459) );
INVx1_ASAP7_75t_L g489 ( .A(n_429), .Y(n_489) );
AND2x4_ASAP7_75t_L g438 ( .A(n_431), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g447 ( .A(n_431), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g457 ( .A(n_431), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_431), .B(n_458), .Y(n_600) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
OR2x2_ASAP7_75t_L g445 ( .A(n_432), .B(n_435), .Y(n_445) );
AND2x2_ASAP7_75t_L g454 ( .A(n_432), .B(n_435), .Y(n_454) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g483 ( .A(n_433), .B(n_435), .Y(n_483) );
AND2x2_ASAP7_75t_L g488 ( .A(n_434), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g501 ( .A(n_434), .Y(n_501) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g468 ( .A(n_435), .Y(n_468) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g1188 ( .A1(n_437), .A2(n_1189), .B1(n_1190), .B2(n_1191), .Y(n_1188) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
BUFx3_ASAP7_75t_L g545 ( .A(n_438), .Y(n_545) );
BUFx3_ASAP7_75t_L g584 ( .A(n_438), .Y(n_584) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_438), .Y(n_611) );
BUFx3_ASAP7_75t_L g941 ( .A(n_438), .Y(n_941) );
INVx1_ASAP7_75t_L g474 ( .A(n_439), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g477 ( .A(n_439), .B(n_454), .Y(n_477) );
AND2x4_ASAP7_75t_L g625 ( .A(n_439), .B(n_444), .Y(n_625) );
AND2x6_ASAP7_75t_L g691 ( .A(n_439), .B(n_454), .Y(n_691) );
INVx4_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_SL g665 ( .A(n_442), .Y(n_665) );
INVx3_ASAP7_75t_L g731 ( .A(n_442), .Y(n_731) );
INVx4_ASAP7_75t_L g838 ( .A(n_442), .Y(n_838) );
OAI21xp33_ASAP7_75t_SL g848 ( .A1(n_442), .A2(n_849), .B(n_850), .Y(n_848) );
INVx11_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx11_ASAP7_75t_L g595 ( .A(n_443), .Y(n_595) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g473 ( .A(n_445), .B(n_474), .Y(n_473) );
INVxp67_ASAP7_75t_L g801 ( .A(n_446), .Y(n_801) );
BUFx3_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx2_ASAP7_75t_L g538 ( .A(n_447), .Y(n_538) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_447), .Y(n_591) );
BUFx3_ASAP7_75t_L g612 ( .A(n_447), .Y(n_612) );
BUFx2_ASAP7_75t_SL g735 ( .A(n_447), .Y(n_735) );
BUFx3_ASAP7_75t_L g757 ( .A(n_447), .Y(n_757) );
BUFx3_ASAP7_75t_L g992 ( .A(n_447), .Y(n_992) );
AND2x2_ASAP7_75t_L g970 ( .A(n_448), .B(n_501), .Y(n_970) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
OR2x6_ASAP7_75t_L g467 ( .A(n_449), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
BUFx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx6_ASAP7_75t_L g542 ( .A(n_453), .Y(n_542) );
BUFx3_ASAP7_75t_L g668 ( .A(n_453), .Y(n_668) );
BUFx3_ASAP7_75t_L g1012 ( .A(n_453), .Y(n_1012) );
AND2x2_ASAP7_75t_L g464 ( .A(n_454), .B(n_458), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g1087 ( .A(n_454), .B(n_458), .Y(n_1087) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g534 ( .A(n_457), .Y(n_534) );
BUFx3_ASAP7_75t_L g616 ( .A(n_457), .Y(n_616) );
BUFx3_ASAP7_75t_L g965 ( .A(n_457), .Y(n_965) );
INVx1_ASAP7_75t_L g508 ( .A(n_459), .Y(n_508) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx2_ASAP7_75t_L g1016 ( .A(n_462), .Y(n_1016) );
INVx5_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx3_ASAP7_75t_L g543 ( .A(n_463), .Y(n_543) );
INVx1_ASAP7_75t_L g582 ( .A(n_463), .Y(n_582) );
INVx2_ASAP7_75t_L g618 ( .A(n_463), .Y(n_618) );
INVx4_ASAP7_75t_L g661 ( .A(n_463), .Y(n_661) );
BUFx3_ASAP7_75t_L g699 ( .A(n_463), .Y(n_699) );
INVx8_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g1214 ( .A(n_465), .Y(n_1214) );
BUFx4f_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
BUFx2_ASAP7_75t_L g546 ( .A(n_466), .Y(n_546) );
BUFx2_ASAP7_75t_L g619 ( .A(n_466), .Y(n_619) );
BUFx2_ASAP7_75t_L g888 ( .A(n_466), .Y(n_888) );
BUFx2_ASAP7_75t_L g942 ( .A(n_466), .Y(n_942) );
INVx6_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g662 ( .A(n_467), .Y(n_662) );
INVx1_ASAP7_75t_SL g700 ( .A(n_467), .Y(n_700) );
INVx1_ASAP7_75t_SL g835 ( .A(n_467), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g851 ( .A1(n_467), .A2(n_505), .B1(n_852), .B2(n_853), .Y(n_851) );
INVx1_ASAP7_75t_L g630 ( .A(n_468), .Y(n_630) );
NOR3xp33_ASAP7_75t_L g469 ( .A(n_470), .B(n_478), .C(n_497), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_475), .B2(n_476), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_472), .A2(n_812), .B1(n_813), .B2(n_814), .Y(n_811) );
INVx1_ASAP7_75t_L g927 ( .A(n_472), .Y(n_927) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx3_ASAP7_75t_L g516 ( .A(n_473), .Y(n_516) );
INVx2_ASAP7_75t_L g562 ( .A(n_473), .Y(n_562) );
INVx2_ASAP7_75t_L g565 ( .A(n_476), .Y(n_565) );
BUFx3_ASAP7_75t_L g1172 ( .A(n_476), .Y(n_1172) );
BUFx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g519 ( .A(n_477), .Y(n_519) );
OAI221xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_484), .B1(n_485), .B2(n_491), .C(n_492), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_479), .A2(n_715), .B(n_716), .Y(n_714) );
OAI221xp5_ASAP7_75t_L g806 ( .A1(n_479), .A2(n_772), .B1(n_807), .B2(n_808), .C(n_809), .Y(n_806) );
OAI221xp5_ASAP7_75t_L g979 ( .A1(n_479), .A2(n_677), .B1(n_980), .B2(n_981), .C(n_982), .Y(n_979) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx4_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI21xp5_ASAP7_75t_SL g520 ( .A1(n_481), .A2(n_521), .B(n_522), .Y(n_520) );
BUFx2_ASAP7_75t_L g645 ( .A(n_481), .Y(n_645) );
INVx4_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx3_ASAP7_75t_L g570 ( .A(n_482), .Y(n_570) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_482), .Y(n_680) );
INVx2_ASAP7_75t_SL g770 ( .A(n_482), .Y(n_770) );
INVx2_ASAP7_75t_L g875 ( .A(n_482), .Y(n_875) );
INVx2_ASAP7_75t_L g1058 ( .A(n_482), .Y(n_1058) );
INVx1_ASAP7_75t_L g506 ( .A(n_483), .Y(n_506) );
AND2x4_ASAP7_75t_L g524 ( .A(n_483), .B(n_508), .Y(n_524) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_487), .Y(n_529) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_487), .Y(n_576) );
BUFx4f_ASAP7_75t_SL g633 ( .A(n_487), .Y(n_633) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_487), .Y(n_648) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g496 ( .A(n_489), .Y(n_496) );
AND2x4_ASAP7_75t_L g495 ( .A(n_490), .B(n_496), .Y(n_495) );
NAND2x1p5_ASAP7_75t_L g500 ( .A(n_490), .B(n_501), .Y(n_500) );
AND2x4_ASAP7_75t_L g629 ( .A(n_490), .B(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g1024 ( .A(n_493), .Y(n_1024) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g776 ( .A(n_494), .Y(n_776) );
BUFx2_ASAP7_75t_L g810 ( .A(n_494), .Y(n_810) );
BUFx6f_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx12f_ASAP7_75t_L g572 ( .A(n_495), .Y(n_572) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_495), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_498), .A2(n_499), .B1(n_502), .B2(n_503), .Y(n_497) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_500), .A2(n_526), .B1(n_527), .B2(n_530), .Y(n_525) );
BUFx3_ASAP7_75t_L g578 ( .A(n_500), .Y(n_578) );
INVx4_ASAP7_75t_L g652 ( .A(n_500), .Y(n_652) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_500), .A2(n_654), .B1(n_804), .B2(n_805), .Y(n_803) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_500), .A2(n_654), .B1(n_1217), .B2(n_1218), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_503), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g1026 ( .A1(n_503), .A2(n_779), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
OAI22xp5_ASAP7_75t_L g1099 ( .A1(n_503), .A2(n_779), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g654 ( .A(n_504), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g986 ( .A(n_505), .Y(n_986) );
OR2x6_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g548 ( .A(n_511), .Y(n_548) );
OA22x2_ASAP7_75t_L g708 ( .A1(n_511), .A2(n_709), .B1(n_710), .B2(n_741), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_511), .Y(n_709) );
XOR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_547), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_513), .B(n_531), .Y(n_512) );
NOR3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_520), .C(n_525), .Y(n_513) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B1(n_517), .B2(n_518), .Y(n_514) );
OAI22xp5_ASAP7_75t_L g845 ( .A1(n_516), .A2(n_768), .B1(n_846), .B2(n_847), .Y(n_845) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_516), .A2(n_564), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
OA211x2_ASAP7_75t_L g620 ( .A1(n_518), .A2(n_621), .B(n_622), .C(n_626), .Y(n_620) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_SL g768 ( .A(n_519), .Y(n_768) );
INVx2_ASAP7_75t_L g814 ( .A(n_519), .Y(n_814) );
BUFx2_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_SL g631 ( .A(n_524), .Y(n_631) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_524), .Y(n_721) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_527), .A2(n_1058), .B1(n_1059), .B2(n_1060), .C(n_1061), .Y(n_1057) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_SL g772 ( .A(n_528), .Y(n_772) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g931 ( .A(n_529), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g531 ( .A(n_532), .B(n_539), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_533), .B(n_535), .Y(n_532) );
BUFx2_ASAP7_75t_L g754 ( .A(n_534), .Y(n_754) );
INVx1_ASAP7_75t_L g1072 ( .A(n_534), .Y(n_1072) );
INVx3_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx3_ASAP7_75t_L g937 ( .A(n_537), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
INVxp67_ASAP7_75t_L g1186 ( .A(n_541), .Y(n_1186) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g607 ( .A(n_542), .Y(n_607) );
INVx2_ASAP7_75t_L g738 ( .A(n_542), .Y(n_738) );
INVx2_ASAP7_75t_L g794 ( .A(n_542), .Y(n_794) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_542), .A2(n_598), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
HB1xp67_ASAP7_75t_L g1006 ( .A(n_545), .Y(n_1006) );
INVx1_ASAP7_75t_L g745 ( .A(n_549), .Y(n_745) );
XOR2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_671), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B1(n_636), .B2(n_670), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B1(n_601), .B2(n_602), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_555), .A2(n_707), .B1(n_708), .B2(n_742), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_555), .Y(n_707) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_579), .Y(n_558) );
NOR3xp33_ASAP7_75t_L g559 ( .A(n_560), .B(n_567), .C(n_573), .Y(n_559) );
OAI22xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_563), .B1(n_564), .B2(n_566), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_SL g641 ( .A(n_562), .Y(n_641) );
INVx2_ASAP7_75t_L g766 ( .A(n_562), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_564), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_564), .A2(n_925), .B1(n_926), .B2(n_928), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g976 ( .A1(n_564), .A2(n_766), .B1(n_977), .B2(n_978), .Y(n_976) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_564), .A2(n_926), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI21xp33_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B(n_571), .Y(n_567) );
OAI21xp5_ASAP7_75t_SL g822 ( .A1(n_569), .A2(n_823), .B(n_824), .Y(n_822) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g718 ( .A(n_572), .Y(n_718) );
BUFx4f_ASAP7_75t_SL g1049 ( .A(n_572), .Y(n_1049) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_575), .B1(n_577), .B2(n_578), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_576), .Y(n_575) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_578), .A2(n_930), .B1(n_931), .B2(n_932), .Y(n_929) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .C(n_592), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_583), .Y(n_580) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_582), .Y(n_790) );
INVx1_ASAP7_75t_L g799 ( .A(n_584), .Y(n_799) );
BUFx2_ASAP7_75t_L g990 ( .A(n_584), .Y(n_990) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_589), .B2(n_590), .Y(n_585) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g590 ( .A(n_591), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_596), .B1(n_597), .B2(n_598), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g606 ( .A(n_595), .Y(n_606) );
INVx5_ASAP7_75t_SL g703 ( .A(n_595), .Y(n_703) );
HB1xp67_ASAP7_75t_L g885 ( .A(n_595), .Y(n_885) );
INVx4_ASAP7_75t_L g964 ( .A(n_595), .Y(n_964) );
INVx2_ASAP7_75t_SL g1093 ( .A(n_595), .Y(n_1093) );
OAI221xp5_ASAP7_75t_SL g1010 ( .A1(n_598), .A2(n_1011), .B1(n_1013), .B2(n_1014), .C(n_1015), .Y(n_1010) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_598), .A2(n_1011), .B1(n_1095), .B2(n_1096), .Y(n_1094) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g796 ( .A(n_599), .Y(n_796) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND4xp75_ASAP7_75t_L g603 ( .A(n_604), .B(n_613), .C(n_620), .D(n_632), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_608), .Y(n_604) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx4_ASAP7_75t_L g666 ( .A(n_610), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_610), .A2(n_1114), .B1(n_1115), .B2(n_1116), .Y(n_1113) );
INVx4_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
HB1xp67_ASAP7_75t_L g1009 ( .A(n_612), .Y(n_1009) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_617), .Y(n_613) );
BUFx4f_ASAP7_75t_SL g732 ( .A(n_616), .Y(n_732) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_618), .Y(n_887) );
INVx1_ASAP7_75t_L g1089 ( .A(n_619), .Y(n_1089) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_623), .Y(n_688) );
INVx5_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx2_ASAP7_75t_L g726 ( .A(n_624), .Y(n_726) );
INVx2_ASAP7_75t_L g881 ( .A(n_624), .Y(n_881) );
INVx2_ASAP7_75t_L g957 ( .A(n_624), .Y(n_957) );
INVx4_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g1128 ( .A(n_628), .Y(n_1128) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
BUFx2_ASAP7_75t_L g686 ( .A(n_629), .Y(n_686) );
BUFx2_ASAP7_75t_L g724 ( .A(n_629), .Y(n_724) );
BUFx3_ASAP7_75t_L g830 ( .A(n_629), .Y(n_830) );
INVx1_ASAP7_75t_L g682 ( .A(n_634), .Y(n_682) );
BUFx4f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g921 ( .A(n_635), .Y(n_921) );
INVx1_ASAP7_75t_L g670 ( .A(n_636), .Y(n_670) );
XOR2x2_ASAP7_75t_L g636 ( .A(n_637), .B(n_669), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_655), .Y(n_637) );
NOR3xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_643), .C(n_649), .Y(n_638) );
OAI21xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_646), .Y(n_643) );
BUFx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g677 ( .A(n_648), .Y(n_677) );
INVx4_ASAP7_75t_L g1125 ( .A(n_648), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_653), .B2(n_654), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_651), .A2(n_986), .B1(n_1063), .B2(n_1064), .Y(n_1062) );
INVx3_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g779 ( .A(n_652), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_663), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_661), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_667), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_706), .B1(n_743), .B2(n_744), .Y(n_671) );
INVx1_ASAP7_75t_L g743 ( .A(n_672), .Y(n_743) );
INVx1_ASAP7_75t_SL g705 ( .A(n_674), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_675), .B(n_692), .Y(n_674) );
NOR2x1_ASAP7_75t_L g675 ( .A(n_676), .B(n_684), .Y(n_675) );
OAI222xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_678), .B1(n_679), .B2(n_681), .C1(n_682), .C2(n_683), .Y(n_676) );
OAI222xp33_ASAP7_75t_L g1021 ( .A1(n_679), .A2(n_772), .B1(n_1022), .B2(n_1023), .C1(n_1024), .C2(n_1025), .Y(n_1021) );
INVx2_ASAP7_75t_SL g679 ( .A(n_680), .Y(n_679) );
INVx2_ASAP7_75t_L g919 ( .A(n_680), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx1_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_SL g827 ( .A(n_690), .Y(n_827) );
INVx1_ASAP7_75t_SL g690 ( .A(n_691), .Y(n_690) );
BUFx2_ASAP7_75t_L g727 ( .A(n_691), .Y(n_727) );
BUFx4f_ASAP7_75t_L g959 ( .A(n_691), .Y(n_959) );
BUFx2_ASAP7_75t_L g1139 ( .A(n_691), .Y(n_1139) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_701), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_694), .B(n_697), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OAI221xp5_ASAP7_75t_SL g1003 ( .A1(n_696), .A2(n_1004), .B1(n_1005), .B2(n_1007), .C(n_1008), .Y(n_1003) );
INVx3_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g1115 ( .A(n_703), .Y(n_1115) );
HB1xp67_ASAP7_75t_L g1182 ( .A(n_703), .Y(n_1182) );
INVx1_ASAP7_75t_L g744 ( .A(n_706), .Y(n_744) );
INVx1_ASAP7_75t_L g742 ( .A(n_708), .Y(n_742) );
INVx1_ASAP7_75t_L g741 ( .A(n_710), .Y(n_741) );
INVx1_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_713), .B(n_728), .Y(n_712) );
NOR2xp33_ASAP7_75t_L g713 ( .A(n_714), .B(n_722), .Y(n_713) );
INVx1_ASAP7_75t_L g1178 ( .A(n_717), .Y(n_1178) );
INVx3_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_723), .B(n_725), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_736), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_737), .B(n_739), .Y(n_736) );
XOR2xp5_ASAP7_75t_L g746 ( .A(n_747), .B(n_866), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_783), .B1(n_864), .B2(n_865), .Y(n_747) );
INVx2_ASAP7_75t_L g864 ( .A(n_748), .Y(n_864) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g782 ( .A(n_750), .Y(n_782) );
AND2x2_ASAP7_75t_SL g750 ( .A(n_751), .B(n_763), .Y(n_750) );
NOR2xp33_ASAP7_75t_SL g751 ( .A(n_752), .B(n_758), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_755), .Y(n_752) );
INVx1_ASAP7_75t_L g1191 ( .A(n_756), .Y(n_1191) );
BUFx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
NOR3xp33_ASAP7_75t_L g763 ( .A(n_764), .B(n_769), .C(n_777), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .B1(n_767), .B2(n_768), .Y(n_764) );
OA211x2_ASAP7_75t_L g1041 ( .A1(n_768), .A2(n_1042), .B(n_1043), .C(n_1044), .Y(n_1041) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_771), .B1(n_772), .B2(n_773), .C(n_774), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_772), .A2(n_1176), .B1(n_1177), .B2(n_1178), .Y(n_1175) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_779), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
INVx2_ASAP7_75t_SL g865 ( .A(n_783), .Y(n_865) );
OA22x2_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_817), .B1(n_862), .B2(n_863), .Y(n_783) );
INVx1_ASAP7_75t_L g862 ( .A(n_784), .Y(n_862) );
INVx1_ASAP7_75t_L g816 ( .A(n_785), .Y(n_816) );
AND2x2_ASAP7_75t_SL g785 ( .A(n_786), .B(n_802), .Y(n_785) );
NOR3xp33_ASAP7_75t_L g786 ( .A(n_787), .B(n_791), .C(n_797), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_793), .B1(n_795), .B2(n_796), .Y(n_791) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g1184 ( .A1(n_796), .A2(n_1185), .B1(n_1186), .B2(n_1187), .Y(n_1184) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_800), .B2(n_801), .Y(n_797) );
INVx1_ASAP7_75t_L g891 ( .A(n_799), .Y(n_891) );
NOR3xp33_ASAP7_75t_SL g802 ( .A(n_803), .B(n_806), .C(n_811), .Y(n_802) );
INVx1_ASAP7_75t_L g863 ( .A(n_817), .Y(n_863) );
XOR2x2_ASAP7_75t_L g817 ( .A(n_818), .B(n_841), .Y(n_817) );
INVx1_ASAP7_75t_L g840 ( .A(n_820), .Y(n_840) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_831), .Y(n_820) );
NOR2xp67_ASAP7_75t_L g821 ( .A(n_822), .B(n_825), .Y(n_821) );
NAND3xp33_ASAP7_75t_L g825 ( .A(n_826), .B(n_828), .C(n_829), .Y(n_825) );
NOR2x1_ASAP7_75t_L g831 ( .A(n_832), .B(n_836), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_839), .Y(n_836) );
INVx2_ASAP7_75t_L g861 ( .A(n_843), .Y(n_861) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_854), .Y(n_843) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_848), .C(n_851), .Y(n_844) );
NOR2xp33_ASAP7_75t_L g854 ( .A(n_855), .B(n_858), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g855 ( .A(n_856), .B(n_857), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g858 ( .A(n_859), .B(n_860), .Y(n_858) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_945), .B1(n_946), .B2(n_997), .Y(n_867) );
INVx1_ASAP7_75t_L g997 ( .A(n_868), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g868 ( .A1(n_869), .A2(n_870), .B1(n_894), .B2(n_895), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_SL g893 ( .A(n_872), .Y(n_893) );
NAND3x1_ASAP7_75t_L g872 ( .A(n_873), .B(n_882), .C(n_889), .Y(n_872) );
NOR2xp33_ASAP7_75t_L g873 ( .A(n_874), .B(n_878), .Y(n_873) );
OAI21xp5_ASAP7_75t_SL g874 ( .A1(n_875), .A2(n_876), .B(n_877), .Y(n_874) );
OAI21xp5_ASAP7_75t_SL g899 ( .A1(n_875), .A2(n_900), .B(n_901), .Y(n_899) );
OAI21xp5_ASAP7_75t_SL g1121 ( .A1(n_875), .A2(n_1122), .B(n_1123), .Y(n_1121) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_881), .Y(n_1098) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_886), .Y(n_882) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
AND2x2_ASAP7_75t_L g889 ( .A(n_890), .B(n_892), .Y(n_889) );
INVx2_ASAP7_75t_SL g894 ( .A(n_895), .Y(n_894) );
AO22x2_ASAP7_75t_SL g895 ( .A1(n_896), .A2(n_914), .B1(n_915), .B2(n_944), .Y(n_895) );
INVx3_ASAP7_75t_L g944 ( .A(n_896), .Y(n_944) );
OAI22x1_ASAP7_75t_L g947 ( .A1(n_896), .A2(n_944), .B1(n_948), .B2(n_949), .Y(n_947) );
XOR2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_913), .Y(n_896) );
NAND2x1_ASAP7_75t_SL g897 ( .A(n_898), .B(n_906), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_902), .Y(n_898) );
NAND3xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_904), .C(n_905), .Y(n_902) );
NOR2x1_ASAP7_75t_L g906 ( .A(n_907), .B(n_910), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_908), .B(n_909), .Y(n_907) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_911), .B(n_912), .Y(n_910) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
XOR2x2_ASAP7_75t_L g915 ( .A(n_916), .B(n_943), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_917), .B(n_933), .Y(n_916) );
NOR3xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_924), .C(n_929), .Y(n_917) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_919), .A2(n_920), .B1(n_921), .B2(n_922), .C(n_923), .Y(n_918) );
OAI21xp5_ASAP7_75t_L g952 ( .A1(n_919), .A2(n_953), .B(n_954), .Y(n_952) );
INVx2_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g933 ( .A(n_934), .B(n_938), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_935), .B(n_936), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_939), .B(n_940), .Y(n_938) );
INVx2_ASAP7_75t_SL g945 ( .A(n_946), .Y(n_945) );
XNOR2x2_ASAP7_75t_L g946 ( .A(n_947), .B(n_972), .Y(n_946) );
INVx3_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
XOR2x2_ASAP7_75t_L g949 ( .A(n_950), .B(n_971), .Y(n_949) );
NAND2xp5_ASAP7_75t_SL g950 ( .A(n_951), .B(n_961), .Y(n_950) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_952), .B(n_955), .Y(n_951) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_958), .C(n_960), .Y(n_955) );
NOR2x1_ASAP7_75t_L g961 ( .A(n_962), .B(n_967), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_963), .B(n_966), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g967 ( .A(n_968), .B(n_969), .Y(n_967) );
INVx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
AND2x2_ASAP7_75t_SL g974 ( .A(n_975), .B(n_987), .Y(n_974) );
NOR3xp33_ASAP7_75t_L g975 ( .A(n_976), .B(n_979), .C(n_983), .Y(n_975) );
NOR2xp33_ASAP7_75t_L g987 ( .A(n_988), .B(n_993), .Y(n_987) );
NAND2xp5_ASAP7_75t_SL g988 ( .A(n_989), .B(n_991), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_995), .Y(n_993) );
INVx1_ASAP7_75t_L g1152 ( .A(n_998), .Y(n_1152) );
AOI22xp5_ASAP7_75t_L g998 ( .A1(n_999), .A2(n_1078), .B1(n_1079), .B2(n_1150), .Y(n_998) );
INVx1_ASAP7_75t_L g1150 ( .A(n_999), .Y(n_1150) );
AOI22xp5_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1031), .B1(n_1032), .B2(n_1077), .Y(n_999) );
INVx2_ASAP7_75t_L g1077 ( .A(n_1000), .Y(n_1077) );
INVx1_ASAP7_75t_SL g1030 ( .A(n_1001), .Y(n_1030) );
AND2x2_ASAP7_75t_SL g1001 ( .A(n_1002), .B(n_1017), .Y(n_1001) );
NOR2xp33_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1010), .Y(n_1002) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx3_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
NOR3xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1021), .C(n_1026), .Y(n_1017) );
INVx1_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
OAI22xp5_ASAP7_75t_SL g1032 ( .A1(n_1033), .A2(n_1034), .B1(n_1051), .B2(n_1076), .Y(n_1032) );
INVx1_ASAP7_75t_SL g1033 ( .A(n_1034), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
INVx2_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
XOR2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1050), .Y(n_1036) );
NAND4xp75_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1041), .C(n_1045), .D(n_1048), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1040), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1047), .Y(n_1045) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1051), .Y(n_1076) );
INVx2_ASAP7_75t_L g1075 ( .A(n_1052), .Y(n_1075) );
AND2x2_ASAP7_75t_SL g1052 ( .A(n_1053), .B(n_1065), .Y(n_1052) );
NOR3xp33_ASAP7_75t_L g1053 ( .A(n_1054), .B(n_1057), .C(n_1062), .Y(n_1053) );
OAI21xp5_ASAP7_75t_SL g1134 ( .A1(n_1058), .A2(n_1135), .B(n_1136), .Y(n_1134) );
NOR2xp33_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1069), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1066 ( .A(n_1067), .B(n_1068), .Y(n_1066) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1073), .Y(n_1069) );
INVx2_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
OAI22xp5_ASAP7_75t_SL g1079 ( .A1(n_1080), .A2(n_1081), .B1(n_1105), .B2(n_1149), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1082), .Y(n_1104) );
AND4x1_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1090), .C(n_1097), .D(n_1102), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1084 ( .A1(n_1085), .A2(n_1086), .B1(n_1088), .B2(n_1089), .Y(n_1084) );
OAI22xp5_ASAP7_75t_L g1211 ( .A1(n_1086), .A2(n_1212), .B1(n_1213), .B2(n_1214), .Y(n_1211) );
BUFx2_ASAP7_75t_R g1086 ( .A(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
INVx1_ASAP7_75t_L g1092 ( .A(n_1093), .Y(n_1092) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1105), .Y(n_1149) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_1106), .A2(n_1107), .B1(n_1130), .B2(n_1131), .Y(n_1105) );
INVx2_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
NAND2xp5_ASAP7_75t_SL g1108 ( .A(n_1109), .B(n_1120), .Y(n_1108) );
NOR3xp33_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1113), .C(n_1117), .Y(n_1109) );
NAND2xp5_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1112), .Y(n_1110) );
NOR2xp33_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1126), .Y(n_1120) );
INVx3_ASAP7_75t_L g1124 ( .A(n_1125), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1129), .Y(n_1126) );
INVx1_ASAP7_75t_L g1130 ( .A(n_1131), .Y(n_1130) );
XOR2x2_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1148), .Y(n_1131) );
NAND3x1_ASAP7_75t_L g1132 ( .A(n_1133), .B(n_1142), .C(n_1145), .Y(n_1132) );
NOR2xp33_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1137), .Y(n_1133) );
NAND3xp33_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1140), .C(n_1141), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1144), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1146), .B(n_1147), .Y(n_1145) );
INVx1_ASAP7_75t_SL g1153 ( .A(n_1154), .Y(n_1153) );
NOR2x1_ASAP7_75t_L g1154 ( .A(n_1155), .B(n_1159), .Y(n_1154) );
OR2x2_ASAP7_75t_SL g1222 ( .A(n_1155), .B(n_1160), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1158), .Y(n_1155) );
CKINVDCx20_ASAP7_75t_R g1195 ( .A(n_1156), .Y(n_1195) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1157), .B(n_1197), .Y(n_1200) );
CKINVDCx16_ASAP7_75t_R g1197 ( .A(n_1158), .Y(n_1197) );
CKINVDCx20_ASAP7_75t_R g1159 ( .A(n_1160), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1162), .Y(n_1160) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1165), .Y(n_1163) );
OAI322xp33_ASAP7_75t_L g1166 ( .A1(n_1167), .A2(n_1194), .A3(n_1196), .B1(n_1198), .B2(n_1201), .C1(n_1202), .C2(n_1220), .Y(n_1166) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1168), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1179), .Y(n_1168) );
OAI211xp5_ASAP7_75t_L g1170 ( .A1(n_1171), .A2(n_1172), .B(n_1173), .C(n_1174), .Y(n_1170) );
NOR3xp33_ASAP7_75t_L g1179 ( .A(n_1180), .B(n_1184), .C(n_1188), .Y(n_1179) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1181), .B(n_1183), .Y(n_1180) );
HB1xp67_ASAP7_75t_L g1194 ( .A(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
CKINVDCx16_ASAP7_75t_R g1198 ( .A(n_1199), .Y(n_1198) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
INVx2_ASAP7_75t_L g1205 ( .A(n_1206), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
AND4x1_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1210), .C(n_1215), .D(n_1219), .Y(n_1207) );
CKINVDCx20_ASAP7_75t_R g1220 ( .A(n_1221), .Y(n_1220) );
CKINVDCx20_ASAP7_75t_R g1221 ( .A(n_1222), .Y(n_1221) );
endmodule