module fake_netlist_1_5388_n_29 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVxp67_ASAP7_75t_SL g13 ( .A(n_7), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
NOR2xp33_ASAP7_75t_L g15 ( .A(n_0), .B(n_11), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_6), .B(n_10), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
INVx4_ASAP7_75t_L g18 ( .A(n_3), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_0), .Y(n_20) );
INVx1_ASAP7_75t_SL g21 ( .A(n_20), .Y(n_21) );
NAND2xp33_ASAP7_75t_R g22 ( .A(n_21), .B(n_20), .Y(n_22) );
AND2x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_20), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AOI321xp33_ASAP7_75t_L g25 ( .A1(n_24), .A2(n_23), .A3(n_19), .B1(n_15), .B2(n_13), .C(n_16), .Y(n_25) );
NAND5xp2_ASAP7_75t_L g26 ( .A(n_25), .B(n_14), .C(n_2), .D(n_3), .E(n_4), .Y(n_26) );
OAI211xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_14), .B(n_17), .C(n_1), .Y(n_27) );
AOI22xp33_ASAP7_75t_R g28 ( .A1(n_26), .A2(n_1), .B1(n_4), .B2(n_5), .Y(n_28) );
AOI22xp33_ASAP7_75t_SL g29 ( .A1(n_28), .A2(n_27), .B1(n_9), .B2(n_12), .Y(n_29) );
endmodule