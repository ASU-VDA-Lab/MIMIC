module fake_jpeg_10700_n_100 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_45),
.B(n_48),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_1),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_2),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

NAND2x1_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_43),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_57),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_42),
.B1(n_36),
.B2(n_35),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_55),
.B1(n_14),
.B2(n_31),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_36),
.B1(n_35),
.B2(n_34),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_44),
.C(n_17),
.Y(n_57)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_59),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_46),
.A2(n_44),
.B1(n_16),
.B2(n_19),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_62),
.A2(n_54),
.B1(n_60),
.B2(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_6),
.Y(n_71)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_9),
.Y(n_76)
);

A2O1A1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_67)
);

AO22x1_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_68),
.B(n_70),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_3),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_73),
.B(n_72),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_61),
.B(n_4),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_71),
.B(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_64),
.B(n_7),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_78),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_73),
.A2(n_11),
.B(n_13),
.Y(n_78)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_79),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_23),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_29),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_91),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_84),
.B(n_80),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_90),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_85),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_96),
.B(n_75),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_87),
.B1(n_88),
.B2(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_76),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g100 ( 
.A(n_99),
.Y(n_100)
);


endmodule