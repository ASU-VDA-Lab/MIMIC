module fake_jpeg_14414_n_633 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_633);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_633;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_18),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx11_ASAP7_75t_SL g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_4),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_14),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_7),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

NAND2x1_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_1),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_62),
.B(n_26),
.C(n_58),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_64),
.Y(n_183)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_66),
.Y(n_158)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_67),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_20),
.B(n_1),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g188 ( 
.A(n_72),
.Y(n_188)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_73),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_76),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_80),
.Y(n_170)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

BUFx4f_ASAP7_75t_SL g176 ( 
.A(n_81),
.Y(n_176)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_21),
.B(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_123),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_84),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_86),
.Y(n_150)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_87),
.Y(n_160)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

BUFx8_ASAP7_75t_L g190 ( 
.A(n_89),
.Y(n_190)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_91),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_92),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_93),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_94),
.Y(n_157)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_96),
.Y(n_186)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_97),
.Y(n_159)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_31),
.Y(n_98)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_98),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

CKINVDCx9p33_ASAP7_75t_R g133 ( 
.A(n_99),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_46),
.Y(n_100)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_102),
.Y(n_210)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_103),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

CKINVDCx11_ASAP7_75t_R g173 ( 
.A(n_105),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_21),
.B(n_1),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_31),
.Y(n_108)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_108),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

BUFx8_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_110),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_111),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_112),
.Y(n_199)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_113),
.Y(n_201)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_114),
.Y(n_200)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_37),
.Y(n_115)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_116),
.Y(n_203)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_117),
.Y(n_205)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_41),
.Y(n_118)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_118),
.Y(n_206)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_120),
.Y(n_211)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_45),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_122),
.Y(n_137)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_30),
.B(n_2),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_49),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_127),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_37),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_48),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_22),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_60),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_61),
.A2(n_33),
.B1(n_28),
.B2(n_49),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_129),
.A2(n_77),
.B1(n_96),
.B2(n_94),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_138),
.B(n_143),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_70),
.B(n_54),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_54),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_148),
.B(n_156),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_127),
.A2(n_60),
.B1(n_33),
.B2(n_28),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_149),
.A2(n_202),
.B1(n_78),
.B2(n_111),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_155),
.B(n_165),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_43),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_61),
.B(n_24),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_163),
.B(n_168),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_109),
.B(n_43),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_109),
.B(n_38),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_172),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_38),
.Y(n_172)
);

BUFx12_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_102),
.B(n_57),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_180),
.B(n_182),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_24),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_34),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_184),
.B(n_185),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_65),
.B(n_34),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_105),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_191),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_82),
.A2(n_58),
.B1(n_56),
.B2(n_51),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_194),
.A2(n_198),
.B1(n_212),
.B2(n_208),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_116),
.B(n_57),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_196),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_63),
.A2(n_26),
.B1(n_19),
.B2(n_53),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_198),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_68),
.A2(n_56),
.B1(n_51),
.B2(n_53),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_97),
.B(n_53),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_204),
.B(n_3),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_74),
.B(n_53),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_207),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_130),
.B(n_2),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_214),
.B(n_225),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_216),
.A2(n_250),
.B1(n_266),
.B2(n_283),
.Y(n_334)
);

CKINVDCx9p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_218),
.Y(n_316)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_133),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_219),
.Y(n_310)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_220),
.Y(n_323)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_159),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_222),
.Y(n_325)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_223),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_224),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_137),
.B(n_2),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_178),
.Y(n_226)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_226),
.Y(n_313)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_178),
.Y(n_227)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_228),
.Y(n_326)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_229),
.Y(n_300)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_162),
.Y(n_230)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_231),
.Y(n_318)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_232),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_131),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_233),
.B(n_237),
.Y(n_333)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_234),
.Y(n_327)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_139),
.Y(n_235)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_235),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_150),
.A2(n_112),
.B1(n_79),
.B2(n_84),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_236),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_131),
.B(n_2),
.Y(n_237)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g343 ( 
.A(n_239),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_139),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g311 ( 
.A(n_241),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_183),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_243),
.B(n_248),
.Y(n_341)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_164),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_246),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_132),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_165),
.B(n_197),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_249),
.B(n_254),
.Y(n_346)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_150),
.A2(n_93),
.B1(n_92),
.B2(n_85),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_166),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_251),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_173),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_253),
.B(n_280),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_140),
.Y(n_254)
);

CKINVDCx12_ASAP7_75t_R g255 ( 
.A(n_174),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_255),
.B(n_257),
.Y(n_296)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_151),
.Y(n_256)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_256),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_174),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_200),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_258),
.B(n_267),
.Y(n_298)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_145),
.Y(n_259)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

INVx3_ASAP7_75t_SL g260 ( 
.A(n_134),
.Y(n_260)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_260),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_209),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_262),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_136),
.B(n_3),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_263),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_151),
.Y(n_264)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_146),
.A2(n_100),
.B1(n_99),
.B2(n_8),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_194),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_147),
.B(n_3),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_268),
.B(n_278),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_271),
.A2(n_176),
.B(n_158),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_152),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_272),
.B(n_273),
.Y(n_317)
);

CKINVDCx12_ASAP7_75t_R g273 ( 
.A(n_141),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_142),
.Y(n_274)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_142),
.Y(n_275)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_275),
.Y(n_328)
);

CKINVDCx9p33_ASAP7_75t_R g276 ( 
.A(n_141),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g347 ( 
.A(n_276),
.B(n_188),
.Y(n_347)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_190),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_279),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_170),
.B(n_3),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_201),
.Y(n_280)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_210),
.B(n_213),
.Y(n_281)
);

NAND2xp33_ASAP7_75t_SL g301 ( 
.A(n_281),
.B(n_285),
.Y(n_301)
);

CKINVDCx12_ASAP7_75t_R g282 ( 
.A(n_187),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_282),
.B(n_176),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_129),
.A2(n_167),
.B1(n_169),
.B2(n_177),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_179),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_284),
.A2(n_286),
.B1(n_288),
.B2(n_187),
.Y(n_291)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_181),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_167),
.A2(n_169),
.B1(n_177),
.B2(n_210),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_287),
.A2(n_153),
.B1(n_186),
.B2(n_157),
.Y(n_307)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_179),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_291),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_271),
.A2(n_242),
.B1(n_218),
.B2(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_302),
.A2(n_260),
.B1(n_222),
.B2(n_277),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_215),
.A2(n_189),
.B1(n_153),
.B2(n_186),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_303),
.A2(n_307),
.B1(n_314),
.B2(n_337),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_249),
.A2(n_144),
.B1(n_189),
.B2(n_134),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_304),
.A2(n_340),
.B1(n_345),
.B2(n_234),
.Y(n_382)
);

NAND2xp33_ASAP7_75t_SL g309 ( 
.A(n_281),
.B(n_157),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g360 ( 
.A1(n_309),
.A2(n_278),
.B(n_240),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_221),
.A2(n_135),
.B1(n_144),
.B2(n_212),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_319),
.B(n_253),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_320),
.B(n_276),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_252),
.B(n_145),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_322),
.B(n_347),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_233),
.A2(n_5),
.B(n_9),
.Y(n_331)
);

OAI21xp33_ASAP7_75t_L g352 ( 
.A1(n_331),
.A2(n_262),
.B(n_268),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_221),
.B(n_175),
.C(n_208),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_335),
.B(n_338),
.C(n_342),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_221),
.A2(n_135),
.B1(n_175),
.B2(n_154),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_237),
.B(n_225),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_270),
.A2(n_154),
.B1(n_188),
.B2(n_176),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_245),
.B(n_261),
.C(n_214),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_269),
.A2(n_188),
.B1(n_190),
.B2(n_10),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_349),
.Y(n_411)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_346),
.B(n_238),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_366),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_351),
.B(n_353),
.Y(n_413)
);

NAND2xp67_ASAP7_75t_SL g394 ( 
.A(n_352),
.B(n_360),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_333),
.B(n_342),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_337),
.B(n_247),
.Y(n_354)
);

XNOR2x1_ASAP7_75t_L g397 ( 
.A(n_354),
.B(n_371),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_301),
.A2(n_217),
.B(n_219),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_356),
.A2(n_358),
.B(n_380),
.Y(n_399)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_299),
.Y(n_357)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_301),
.A2(n_230),
.B(n_227),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_323),
.Y(n_359)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_359),
.Y(n_426)
);

INVx8_ASAP7_75t_L g361 ( 
.A(n_316),
.Y(n_361)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_294),
.B(n_246),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_362),
.B(n_363),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_294),
.B(n_251),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_298),
.A2(n_321),
.B1(n_307),
.B2(n_335),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_364),
.A2(n_334),
.B1(n_289),
.B2(n_345),
.Y(n_407)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_324),
.Y(n_365)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_365),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_332),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_326),
.Y(n_367)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_367),
.Y(n_415)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_312),
.Y(n_368)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_368),
.Y(n_422)
);

INVx8_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_292),
.B(n_226),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_370),
.B(n_374),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_314),
.B(n_285),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_300),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_372),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_292),
.B(n_220),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_300),
.Y(n_375)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_375),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_306),
.B(n_228),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_374),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_341),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_378),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g378 ( 
.A1(n_309),
.A2(n_231),
.A3(n_239),
.B1(n_259),
.B2(n_264),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_229),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_379),
.B(n_385),
.C(n_340),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_347),
.A2(n_321),
.B(n_296),
.Y(n_380)
);

INVx13_ASAP7_75t_L g381 ( 
.A(n_310),
.Y(n_381)
);

INVx2_ASAP7_75t_SL g412 ( 
.A(n_381),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_382),
.A2(n_384),
.B1(n_325),
.B2(n_318),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_304),
.B(n_288),
.C(n_284),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_290),
.B(n_275),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_388),
.Y(n_409)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_387),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_295),
.B(n_265),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_297),
.B(n_274),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_389),
.Y(n_425)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g398 ( 
.A1(n_390),
.A2(n_392),
.B1(n_343),
.B2(n_318),
.Y(n_398)
);

OR2x2_ASAP7_75t_SL g391 ( 
.A(n_331),
.B(n_277),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_391),
.A2(n_327),
.B(n_315),
.Y(n_424)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_343),
.Y(n_392)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_393),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_395),
.B(n_427),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_398),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_353),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_339),
.C(n_305),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_404),
.B(n_408),
.C(n_419),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_407),
.A2(n_410),
.B1(n_428),
.B2(n_384),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_383),
.B(n_339),
.C(n_329),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_336),
.B1(n_330),
.B2(n_308),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_325),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_416),
.A2(n_424),
.B(n_361),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_339),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_363),
.B(n_291),
.C(n_327),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_420),
.B(n_431),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_421),
.A2(n_348),
.B1(n_371),
.B2(n_378),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_362),
.B(n_293),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_354),
.A2(n_336),
.B1(n_330),
.B2(n_256),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_360),
.B(n_376),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_432),
.B(n_441),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_425),
.B(n_366),
.Y(n_433)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_433),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_434),
.A2(n_437),
.B1(n_440),
.B2(n_449),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_413),
.B(n_389),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g471 ( 
.A(n_435),
.B(n_438),
.Y(n_471)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_422),
.Y(n_436)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_436),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_407),
.A2(n_382),
.B1(n_355),
.B2(n_385),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_411),
.B(n_357),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_401),
.B(n_390),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_439),
.B(n_442),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_406),
.A2(n_356),
.B1(n_350),
.B2(n_373),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_SL g441 ( 
.A(n_394),
.B(n_354),
.C(n_373),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_409),
.B(n_368),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g443 ( 
.A1(n_399),
.A2(n_380),
.B(n_349),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_443),
.A2(n_458),
.B(n_416),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_431),
.B(n_370),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_445),
.B(n_461),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_446),
.A2(n_460),
.B1(n_428),
.B2(n_429),
.Y(n_487)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_447),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_400),
.A2(n_371),
.B1(n_369),
.B2(n_361),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_448),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_395),
.A2(n_348),
.B1(n_391),
.B2(n_386),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_365),
.Y(n_450)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

INVx8_ASAP7_75t_L g452 ( 
.A(n_396),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g494 ( 
.A(n_452),
.Y(n_494)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_405),
.Y(n_453)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_453),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_414),
.B(n_375),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_454),
.B(n_455),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_414),
.B(n_372),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_420),
.A2(n_387),
.B1(n_392),
.B2(n_315),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_457),
.A2(n_416),
.B(n_429),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_416),
.A2(n_369),
.B1(n_359),
.B2(n_367),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_415),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_313),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_462),
.B(n_464),
.Y(n_476)
);

NAND3xp33_ASAP7_75t_L g463 ( 
.A(n_394),
.B(n_293),
.C(n_344),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_466),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_313),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_410),
.A2(n_235),
.B1(n_241),
.B2(n_311),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_465),
.A2(n_393),
.B1(n_381),
.B2(n_190),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_418),
.B(n_344),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_404),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_467),
.B(n_472),
.Y(n_523)
);

A2O1A1O1Ixp25_ASAP7_75t_L g468 ( 
.A1(n_432),
.A2(n_399),
.B(n_424),
.C(n_408),
.D(n_397),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_468),
.B(n_470),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_459),
.B(n_419),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_397),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_475),
.B(n_491),
.C(n_499),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_415),
.Y(n_478)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_478),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_479),
.A2(n_481),
.B(n_489),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_454),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_484),
.B(n_486),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_455),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_487),
.A2(n_440),
.B1(n_466),
.B2(n_462),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_458),
.A2(n_400),
.B(n_423),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_444),
.B(n_426),
.C(n_402),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_430),
.Y(n_492)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_492),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_446),
.A2(n_430),
.B1(n_396),
.B2(n_412),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_493),
.A2(n_434),
.B1(n_465),
.B2(n_437),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_464),
.B(n_412),
.Y(n_495)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_495),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_435),
.B(n_412),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g506 ( 
.A(n_496),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_498),
.A2(n_451),
.B1(n_460),
.B2(n_457),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_444),
.B(n_393),
.C(n_381),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_501),
.A2(n_516),
.B1(n_486),
.B2(n_471),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_439),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_502),
.B(n_518),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_450),
.Y(n_504)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_505),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_481),
.B(n_451),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_507),
.A2(n_479),
.B(n_489),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_478),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_509),
.B(n_522),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_467),
.B(n_456),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_510),
.B(n_512),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_472),
.B(n_449),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g539 ( 
.A1(n_513),
.A2(n_514),
.B1(n_517),
.B2(n_520),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_490),
.A2(n_443),
.B1(n_445),
.B2(n_442),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_487),
.A2(n_447),
.B1(n_436),
.B2(n_461),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_497),
.B(n_453),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_493),
.A2(n_473),
.B1(n_469),
.B2(n_484),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_499),
.C(n_475),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_521),
.B(n_524),
.C(n_485),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_492),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_469),
.B(n_441),
.C(n_452),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_480),
.A2(n_452),
.B1(n_9),
.B2(n_10),
.Y(n_525)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_525),
.Y(n_551)
);

INVx4_ASAP7_75t_L g526 ( 
.A(n_494),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_482),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_473),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_527),
.A2(n_498),
.B1(n_488),
.B2(n_477),
.Y(n_553)
);

INVx1_ASAP7_75t_SL g528 ( 
.A(n_474),
.Y(n_528)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_528),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_SL g548 ( 
.A(n_529),
.B(n_468),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_SL g530 ( 
.A(n_512),
.B(n_483),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_530),
.B(n_533),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_531),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_SL g533 ( 
.A(n_516),
.B(n_483),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_535),
.B(n_542),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_503),
.Y(n_536)
);

NOR3xp33_ASAP7_75t_L g570 ( 
.A(n_536),
.B(n_508),
.C(n_515),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_537),
.A2(n_505),
.B1(n_500),
.B2(n_515),
.Y(n_564)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_524),
.A2(n_511),
.B(n_507),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_538),
.A2(n_511),
.B(n_507),
.Y(n_560)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_540),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_510),
.B(n_476),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_519),
.B(n_476),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_543),
.B(n_545),
.C(n_549),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_519),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_SL g556 ( 
.A(n_544),
.B(n_547),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_521),
.B(n_485),
.C(n_495),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_523),
.B(n_514),
.Y(n_547)
);

XOR2x2_ASAP7_75t_L g563 ( 
.A(n_548),
.B(n_554),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_503),
.B(n_482),
.Y(n_549)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_553),
.Y(n_562)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_520),
.B(n_477),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_534),
.Y(n_555)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_555),
.Y(n_577)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_546),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_559),
.B(n_561),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_560),
.B(n_547),
.Y(n_581)
);

BUFx12_ASAP7_75t_L g561 ( 
.A(n_531),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_564),
.A2(n_526),
.B1(n_474),
.B2(n_488),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_537),
.A2(n_551),
.B1(n_513),
.B2(n_532),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_567),
.Y(n_575)
);

OA21x2_ASAP7_75t_SL g568 ( 
.A1(n_548),
.A2(n_504),
.B(n_471),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g582 ( 
.A1(n_568),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.Y(n_582)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_552),
.Y(n_569)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_550),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_549),
.B(n_528),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_572),
.B(n_542),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_533),
.A2(n_517),
.B1(n_506),
.B2(n_527),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_574),
.B(n_554),
.Y(n_576)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_576),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_573),
.A2(n_539),
.B(n_535),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_579),
.Y(n_597)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_581),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_566),
.B(n_543),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_583),
.B(n_587),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_566),
.B(n_545),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g602 ( 
.A(n_584),
.B(n_586),
.Y(n_602)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_585),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_555),
.B(n_541),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_558),
.B(n_541),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g588 ( 
.A1(n_562),
.A2(n_530),
.B1(n_544),
.B2(n_265),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_588),
.B(n_560),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_564),
.A2(n_265),
.B1(n_12),
.B2(n_13),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_589),
.A2(n_561),
.B1(n_12),
.B2(n_13),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_557),
.B(n_15),
.C(n_12),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_590),
.B(n_573),
.C(n_572),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_565),
.B(n_11),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_591),
.B(n_565),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_592),
.B(n_593),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_562),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_599),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g596 ( 
.A(n_588),
.B(n_563),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_596),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_577),
.B(n_563),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g612 ( 
.A(n_600),
.B(n_579),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g606 ( 
.A1(n_603),
.A2(n_575),
.B1(n_590),
.B2(n_581),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_580),
.B(n_556),
.Y(n_605)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_605),
.Y(n_614)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_606),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_602),
.B(n_582),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_607),
.B(n_610),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_598),
.C(n_578),
.Y(n_610)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_613),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g613 ( 
.A1(n_601),
.A2(n_585),
.B(n_561),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g615 ( 
.A(n_598),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_615),
.B(n_595),
.Y(n_617)
);

INVxp33_ASAP7_75t_SL g616 ( 
.A(n_611),
.Y(n_616)
);

NOR3xp33_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_617),
.C(n_604),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_610),
.B(n_597),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_618),
.B(n_620),
.Y(n_623)
);

CKINVDCx14_ASAP7_75t_R g620 ( 
.A(n_608),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_616),
.B(n_614),
.C(n_615),
.Y(n_624)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_624),
.B(n_625),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_621),
.A2(n_622),
.B(n_609),
.Y(n_625)
);

AOI322xp5_ASAP7_75t_L g628 ( 
.A1(n_626),
.A2(n_609),
.A3(n_619),
.B1(n_594),
.B2(n_600),
.C1(n_596),
.C2(n_589),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g629 ( 
.A(n_628),
.B(n_623),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_629),
.Y(n_630)
);

OAI21xp5_ASAP7_75t_L g631 ( 
.A1(n_630),
.A2(n_627),
.B(n_556),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_631),
.B(n_11),
.C(n_14),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_632),
.B(n_14),
.C(n_15),
.Y(n_633)
);


endmodule