module fake_jpeg_31004_n_152 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_152);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_152;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_39),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_9),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_27),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_12),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_2),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_56),
.Y(n_74)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_48),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_74),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_57),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_52),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_60),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_80),
.B(n_61),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_73),
.A2(n_64),
.B(n_59),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_94),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_55),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_7),
.C(n_8),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_84),
.A2(n_65),
.B1(n_56),
.B2(n_60),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_89),
.B(n_23),
.C(n_45),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_63),
.B1(n_49),
.B2(n_58),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_97),
.Y(n_105)
);

CKINVDCx10_ASAP7_75t_R g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_96),
.Y(n_102)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_54),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_95),
.B(n_101),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g96 ( 
.A(n_81),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_53),
.B1(n_62),
.B2(n_46),
.Y(n_97)
);

INVx13_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_99),
.B(n_100),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_3),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_116),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_111),
.B(n_19),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_91),
.A2(n_4),
.B(n_5),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_117),
.Y(n_125)
);

XOR2x1_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_5),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_113),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_6),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_7),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_119),
.Y(n_127)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_26),
.C(n_44),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_29),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_8),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_9),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_33),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_128),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_122),
.B(n_124),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_107),
.A2(n_10),
.B1(n_14),
.B2(n_15),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_133),
.Y(n_139)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_130),
.A2(n_134),
.B(n_110),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_103),
.A2(n_24),
.B1(n_30),
.B2(n_32),
.Y(n_131)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_102),
.B(n_36),
.Y(n_134)
);

NOR4xp25_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_137),
.C(n_140),
.D(n_138),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_123),
.A2(n_111),
.B(n_104),
.C(n_126),
.D(n_125),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_117),
.C(n_118),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_142),
.A2(n_144),
.B(n_141),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_136),
.A2(n_122),
.B1(n_131),
.B2(n_128),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_141),
.A2(n_127),
.B1(n_132),
.B2(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_146),
.B(n_139),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_147),
.B(n_145),
.Y(n_148)
);

FAx1_ASAP7_75t_SL g149 ( 
.A(n_148),
.B(n_38),
.CI(n_40),
.CON(n_149),
.SN(n_149)
);

NAND3xp33_ASAP7_75t_SL g150 ( 
.A(n_149),
.B(n_42),
.C(n_43),
.Y(n_150)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_150),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_149),
.Y(n_152)
);


endmodule