module fake_netlist_5_2479_n_1689 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1689);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1689;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_155;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_150;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_156;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_157;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_154;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_368;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_151;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1685;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1543;
wire n_1399;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_158;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_36),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_106),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_102),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_18),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_30),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_94),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_66),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_31),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_7),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_85),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_73),
.Y(n_164)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_36),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_77),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_39),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_22),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_3),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_130),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_129),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_5),
.Y(n_175)
);

BUFx3_ASAP7_75t_L g176 ( 
.A(n_62),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_59),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_88),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_72),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_90),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_80),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_7),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_149),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_61),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_30),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_74),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g188 ( 
.A(n_49),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_17),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_44),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_10),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_20),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_112),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_59),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_10),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_34),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_39),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_126),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_52),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_69),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_52),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_25),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_116),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_101),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_131),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_15),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_87),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_137),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_114),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_43),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_8),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_92),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_135),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_45),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_18),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_51),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_144),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_98),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_67),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_120),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_45),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_125),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_145),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_26),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_89),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_19),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_82),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_140),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_23),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_23),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_0),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_111),
.Y(n_236)
);

BUFx8_ASAP7_75t_SL g237 ( 
.A(n_8),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_33),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_96),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_60),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_79),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_148),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_42),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_0),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_124),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_49),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_81),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_86),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_55),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_20),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_53),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_38),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_105),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_29),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_34),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_76),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_14),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_103),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_2),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_57),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_63),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_65),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_113),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_38),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_35),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_91),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_21),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_128),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_1),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_19),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_141),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_46),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_61),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_136),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_31),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_26),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_75),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_47),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_110),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_4),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_108),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_55),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_56),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_93),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_147),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_146),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_193),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g296 ( 
.A(n_157),
.B(n_1),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_193),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_193),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_179),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g300 ( 
.A(n_240),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_205),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_193),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_193),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_212),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_193),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_281),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_259),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_259),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_224),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_259),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_259),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_237),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_150),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_242),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_280),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_153),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_291),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_271),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_271),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_154),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_277),
.B(n_2),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_158),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_163),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_164),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_271),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_166),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_271),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_271),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_168),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_162),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_287),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_180),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_160),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_287),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_160),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_181),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_183),
.Y(n_344)
);

NOR2xp67_ASAP7_75t_L g345 ( 
.A(n_188),
.B(n_4),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_162),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_170),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_287),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_277),
.B(n_5),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_170),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_194),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_209),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_241),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_202),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_209),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_229),
.B(n_6),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_241),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_209),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_151),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_157),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_211),
.B(n_9),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_152),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_261),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_207),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_208),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_161),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_328),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_178),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_331),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_295),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_295),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_297),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_297),
.B(n_176),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_298),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_349),
.B(n_324),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_298),
.B(n_232),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_302),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_302),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_303),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_346),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_167),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_303),
.Y(n_385)
);

CKINVDCx6p67_ASAP7_75t_R g386 ( 
.A(n_362),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_357),
.B(n_206),
.Y(n_387)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_305),
.B(n_176),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_305),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_307),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_308),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_308),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_310),
.B(n_176),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_310),
.B(n_211),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_311),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_300),
.B(n_233),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_311),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_357),
.B(n_206),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_312),
.Y(n_400)
);

AND2x4_ASAP7_75t_SL g401 ( 
.A(n_359),
.B(n_206),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_312),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_345),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_316),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_345),
.B(n_206),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_316),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_321),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_321),
.B(n_322),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_322),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_330),
.Y(n_411)
);

BUFx8_ASAP7_75t_L g412 ( 
.A(n_306),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_330),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_350),
.A2(n_294),
.B1(n_276),
.B2(n_182),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_332),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_335),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_306),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_356),
.B(n_173),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_337),
.B(n_213),
.Y(n_421)
);

BUFx2_ASAP7_75t_L g422 ( 
.A(n_353),
.Y(n_422)
);

BUFx8_ASAP7_75t_L g423 ( 
.A(n_296),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_337),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_339),
.B(n_341),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_339),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_341),
.B(n_216),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_343),
.B(n_221),
.Y(n_428)
);

CKINVDCx8_ASAP7_75t_R g429 ( 
.A(n_334),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_343),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_255),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_314),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_348),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_409),
.Y(n_436)
);

INVxp33_ASAP7_75t_SL g437 ( 
.A(n_384),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_409),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_403),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_392),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_378),
.B(n_355),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_409),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_384),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_432),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_419),
.B(n_378),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g450 ( 
.A(n_419),
.B(n_319),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_367),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_401),
.B(n_323),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_403),
.B(n_325),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_367),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_370),
.B(n_326),
.Y(n_456)
);

BUFx10_ASAP7_75t_L g457 ( 
.A(n_397),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_374),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_397),
.A2(n_399),
.B1(n_387),
.B2(n_165),
.Y(n_459)
);

INVx2_ASAP7_75t_SL g460 ( 
.A(n_423),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_376),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_386),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_401),
.B(n_327),
.Y(n_464)
);

BUFx3_ASAP7_75t_L g465 ( 
.A(n_376),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_370),
.B(n_329),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_401),
.B(n_333),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g468 ( 
.A(n_423),
.Y(n_468)
);

OAI22xp33_ASAP7_75t_L g469 ( 
.A1(n_387),
.A2(n_399),
.B1(n_334),
.B2(n_318),
.Y(n_469)
);

AND2x6_ASAP7_75t_L g470 ( 
.A(n_376),
.B(n_200),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_405),
.B(n_336),
.Y(n_471)
);

NOR3xp33_ASAP7_75t_L g472 ( 
.A(n_418),
.B(n_196),
.C(n_268),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_380),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_367),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_380),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_423),
.B(n_342),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_388),
.B(n_355),
.Y(n_480)
);

NOR3xp33_ASAP7_75t_L g481 ( 
.A(n_418),
.B(n_296),
.C(n_360),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_405),
.B(n_344),
.Y(n_482)
);

INVxp67_ASAP7_75t_SL g483 ( 
.A(n_421),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_367),
.Y(n_485)
);

AOI21x1_ASAP7_75t_L g486 ( 
.A1(n_395),
.A2(n_358),
.B(n_200),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_383),
.A2(n_228),
.B1(n_230),
.B2(n_218),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_379),
.B(n_351),
.Y(n_488)
);

BUFx6f_ASAP7_75t_SL g489 ( 
.A(n_429),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_429),
.B(n_354),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_429),
.B(n_364),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_375),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_375),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_372),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_372),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_375),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_379),
.B(n_365),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_372),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_367),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_421),
.B(n_255),
.Y(n_501)
);

OAI22xp33_ASAP7_75t_L g502 ( 
.A1(n_383),
.A2(n_171),
.B1(n_290),
.B2(n_289),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_427),
.B(n_255),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_382),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_382),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_388),
.A2(n_366),
.B(n_200),
.C(n_159),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_367),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_394),
.B(n_156),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_427),
.B(n_222),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_394),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_375),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_367),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_377),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_394),
.B(n_159),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_377),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_428),
.B(n_223),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_392),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_428),
.B(n_227),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_367),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_392),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_431),
.B(n_156),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_412),
.B(n_313),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_382),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_431),
.B(n_174),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_377),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_389),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_389),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_389),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_412),
.B(n_231),
.Y(n_529)
);

BUFx4f_ASAP7_75t_L g530 ( 
.A(n_392),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_390),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_412),
.B(n_236),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_377),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_412),
.B(n_239),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_433),
.B(n_299),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_431),
.Y(n_536)
);

OA22x2_ASAP7_75t_L g537 ( 
.A1(n_414),
.A2(n_247),
.B1(n_169),
.B2(n_177),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_412),
.B(n_245),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_386),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_390),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_412),
.B(n_248),
.Y(n_541)
);

NOR2x1p5_ASAP7_75t_L g542 ( 
.A(n_386),
.B(n_198),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_433),
.B(n_301),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_381),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_390),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_392),
.Y(n_546)
);

BUFx4f_ASAP7_75t_L g547 ( 
.A(n_392),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_433),
.A2(n_188),
.B1(n_261),
.B2(n_283),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_392),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_414),
.B(n_249),
.Y(n_550)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_368),
.B(n_198),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_381),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_381),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_393),
.Y(n_554)
);

OR2x6_ASAP7_75t_L g555 ( 
.A(n_368),
.B(n_174),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_381),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_433),
.B(n_253),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_433),
.B(n_304),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_393),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_393),
.Y(n_560)
);

NOR2x1p5_ASAP7_75t_L g561 ( 
.A(n_433),
.B(n_198),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_368),
.B(n_258),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_396),
.B(n_260),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_385),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_385),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_396),
.A2(n_283),
.B1(n_161),
.B2(n_250),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_396),
.Y(n_567)
);

INVx3_ASAP7_75t_L g568 ( 
.A(n_392),
.Y(n_568)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_402),
.Y(n_569)
);

INVx1_ASAP7_75t_SL g570 ( 
.A(n_384),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_407),
.A2(n_192),
.B1(n_203),
.B2(n_201),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_385),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_385),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_402),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_402),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_391),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_413),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_404),
.B(n_262),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_391),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_404),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_461),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_461),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_448),
.B(n_440),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_496),
.Y(n_585)
);

AND2x4_ASAP7_75t_SL g586 ( 
.A(n_555),
.B(n_309),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_471),
.B(n_315),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_440),
.B(n_155),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_483),
.B(n_514),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_461),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_465),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_536),
.B(n_186),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_514),
.B(n_404),
.Y(n_593)
);

NAND2xp33_ASAP7_75t_L g594 ( 
.A(n_470),
.B(n_264),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_496),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_L g596 ( 
.A(n_464),
.B(n_267),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_536),
.B(n_317),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_514),
.B(n_406),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_496),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_465),
.B(n_186),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_450),
.B(n_172),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_442),
.B(n_320),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_442),
.B(n_407),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_553),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_456),
.B(n_175),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_465),
.B(n_406),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_476),
.B(n_210),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_466),
.B(n_185),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_553),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_488),
.B(n_497),
.Y(n_610)
);

O2A1O1Ixp33_ASAP7_75t_L g611 ( 
.A1(n_506),
.A2(n_219),
.B(n_247),
.C(n_234),
.Y(n_611)
);

INVxp33_ASAP7_75t_SL g612 ( 
.A(n_445),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_476),
.B(n_210),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_553),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_436),
.A2(n_219),
.B1(n_184),
.B2(n_177),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_551),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_437),
.B(n_407),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_476),
.A2(n_265),
.B1(n_226),
.B2(n_292),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_510),
.B(n_210),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_470),
.B(n_270),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_510),
.B(n_406),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_454),
.B(n_190),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_459),
.B(n_191),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_457),
.B(n_422),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_557),
.A2(n_411),
.B(n_408),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_535),
.B(n_195),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_510),
.B(n_408),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_573),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_436),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_569),
.B(n_408),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_457),
.B(n_422),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_569),
.B(n_411),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_543),
.B(n_197),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_439),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_439),
.B(n_411),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_469),
.B(n_210),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_457),
.B(n_422),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_443),
.B(n_210),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_443),
.B(n_210),
.Y(n_639)
);

OAI221xp5_ASAP7_75t_L g640 ( 
.A1(n_566),
.A2(n_214),
.B1(n_184),
.B2(n_169),
.C(n_220),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_558),
.A2(n_288),
.B1(n_187),
.B2(n_272),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_446),
.B(n_187),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_446),
.B(n_189),
.Y(n_643)
);

OR2x6_ASAP7_75t_L g644 ( 
.A(n_542),
.B(n_214),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_447),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_551),
.Y(n_646)
);

INVxp67_ASAP7_75t_L g647 ( 
.A(n_457),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_447),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_449),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_573),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_561),
.A2(n_479),
.B1(n_482),
.B2(n_508),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_573),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_449),
.B(n_416),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_562),
.Y(n_654)
);

BUFx8_ASAP7_75t_L g655 ( 
.A(n_489),
.Y(n_655)
);

NAND2x1p5_ASAP7_75t_L g656 ( 
.A(n_438),
.B(n_217),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_555),
.Y(n_657)
);

NAND3xp33_ASAP7_75t_L g658 ( 
.A(n_481),
.B(n_273),
.C(n_215),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_487),
.B(n_204),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_509),
.B(n_416),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_516),
.B(n_416),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_518),
.B(n_417),
.Y(n_662)
);

NOR3xp33_ASAP7_75t_L g663 ( 
.A(n_550),
.B(n_199),
.C(n_235),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_572),
.B(n_238),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_480),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_501),
.B(n_243),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_503),
.B(n_417),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_502),
.B(n_453),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_480),
.B(n_508),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_473),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_561),
.A2(n_292),
.B1(n_284),
.B2(n_286),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_508),
.A2(n_286),
.B1(n_284),
.B2(n_293),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_467),
.B(n_244),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_563),
.B(n_251),
.Y(n_674)
);

AND2x6_ASAP7_75t_L g675 ( 
.A(n_508),
.B(n_275),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_521),
.A2(n_293),
.B1(n_275),
.B2(n_426),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_473),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_521),
.B(n_417),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_487),
.B(n_256),
.Y(n_679)
);

A2O1A1Ixp33_ASAP7_75t_L g680 ( 
.A1(n_521),
.A2(n_420),
.B(n_424),
.C(n_426),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_L g681 ( 
.A(n_470),
.B(n_257),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_521),
.B(n_420),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_555),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_555),
.B(n_204),
.Y(n_684)
);

AOI221xp5_ASAP7_75t_L g685 ( 
.A1(n_472),
.A2(n_225),
.B1(n_220),
.B2(n_234),
.C(n_250),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_478),
.B(n_420),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_478),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_494),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_524),
.B(n_363),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_460),
.B(n_434),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_579),
.B(n_424),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_580),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_494),
.B(n_424),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_460),
.B(n_434),
.Y(n_694)
);

BUFx5_ASAP7_75t_L g695 ( 
.A(n_470),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_468),
.B(n_434),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_468),
.B(n_434),
.Y(n_697)
);

NOR2x1p5_ASAP7_75t_L g698 ( 
.A(n_462),
.B(n_263),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_495),
.A2(n_426),
.B(n_398),
.C(n_279),
.Y(n_699)
);

AOI221xp5_ASAP7_75t_L g700 ( 
.A1(n_548),
.A2(n_279),
.B1(n_225),
.B2(n_252),
.C(n_254),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_495),
.B(n_398),
.Y(n_701)
);

BUFx8_ASAP7_75t_L g702 ( 
.A(n_489),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_498),
.B(n_398),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_580),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_498),
.B(n_398),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_504),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_505),
.B(n_523),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_505),
.B(n_434),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_444),
.B(n_269),
.Y(n_709)
);

INVx1_ASAP7_75t_SL g710 ( 
.A(n_570),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_580),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_523),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_458),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_490),
.B(n_491),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_SL g715 ( 
.A1(n_489),
.A2(n_204),
.B1(n_246),
.B2(n_285),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_526),
.B(n_398),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_524),
.B(n_274),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_524),
.B(n_282),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_527),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_524),
.B(n_204),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_458),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_475),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_527),
.B(n_398),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_475),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_528),
.B(n_435),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_524),
.A2(n_252),
.B(n_254),
.C(n_278),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_539),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_528),
.B(n_413),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_531),
.B(n_413),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_555),
.B(n_246),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_477),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_438),
.B(n_246),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_531),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_542),
.B(n_540),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_529),
.B(n_278),
.C(n_363),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_540),
.B(n_246),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_545),
.B(n_435),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_545),
.B(n_413),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_537),
.A2(n_285),
.B1(n_358),
.B2(n_435),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_554),
.B(n_435),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_554),
.B(n_413),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_559),
.B(n_413),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_559),
.B(n_413),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_560),
.B(n_64),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_560),
.B(n_285),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_L g746 ( 
.A(n_470),
.B(n_413),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_567),
.B(n_400),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_584),
.B(n_522),
.Y(n_748)
);

AOI21xp5_ASAP7_75t_L g749 ( 
.A1(n_669),
.A2(n_547),
.B(n_530),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_695),
.B(n_589),
.Y(n_750)
);

AOI21xp5_ASAP7_75t_L g751 ( 
.A1(n_593),
.A2(n_547),
.B(n_530),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_610),
.B(n_470),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_598),
.A2(n_682),
.B(n_678),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_660),
.A2(n_547),
.B(n_530),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_661),
.A2(n_662),
.B(n_691),
.Y(n_755)
);

AND2x4_ASAP7_75t_L g756 ( 
.A(n_734),
.B(n_451),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_690),
.A2(n_578),
.B(n_441),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_690),
.A2(n_578),
.B(n_441),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_744),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_734),
.B(n_451),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_694),
.A2(n_578),
.B(n_441),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_694),
.A2(n_697),
.B(n_696),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_610),
.B(n_470),
.Y(n_763)
);

NAND2xp33_ASAP7_75t_L g764 ( 
.A(n_695),
.B(n_567),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_L g765 ( 
.A1(n_625),
.A2(n_581),
.B(n_575),
.Y(n_765)
);

NOR2x1p5_ASAP7_75t_SL g766 ( 
.A(n_695),
.B(n_486),
.Y(n_766)
);

NAND2x1p5_ASAP7_75t_L g767 ( 
.A(n_744),
.B(n_575),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_696),
.A2(n_578),
.B(n_441),
.Y(n_768)
);

AOI21xp5_ASAP7_75t_L g769 ( 
.A1(n_697),
.A2(n_463),
.B(n_519),
.Y(n_769)
);

OAI21xp5_ASAP7_75t_L g770 ( 
.A1(n_701),
.A2(n_581),
.B(n_576),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_667),
.A2(n_463),
.B(n_519),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_606),
.A2(n_463),
.B(n_519),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_584),
.B(n_576),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_621),
.A2(n_627),
.B(n_746),
.Y(n_774)
);

O2A1O1Ixp33_ASAP7_75t_L g775 ( 
.A1(n_636),
.A2(n_532),
.B(n_534),
.C(n_538),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_612),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_582),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_666),
.B(n_452),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_583),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_623),
.A2(n_541),
.B(n_452),
.C(n_507),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_590),
.Y(n_781)
);

AOI21x1_ASAP7_75t_L g782 ( 
.A1(n_708),
.A2(n_486),
.B(n_574),
.Y(n_782)
);

O2A1O1Ixp33_ASAP7_75t_L g783 ( 
.A1(n_623),
.A2(n_577),
.B(n_574),
.C(n_484),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_591),
.Y(n_784)
);

AOI21x1_ASAP7_75t_L g785 ( 
.A1(n_708),
.A2(n_577),
.B(n_493),
.Y(n_785)
);

O2A1O1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_642),
.A2(n_552),
.B(n_493),
.C(n_492),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_707),
.A2(n_463),
.B(n_519),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_688),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_594),
.A2(n_519),
.B(n_507),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_620),
.A2(n_500),
.B(n_512),
.Y(n_790)
);

CKINVDCx20_ASAP7_75t_R g791 ( 
.A(n_727),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_666),
.B(n_605),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_695),
.B(n_452),
.Y(n_793)
);

AO21x1_ASAP7_75t_L g794 ( 
.A1(n_626),
.A2(n_556),
.B(n_492),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_706),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_607),
.A2(n_507),
.B(n_512),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_668),
.A2(n_477),
.B(n_484),
.C(n_565),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_607),
.A2(n_512),
.B(n_507),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_613),
.A2(n_512),
.B(n_500),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_613),
.A2(n_500),
.B(n_499),
.Y(n_800)
);

INVx3_ASAP7_75t_L g801 ( 
.A(n_712),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_703),
.A2(n_511),
.B(n_513),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_603),
.B(n_537),
.Y(n_803)
);

INVx8_ASAP7_75t_L g804 ( 
.A(n_675),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_719),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_695),
.B(n_452),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_619),
.A2(n_499),
.B(n_500),
.Y(n_807)
);

AOI21x1_ASAP7_75t_L g808 ( 
.A1(n_725),
.A2(n_513),
.B(n_511),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_605),
.B(n_455),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_733),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_629),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_705),
.A2(n_515),
.B(n_525),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_SL g813 ( 
.A(n_602),
.B(n_285),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_668),
.A2(n_525),
.B(n_515),
.C(n_565),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_585),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_SL g816 ( 
.A(n_655),
.B(n_533),
.Y(n_816)
);

OAI21xp5_ASAP7_75t_L g817 ( 
.A1(n_716),
.A2(n_552),
.B(n_544),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_695),
.B(n_455),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_619),
.A2(n_653),
.B(n_635),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_608),
.B(n_455),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_608),
.B(n_455),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_651),
.A2(n_474),
.B1(n_485),
.B2(n_499),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_723),
.A2(n_564),
.B(n_556),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_626),
.B(n_474),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_630),
.A2(n_474),
.B(n_485),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_689),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_642),
.A2(n_564),
.B(n_544),
.C(n_410),
.Y(n_827)
);

NOR2xp67_ASAP7_75t_L g828 ( 
.A(n_654),
.B(n_474),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_646),
.B(n_485),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_632),
.A2(n_485),
.B(n_499),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_634),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_633),
.B(n_568),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_595),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_633),
.B(n_568),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_728),
.A2(n_738),
.B(n_729),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_680),
.A2(n_520),
.B(n_568),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_645),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_741),
.A2(n_568),
.B(n_549),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_742),
.A2(n_549),
.B(n_546),
.Y(n_839)
);

AOI21x1_ASAP7_75t_L g840 ( 
.A1(n_725),
.A2(n_369),
.B(n_371),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_SL g841 ( 
.A(n_655),
.B(n_430),
.Y(n_841)
);

BUFx4f_ASAP7_75t_L g842 ( 
.A(n_644),
.Y(n_842)
);

NOR2xp33_ASAP7_75t_L g843 ( 
.A(n_616),
.B(n_549),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_648),
.B(n_549),
.Y(n_844)
);

A2O1A1Ixp33_ASAP7_75t_L g845 ( 
.A1(n_622),
.A2(n_546),
.B(n_520),
.C(n_415),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_649),
.A2(n_641),
.B1(n_714),
.B2(n_657),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_670),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_615),
.A2(n_435),
.B1(n_434),
.B2(n_415),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_743),
.A2(n_546),
.B(n_520),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_747),
.A2(n_693),
.B(n_681),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_714),
.A2(n_546),
.B1(n_520),
.B2(n_571),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_599),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_638),
.A2(n_410),
.B(n_391),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_674),
.B(n_677),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_674),
.B(n_571),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_686),
.A2(n_571),
.B(n_517),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_687),
.B(n_571),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_638),
.A2(n_410),
.B(n_391),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_665),
.B(n_571),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_647),
.B(n_9),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_600),
.A2(n_517),
.B(n_369),
.Y(n_861)
);

O2A1O1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_643),
.A2(n_430),
.B(n_415),
.C(n_410),
.Y(n_862)
);

O2A1O1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_643),
.A2(n_430),
.B(n_415),
.C(n_400),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_713),
.Y(n_864)
);

OAI21xp33_ASAP7_75t_L g865 ( 
.A1(n_664),
.A2(n_430),
.B(n_400),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_739),
.B(n_435),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_656),
.A2(n_601),
.B1(n_600),
.B2(n_683),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_592),
.B(n_400),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_639),
.A2(n_517),
.B(n_373),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_639),
.A2(n_517),
.B(n_373),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_721),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_722),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_592),
.B(n_373),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_737),
.A2(n_517),
.B(n_373),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_702),
.Y(n_875)
);

AOI21x1_ASAP7_75t_L g876 ( 
.A1(n_737),
.A2(n_371),
.B(n_369),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_740),
.A2(n_517),
.B(n_371),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_588),
.B(n_371),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_587),
.B(n_11),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_689),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_588),
.B(n_369),
.Y(n_881)
);

O2A1O1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_618),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_624),
.Y(n_883)
);

BUFx12f_ASAP7_75t_L g884 ( 
.A(n_702),
.Y(n_884)
);

BUFx3_ASAP7_75t_L g885 ( 
.A(n_586),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_740),
.A2(n_435),
.B(n_434),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_736),
.B(n_435),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_656),
.A2(n_435),
.B1(n_434),
.B2(n_143),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_664),
.A2(n_434),
.B(n_13),
.C(n_14),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_736),
.B(n_12),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_724),
.A2(n_138),
.B(n_133),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_731),
.A2(n_127),
.B(n_123),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_597),
.B(n_16),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_604),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_739),
.B(n_119),
.Y(n_895)
);

AOI21xp5_ASAP7_75t_L g896 ( 
.A1(n_609),
.A2(n_115),
.B(n_107),
.Y(n_896)
);

OAI21xp33_ASAP7_75t_SL g897 ( 
.A1(n_601),
.A2(n_17),
.B(n_21),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_745),
.B(n_24),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_614),
.A2(n_104),
.B(n_100),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_628),
.A2(n_99),
.B(n_97),
.Y(n_900)
);

O2A1O1Ixp5_ASAP7_75t_L g901 ( 
.A1(n_745),
.A2(n_24),
.B(n_27),
.C(n_28),
.Y(n_901)
);

AND2x6_ASAP7_75t_L g902 ( 
.A(n_684),
.B(n_78),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_650),
.Y(n_903)
);

OAI21xp33_ASAP7_75t_L g904 ( 
.A1(n_673),
.A2(n_27),
.B(n_28),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_659),
.B(n_32),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_652),
.A2(n_71),
.B(n_68),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_692),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_735),
.B(n_32),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_704),
.A2(n_33),
.B(n_35),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_615),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_596),
.B(n_671),
.Y(n_911)
);

AOI22x1_ASAP7_75t_L g912 ( 
.A1(n_711),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_912)
);

AND2x6_ASAP7_75t_L g913 ( 
.A(n_720),
.B(n_730),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_720),
.B(n_42),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_710),
.B(n_43),
.Y(n_915)
);

OAI21xp5_ASAP7_75t_L g916 ( 
.A1(n_717),
.A2(n_718),
.B(n_699),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_717),
.B(n_44),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_718),
.B(n_46),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_676),
.B(n_675),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_675),
.B(n_48),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_675),
.A2(n_50),
.B(n_54),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_673),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_732),
.A2(n_58),
.B(n_60),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_672),
.A2(n_730),
.B1(n_658),
.B2(n_679),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_L g925 ( 
.A1(n_675),
.A2(n_726),
.B(n_611),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_644),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_663),
.A2(n_700),
.B(n_709),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_631),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_637),
.B(n_586),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_640),
.A2(n_685),
.B(n_715),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_698),
.B(n_617),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_669),
.A2(n_536),
.B(n_514),
.Y(n_932)
);

OAI22xp5_ASAP7_75t_L g933 ( 
.A1(n_792),
.A2(n_767),
.B1(n_759),
.B2(n_854),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_755),
.B(n_748),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_748),
.B(n_773),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_826),
.B(n_756),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_883),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_752),
.A2(n_763),
.B(n_850),
.Y(n_938)
);

OAI22xp5_ASAP7_75t_L g939 ( 
.A1(n_767),
.A2(n_759),
.B1(n_916),
.B2(n_867),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_913),
.A2(n_924),
.B1(n_905),
.B2(n_759),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_847),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_815),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_759),
.A2(n_810),
.B1(n_788),
.B2(n_801),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_811),
.B(n_831),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_833),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_913),
.A2(n_905),
.B1(n_879),
.B2(n_929),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_774),
.A2(n_855),
.B(n_819),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_753),
.A2(n_750),
.B(n_809),
.Y(n_948)
);

INVx1_ASAP7_75t_SL g949 ( 
.A(n_915),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_803),
.B(n_928),
.Y(n_950)
);

OAI22xp5_ASAP7_75t_L g951 ( 
.A1(n_788),
.A2(n_810),
.B1(n_801),
.B2(n_932),
.Y(n_951)
);

OAI21xp33_ASAP7_75t_L g952 ( 
.A1(n_879),
.A2(n_893),
.B(n_813),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_826),
.B(n_756),
.Y(n_953)
);

A2O1A1Ixp33_ASAP7_75t_SL g954 ( 
.A1(n_860),
.A2(n_775),
.B(n_765),
.C(n_927),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_852),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_928),
.B(n_929),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_837),
.B(n_913),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_889),
.A2(n_918),
.B(n_917),
.C(n_898),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_846),
.A2(n_880),
.B1(n_762),
.B2(n_919),
.Y(n_959)
);

HB1xp67_ASAP7_75t_L g960 ( 
.A(n_928),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_928),
.Y(n_961)
);

OAI21xp33_ASAP7_75t_L g962 ( 
.A1(n_893),
.A2(n_904),
.B(n_890),
.Y(n_962)
);

NAND2x1p5_ASAP7_75t_L g963 ( 
.A(n_880),
.B(n_760),
.Y(n_963)
);

OAI22xp33_ASAP7_75t_L g964 ( 
.A1(n_921),
.A2(n_930),
.B1(n_914),
.B2(n_918),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_913),
.B(n_795),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_860),
.B(n_776),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_781),
.Y(n_967)
);

NOR3xp33_ASAP7_75t_SL g968 ( 
.A(n_922),
.B(n_897),
.C(n_917),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_750),
.A2(n_821),
.B(n_820),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_781),
.Y(n_970)
);

AOI21x1_ASAP7_75t_L g971 ( 
.A1(n_824),
.A2(n_834),
.B(n_832),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_778),
.A2(n_764),
.B(n_751),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_760),
.B(n_842),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_885),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_842),
.B(n_805),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_913),
.B(n_829),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_754),
.A2(n_787),
.B(n_771),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_777),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_895),
.A2(n_780),
.B(n_925),
.C(n_923),
.Y(n_979)
);

AOI21x1_ASAP7_75t_L g980 ( 
.A1(n_887),
.A2(n_782),
.B(n_881),
.Y(n_980)
);

O2A1O1Ixp33_ASAP7_75t_L g981 ( 
.A1(n_889),
.A2(n_901),
.B(n_797),
.C(n_814),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_851),
.A2(n_911),
.B1(n_859),
.B2(n_910),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_931),
.B(n_779),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_911),
.A2(n_749),
.B(n_784),
.C(n_783),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_926),
.B(n_791),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_843),
.B(n_828),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_843),
.B(n_868),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_878),
.B(n_873),
.Y(n_988)
);

A2O1A1Ixp33_ASAP7_75t_SL g989 ( 
.A1(n_770),
.A2(n_836),
.B(n_817),
.C(n_812),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_772),
.A2(n_790),
.B(n_789),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_894),
.Y(n_991)
);

NAND2x1_ASAP7_75t_L g992 ( 
.A(n_903),
.B(n_907),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_804),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_804),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_864),
.B(n_871),
.Y(n_995)
);

CKINVDCx20_ASAP7_75t_R g996 ( 
.A(n_884),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_841),
.B(n_910),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_872),
.Y(n_998)
);

NOR3xp33_ASAP7_75t_L g999 ( 
.A(n_908),
.B(n_920),
.C(n_882),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_816),
.B(n_857),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_835),
.A2(n_866),
.B(n_758),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_875),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_902),
.Y(n_1003)
);

O2A1O1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_901),
.A2(n_797),
.B(n_814),
.C(n_908),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_844),
.B(n_804),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_865),
.B(n_902),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_902),
.Y(n_1007)
);

OA21x2_ASAP7_75t_L g1008 ( 
.A1(n_794),
.A2(n_845),
.B(n_823),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_902),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_902),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_825),
.B(n_830),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_866),
.A2(n_757),
.B(n_761),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_785),
.Y(n_1013)
);

A2O1A1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_766),
.A2(n_786),
.B(n_807),
.C(n_798),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_888),
.B(n_822),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_838),
.B(n_839),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_849),
.B(n_802),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_912),
.Y(n_1018)
);

NOR2x1_ASAP7_75t_SL g1019 ( 
.A(n_793),
.B(n_806),
.Y(n_1019)
);

OR2x6_ASAP7_75t_SL g1020 ( 
.A(n_909),
.B(n_906),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_768),
.A2(n_818),
.B(n_793),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_SL g1022 ( 
.A(n_769),
.B(n_861),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_806),
.B(n_818),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_796),
.B(n_799),
.Y(n_1024)
);

A2O1A1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_800),
.A2(n_827),
.B(n_856),
.C(n_863),
.Y(n_1025)
);

AOI21x1_ASAP7_75t_L g1026 ( 
.A1(n_808),
.A2(n_840),
.B(n_876),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_848),
.B(n_877),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_874),
.B(n_886),
.Y(n_1028)
);

INVx4_ASAP7_75t_L g1029 ( 
.A(n_848),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_869),
.B(n_870),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_853),
.A2(n_858),
.B(n_862),
.Y(n_1031)
);

O2A1O1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_891),
.A2(n_892),
.B(n_896),
.C(n_899),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_900),
.B(n_748),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_915),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_752),
.A2(n_763),
.B(n_755),
.Y(n_1035)
);

OAI22x1_ASAP7_75t_L g1036 ( 
.A1(n_905),
.A2(n_459),
.B1(n_668),
.B2(n_414),
.Y(n_1036)
);

NOR2x1_ASAP7_75t_L g1037 ( 
.A(n_776),
.B(n_791),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_855),
.A2(n_824),
.B(n_820),
.Y(n_1038)
);

O2A1O1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_792),
.A2(n_448),
.B(n_636),
.C(n_889),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_SL g1040 ( 
.A1(n_792),
.A2(n_895),
.B(n_636),
.C(n_917),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_815),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_792),
.A2(n_448),
.B(n_636),
.C(n_889),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_752),
.A2(n_763),
.B(n_755),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_792),
.B(n_610),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_792),
.B(n_610),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_752),
.A2(n_763),
.B(n_755),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_792),
.B(n_610),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_776),
.B(n_804),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_748),
.B(n_792),
.Y(n_1049)
);

NOR3xp33_ASAP7_75t_L g1050 ( 
.A(n_792),
.B(n_668),
.C(n_448),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_792),
.B(n_610),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_815),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_826),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_792),
.B(n_610),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_SL g1055 ( 
.A(n_791),
.B(n_612),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_792),
.B(n_610),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_883),
.Y(n_1057)
);

OAI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_792),
.A2(n_932),
.B(n_755),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_815),
.Y(n_1059)
);

O2A1O1Ixp5_ASAP7_75t_L g1060 ( 
.A1(n_792),
.A2(n_794),
.B(n_636),
.C(n_916),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_R g1061 ( 
.A(n_791),
.B(n_445),
.Y(n_1061)
);

INVxp67_ASAP7_75t_L g1062 ( 
.A(n_883),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_792),
.A2(n_610),
.B1(n_748),
.B2(n_668),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_792),
.B(n_610),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_792),
.B(n_610),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_847),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_791),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_883),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_815),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_883),
.B(n_603),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_792),
.A2(n_610),
.B1(n_748),
.B2(n_668),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_748),
.B(n_792),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_815),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_804),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_826),
.B(n_756),
.Y(n_1075)
);

CKINVDCx8_ASAP7_75t_R g1076 ( 
.A(n_883),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_815),
.Y(n_1077)
);

AO21x2_ASAP7_75t_L g1078 ( 
.A1(n_1058),
.A2(n_947),
.B(n_938),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_934),
.A2(n_947),
.B(n_1035),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_937),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1063),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1035),
.A2(n_1046),
.B(n_1043),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_1044),
.B(n_1051),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_977),
.A2(n_990),
.B(n_1012),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1043),
.A2(n_1046),
.B(n_989),
.Y(n_1085)
);

AOI221x1_ASAP7_75t_L g1086 ( 
.A1(n_952),
.A2(n_1036),
.B1(n_1050),
.B2(n_962),
.C(n_979),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_1012),
.A2(n_1021),
.B(n_1001),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_1070),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_938),
.A2(n_1001),
.B(n_972),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_974),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_972),
.A2(n_1017),
.B(n_1033),
.Y(n_1091)
);

O2A1O1Ixp5_ASAP7_75t_L g1092 ( 
.A1(n_1045),
.A2(n_1056),
.B(n_1047),
.C(n_964),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1054),
.B(n_1064),
.Y(n_1093)
);

NAND3xp33_ASAP7_75t_L g1094 ( 
.A(n_1050),
.B(n_1065),
.C(n_1049),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_958),
.A2(n_1039),
.B(n_1042),
.C(n_940),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_983),
.B(n_1062),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_993),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_948),
.A2(n_969),
.A3(n_959),
.B(n_939),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_1060),
.A2(n_964),
.B(n_1072),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_SL g1100 ( 
.A(n_1055),
.B(n_966),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_1057),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1066),
.Y(n_1102)
);

OAI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_1015),
.A2(n_935),
.B(n_1004),
.Y(n_1103)
);

HB1xp67_ASAP7_75t_L g1104 ( 
.A(n_1068),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_1062),
.Y(n_1105)
);

AO32x2_ASAP7_75t_L g1106 ( 
.A1(n_982),
.A2(n_933),
.A3(n_951),
.B1(n_1029),
.B2(n_943),
.Y(n_1106)
);

AOI221x1_ASAP7_75t_L g1107 ( 
.A1(n_999),
.A2(n_1006),
.B1(n_1025),
.B2(n_1014),
.C(n_1011),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1029),
.B(n_950),
.Y(n_1108)
);

BUFx4f_ASAP7_75t_SL g1109 ( 
.A(n_1002),
.Y(n_1109)
);

OR2x2_ASAP7_75t_L g1110 ( 
.A(n_949),
.B(n_1034),
.Y(n_1110)
);

AO21x2_ASAP7_75t_L g1111 ( 
.A1(n_971),
.A2(n_1038),
.B(n_1040),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_1021),
.A2(n_1016),
.B(n_1013),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_988),
.A2(n_1022),
.B(n_1032),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_936),
.B(n_953),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_987),
.A2(n_986),
.B(n_1032),
.Y(n_1115)
);

NOR2xp67_ASAP7_75t_L g1116 ( 
.A(n_985),
.B(n_998),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_980),
.A2(n_1031),
.B(n_976),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_944),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_956),
.B(n_946),
.Y(n_1119)
);

NAND3xp33_ASAP7_75t_L g1120 ( 
.A(n_968),
.B(n_999),
.C(n_997),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1030),
.A2(n_1004),
.B(n_1027),
.Y(n_1121)
);

INVx3_ASAP7_75t_SL g1122 ( 
.A(n_996),
.Y(n_1122)
);

AOI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1031),
.A2(n_957),
.B(n_965),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_973),
.A2(n_1018),
.B1(n_960),
.B2(n_975),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_978),
.B(n_960),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_968),
.A2(n_981),
.B(n_1000),
.C(n_1023),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1024),
.A2(n_1005),
.B(n_981),
.Y(n_1127)
);

BUFx2_ASAP7_75t_SL g1128 ( 
.A(n_1076),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1024),
.A2(n_1028),
.B(n_995),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_967),
.B(n_970),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_942),
.B(n_1077),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_992),
.A2(n_1008),
.B(n_991),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_945),
.B(n_1073),
.Y(n_1133)
);

AO31x2_ASAP7_75t_L g1134 ( 
.A1(n_1019),
.A2(n_1020),
.A3(n_1008),
.B(n_955),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1041),
.A2(n_1069),
.A3(n_1052),
.B(n_1059),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1003),
.B(n_1037),
.C(n_953),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_963),
.A2(n_1028),
.B(n_1074),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_963),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1007),
.A2(n_1010),
.B(n_1074),
.Y(n_1139)
);

AO31x2_ASAP7_75t_L g1140 ( 
.A1(n_994),
.A2(n_1053),
.A3(n_1009),
.B(n_961),
.Y(n_1140)
);

OR2x2_ASAP7_75t_L g1141 ( 
.A(n_1067),
.B(n_1075),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_961),
.B(n_936),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1074),
.A2(n_1009),
.B(n_994),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1074),
.A2(n_1009),
.B(n_1075),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_961),
.A2(n_1053),
.B(n_1048),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1048),
.B(n_1061),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_1048),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_974),
.Y(n_1148)
);

INVx5_ASAP7_75t_L g1149 ( 
.A(n_1074),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_934),
.A2(n_1058),
.B(n_792),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1045),
.B(n_1047),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_941),
.Y(n_1152)
);

A2O1A1Ixp33_ASAP7_75t_L g1153 ( 
.A1(n_1045),
.A2(n_1056),
.B(n_1047),
.C(n_1063),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1063),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_934),
.A2(n_1058),
.B(n_792),
.Y(n_1155)
);

O2A1O1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_952),
.A2(n_792),
.B(n_448),
.C(n_1045),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_934),
.A2(n_1058),
.B(n_792),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_934),
.A2(n_1058),
.B(n_792),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_941),
.Y(n_1159)
);

O2A1O1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_954),
.A2(n_792),
.B(n_964),
.C(n_918),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_934),
.A2(n_1058),
.B(n_792),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_952),
.A2(n_792),
.B(n_448),
.C(n_1045),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1026),
.A2(n_977),
.B(n_990),
.Y(n_1163)
);

AND2x2_ASAP7_75t_SL g1164 ( 
.A(n_1045),
.B(n_1047),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_934),
.A2(n_1058),
.B(n_792),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_934),
.A2(n_1058),
.B(n_1043),
.Y(n_1166)
);

AO21x1_ASAP7_75t_L g1167 ( 
.A1(n_964),
.A2(n_792),
.B(n_1063),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_954),
.A2(n_792),
.B(n_964),
.C(n_918),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_941),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_937),
.Y(n_1170)
);

NOR4xp25_ASAP7_75t_L g1171 ( 
.A(n_952),
.B(n_792),
.C(n_1047),
.D(n_1045),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_941),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_952),
.A2(n_792),
.B(n_448),
.C(n_1045),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_934),
.A2(n_1058),
.B(n_1043),
.Y(n_1174)
);

INVxp67_ASAP7_75t_SL g1175 ( 
.A(n_1045),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_1045),
.A2(n_1056),
.B(n_1047),
.C(n_1063),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_979),
.A2(n_794),
.A3(n_984),
.B(n_1001),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_934),
.A2(n_1058),
.B(n_1043),
.Y(n_1178)
);

OA21x2_ASAP7_75t_L g1179 ( 
.A1(n_1060),
.A2(n_1058),
.B(n_969),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1070),
.B(n_602),
.Y(n_1180)
);

NOR2x1_ASAP7_75t_SL g1181 ( 
.A(n_1074),
.B(n_1009),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_941),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1045),
.B(n_1047),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_974),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1045),
.A2(n_1056),
.B(n_1047),
.C(n_1063),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_979),
.A2(n_794),
.A3(n_984),
.B(n_1001),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1045),
.B(n_1047),
.Y(n_1187)
);

OAI22x1_ASAP7_75t_L g1188 ( 
.A1(n_1063),
.A2(n_1071),
.B1(n_459),
.B2(n_905),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_941),
.Y(n_1189)
);

A2O1A1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1045),
.A2(n_1056),
.B(n_1047),
.C(n_1063),
.Y(n_1190)
);

BUFx3_ASAP7_75t_L g1191 ( 
.A(n_974),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1026),
.A2(n_977),
.B(n_990),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_934),
.A2(n_1058),
.B(n_792),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_941),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_SL g1195 ( 
.A1(n_1019),
.A2(n_921),
.B(n_958),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1045),
.A2(n_1056),
.B1(n_1047),
.B2(n_792),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_941),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1044),
.B(n_710),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1045),
.B(n_1047),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1045),
.A2(n_1056),
.B(n_1047),
.C(n_1063),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_941),
.Y(n_1201)
);

AO22x2_ASAP7_75t_L g1202 ( 
.A1(n_997),
.A2(n_939),
.B1(n_917),
.B2(n_918),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_SL g1203 ( 
.A1(n_934),
.A2(n_982),
.B(n_939),
.Y(n_1203)
);

O2A1O1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_952),
.A2(n_792),
.B(n_448),
.C(n_1045),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_934),
.A2(n_1058),
.B(n_1043),
.Y(n_1205)
);

AND2x4_ASAP7_75t_L g1206 ( 
.A(n_936),
.B(n_953),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_941),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1045),
.B(n_1047),
.Y(n_1208)
);

NAND3xp33_ASAP7_75t_SL g1209 ( 
.A(n_1063),
.B(n_1071),
.C(n_952),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_979),
.A2(n_794),
.A3(n_984),
.B(n_1001),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_941),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1060),
.A2(n_1071),
.B(n_1063),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1196),
.A2(n_1208),
.B1(n_1183),
.B2(n_1199),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1164),
.B(n_1180),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_L g1215 ( 
.A(n_1136),
.B(n_1141),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1122),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1209),
.A2(n_1188),
.B1(n_1120),
.B2(n_1167),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_1146),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1102),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1202),
.A2(n_1119),
.B1(n_1094),
.B2(n_1154),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1153),
.A2(n_1200),
.B1(n_1190),
.B2(n_1185),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1202),
.A2(n_1175),
.B1(n_1151),
.B2(n_1208),
.Y(n_1222)
);

OAI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1176),
.A2(n_1199),
.B1(n_1187),
.B2(n_1183),
.Y(n_1223)
);

AOI22xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1202),
.A2(n_1187),
.B1(n_1151),
.B2(n_1154),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1081),
.A2(n_1212),
.B1(n_1103),
.B2(n_1119),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1083),
.B(n_1093),
.Y(n_1226)
);

BUFx3_ASAP7_75t_L g1227 ( 
.A(n_1090),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1172),
.Y(n_1228)
);

BUFx2_ASAP7_75t_L g1229 ( 
.A(n_1080),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_L g1230 ( 
.A1(n_1081),
.A2(n_1212),
.B1(n_1103),
.B2(n_1099),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1093),
.A2(n_1086),
.B1(n_1118),
.B2(n_1198),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_L g1232 ( 
.A1(n_1099),
.A2(n_1195),
.B1(n_1100),
.B2(n_1121),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1110),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1171),
.B(n_1088),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_L g1235 ( 
.A(n_1170),
.Y(n_1235)
);

OAI22xp33_ASAP7_75t_L g1236 ( 
.A1(n_1088),
.A2(n_1108),
.B1(n_1116),
.B2(n_1125),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_SL g1237 ( 
.A1(n_1121),
.A2(n_1128),
.B1(n_1108),
.B2(n_1179),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1152),
.Y(n_1238)
);

BUFx2_ASAP7_75t_SL g1239 ( 
.A(n_1096),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1159),
.Y(n_1240)
);

BUFx4f_ASAP7_75t_L g1241 ( 
.A(n_1114),
.Y(n_1241)
);

OAI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1124),
.A2(n_1126),
.B1(n_1095),
.B2(n_1105),
.Y(n_1242)
);

AOI22xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1147),
.A2(n_1114),
.B1(n_1206),
.B2(n_1104),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1169),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_1109),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1182),
.Y(n_1246)
);

BUFx4_ASAP7_75t_SL g1247 ( 
.A(n_1148),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1101),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1129),
.Y(n_1249)
);

INVx6_ASAP7_75t_L g1250 ( 
.A(n_1206),
.Y(n_1250)
);

BUFx2_ASAP7_75t_L g1251 ( 
.A(n_1191),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1138),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_1160),
.A2(n_1168),
.B1(n_1142),
.B2(n_1129),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1189),
.Y(n_1254)
);

BUFx8_ASAP7_75t_L g1255 ( 
.A(n_1184),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1145),
.Y(n_1256)
);

BUFx8_ASAP7_75t_L g1257 ( 
.A(n_1194),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1211),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1150),
.A2(n_1155),
.B1(n_1157),
.B2(n_1193),
.Y(n_1259)
);

INVx2_ASAP7_75t_SL g1260 ( 
.A(n_1140),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1181),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1140),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1144),
.Y(n_1263)
);

CKINVDCx11_ASAP7_75t_R g1264 ( 
.A(n_1197),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1092),
.A2(n_1173),
.B(n_1204),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1139),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_SL g1267 ( 
.A1(n_1179),
.A2(n_1157),
.B1(n_1165),
.B2(n_1150),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1156),
.B(n_1162),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1201),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1155),
.A2(n_1161),
.B1(n_1165),
.B2(n_1158),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1207),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1135),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1158),
.A2(n_1193),
.B1(n_1161),
.B2(n_1127),
.Y(n_1273)
);

OAI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1107),
.A2(n_1131),
.B1(n_1133),
.B2(n_1130),
.Y(n_1274)
);

OAI22xp33_ASAP7_75t_R g1275 ( 
.A1(n_1203),
.A2(n_1106),
.B1(n_1135),
.B2(n_1131),
.Y(n_1275)
);

OAI22xp5_ASAP7_75t_L g1276 ( 
.A1(n_1139),
.A2(n_1133),
.B1(n_1130),
.B2(n_1097),
.Y(n_1276)
);

CKINVDCx11_ASAP7_75t_R g1277 ( 
.A(n_1143),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1132),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1078),
.A2(n_1115),
.B1(n_1205),
.B2(n_1178),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1097),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1166),
.A2(n_1174),
.B1(n_1113),
.B2(n_1123),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1134),
.Y(n_1282)
);

INVx5_ASAP7_75t_L g1283 ( 
.A(n_1137),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1106),
.B(n_1134),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1113),
.A2(n_1091),
.B1(n_1085),
.B2(n_1079),
.Y(n_1285)
);

CKINVDCx11_ASAP7_75t_R g1286 ( 
.A(n_1106),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1112),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1117),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1091),
.Y(n_1289)
);

NAND2x1p5_ASAP7_75t_L g1290 ( 
.A(n_1087),
.B(n_1084),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1079),
.A2(n_1089),
.B1(n_1111),
.B2(n_1082),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1177),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_1089),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1177),
.Y(n_1294)
);

BUFx8_ASAP7_75t_L g1295 ( 
.A(n_1098),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1098),
.Y(n_1296)
);

AOI22x1_ASAP7_75t_SL g1297 ( 
.A1(n_1186),
.A2(n_1210),
.B1(n_1163),
.B2(n_1192),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1186),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1210),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1149),
.Y(n_1300)
);

INVxp67_ASAP7_75t_SL g1301 ( 
.A(n_1121),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1164),
.A2(n_952),
.B1(n_301),
.B2(n_304),
.Y(n_1302)
);

OR2x2_ASAP7_75t_L g1303 ( 
.A(n_1088),
.B(n_1175),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1209),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1109),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1209),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1196),
.A2(n_1071),
.B1(n_1063),
.B2(n_1047),
.Y(n_1307)
);

OAI22xp5_ASAP7_75t_L g1308 ( 
.A1(n_1196),
.A2(n_1071),
.B1(n_1063),
.B2(n_1047),
.Y(n_1308)
);

CKINVDCx11_ASAP7_75t_R g1309 ( 
.A(n_1122),
.Y(n_1309)
);

BUFx12f_ASAP7_75t_L g1310 ( 
.A(n_1080),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1164),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1164),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1209),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1164),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_SL g1316 ( 
.A1(n_1188),
.A2(n_1036),
.B1(n_905),
.B2(n_623),
.Y(n_1316)
);

INVx6_ASAP7_75t_L g1317 ( 
.A(n_1149),
.Y(n_1317)
);

BUFx8_ASAP7_75t_L g1318 ( 
.A(n_1080),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1209),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1319)
);

INVx1_ASAP7_75t_SL g1320 ( 
.A(n_1110),
.Y(n_1320)
);

BUFx12f_ASAP7_75t_L g1321 ( 
.A(n_1080),
.Y(n_1321)
);

INVx6_ASAP7_75t_L g1322 ( 
.A(n_1149),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1164),
.A2(n_1045),
.B1(n_1056),
.B2(n_1047),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1080),
.Y(n_1324)
);

INVx1_ASAP7_75t_SL g1325 ( 
.A(n_1303),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1291),
.A2(n_1285),
.B(n_1279),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1272),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_L g1328 ( 
.A1(n_1291),
.A2(n_1285),
.B(n_1279),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1292),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1289),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1286),
.B(n_1224),
.Y(n_1331)
);

AO21x1_ASAP7_75t_SL g1332 ( 
.A1(n_1230),
.A2(n_1268),
.B(n_1265),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1294),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1259),
.A2(n_1273),
.B(n_1230),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1259),
.A2(n_1273),
.B(n_1249),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1290),
.A2(n_1278),
.B(n_1287),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1301),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1282),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1213),
.B(n_1223),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1301),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1213),
.B(n_1299),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1249),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1284),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1296),
.B(n_1234),
.Y(n_1344)
);

INVx2_ASAP7_75t_SL g1345 ( 
.A(n_1283),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1221),
.A2(n_1307),
.B1(n_1308),
.B2(n_1313),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1232),
.A2(n_1253),
.B(n_1225),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1232),
.A2(n_1225),
.B(n_1220),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_SL g1349 ( 
.A1(n_1260),
.A2(n_1217),
.B(n_1242),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1304),
.A2(n_1319),
.B1(n_1315),
.B2(n_1306),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1276),
.A2(n_1215),
.B(n_1238),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1293),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1298),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1295),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1295),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1275),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1297),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1288),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1248),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1288),
.Y(n_1360)
);

BUFx2_ASAP7_75t_L g1361 ( 
.A(n_1262),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_SL g1362 ( 
.A1(n_1217),
.A2(n_1299),
.B(n_1269),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1244),
.A2(n_1254),
.B(n_1246),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1240),
.A2(n_1228),
.B(n_1219),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1256),
.Y(n_1365)
);

INVx1_ASAP7_75t_SL g1366 ( 
.A(n_1233),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1270),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1316),
.B(n_1222),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1304),
.A2(n_1315),
.B(n_1313),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1270),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1320),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1222),
.B(n_1237),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1281),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1267),
.Y(n_1374)
);

AO21x2_ASAP7_75t_L g1375 ( 
.A1(n_1274),
.A2(n_1231),
.B(n_1236),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1267),
.Y(n_1376)
);

OA21x2_ASAP7_75t_L g1377 ( 
.A1(n_1306),
.A2(n_1319),
.B(n_1226),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_1300),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1237),
.Y(n_1379)
);

INVxp67_ASAP7_75t_L g1380 ( 
.A(n_1239),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1274),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1311),
.A2(n_1314),
.B1(n_1323),
.B2(n_1312),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1214),
.A2(n_1251),
.B(n_1324),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1277),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1231),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1236),
.A2(n_1322),
.B(n_1317),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1311),
.B(n_1323),
.Y(n_1387)
);

OA21x2_ASAP7_75t_L g1388 ( 
.A1(n_1271),
.A2(n_1302),
.B(n_1280),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1312),
.A2(n_1314),
.B(n_1266),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1216),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1325),
.B(n_1229),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1346),
.A2(n_1243),
.B(n_1241),
.C(n_1257),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1325),
.B(n_1318),
.Y(n_1393)
);

BUFx8_ASAP7_75t_SL g1394 ( 
.A(n_1390),
.Y(n_1394)
);

AOI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1339),
.A2(n_1241),
.B(n_1317),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1363),
.Y(n_1396)
);

AO32x2_ASAP7_75t_L g1397 ( 
.A1(n_1345),
.A2(n_1378),
.A3(n_1344),
.B1(n_1356),
.B2(n_1343),
.Y(n_1397)
);

NOR2xp33_ASAP7_75t_L g1398 ( 
.A(n_1352),
.B(n_1321),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1353),
.B(n_1218),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1363),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1339),
.A2(n_1263),
.B(n_1261),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1379),
.B(n_1218),
.Y(n_1402)
);

OR2x2_ASAP7_75t_L g1403 ( 
.A(n_1344),
.B(n_1227),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1365),
.B(n_1305),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1334),
.A2(n_1250),
.B(n_1252),
.Y(n_1405)
);

AOI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1382),
.A2(n_1245),
.B1(n_1264),
.B2(n_1258),
.C(n_1257),
.Y(n_1406)
);

AOI221xp5_ASAP7_75t_L g1407 ( 
.A1(n_1350),
.A2(n_1247),
.B1(n_1318),
.B2(n_1310),
.C(n_1235),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1352),
.A2(n_1250),
.B1(n_1247),
.B2(n_1255),
.Y(n_1408)
);

AND2x2_ASAP7_75t_SL g1409 ( 
.A(n_1334),
.B(n_1309),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1389),
.A2(n_1255),
.B1(n_1387),
.B2(n_1380),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1389),
.A2(n_1387),
.B1(n_1380),
.B2(n_1369),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1369),
.A2(n_1368),
.B1(n_1332),
.B2(n_1356),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1366),
.B(n_1371),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1369),
.A2(n_1368),
.B1(n_1332),
.B2(n_1388),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1415)
);

AND2x2_ASAP7_75t_L g1416 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1416)
);

A2O1A1Ixp33_ASAP7_75t_L g1417 ( 
.A1(n_1347),
.A2(n_1348),
.B(n_1372),
.C(n_1341),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1366),
.B(n_1371),
.Y(n_1418)
);

AOI221xp5_ASAP7_75t_L g1419 ( 
.A1(n_1385),
.A2(n_1381),
.B1(n_1370),
.B2(n_1367),
.C(n_1341),
.Y(n_1419)
);

AO32x1_ASAP7_75t_L g1420 ( 
.A1(n_1385),
.A2(n_1381),
.A3(n_1372),
.B1(n_1329),
.B2(n_1333),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1348),
.A2(n_1369),
.B(n_1347),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1330),
.B(n_1359),
.Y(n_1422)
);

OR2x2_ASAP7_75t_L g1423 ( 
.A(n_1342),
.B(n_1373),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1365),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1334),
.B(n_1358),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1377),
.B(n_1388),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1369),
.A2(n_1388),
.B1(n_1330),
.B2(n_1331),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1334),
.B(n_1360),
.Y(n_1428)
);

NOR2xp67_ASAP7_75t_SL g1429 ( 
.A(n_1384),
.B(n_1388),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1377),
.B(n_1364),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1384),
.Y(n_1431)
);

AO21x2_ASAP7_75t_L g1432 ( 
.A1(n_1349),
.A2(n_1328),
.B(n_1326),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1331),
.B(n_1337),
.Y(n_1433)
);

AOI211xp5_ASAP7_75t_L g1434 ( 
.A1(n_1357),
.A2(n_1355),
.B(n_1354),
.C(n_1384),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1377),
.A2(n_1375),
.B1(n_1384),
.B2(n_1362),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1326),
.A2(n_1328),
.B(n_1386),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1384),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1340),
.B(n_1335),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1364),
.B(n_1354),
.Y(n_1439)
);

OR2x2_ASAP7_75t_L g1440 ( 
.A(n_1338),
.B(n_1335),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1402),
.B(n_1383),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1396),
.Y(n_1442)
);

OAI221xp5_ASAP7_75t_SL g1443 ( 
.A1(n_1414),
.A2(n_1357),
.B1(n_1355),
.B2(n_1375),
.C(n_1362),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1438),
.B(n_1335),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1400),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1425),
.B(n_1375),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1438),
.B(n_1335),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1430),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1425),
.B(n_1428),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1436),
.B(n_1421),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1439),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1397),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1432),
.B(n_1335),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1432),
.B(n_1326),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1428),
.B(n_1375),
.Y(n_1455)
);

INVxp67_ASAP7_75t_SL g1456 ( 
.A(n_1440),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1432),
.B(n_1328),
.Y(n_1457)
);

OR2x2_ASAP7_75t_L g1458 ( 
.A(n_1426),
.B(n_1338),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1411),
.A2(n_1349),
.B1(n_1384),
.B2(n_1386),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1397),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1420),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1424),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1397),
.Y(n_1463)
);

AND2x2_ASAP7_75t_SL g1464 ( 
.A(n_1409),
.B(n_1361),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1442),
.Y(n_1465)
);

INVxp67_ASAP7_75t_SL g1466 ( 
.A(n_1456),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1444),
.B(n_1417),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1449),
.B(n_1417),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1444),
.B(n_1447),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1442),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1462),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1442),
.Y(n_1472)
);

OAI21xp33_ASAP7_75t_L g1473 ( 
.A1(n_1459),
.A2(n_1412),
.B(n_1427),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1445),
.Y(n_1474)
);

AOI211xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1443),
.A2(n_1410),
.B(n_1434),
.C(n_1405),
.Y(n_1475)
);

INVx3_ASAP7_75t_SL g1476 ( 
.A(n_1464),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1451),
.B(n_1415),
.Y(n_1477)
);

NOR2xp33_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1393),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1444),
.B(n_1415),
.Y(n_1479)
);

NAND3xp33_ASAP7_75t_L g1480 ( 
.A(n_1443),
.B(n_1419),
.C(n_1429),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1458),
.B(n_1446),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1447),
.B(n_1416),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1445),
.A2(n_1351),
.B(n_1336),
.Y(n_1483)
);

NOR2xp67_ASAP7_75t_L g1484 ( 
.A(n_1446),
.B(n_1401),
.Y(n_1484)
);

AOI31xp33_ASAP7_75t_L g1485 ( 
.A1(n_1459),
.A2(n_1406),
.A3(n_1408),
.B(n_1407),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1447),
.B(n_1416),
.Y(n_1486)
);

INVxp67_ASAP7_75t_SL g1487 ( 
.A(n_1456),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1458),
.B(n_1446),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1447),
.B(n_1433),
.Y(n_1489)
);

OAI33xp33_ASAP7_75t_L g1490 ( 
.A1(n_1461),
.A2(n_1413),
.A3(n_1391),
.B1(n_1403),
.B2(n_1423),
.B3(n_1327),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1452),
.B(n_1433),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1469),
.B(n_1452),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1469),
.B(n_1452),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1465),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1465),
.Y(n_1495)
);

NAND2x1p5_ASAP7_75t_L g1496 ( 
.A(n_1483),
.B(n_1453),
.Y(n_1496)
);

BUFx4f_ASAP7_75t_SL g1497 ( 
.A(n_1476),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1481),
.B(n_1463),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1483),
.A2(n_1457),
.B(n_1454),
.Y(n_1499)
);

INVx4_ASAP7_75t_L g1500 ( 
.A(n_1476),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1467),
.B(n_1460),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1467),
.B(n_1460),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1470),
.Y(n_1503)
);

INVx2_ASAP7_75t_L g1504 ( 
.A(n_1474),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1470),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1467),
.B(n_1463),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1472),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1466),
.B(n_1448),
.Y(n_1508)
);

BUFx2_ASAP7_75t_L g1509 ( 
.A(n_1476),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1480),
.B(n_1435),
.C(n_1450),
.Y(n_1510)
);

NAND2x1p5_ASAP7_75t_L g1511 ( 
.A(n_1483),
.B(n_1453),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1471),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1491),
.B(n_1489),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1466),
.B(n_1448),
.Y(n_1514)
);

NOR2xp67_ASAP7_75t_L g1515 ( 
.A(n_1468),
.B(n_1480),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1494),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1494),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1509),
.B(n_1489),
.Y(n_1518)
);

INVxp67_ASAP7_75t_L g1519 ( 
.A(n_1515),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1513),
.Y(n_1520)
);

AO21x1_ASAP7_75t_L g1521 ( 
.A1(n_1501),
.A2(n_1485),
.B(n_1487),
.Y(n_1521)
);

AND2x4_ASAP7_75t_L g1522 ( 
.A(n_1500),
.B(n_1509),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1509),
.B(n_1479),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1513),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1494),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1510),
.B(n_1394),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1515),
.B(n_1468),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1508),
.B(n_1481),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1500),
.B(n_1484),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1495),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1495),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1495),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1503),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1510),
.B(n_1484),
.Y(n_1534)
);

INVx2_ASAP7_75t_SL g1535 ( 
.A(n_1512),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1501),
.B(n_1479),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1513),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1508),
.B(n_1478),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1514),
.B(n_1477),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1503),
.Y(n_1540)
);

OAI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1501),
.A2(n_1473),
.B(n_1475),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1514),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1500),
.B(n_1464),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1498),
.B(n_1488),
.Y(n_1544)
);

NAND4xp25_ASAP7_75t_L g1545 ( 
.A(n_1500),
.B(n_1475),
.C(n_1473),
.D(n_1422),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1503),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1505),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1502),
.B(n_1479),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1502),
.B(n_1482),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1482),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1506),
.B(n_1477),
.Y(n_1552)
);

INVxp67_ASAP7_75t_SL g1553 ( 
.A(n_1512),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1505),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1505),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1507),
.Y(n_1556)
);

OR2x2_ASAP7_75t_L g1557 ( 
.A(n_1498),
.B(n_1488),
.Y(n_1557)
);

INVxp67_ASAP7_75t_L g1558 ( 
.A(n_1527),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1519),
.B(n_1482),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1521),
.A2(n_1409),
.B1(n_1450),
.B2(n_1464),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1541),
.A2(n_1500),
.B1(n_1497),
.B2(n_1450),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1536),
.B(n_1506),
.Y(n_1562)
);

INVx1_ASAP7_75t_SL g1563 ( 
.A(n_1522),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1516),
.Y(n_1564)
);

HB1xp67_ASAP7_75t_L g1565 ( 
.A(n_1518),
.Y(n_1565)
);

NOR2x1_ASAP7_75t_L g1566 ( 
.A(n_1545),
.B(n_1512),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1521),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1538),
.B(n_1486),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1522),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1552),
.B(n_1498),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1543),
.Y(n_1571)
);

NAND2x1_ASAP7_75t_SL g1572 ( 
.A(n_1522),
.B(n_1512),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1516),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1543),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1536),
.B(n_1506),
.Y(n_1575)
);

NAND4xp25_ASAP7_75t_L g1576 ( 
.A(n_1526),
.B(n_1418),
.C(n_1398),
.D(n_1450),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1548),
.B(n_1492),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1534),
.A2(n_1485),
.B(n_1499),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1548),
.Y(n_1579)
);

NOR2xp67_ASAP7_75t_L g1580 ( 
.A(n_1535),
.B(n_1518),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1549),
.B(n_1492),
.Y(n_1581)
);

INVx1_ASAP7_75t_SL g1582 ( 
.A(n_1523),
.Y(n_1582)
);

NOR2xp33_ASAP7_75t_L g1583 ( 
.A(n_1542),
.B(n_1394),
.Y(n_1583)
);

NAND3xp33_ASAP7_75t_L g1584 ( 
.A(n_1529),
.B(n_1457),
.C(n_1454),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1523),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1539),
.B(n_1486),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1587)
);

INVx2_ASAP7_75t_SL g1588 ( 
.A(n_1535),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1549),
.B(n_1493),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1528),
.B(n_1520),
.Y(n_1590)
);

OAI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1543),
.A2(n_1497),
.B1(n_1455),
.B2(n_1437),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1551),
.B(n_1493),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1564),
.Y(n_1593)
);

INVx1_ASAP7_75t_SL g1594 ( 
.A(n_1563),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

NAND2x1p5_ASAP7_75t_L g1596 ( 
.A(n_1566),
.B(n_1529),
.Y(n_1596)
);

AOI21xp33_ASAP7_75t_L g1597 ( 
.A1(n_1567),
.A2(n_1529),
.B(n_1553),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1566),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1558),
.B(n_1551),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1560),
.A2(n_1457),
.B1(n_1454),
.B2(n_1464),
.Y(n_1600)
);

AOI322xp5_ASAP7_75t_L g1601 ( 
.A1(n_1560),
.A2(n_1561),
.A3(n_1583),
.B1(n_1582),
.B2(n_1562),
.C1(n_1575),
.C2(n_1585),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1569),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1573),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1576),
.B(n_1520),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1573),
.Y(n_1605)
);

NOR2xp33_ASAP7_75t_L g1606 ( 
.A(n_1576),
.B(n_1524),
.Y(n_1606)
);

NOR2x1_ASAP7_75t_L g1607 ( 
.A(n_1578),
.B(n_1556),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1574),
.B(n_1464),
.Y(n_1608)
);

OAI31xp33_ASAP7_75t_SL g1609 ( 
.A1(n_1584),
.A2(n_1499),
.A3(n_1524),
.B(n_1537),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1565),
.Y(n_1610)
);

O2A1O1Ixp33_ASAP7_75t_L g1611 ( 
.A1(n_1571),
.A2(n_1511),
.B(n_1496),
.C(n_1392),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1584),
.A2(n_1580),
.B1(n_1571),
.B2(n_1574),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1590),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1590),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1562),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1575),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1579),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1596),
.B(n_1572),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1593),
.Y(n_1619)
);

OAI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1607),
.A2(n_1574),
.B1(n_1572),
.B2(n_1580),
.C(n_1559),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1595),
.Y(n_1621)
);

INVxp67_ASAP7_75t_SL g1622 ( 
.A(n_1596),
.Y(n_1622)
);

NAND3xp33_ASAP7_75t_L g1623 ( 
.A(n_1601),
.B(n_1588),
.C(n_1591),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1594),
.B(n_1568),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1602),
.B(n_1610),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1613),
.B(n_1588),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1599),
.B(n_1579),
.Y(n_1627)
);

AOI21xp33_ASAP7_75t_SL g1628 ( 
.A1(n_1609),
.A2(n_1587),
.B(n_1570),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1614),
.B(n_1577),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1603),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1597),
.Y(n_1631)
);

INVx3_ASAP7_75t_L g1632 ( 
.A(n_1615),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1604),
.B(n_1577),
.Y(n_1633)
);

INVx2_ASAP7_75t_L g1634 ( 
.A(n_1616),
.Y(n_1634)
);

NOR2xp33_ASAP7_75t_L g1635 ( 
.A(n_1604),
.B(n_1586),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1605),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1632),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1625),
.B(n_1598),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1631),
.A2(n_1598),
.B(n_1612),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1618),
.Y(n_1640)
);

INVx2_ASAP7_75t_L g1641 ( 
.A(n_1618),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1632),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1625),
.B(n_1606),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_SL g1644 ( 
.A1(n_1623),
.A2(n_1606),
.B1(n_1617),
.B2(n_1600),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1629),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1626),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1626),
.Y(n_1647)
);

NAND3x1_ASAP7_75t_L g1648 ( 
.A(n_1638),
.B(n_1621),
.C(n_1619),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1643),
.B(n_1631),
.Y(n_1649)
);

NOR2x1_ASAP7_75t_L g1650 ( 
.A(n_1642),
.B(n_1618),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1646),
.B(n_1635),
.Y(n_1651)
);

NAND4xp25_ASAP7_75t_L g1652 ( 
.A(n_1644),
.B(n_1623),
.C(n_1633),
.D(n_1624),
.Y(n_1652)
);

NAND4xp25_ASAP7_75t_L g1653 ( 
.A(n_1643),
.B(n_1620),
.C(n_1634),
.D(n_1627),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1642),
.B(n_1630),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_L g1655 ( 
.A(n_1637),
.B(n_1636),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1639),
.A2(n_1628),
.B(n_1622),
.C(n_1611),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1647),
.B(n_1608),
.Y(n_1657)
);

AOI221xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1656),
.A2(n_1641),
.B1(n_1645),
.B2(n_1640),
.C(n_1587),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_L g1659 ( 
.A(n_1649),
.B(n_1641),
.Y(n_1659)
);

INVx1_ASAP7_75t_SL g1660 ( 
.A(n_1650),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1657),
.B(n_1592),
.Y(n_1661)
);

AND5x1_ASAP7_75t_L g1662 ( 
.A(n_1652),
.B(n_1490),
.C(n_1441),
.D(n_1392),
.E(n_1395),
.Y(n_1662)
);

O2A1O1Ixp33_ASAP7_75t_L g1663 ( 
.A1(n_1660),
.A2(n_1659),
.B(n_1651),
.C(n_1654),
.Y(n_1663)
);

AOI211xp5_ASAP7_75t_L g1664 ( 
.A1(n_1658),
.A2(n_1653),
.B(n_1648),
.C(n_1655),
.Y(n_1664)
);

AOI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1661),
.A2(n_1592),
.B1(n_1589),
.B2(n_1581),
.Y(n_1665)
);

OAI21xp33_ASAP7_75t_L g1666 ( 
.A1(n_1662),
.A2(n_1589),
.B(n_1581),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1659),
.B(n_1537),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1659),
.A2(n_1570),
.B1(n_1437),
.B2(n_1431),
.Y(n_1668)
);

INVx1_ASAP7_75t_SL g1669 ( 
.A(n_1667),
.Y(n_1669)
);

AOI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1664),
.A2(n_1556),
.B1(n_1530),
.B2(n_1517),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1665),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1663),
.Y(n_1672)
);

NOR2xp67_ASAP7_75t_L g1673 ( 
.A(n_1668),
.B(n_1540),
.Y(n_1673)
);

XOR2xp5_ASAP7_75t_L g1674 ( 
.A(n_1671),
.B(n_1399),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_L g1675 ( 
.A(n_1672),
.B(n_1666),
.C(n_1399),
.Y(n_1675)
);

OAI21xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1670),
.A2(n_1437),
.B(n_1404),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1675),
.B(n_1669),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1677),
.A2(n_1674),
.B1(n_1676),
.B2(n_1673),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1550),
.B1(n_1525),
.B2(n_1533),
.Y(n_1679)
);

BUFx2_ASAP7_75t_SL g1680 ( 
.A(n_1678),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_SL g1681 ( 
.A1(n_1680),
.A2(n_1437),
.B1(n_1517),
.B2(n_1525),
.Y(n_1681)
);

OAI22x1_ASAP7_75t_L g1682 ( 
.A1(n_1679),
.A2(n_1550),
.B1(n_1547),
.B2(n_1532),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1681),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1682),
.A2(n_1531),
.B(n_1530),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1683),
.A2(n_1532),
.B1(n_1533),
.B2(n_1531),
.C(n_1547),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1685),
.A2(n_1684),
.B1(n_1555),
.B2(n_1554),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1686),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_R g1688 ( 
.A1(n_1687),
.A2(n_1546),
.B1(n_1512),
.B2(n_1544),
.C(n_1557),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1557),
.B(n_1544),
.C(n_1404),
.Y(n_1689)
);


endmodule