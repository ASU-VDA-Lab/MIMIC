module fake_ariane_3106_n_1141 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1141);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1141;

wire n_295;
wire n_356;
wire n_556;
wire n_1127;
wire n_698;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_423;
wire n_347;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_220;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_819;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_214;
wire n_1138;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_945;
wire n_958;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_779;
wire n_754;
wire n_871;
wire n_315;
wire n_903;
wire n_1073;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_1052;
wire n_1068;
wire n_272;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_1018;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_1047;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_1134;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_253;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_1099;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_997;
wire n_635;
wire n_707;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_1080;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_977;
wire n_957;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_1140;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_260;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_888;
wire n_845;
wire n_1135;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_1043;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_933;
wire n_872;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_213;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_1083;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_275;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_1139;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_1051;
wire n_494;
wire n_959;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_854;
wire n_841;
wire n_471;
wire n_351;
wire n_1069;
wire n_965;
wire n_393;
wire n_886;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_58),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_15),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_11),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_110),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_82),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_131),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_211),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_98),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_111),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_205),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_132),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_16),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_90),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_118),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_96),
.Y(n_230)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_151),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_25),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_158),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_44),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_19),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_91),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_67),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_17),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_84),
.Y(n_241)
);

BUFx8_ASAP7_75t_SL g242 ( 
.A(n_42),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_0),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_105),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_26),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_125),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_197),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_134),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_50),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_34),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_165),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_19),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_187),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_206),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_11),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_38),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_178),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_107),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_160),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_194),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_15),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_49),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_182),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_169),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_166),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_14),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_92),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_14),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_37),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_24),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_17),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_33),
.Y(n_273)
);

INVxp33_ASAP7_75t_SL g274 ( 
.A(n_12),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_135),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_49),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_12),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_168),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_72),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_13),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_62),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_139),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_177),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_255),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g289 ( 
.A(n_267),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_264),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_277),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_282),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_213),
.Y(n_297)
);

INVxp67_ASAP7_75t_SL g298 ( 
.A(n_231),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_217),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_224),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_231),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_279),
.Y(n_304)
);

INVxp67_ASAP7_75t_SL g305 ( 
.A(n_246),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_256),
.Y(n_307)
);

BUFx2_ASAP7_75t_SL g308 ( 
.A(n_282),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_246),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_238),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_274),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_249),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_226),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_254),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_265),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_233),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_269),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_223),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_223),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_237),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_237),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_237),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_237),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_237),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_236),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_218),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_280),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_218),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_326),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_239),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_326),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_220),
.Y(n_341)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_323),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_290),
.Y(n_347)
);

AND2x4_ASAP7_75t_L g348 ( 
.A(n_303),
.B(n_225),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_292),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_311),
.A2(n_274),
.B1(n_280),
.B2(n_235),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_299),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_309),
.B(n_219),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_325),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_312),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_289),
.B(n_243),
.Y(n_358)
);

NOR2x1_ASAP7_75t_L g359 ( 
.A(n_308),
.B(n_268),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

AND2x4_ASAP7_75t_L g361 ( 
.A(n_303),
.B(n_297),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_327),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_309),
.B(n_219),
.Y(n_363)
);

OA21x2_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_250),
.B(n_245),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_313),
.B(n_317),
.Y(n_366)
);

BUFx2_ASAP7_75t_L g367 ( 
.A(n_312),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_329),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_308),
.Y(n_369)
);

OAI22x1_ASAP7_75t_SL g370 ( 
.A1(n_307),
.A2(n_252),
.B1(n_270),
.B2(n_262),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_297),
.B(n_248),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_248),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_301),
.B(n_278),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_301),
.B(n_278),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_302),
.B(n_281),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_330),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_330),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_304),
.A2(n_273),
.B1(n_276),
.B2(n_271),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_332),
.B(n_281),
.Y(n_380)
);

BUFx8_ASAP7_75t_L g381 ( 
.A(n_320),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_331),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_302),
.B(n_212),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_306),
.B(n_221),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_306),
.B(n_222),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_291),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_331),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_324),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_314),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_310),
.B(n_227),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_322),
.A2(n_251),
.B1(n_275),
.B2(n_263),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_369),
.B(n_320),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_341),
.B(n_296),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_349),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_369),
.A2(n_333),
.B1(n_335),
.B2(n_318),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_356),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_379),
.A2(n_322),
.B1(n_286),
.B2(n_300),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_356),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_371),
.A2(n_335),
.B1(n_284),
.B2(n_305),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_357),
.A2(n_315),
.B1(n_319),
.B2(n_316),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_388),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_365),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_341),
.B(n_298),
.Y(n_408)
);

BUFx6f_ASAP7_75t_SL g409 ( 
.A(n_341),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_365),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_354),
.B(n_315),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_374),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_374),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_336),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_382),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_371),
.A2(n_319),
.B1(n_316),
.B2(n_294),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_387),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_341),
.B(n_293),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_339),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_349),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_349),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_336),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_359),
.B(n_229),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_389),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_371),
.B(n_293),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_375),
.A2(n_295),
.B1(n_294),
.B2(n_258),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_338),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_338),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_348),
.B(n_383),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_380),
.B(n_295),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_340),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_389),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_340),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_338),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_340),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_379),
.A2(n_285),
.B1(n_288),
.B2(n_287),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_381),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_345),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_345),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_346),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g450 ( 
.A(n_392),
.B(n_230),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_367),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_346),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_346),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_375),
.B(n_287),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_392),
.A2(n_285),
.B1(n_288),
.B2(n_283),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_352),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_342),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_352),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_348),
.B(n_232),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_352),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_360),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_360),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_357),
.A2(n_386),
.B1(n_375),
.B2(n_353),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_386),
.A2(n_247),
.B1(n_259),
.B2(n_257),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_360),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_383),
.B(n_234),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_368),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_368),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_414),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_436),
.B(n_359),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_451),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_408),
.B(n_366),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_438),
.B(n_383),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_457),
.Y(n_475)
);

INVx8_ASAP7_75t_L g476 ( 
.A(n_409),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_414),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_411),
.B(n_381),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_L g479 ( 
.A(n_445),
.B(n_395),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_421),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_342),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_398),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_400),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_432),
.B(n_348),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_432),
.B(n_348),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_445),
.B(n_370),
.Y(n_486)
);

NOR3xp33_ASAP7_75t_L g487 ( 
.A(n_463),
.B(n_353),
.C(n_337),
.Y(n_487)
);

NAND2xp33_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_373),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_466),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_419),
.B(n_361),
.Y(n_490)
);

NAND3xp33_ASAP7_75t_SL g491 ( 
.A(n_423),
.B(n_376),
.C(n_373),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_394),
.B(n_381),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_409),
.B(n_381),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_400),
.Y(n_494)
);

NAND3xp33_ASAP7_75t_L g495 ( 
.A(n_397),
.B(n_358),
.C(n_376),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_402),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_405),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_409),
.B(n_384),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_454),
.B(n_361),
.Y(n_500)
);

AO221x1_ASAP7_75t_L g501 ( 
.A1(n_399),
.A2(n_370),
.B1(n_393),
.B2(n_344),
.C(n_351),
.Y(n_501)
);

NOR3xp33_ASAP7_75t_L g502 ( 
.A(n_455),
.B(n_450),
.C(n_464),
.Y(n_502)
);

INVxp33_ASAP7_75t_L g503 ( 
.A(n_454),
.Y(n_503)
);

AO221x1_ASAP7_75t_L g504 ( 
.A1(n_444),
.A2(n_393),
.B1(n_344),
.B2(n_351),
.C(n_347),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_417),
.B(n_361),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_421),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_361),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_459),
.B(n_391),
.Y(n_508)
);

NOR3xp33_ASAP7_75t_L g509 ( 
.A(n_403),
.B(n_385),
.C(n_384),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_396),
.B(n_385),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_401),
.B(n_358),
.Y(n_511)
);

NOR3xp33_ASAP7_75t_L g512 ( 
.A(n_430),
.B(n_391),
.C(n_363),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_431),
.Y(n_513)
);

NOR2xp67_ASAP7_75t_L g514 ( 
.A(n_406),
.B(n_390),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_396),
.B(n_355),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_396),
.B(n_355),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_425),
.B(n_363),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_429),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_407),
.B(n_390),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_425),
.B(n_372),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_425),
.B(n_372),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_428),
.B(n_390),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_429),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_428),
.B(n_390),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_407),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g530 ( 
.A(n_431),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_434),
.Y(n_531)
);

BUFx8_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_428),
.B(n_389),
.Y(n_533)
);

AND2x2_ASAP7_75t_L g534 ( 
.A(n_412),
.B(n_347),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_412),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_413),
.Y(n_536)
);

BUFx6f_ASAP7_75t_SL g537 ( 
.A(n_413),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_415),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_415),
.B(n_350),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_416),
.B(n_350),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_404),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_431),
.B(n_440),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_435),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_418),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_418),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_440),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_420),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_420),
.B(n_364),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_435),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_422),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_440),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_487),
.A2(n_422),
.B1(n_437),
.B2(n_424),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_489),
.B(n_424),
.Y(n_554)
);

OR2x6_ASAP7_75t_L g555 ( 
.A(n_476),
.B(n_447),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_471),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_L g557 ( 
.A(n_509),
.B(n_404),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_479),
.B(n_437),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_469),
.Y(n_559)
);

OAI221xp5_ASAP7_75t_L g560 ( 
.A1(n_502),
.A2(n_443),
.B1(n_467),
.B2(n_465),
.C(n_446),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_469),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_477),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_482),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_483),
.Y(n_564)
);

OAI221xp5_ASAP7_75t_L g565 ( 
.A1(n_472),
.A2(n_443),
.B1(n_467),
.B2(n_465),
.C(n_446),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_475),
.B(n_404),
.Y(n_566)
);

AOI22x1_ASAP7_75t_L g567 ( 
.A1(n_494),
.A2(n_441),
.B1(n_449),
.B2(n_439),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_478),
.B(n_439),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

OAI221xp5_ASAP7_75t_L g570 ( 
.A1(n_511),
.A2(n_441),
.B1(n_461),
.B2(n_449),
.C(n_458),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_481),
.Y(n_571)
);

BUFx8_ASAP7_75t_L g572 ( 
.A(n_537),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_496),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_551),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_478),
.B(n_452),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_497),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_473),
.Y(n_577)
);

BUFx8_ASAP7_75t_L g578 ( 
.A(n_537),
.Y(n_578)
);

NAND2x1p5_ASAP7_75t_L g579 ( 
.A(n_529),
.B(n_493),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_551),
.B(n_452),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_474),
.B(n_453),
.Y(n_581)
);

BUFx6f_ASAP7_75t_SL g582 ( 
.A(n_532),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_516),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_526),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_473),
.B(n_404),
.Y(n_585)
);

AO22x2_ASAP7_75t_L g586 ( 
.A1(n_486),
.A2(n_495),
.B1(n_507),
.B2(n_485),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_539),
.A2(n_458),
.B1(n_461),
.B2(n_453),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_484),
.A2(n_468),
.B1(n_462),
.B2(n_460),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_527),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_535),
.Y(n_590)
);

AO22x2_ASAP7_75t_L g591 ( 
.A1(n_505),
.A2(n_468),
.B1(n_462),
.B2(n_460),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_488),
.A2(n_456),
.B1(n_448),
.B2(n_447),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_492),
.B(n_508),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_536),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_508),
.B(n_448),
.Y(n_595)
);

AO22x2_ASAP7_75t_L g596 ( 
.A1(n_504),
.A2(n_456),
.B1(n_364),
.B2(n_442),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_532),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_488),
.B(n_364),
.C(n_404),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_538),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_532),
.Y(n_600)
);

AO22x2_ASAP7_75t_L g601 ( 
.A1(n_540),
.A2(n_364),
.B1(n_442),
.B2(n_377),
.Y(n_601)
);

AOI22xp5_ASAP7_75t_L g602 ( 
.A1(n_492),
.A2(n_364),
.B1(n_426),
.B2(n_427),
.Y(n_602)
);

BUFx6f_ASAP7_75t_SL g603 ( 
.A(n_529),
.Y(n_603)
);

AO22x2_ASAP7_75t_L g604 ( 
.A1(n_545),
.A2(n_368),
.B1(n_377),
.B2(n_378),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_546),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_477),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_480),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_548),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_534),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_541),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_541),
.Y(n_611)
);

NAND2x1p5_ASAP7_75t_L g612 ( 
.A(n_493),
.B(n_426),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_470),
.B(n_426),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_500),
.B(n_498),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_520),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_498),
.B(n_426),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_470),
.Y(n_617)
);

AOI22x1_ASAP7_75t_L g618 ( 
.A1(n_498),
.A2(n_542),
.B1(n_530),
.B2(n_513),
.Y(n_618)
);

AO22x2_ASAP7_75t_L g619 ( 
.A1(n_501),
.A2(n_377),
.B1(n_378),
.B2(n_2),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_480),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_506),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_595),
.A2(n_510),
.B(n_522),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_593),
.A2(n_499),
.B1(n_503),
.B2(n_491),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_559),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_577),
.B(n_503),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_561),
.Y(n_626)
);

AO21x1_ASAP7_75t_L g627 ( 
.A1(n_585),
.A2(n_549),
.B(n_499),
.Y(n_627)
);

BUFx6f_ASAP7_75t_SL g628 ( 
.A(n_597),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_617),
.B(n_490),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_609),
.B(n_566),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_615),
.B(n_476),
.Y(n_632)
);

AO22x1_ASAP7_75t_L g633 ( 
.A1(n_600),
.A2(n_476),
.B1(n_512),
.B2(n_549),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_610),
.A2(n_522),
.B(n_510),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_580),
.B(n_476),
.Y(n_635)
);

O2A1O1Ixp5_ASAP7_75t_L g636 ( 
.A1(n_598),
.A2(n_542),
.B(n_517),
.C(n_518),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_580),
.B(n_547),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_556),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_563),
.B(n_515),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_574),
.B(n_506),
.Y(n_640)
);

AOI21xp5_ASAP7_75t_L g641 ( 
.A1(n_557),
.A2(n_521),
.B(n_533),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_564),
.B(n_514),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_573),
.B(n_552),
.Y(n_643)
);

OA22x2_ASAP7_75t_L g644 ( 
.A1(n_569),
.A2(n_550),
.B1(n_544),
.B2(n_519),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_576),
.B(n_519),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_571),
.A2(n_603),
.B1(n_554),
.B2(n_586),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_583),
.B(n_524),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_614),
.B(n_523),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_581),
.A2(n_543),
.B(n_525),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_614),
.B(n_542),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_584),
.A2(n_550),
.B1(n_544),
.B2(n_531),
.Y(n_651)
);

AOI21xp5_ASAP7_75t_L g652 ( 
.A1(n_613),
.A2(n_528),
.B(n_524),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_582),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_589),
.B(n_590),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_L g655 ( 
.A1(n_611),
.A2(n_528),
.B(n_531),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_594),
.B(n_599),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_605),
.B(n_426),
.Y(n_657)
);

OAI22xp5_ASAP7_75t_L g658 ( 
.A1(n_608),
.A2(n_427),
.B1(n_260),
.B2(n_253),
.Y(n_658)
);

NOR2x1p5_ASAP7_75t_SL g659 ( 
.A(n_562),
.B(n_378),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_554),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_603),
.A2(n_427),
.B1(n_244),
.B2(n_240),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_SL g662 ( 
.A1(n_560),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_616),
.A2(n_427),
.B(n_343),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_586),
.B(n_427),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_568),
.A2(n_343),
.B1(n_3),
.B2(n_4),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_616),
.A2(n_343),
.B(n_54),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_619),
.B(n_1),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_587),
.B(n_343),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_582),
.B(n_343),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_579),
.B(n_3),
.Y(n_670)
);

INVx3_ASAP7_75t_L g671 ( 
.A(n_555),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_565),
.A2(n_343),
.B(n_55),
.Y(n_672)
);

OAI21xp5_ASAP7_75t_L g673 ( 
.A1(n_592),
.A2(n_343),
.B(n_4),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_568),
.B(n_5),
.Y(n_674)
);

O2A1O1Ixp33_ASAP7_75t_SL g675 ( 
.A1(n_570),
.A2(n_5),
.B(n_6),
.C(n_7),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_606),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_575),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_677)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_575),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_620),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_567),
.A2(n_56),
.B(n_53),
.Y(n_680)
);

OAI22xp5_ASAP7_75t_L g681 ( 
.A1(n_567),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_618),
.A2(n_553),
.B(n_602),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_612),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_621),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_629),
.B(n_558),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_630),
.B(n_558),
.Y(n_686)
);

BUFx12f_ASAP7_75t_L g687 ( 
.A(n_653),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_673),
.A2(n_607),
.B(n_553),
.C(n_619),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_679),
.Y(n_689)
);

BUFx2_ASAP7_75t_L g690 ( 
.A(n_644),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_684),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_636),
.Y(n_692)
);

BUFx2_ASAP7_75t_SL g693 ( 
.A(n_628),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_644),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_645),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_667),
.A2(n_572),
.B1(n_578),
.B2(n_596),
.Y(n_696)
);

INVxp33_ASAP7_75t_SL g697 ( 
.A(n_637),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_623),
.B(n_572),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_647),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_674),
.B(n_660),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_636),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_655),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_631),
.B(n_578),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_624),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_625),
.B(n_596),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_626),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_646),
.A2(n_591),
.B1(n_588),
.B2(n_604),
.Y(n_707)
);

CKINVDCx20_ASAP7_75t_R g708 ( 
.A(n_640),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_676),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g710 ( 
.A(n_628),
.B(n_618),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_635),
.Y(n_711)
);

AND2x2_ASAP7_75t_L g712 ( 
.A(n_674),
.B(n_604),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_632),
.B(n_16),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_638),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g715 ( 
.A1(n_641),
.A2(n_649),
.B(n_622),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_648),
.B(n_588),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_661),
.Y(n_717)
);

AND2x2_ASAP7_75t_L g718 ( 
.A(n_639),
.B(n_650),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_650),
.B(n_601),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_634),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_648),
.B(n_591),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_683),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_657),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_654),
.B(n_601),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_656),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_670),
.B(n_18),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_629),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_633),
.B(n_18),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_664),
.A2(n_677),
.B1(n_642),
.B2(n_665),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_683),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_643),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_671),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_671),
.Y(n_733)
);

BUFx2_ASAP7_75t_R g734 ( 
.A(n_668),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_678),
.A2(n_681),
.B1(n_651),
.B2(n_672),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_678),
.B(n_627),
.Y(n_736)
);

BUFx12f_ASAP7_75t_L g737 ( 
.A(n_669),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_651),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_658),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_739)
);

BUFx6f_ASAP7_75t_L g740 ( 
.A(n_668),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_682),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_652),
.B(n_20),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_659),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_663),
.B(n_21),
.Y(n_744)
);

BUFx2_ASAP7_75t_L g745 ( 
.A(n_662),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_666),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_L g747 ( 
.A1(n_715),
.A2(n_680),
.B(n_675),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_735),
.A2(n_675),
.B(n_662),
.Y(n_748)
);

AO21x2_ASAP7_75t_L g749 ( 
.A1(n_736),
.A2(n_59),
.B(n_57),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_714),
.Y(n_750)
);

INVx1_ASAP7_75t_SL g751 ( 
.A(n_733),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_706),
.Y(n_752)
);

INVxp67_ASAP7_75t_L g753 ( 
.A(n_703),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_735),
.A2(n_22),
.B(n_23),
.Y(n_754)
);

INVx1_ASAP7_75t_SL g755 ( 
.A(n_733),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_694),
.B(n_60),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_SL g757 ( 
.A1(n_698),
.A2(n_23),
.B(n_24),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_714),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_685),
.B(n_733),
.Y(n_759)
);

OR2x2_ASAP7_75t_SL g760 ( 
.A(n_728),
.B(n_25),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_727),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_689),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_734),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_685),
.B(n_26),
.Y(n_764)
);

NAND2x1p5_ASAP7_75t_L g765 ( 
.A(n_685),
.B(n_61),
.Y(n_765)
);

BUFx2_ASAP7_75t_L g766 ( 
.A(n_708),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_687),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_746),
.A2(n_27),
.B(n_28),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_718),
.B(n_27),
.Y(n_769)
);

BUFx5_ASAP7_75t_L g770 ( 
.A(n_702),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_718),
.B(n_28),
.Y(n_771)
);

INVx5_ASAP7_75t_L g772 ( 
.A(n_737),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_685),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_700),
.B(n_29),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_689),
.Y(n_775)
);

NAND2x1p5_ASAP7_75t_L g776 ( 
.A(n_722),
.B(n_63),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_687),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_722),
.B(n_29),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_687),
.Y(n_779)
);

INVx3_ASAP7_75t_L g780 ( 
.A(n_737),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_745),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_697),
.B(n_30),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_691),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_691),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_704),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_692),
.A2(n_31),
.B(n_32),
.Y(n_786)
);

AND2x4_ASAP7_75t_L g787 ( 
.A(n_722),
.B(n_33),
.Y(n_787)
);

AOI21xp5_ASAP7_75t_L g788 ( 
.A1(n_692),
.A2(n_34),
.B(n_35),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_700),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_732),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_725),
.B(n_35),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_717),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_692),
.A2(n_36),
.B(n_39),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_712),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_725),
.B(n_40),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_745),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_796)
);

AOI21xp5_ASAP7_75t_L g797 ( 
.A1(n_701),
.A2(n_43),
.B(n_44),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_739),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_798)
);

INVxp67_ASAP7_75t_SL g799 ( 
.A(n_731),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_737),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_710),
.B(n_45),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_731),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_732),
.Y(n_803)
);

INVx1_ASAP7_75t_SL g804 ( 
.A(n_732),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_701),
.A2(n_46),
.B(n_47),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_704),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_722),
.B(n_48),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_706),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_706),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_711),
.Y(n_810)
);

INVx3_ASAP7_75t_SL g811 ( 
.A(n_726),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_709),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_729),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_710),
.B(n_51),
.Y(n_814)
);

INVx5_ASAP7_75t_L g815 ( 
.A(n_711),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_701),
.A2(n_52),
.B(n_210),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_686),
.B(n_52),
.Y(n_817)
);

AND2x2_ASAP7_75t_SL g818 ( 
.A(n_764),
.B(n_690),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_789),
.B(n_731),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_771),
.B(n_695),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_750),
.Y(n_821)
);

O2A1O1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_813),
.A2(n_728),
.B(n_688),
.C(n_713),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_774),
.B(n_712),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_772),
.Y(n_824)
);

OA21x2_ASAP7_75t_L g825 ( 
.A1(n_747),
.A2(n_741),
.B(n_707),
.Y(n_825)
);

NOR2x1_ASAP7_75t_L g826 ( 
.A(n_780),
.B(n_693),
.Y(n_826)
);

CKINVDCx20_ASAP7_75t_R g827 ( 
.A(n_779),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_773),
.B(n_719),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_759),
.B(n_719),
.Y(n_829)
);

AND2x4_ASAP7_75t_L g830 ( 
.A(n_759),
.B(n_690),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_794),
.A2(n_813),
.B1(n_748),
.B2(n_760),
.Y(n_831)
);

O2A1O1Ixp5_ASAP7_75t_L g832 ( 
.A1(n_754),
.A2(n_744),
.B(n_742),
.C(n_705),
.Y(n_832)
);

OR2x6_ASAP7_75t_L g833 ( 
.A(n_810),
.B(n_721),
.Y(n_833)
);

O2A1O1Ixp5_ASAP7_75t_L g834 ( 
.A1(n_798),
.A2(n_742),
.B(n_716),
.C(n_720),
.Y(n_834)
);

A2O1A1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_768),
.A2(n_696),
.B(n_738),
.C(n_721),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_764),
.B(n_694),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_758),
.B(n_695),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_751),
.A2(n_720),
.B(n_724),
.Y(n_838)
);

NOR2x2_ASAP7_75t_L g839 ( 
.A(n_767),
.B(n_693),
.Y(n_839)
);

OR2x6_ASAP7_75t_L g840 ( 
.A(n_765),
.B(n_740),
.Y(n_840)
);

AOI21x1_ASAP7_75t_SL g841 ( 
.A1(n_778),
.A2(n_724),
.B(n_740),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_751),
.A2(n_755),
.B(n_816),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_755),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_762),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_775),
.B(n_738),
.Y(n_845)
);

NAND2x1p5_ASAP7_75t_L g846 ( 
.A(n_772),
.B(n_711),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_SL g847 ( 
.A1(n_782),
.A2(n_743),
.B(n_730),
.C(n_723),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_749),
.A2(n_723),
.B(n_740),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_803),
.B(n_740),
.Y(n_849)
);

OR2x2_ASAP7_75t_L g850 ( 
.A(n_783),
.B(n_699),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_802),
.B(n_699),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_766),
.B(n_711),
.Y(n_852)
);

AND2x4_ASAP7_75t_L g853 ( 
.A(n_772),
.B(n_740),
.Y(n_853)
);

OA21x2_ASAP7_75t_L g854 ( 
.A1(n_786),
.A2(n_702),
.B(n_743),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_795),
.B(n_711),
.Y(n_855)
);

AOI211xp5_ASAP7_75t_L g856 ( 
.A1(n_781),
.A2(n_711),
.B(n_740),
.C(n_730),
.Y(n_856)
);

OR2x6_ASAP7_75t_SL g857 ( 
.A(n_769),
.B(n_730),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_784),
.B(n_723),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_794),
.A2(n_792),
.B1(n_798),
.B2(n_817),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_790),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_785),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_SL g862 ( 
.A1(n_788),
.A2(n_797),
.B(n_793),
.C(n_805),
.Y(n_862)
);

NAND2x1p5_ASAP7_75t_L g863 ( 
.A(n_780),
.B(n_709),
.Y(n_863)
);

INVx3_ASAP7_75t_SL g864 ( 
.A(n_761),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_L g865 ( 
.A1(n_801),
.A2(n_743),
.B(n_709),
.C(n_66),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_814),
.A2(n_64),
.B(n_65),
.C(n_68),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_799),
.B(n_209),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_790),
.B(n_69),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_778),
.B(n_70),
.Y(n_869)
);

O2A1O1Ixp5_ASAP7_75t_L g870 ( 
.A1(n_796),
.A2(n_71),
.B(n_73),
.C(n_74),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_806),
.Y(n_871)
);

O2A1O1Ixp5_ASAP7_75t_L g872 ( 
.A1(n_791),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_872)
);

AOI221xp5_ASAP7_75t_L g873 ( 
.A1(n_757),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_873)
);

AND2x2_ASAP7_75t_SL g874 ( 
.A(n_800),
.B(n_787),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_753),
.A2(n_83),
.B(n_85),
.C(n_86),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_804),
.B(n_770),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_752),
.Y(n_877)
);

OR2x2_ASAP7_75t_L g878 ( 
.A(n_804),
.B(n_763),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_815),
.B(n_87),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_787),
.B(n_88),
.Y(n_880)
);

HB1xp67_ASAP7_75t_L g881 ( 
.A(n_815),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_808),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_812),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_763),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_807),
.A2(n_89),
.B(n_93),
.C(n_94),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_809),
.B(n_95),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_SL g887 ( 
.A1(n_831),
.A2(n_756),
.B1(n_749),
.B2(n_815),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_831),
.A2(n_811),
.B1(n_807),
.B2(n_777),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_821),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_820),
.B(n_770),
.Y(n_890)
);

INVx5_ASAP7_75t_SL g891 ( 
.A(n_840),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_SL g892 ( 
.A1(n_859),
.A2(n_756),
.B1(n_770),
.B2(n_776),
.Y(n_892)
);

HB1xp67_ASAP7_75t_L g893 ( 
.A(n_843),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_859),
.A2(n_756),
.B1(n_770),
.B2(n_100),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_823),
.A2(n_756),
.B1(n_770),
.B2(n_101),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_819),
.B(n_208),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_878),
.B(n_844),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_877),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_L g899 ( 
.A1(n_836),
.A2(n_97),
.B1(n_99),
.B2(n_102),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_822),
.A2(n_103),
.B(n_104),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_852),
.B(n_829),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_824),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_828),
.B(n_207),
.Y(n_903)
);

AOI22xp33_ASAP7_75t_L g904 ( 
.A1(n_818),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_825),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_905)
);

INVx6_ASAP7_75t_L g906 ( 
.A(n_824),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_882),
.Y(n_907)
);

OR2x2_ASAP7_75t_SL g908 ( 
.A(n_839),
.B(n_115),
.Y(n_908)
);

BUFx3_ASAP7_75t_L g909 ( 
.A(n_824),
.Y(n_909)
);

INVx4_ASAP7_75t_L g910 ( 
.A(n_874),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_834),
.B(n_116),
.C(n_117),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_883),
.Y(n_912)
);

AOI22xp33_ASAP7_75t_L g913 ( 
.A1(n_825),
.A2(n_884),
.B1(n_873),
.B2(n_855),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_827),
.Y(n_914)
);

INVx3_ASAP7_75t_L g915 ( 
.A(n_849),
.Y(n_915)
);

AOI22xp33_ASAP7_75t_L g916 ( 
.A1(n_838),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_861),
.Y(n_917)
);

BUFx5_ASAP7_75t_L g918 ( 
.A(n_853),
.Y(n_918)
);

NOR3xp33_ASAP7_75t_SL g919 ( 
.A(n_880),
.B(n_122),
.C(n_123),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_830),
.B(n_124),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_871),
.Y(n_921)
);

AOI22xp33_ASAP7_75t_L g922 ( 
.A1(n_854),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_850),
.Y(n_923)
);

INVx1_ASAP7_75t_SL g924 ( 
.A(n_864),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_830),
.B(n_129),
.Y(n_925)
);

OAI22xp5_ASAP7_75t_L g926 ( 
.A1(n_835),
.A2(n_130),
.B1(n_133),
.B2(n_136),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_851),
.Y(n_927)
);

INVx8_ASAP7_75t_L g928 ( 
.A(n_840),
.Y(n_928)
);

BUFx2_ASAP7_75t_L g929 ( 
.A(n_881),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_851),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_837),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_858),
.Y(n_932)
);

OAI21xp5_ASAP7_75t_SL g933 ( 
.A1(n_869),
.A2(n_137),
.B(n_140),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_856),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_SL g935 ( 
.A1(n_856),
.A2(n_826),
.B1(n_840),
.B2(n_857),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_901),
.B(n_876),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_907),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_915),
.B(n_876),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_893),
.B(n_860),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_924),
.B(n_863),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_907),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_912),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_912),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_933),
.A2(n_900),
.B(n_913),
.C(n_887),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_909),
.Y(n_945)
);

AO32x1_ASAP7_75t_L g946 ( 
.A1(n_888),
.A2(n_847),
.A3(n_841),
.B1(n_833),
.B2(n_848),
.Y(n_946)
);

AND2x4_ASAP7_75t_L g947 ( 
.A(n_915),
.B(n_849),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_929),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_889),
.Y(n_949)
);

NAND2x1_ASAP7_75t_L g950 ( 
.A(n_910),
.B(n_906),
.Y(n_950)
);

NOR2x1_ASAP7_75t_SL g951 ( 
.A(n_910),
.B(n_833),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_913),
.A2(n_865),
.B(n_862),
.C(n_875),
.Y(n_952)
);

AO21x2_ASAP7_75t_L g953 ( 
.A1(n_911),
.A2(n_842),
.B(n_867),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_898),
.Y(n_954)
);

OR2x2_ASAP7_75t_L g955 ( 
.A(n_897),
.B(n_923),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_894),
.A2(n_885),
.B(n_870),
.C(n_872),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_890),
.A2(n_867),
.B(n_868),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_915),
.B(n_833),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_928),
.B(n_853),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_898),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_909),
.B(n_845),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_927),
.B(n_854),
.Y(n_962)
);

OR2x2_ASAP7_75t_L g963 ( 
.A(n_930),
.B(n_868),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_917),
.B(n_832),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_931),
.B(n_910),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_894),
.A2(n_866),
.B(n_879),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_951),
.B(n_902),
.Y(n_967)
);

AOI22xp33_ASAP7_75t_L g968 ( 
.A1(n_966),
.A2(n_953),
.B1(n_926),
.B2(n_905),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_962),
.Y(n_969)
);

OR2x2_ASAP7_75t_L g970 ( 
.A(n_955),
.B(n_932),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_966),
.A2(n_905),
.B1(n_892),
.B2(n_895),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_955),
.B(n_921),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_962),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_964),
.B(n_935),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_949),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_948),
.B(n_918),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_951),
.B(n_902),
.Y(n_977)
);

NAND2x1p5_ASAP7_75t_L g978 ( 
.A(n_950),
.B(n_934),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_949),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_953),
.A2(n_895),
.B1(n_899),
.B2(n_904),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_944),
.A2(n_899),
.B1(n_904),
.B2(n_916),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_937),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_937),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_964),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_948),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_942),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_941),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_942),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_984),
.A2(n_974),
.B(n_985),
.Y(n_989)
);

A2O1A1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_981),
.A2(n_968),
.B(n_980),
.C(n_971),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_L g991 ( 
.A(n_984),
.B(n_952),
.C(n_963),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_978),
.A2(n_940),
.B(n_939),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_975),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_979),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_985),
.Y(n_995)
);

NAND4xp25_ASAP7_75t_L g996 ( 
.A(n_976),
.B(n_948),
.C(n_956),
.D(n_965),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_978),
.A2(n_946),
.B(n_950),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_970),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_970),
.B(n_936),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_976),
.B(n_936),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_969),
.A2(n_919),
.B(n_916),
.C(n_922),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_969),
.B(n_965),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_986),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_972),
.Y(n_1004)
);

NAND3xp33_ASAP7_75t_SL g1005 ( 
.A(n_978),
.B(n_963),
.C(n_914),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_993),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_995),
.B(n_967),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_989),
.B(n_967),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_990),
.B(n_973),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_1003),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_994),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_990),
.B(n_973),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_998),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1000),
.B(n_967),
.Y(n_1014)
);

OR2x2_ASAP7_75t_L g1015 ( 
.A(n_1004),
.B(n_972),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_1003),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_991),
.B(n_977),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_1006),
.B(n_999),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_1006),
.B(n_1000),
.Y(n_1019)
);

NOR4xp25_ASAP7_75t_L g1020 ( 
.A(n_1009),
.B(n_996),
.C(n_1005),
.D(n_1001),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_1011),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_1013),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_1012),
.B(n_992),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_1017),
.B(n_997),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_1017),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1014),
.Y(n_1026)
);

AOI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_1023),
.A2(n_1017),
.B1(n_1001),
.B2(n_1008),
.Y(n_1027)
);

OAI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_1020),
.A2(n_1008),
.B(n_1007),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1021),
.Y(n_1029)
);

OAI211xp5_ASAP7_75t_L g1030 ( 
.A1(n_1025),
.A2(n_1014),
.B(n_914),
.C(n_1015),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_1025),
.B(n_1007),
.Y(n_1031)
);

NAND2xp33_ASAP7_75t_SL g1032 ( 
.A(n_1024),
.B(n_1007),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1027),
.A2(n_1026),
.B1(n_1019),
.B2(n_1018),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1030),
.B(n_1022),
.Y(n_1034)
);

AOI22xp33_ASAP7_75t_L g1035 ( 
.A1(n_1028),
.A2(n_953),
.B1(n_1016),
.B2(n_1010),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_1031),
.B(n_1015),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_1029),
.B(n_1002),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1032),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_1032),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1031),
.B(n_977),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_1029),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_1029),
.Y(n_1042)
);

XNOR2x1_ASAP7_75t_L g1043 ( 
.A(n_1039),
.B(n_920),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1036),
.B(n_1016),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_1041),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1041),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_1042),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1042),
.B(n_1010),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_1038),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_1037),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1050),
.B(n_1049),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_1044),
.B(n_1033),
.Y(n_1052)
);

AOI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1043),
.A2(n_1035),
.B1(n_1034),
.B2(n_1040),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1049),
.B(n_982),
.Y(n_1054)
);

CKINVDCx14_ASAP7_75t_R g1055 ( 
.A(n_1049),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1047),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1045),
.B(n_983),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_1055),
.B(n_1046),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_SL g1059 ( 
.A(n_1052),
.B(n_1056),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1051),
.Y(n_1060)
);

NAND3xp33_ASAP7_75t_L g1061 ( 
.A(n_1053),
.B(n_1048),
.C(n_922),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1054),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1059),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1058),
.B(n_1057),
.Y(n_1064)
);

INVx1_ASAP7_75t_SL g1065 ( 
.A(n_1060),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1062),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_1061),
.B(n_908),
.Y(n_1067)
);

INVxp67_ASAP7_75t_SL g1068 ( 
.A(n_1059),
.Y(n_1068)
);

AND2x2_ASAP7_75t_L g1069 ( 
.A(n_1068),
.B(n_977),
.Y(n_1069)
);

AOI221xp5_ASAP7_75t_L g1070 ( 
.A1(n_1067),
.A2(n_953),
.B1(n_987),
.B2(n_896),
.C(n_903),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_1063),
.B(n_945),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1066),
.A2(n_957),
.B1(n_925),
.B2(n_986),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1065),
.A2(n_957),
.B1(n_988),
.B2(n_945),
.Y(n_1073)
);

AOI211xp5_ASAP7_75t_L g1074 ( 
.A1(n_1064),
.A2(n_879),
.B(n_945),
.C(n_946),
.Y(n_1074)
);

AOI221xp5_ASAP7_75t_L g1075 ( 
.A1(n_1069),
.A2(n_988),
.B1(n_946),
.B2(n_943),
.C(n_941),
.Y(n_1075)
);

AOI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_1071),
.A2(n_957),
.B(n_886),
.Y(n_1076)
);

BUFx4f_ASAP7_75t_L g1077 ( 
.A(n_1070),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_1073),
.B(n_945),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1072),
.B(n_957),
.Y(n_1079)
);

INVx1_ASAP7_75t_SL g1080 ( 
.A(n_1074),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1069),
.B(n_945),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1069),
.B(n_961),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_1080),
.B(n_961),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1082),
.Y(n_1084)
);

OAI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_1081),
.A2(n_945),
.B(n_938),
.Y(n_1085)
);

NOR2x1_ASAP7_75t_L g1086 ( 
.A(n_1078),
.B(n_961),
.Y(n_1086)
);

NOR2x1_ASAP7_75t_L g1087 ( 
.A(n_1079),
.B(n_1077),
.Y(n_1087)
);

NOR4xp75_ASAP7_75t_L g1088 ( 
.A(n_1075),
.B(n_938),
.C(n_946),
.D(n_958),
.Y(n_1088)
);

NAND4xp25_ASAP7_75t_L g1089 ( 
.A(n_1076),
.B(n_961),
.C(n_958),
.D(n_947),
.Y(n_1089)
);

XNOR2xp5_ASAP7_75t_L g1090 ( 
.A(n_1080),
.B(n_846),
.Y(n_1090)
);

XNOR2xp5_ASAP7_75t_L g1091 ( 
.A(n_1090),
.B(n_959),
.Y(n_1091)
);

NOR2x1_ASAP7_75t_L g1092 ( 
.A(n_1084),
.B(n_959),
.Y(n_1092)
);

OAI211xp5_ASAP7_75t_SL g1093 ( 
.A1(n_1087),
.A2(n_946),
.B(n_943),
.C(n_146),
.Y(n_1093)
);

NOR3x1_ASAP7_75t_L g1094 ( 
.A(n_1083),
.B(n_906),
.C(n_145),
.Y(n_1094)
);

NAND4xp25_ASAP7_75t_L g1095 ( 
.A(n_1086),
.B(n_947),
.C(n_906),
.D(n_148),
.Y(n_1095)
);

NOR2x1_ASAP7_75t_L g1096 ( 
.A(n_1089),
.B(n_959),
.Y(n_1096)
);

NAND4xp75_ASAP7_75t_L g1097 ( 
.A(n_1088),
.B(n_942),
.C(n_147),
.D(n_149),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1085),
.A2(n_947),
.B1(n_954),
.B2(n_960),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1086),
.B(n_947),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_1094),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_1099),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1097),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1092),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1095),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1096),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_1091),
.B(n_918),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_1098),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1093),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1097),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1097),
.Y(n_1110)
);

NOR2xp67_ASAP7_75t_L g1111 ( 
.A(n_1095),
.B(n_144),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1094),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1100),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1108),
.A2(n_960),
.B1(n_954),
.B2(n_959),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1112),
.B(n_1111),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_1112),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1103),
.Y(n_1117)
);

OAI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1104),
.A2(n_959),
.B1(n_954),
.B2(n_960),
.C(n_154),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1101),
.A2(n_891),
.B1(n_928),
.B2(n_918),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_1105),
.B(n_150),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1102),
.B(n_152),
.Y(n_1121)
);

OAI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1116),
.A2(n_1110),
.B1(n_1109),
.B2(n_1107),
.C(n_1106),
.Y(n_1122)
);

AOI211xp5_ASAP7_75t_L g1123 ( 
.A1(n_1117),
.A2(n_153),
.B(n_155),
.C(n_156),
.Y(n_1123)
);

NAND2x1_ASAP7_75t_L g1124 ( 
.A(n_1113),
.B(n_159),
.Y(n_1124)
);

OAI211xp5_ASAP7_75t_L g1125 ( 
.A1(n_1115),
.A2(n_161),
.B(n_162),
.C(n_163),
.Y(n_1125)
);

XOR2x2_ASAP7_75t_L g1126 ( 
.A(n_1121),
.B(n_164),
.Y(n_1126)
);

AOI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_1120),
.A2(n_167),
.B(n_170),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1122),
.A2(n_1118),
.B1(n_1119),
.B2(n_1114),
.Y(n_1128)
);

AOI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1126),
.A2(n_918),
.B1(n_928),
.B2(n_891),
.Y(n_1129)
);

NAND5xp2_ASAP7_75t_L g1130 ( 
.A(n_1123),
.B(n_171),
.C(n_172),
.D(n_173),
.E(n_174),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_SL g1131 ( 
.A1(n_1128),
.A2(n_1124),
.B1(n_1127),
.B2(n_1125),
.Y(n_1131)
);

OAI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_1131),
.A2(n_1129),
.B1(n_1130),
.B2(n_891),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1132),
.A2(n_175),
.B(n_176),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1132),
.B(n_181),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1134),
.Y(n_1135)
);

OAI222xp33_ASAP7_75t_L g1136 ( 
.A1(n_1133),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.C1(n_186),
.C2(n_188),
.Y(n_1136)
);

OAI322xp33_ASAP7_75t_L g1137 ( 
.A1(n_1134),
.A2(n_189),
.A3(n_190),
.B1(n_191),
.B2(n_192),
.C1(n_195),
.C2(n_196),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1135),
.B(n_928),
.Y(n_1138)
);

INVxp33_ASAP7_75t_L g1139 ( 
.A(n_1136),
.Y(n_1139)
);

AOI221xp5_ASAP7_75t_L g1140 ( 
.A1(n_1139),
.A2(n_1137),
.B1(n_198),
.B2(n_199),
.C(n_200),
.Y(n_1140)
);

AOI211xp5_ASAP7_75t_L g1141 ( 
.A1(n_1140),
.A2(n_1138),
.B(n_201),
.C(n_203),
.Y(n_1141)
);


endmodule