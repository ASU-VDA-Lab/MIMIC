module fake_jpeg_8619_n_314 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_314);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx5_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_38),
.Y(n_45)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_19),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_24),
.Y(n_50)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_16),
.B1(n_31),
.B2(n_17),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_51),
.B1(n_67),
.B2(n_19),
.Y(n_80)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_59),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_39),
.A2(n_30),
.B1(n_17),
.B2(n_27),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_R g53 ( 
.A(n_35),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_20),
.Y(n_73)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_19),
.B1(n_20),
.B2(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_25),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_68),
.Y(n_87)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_42),
.A2(n_31),
.B1(n_24),
.B2(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_69),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_61),
.A2(n_38),
.B1(n_42),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_74),
.A2(n_62),
.B1(n_52),
.B2(n_48),
.Y(n_104)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_77),
.B(n_93),
.Y(n_109)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_78),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_79),
.A2(n_81),
.B1(n_22),
.B2(n_24),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_80),
.A2(n_68),
.B1(n_29),
.B2(n_21),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_50),
.A2(n_42),
.B1(n_38),
.B2(n_20),
.Y(n_81)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_64),
.A2(n_28),
.B(n_32),
.C(n_34),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g121 ( 
.A1(n_88),
.A2(n_28),
.B(n_32),
.C(n_47),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_90),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_21),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_45),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_65),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_96),
.A2(n_115),
.B1(n_22),
.B2(n_26),
.Y(n_132)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_101),
.B(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_104),
.A2(n_111),
.B1(n_71),
.B2(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_51),
.B(n_53),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_105),
.A2(n_113),
.B(n_36),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_106),
.B(n_119),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_91),
.A2(n_49),
.B1(n_46),
.B2(n_54),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_38),
.B1(n_48),
.B2(n_52),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_57),
.B1(n_55),
.B2(n_36),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_46),
.B1(n_60),
.B2(n_58),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_117),
.B(n_85),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_62),
.B1(n_44),
.B2(n_40),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_45),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_116),
.Y(n_124)
);

AO21x2_ASAP7_75t_SL g113 ( 
.A1(n_73),
.A2(n_40),
.B(n_38),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_44),
.B1(n_21),
.B2(n_26),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_56),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_56),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_60),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_85),
.C(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_127),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_135),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_147),
.B1(n_139),
.B2(n_131),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_128),
.B(n_136),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_90),
.A3(n_70),
.B1(n_86),
.B2(n_36),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_131),
.B(n_120),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g130 ( 
.A(n_113),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_130),
.Y(n_153)
);

AOI221xp5_ASAP7_75t_L g158 ( 
.A1(n_132),
.A2(n_145),
.B1(n_103),
.B2(n_141),
.C(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_139),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_71),
.B1(n_48),
.B2(n_84),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_134),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_75),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_75),
.C(n_89),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_78),
.B1(n_72),
.B2(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_69),
.B1(n_40),
.B2(n_82),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_113),
.A2(n_94),
.B1(n_72),
.B2(n_22),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_116),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_133),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_140),
.B(n_146),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_70),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_120),
.Y(n_167)
);

AND2x6_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_114),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_151),
.B1(n_160),
.B2(n_123),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_111),
.B1(n_115),
.B2(n_104),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_111),
.B1(n_122),
.B2(n_121),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_158),
.B1(n_165),
.B2(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_154),
.B(n_161),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_114),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_156),
.B(n_164),
.Y(n_176)
);

OAI22x1_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_117),
.B1(n_114),
.B2(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_138),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_170),
.B(n_173),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_130),
.A2(n_111),
.B1(n_96),
.B2(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_166),
.B(n_168),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_118),
.B1(n_97),
.B2(n_98),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_127),
.B(n_99),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_171),
.B(n_174),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_143),
.A2(n_145),
.B(n_144),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_99),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_136),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_180),
.C(n_200),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_167),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_190),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_128),
.C(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_163),
.A2(n_142),
.B1(n_132),
.B2(n_144),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_187),
.A2(n_188),
.B1(n_153),
.B2(n_156),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_163),
.A2(n_123),
.B1(n_98),
.B2(n_147),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_165),
.B1(n_151),
.B2(n_152),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_153),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_192),
.Y(n_207)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_97),
.B(n_118),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_154),
.B(n_127),
.Y(n_194)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_195),
.B(n_197),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_102),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_196),
.B(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_102),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_55),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_162),
.B(n_94),
.C(n_57),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_201),
.Y(n_242)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_149),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_215),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_213),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_151),
.B1(n_153),
.B2(n_57),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_192),
.B1(n_176),
.B2(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_211),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_151),
.C(n_55),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_218),
.C(n_219),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_214),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_184),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_23),
.C(n_1),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_23),
.C(n_1),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_184),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_220),
.B(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_23),
.C(n_2),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_191),
.B(n_23),
.Y(n_224)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_224),
.Y(n_230)
);

INVxp33_ASAP7_75t_SL g225 ( 
.A(n_223),
.Y(n_225)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_225),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_193),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_226),
.B(n_234),
.Y(n_253)
);

NOR2x1_ASAP7_75t_L g228 ( 
.A(n_205),
.B(n_199),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_240),
.C(n_244),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_183),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_215),
.B(n_189),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_212),
.C(n_210),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_185),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_238),
.B(n_239),
.Y(n_248)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_204),
.A2(n_189),
.B(n_197),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_208),
.A2(n_189),
.B(n_190),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_241),
.A2(n_206),
.B(n_216),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_188),
.B1(n_187),
.B2(n_198),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_243),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_23),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_258),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_214),
.Y(n_247)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_249),
.A2(n_255),
.B(n_237),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_217),
.B(n_216),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_251),
.A2(n_229),
.B(n_244),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_230),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_252),
.Y(n_262)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_228),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_259),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_241),
.A2(n_210),
.B(n_221),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_231),
.B(n_219),
.C(n_218),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_260),
.C(n_237),
.Y(n_271)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_257),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_226),
.B(n_14),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_15),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_261),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_231),
.C(n_234),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_SL g278 ( 
.A(n_263),
.B(n_256),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_243),
.B1(n_240),
.B2(n_235),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_251),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_249),
.Y(n_277)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_273),
.C(n_260),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_233),
.C(n_13),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_258),
.C(n_250),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_253),
.B(n_255),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_261),
.Y(n_281)
);

NOR2xp67_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_246),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_277),
.B(n_278),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_248),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_279),
.B(n_281),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_0),
.C(n_3),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_11),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_0),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_270),
.C(n_273),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_290),
.B(n_294),
.C(n_7),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_264),
.A3(n_267),
.B1(n_265),
.B2(n_263),
.C1(n_270),
.C2(n_266),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_291),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

INVxp33_ASAP7_75t_SL g292 ( 
.A(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_283),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_7),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_266),
.C(n_4),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_296),
.B(n_6),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_288),
.A2(n_283),
.B(n_285),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_300),
.C(n_303),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_295),
.B(n_291),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_298),
.A2(n_7),
.B(n_8),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_299),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_288),
.A2(n_5),
.B(n_6),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_302),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_302),
.B(n_304),
.Y(n_307)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_10),
.B(n_8),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_309),
.A2(n_8),
.B(n_9),
.Y(n_310)
);

A2O1A1Ixp33_ASAP7_75t_SL g312 ( 
.A1(n_310),
.A2(n_311),
.B(n_9),
.C(n_10),
.Y(n_312)
);

O2A1O1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_312),
.A2(n_308),
.B(n_305),
.C(n_306),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_10),
.Y(n_314)
);


endmodule