module fake_jpeg_29633_n_247 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_7),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_31),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_40),
.B(n_42),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_20),
.B(n_15),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_13),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_49),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_25),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_32),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_22),
.B(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_57),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_36),
.Y(n_73)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_22),
.B(n_12),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_12),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_63),
.Y(n_91)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

AO22x1_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_17),
.B1(n_32),
.B2(n_24),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_93),
.B(n_62),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_90),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_18),
.C(n_34),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_75),
.B(n_3),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_78),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_63),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_40),
.A2(n_18),
.B1(n_34),
.B2(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_82),
.A2(n_85),
.B1(n_87),
.B2(n_3),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_83),
.B(n_98),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_27),
.B1(n_24),
.B2(n_29),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_38),
.A2(n_37),
.B1(n_33),
.B2(n_29),
.Y(n_87)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_28),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_49),
.A2(n_28),
.B(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_45),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_27),
.B1(n_1),
.B2(n_2),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_97),
.A2(n_61),
.B1(n_56),
.B2(n_45),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_41),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_7),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_101),
.B(n_105),
.Y(n_153)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

INVx2_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_53),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_106),
.B(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_109),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_27),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

BUFx4f_ASAP7_75t_SL g113 ( 
.A(n_66),
.Y(n_113)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_47),
.B1(n_43),
.B2(n_4),
.Y(n_114)
);

AO22x1_ASAP7_75t_L g133 ( 
.A1(n_114),
.A2(n_87),
.B1(n_70),
.B2(n_69),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_0),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_124),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_91),
.B(n_0),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_116),
.B(n_118),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_117),
.A2(n_126),
.B1(n_71),
.B2(n_99),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_120),
.Y(n_148)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_6),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_74),
.B(n_92),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_8),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_97),
.A2(n_85),
.B1(n_68),
.B2(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_129),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_79),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_133),
.A2(n_137),
.B1(n_129),
.B2(n_123),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_143),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_115),
.B(n_70),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_65),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_104),
.A2(n_92),
.B1(n_74),
.B2(n_65),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_127),
.B1(n_123),
.B2(n_108),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_154),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_126),
.A2(n_118),
.B(n_101),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_122),
.B(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_114),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_155),
.B(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_142),
.B(n_102),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_163),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g159 ( 
.A1(n_133),
.A2(n_105),
.B1(n_114),
.B2(n_103),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_159),
.A2(n_161),
.B1(n_157),
.B2(n_156),
.Y(n_195)
);

XNOR2x1_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_105),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_160),
.B(n_165),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_178),
.B(n_137),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_176),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_135),
.B(n_131),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_149),
.B(n_128),
.C(n_121),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_173),
.C(n_156),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_167),
.B(n_141),
.Y(n_180)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_136),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_170),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_113),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g172 ( 
.A(n_157),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_113),
.C(n_151),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_155),
.A2(n_140),
.B1(n_133),
.B2(n_153),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g177 ( 
.A(n_153),
.B(n_138),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_148),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_145),
.A2(n_144),
.B(n_141),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_132),
.Y(n_179)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_179),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_180),
.A2(n_195),
.B1(n_167),
.B2(n_152),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_186),
.B(n_174),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_194),
.Y(n_208)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_189),
.Y(n_205)
);

OR2x2_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_150),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_190),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_177),
.B(n_147),
.Y(n_210)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_173),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_204),
.C(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_200),
.B(n_202),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_185),
.B(n_134),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_183),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_197),
.A2(n_170),
.B1(n_160),
.B2(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_203),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_165),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_178),
.C(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_162),
.Y(n_207)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_209),
.B(n_210),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_193),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_212),
.B(n_219),
.C(n_204),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_209),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_188),
.C(n_190),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_208),
.B(n_181),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_221),
.B(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_223),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_203),
.B1(n_191),
.B2(n_182),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_181),
.B1(n_210),
.B2(n_197),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_224),
.B(n_215),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_207),
.B(n_182),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_225),
.A2(n_226),
.B(n_213),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_218),
.A2(n_211),
.B(n_205),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_219),
.A2(n_180),
.B(n_200),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_214),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_212),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_233),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_232),
.A2(n_234),
.A3(n_225),
.B1(n_223),
.B2(n_228),
.C1(n_216),
.C2(n_184),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_214),
.C(n_187),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_235),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_139),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_232),
.A2(n_172),
.B1(n_180),
.B2(n_184),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_238),
.A2(n_230),
.B(n_147),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_139),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_189),
.B(n_172),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_243),
.A2(n_238),
.B(n_236),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g246 ( 
.A(n_245),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_244),
.Y(n_247)
);


endmodule