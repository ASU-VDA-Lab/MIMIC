module fake_jpeg_27420_n_129 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_129);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_129;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

OAI21xp33_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_30),
.B(n_4),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_18),
.B(n_1),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_21),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_15),
.A2(n_2),
.B1(n_4),
.B2(n_8),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_24),
.B1(n_20),
.B2(n_23),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

OA22x2_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_22),
.B1(n_17),
.B2(n_27),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_45),
.A2(n_46),
.B1(n_35),
.B2(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_47),
.B(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_48),
.B(n_13),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_24),
.B1(n_23),
.B2(n_21),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_19),
.B(n_13),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_20),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_8),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_25),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_54),
.B(n_19),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_SL g77 ( 
.A(n_56),
.B(n_57),
.C(n_67),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_16),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_17),
.B1(n_26),
.B2(n_27),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_45),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_17),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_62),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_52),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_65),
.Y(n_82)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_69),
.Y(n_85)
);

OR2x2_ASAP7_75t_SL g67 ( 
.A(n_48),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_25),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_74),
.B(n_57),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_81),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_80),
.B(n_56),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_54),
.B(n_43),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_44),
.C(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_44),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_77),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_80),
.B(n_71),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_92),
.B(n_95),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_85),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_71),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_58),
.B1(n_77),
.B2(n_74),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_100),
.A2(n_103),
.B(n_104),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_76),
.B(n_41),
.Y(n_103)
);

XNOR2x1_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_45),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_84),
.B(n_45),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_105),
.A2(n_92),
.B(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_111),
.Y(n_118)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_114),
.B(n_75),
.Y(n_117)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_93),
.A3(n_96),
.B1(n_86),
.B2(n_26),
.C(n_9),
.Y(n_112)
);

AOI221xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_41),
.B1(n_26),
.B2(n_11),
.C(n_9),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_113),
.A2(n_102),
.B1(n_101),
.B2(n_68),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_94),
.B(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_117),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_11),
.B(n_4),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_119),
.B(n_31),
.C(n_40),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_119),
.B(n_40),
.C(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_120),
.B(n_122),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_118),
.B(n_117),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

OAI31xp33_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_68),
.A3(n_49),
.B(n_40),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_SL g128 ( 
.A1(n_126),
.A2(n_49),
.B(n_68),
.C(n_125),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_128),
.B(n_127),
.Y(n_129)
);


endmodule