module fake_jpeg_30066_n_63 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_16),
.A2(n_21),
.B(n_25),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_24),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_28),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_27),
.B(n_30),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_31),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_9),
.B1(n_22),
.B2(n_19),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_26),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_1),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_43),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_13),
.B(n_23),
.Y(n_54)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_34),
.A2(n_8),
.B1(n_17),
.B2(n_15),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_3),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_11),
.C(n_14),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_50),
.C(n_46),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_54),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_42),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_40),
.B1(n_44),
.B2(n_49),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_51),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_60),
.A2(n_58),
.B1(n_55),
.B2(n_50),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_59),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_61),
.Y(n_63)
);


endmodule