module fake_jpeg_14330_n_131 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_131);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_131;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_1),
.B(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_8),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_28),
.B(n_34),
.Y(n_57)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_19),
.B(n_9),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_0),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_13),
.B(n_17),
.C(n_25),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_4),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_38),
.A2(n_18),
.B1(n_27),
.B2(n_16),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_41),
.A2(n_55),
.B1(n_51),
.B2(n_53),
.Y(n_62)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_16),
.B(n_26),
.C(n_17),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_51),
.Y(n_68)
);

AOI32xp33_ASAP7_75t_L g45 ( 
.A1(n_30),
.A2(n_22),
.A3(n_26),
.B1(n_13),
.B2(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_45),
.B(n_49),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_41),
.Y(n_69)
);

OA21x2_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_31),
.B(n_30),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_35),
.B1(n_11),
.B2(n_12),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_24),
.B(n_21),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_21),
.C(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_22),
.B1(n_2),
.B2(n_1),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_55),
.B1(n_31),
.B2(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_30),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_1),
.B1(n_4),
.B2(n_10),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_58),
.B(n_59),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_11),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_60),
.B(n_64),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_12),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_62),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_43),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_52),
.A2(n_44),
.B1(n_48),
.B2(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_67),
.B(n_69),
.Y(n_88)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_74),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_83),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_79),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_65),
.C(n_63),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_54),
.Y(n_83)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_63),
.B1(n_72),
.B2(n_61),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2x1_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_58),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_92),
.B(n_95),
.Y(n_103)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_84),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_97),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_59),
.B1(n_66),
.B2(n_82),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_59),
.B1(n_81),
.B2(n_75),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_59),
.B(n_78),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_86),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_102),
.A2(n_87),
.B(n_99),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_108),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_104),
.A2(n_97),
.B1(n_95),
.B2(n_100),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_94),
.C(n_98),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_115),
.C(n_109),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_92),
.B(n_94),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_87),
.B(n_105),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_109),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_104),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_117),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_118),
.B(n_119),
.Y(n_121)
);

BUFx24_ASAP7_75t_SL g119 ( 
.A(n_113),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_122),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_111),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_96),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_115),
.B1(n_106),
.B2(n_90),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_106),
.C(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_127),
.B(n_121),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_125),
.Y(n_131)
);


endmodule