module fake_netlist_1_12461_n_726 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_726);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_726;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g101 ( .A(n_73), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_77), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_51), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_21), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_89), .Y(n_105) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_25), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_4), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_45), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_47), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_1), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_85), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_39), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_61), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_90), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_33), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_30), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_19), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_84), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_10), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_78), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_34), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_46), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_7), .Y(n_124) );
BUFx10_ASAP7_75t_L g125 ( .A(n_53), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_62), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_8), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_43), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_97), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_23), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_36), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_48), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_86), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_60), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_68), .Y(n_136) );
BUFx2_ASAP7_75t_SL g137 ( .A(n_72), .Y(n_137) );
INVxp67_ASAP7_75t_SL g138 ( .A(n_69), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_76), .Y(n_139) );
INVx2_ASAP7_75t_SL g140 ( .A(n_44), .Y(n_140) );
INVx1_ASAP7_75t_SL g141 ( .A(n_13), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_106), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_106), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_108), .B(n_125), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_124), .Y(n_145) );
OA21x2_ASAP7_75t_L g146 ( .A1(n_101), .A2(n_0), .B(n_1), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_121), .B(n_0), .Y(n_148) );
AND2x2_ASAP7_75t_SL g149 ( .A(n_102), .B(n_18), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_125), .B(n_2), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_124), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_121), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_125), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_107), .B(n_2), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_106), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_140), .B(n_3), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_106), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_109), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_140), .Y(n_159) );
INVxp67_ASAP7_75t_L g160 ( .A(n_120), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_112), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_153), .B(n_105), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_153), .B(n_111), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_161), .Y(n_164) );
BUFx3_ASAP7_75t_L g165 ( .A(n_156), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_161), .Y(n_166) );
INVxp67_ASAP7_75t_SL g167 ( .A(n_147), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_144), .B(n_110), .Y(n_168) );
OA22x2_ASAP7_75t_L g169 ( .A1(n_148), .A2(n_128), .B1(n_110), .B2(n_141), .Y(n_169) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_149), .B(n_113), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_148), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_148), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_148), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_161), .Y(n_174) );
INVx2_ASAP7_75t_SL g175 ( .A(n_153), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_149), .A2(n_131), .B1(n_117), .B2(n_116), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
OR2x6_ASAP7_75t_L g179 ( .A(n_150), .B(n_137), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_147), .Y(n_180) );
INVxp67_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_153), .B(n_111), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_144), .B(n_116), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_143), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_161), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_147), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_150), .Y(n_189) );
NAND3xp33_ASAP7_75t_L g190 ( .A(n_146), .B(n_139), .C(n_127), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_184), .B(n_153), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_163), .B(n_160), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_176), .B(n_149), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_179), .B(n_150), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_172), .A2(n_156), .B(n_149), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_168), .B(n_160), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g197 ( .A1(n_170), .A2(n_156), .B1(n_154), .B2(n_131), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_184), .B(n_158), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_176), .B(n_156), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_182), .B(n_158), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_176), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_167), .B(n_156), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_176), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_170), .A2(n_154), .B1(n_146), .B2(n_156), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_168), .B(n_147), .Y(n_205) );
AND2x4_ASAP7_75t_L g206 ( .A(n_179), .B(n_154), .Y(n_206) );
O2A1O1Ixp5_ASAP7_75t_L g207 ( .A1(n_178), .A2(n_159), .B(n_152), .C(n_138), .Y(n_207) );
INVx5_ASAP7_75t_L g208 ( .A(n_178), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_170), .A2(n_117), .B1(n_159), .B2(n_152), .Y(n_209) );
BUFx2_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
NAND3xp33_ASAP7_75t_L g211 ( .A(n_181), .B(n_146), .C(n_159), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_178), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_178), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_180), .Y(n_214) );
INVx2_ASAP7_75t_SL g215 ( .A(n_179), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_162), .B(n_159), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_171), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_175), .B(n_152), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_175), .B(n_118), .Y(n_219) );
OR2x2_ASAP7_75t_L g220 ( .A(n_179), .B(n_151), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_172), .B(n_151), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_171), .B(n_161), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_173), .B(n_133), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_177), .A2(n_146), .B1(n_132), .B2(n_118), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_179), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_169), .Y(n_226) );
AOI22xp33_ASAP7_75t_L g227 ( .A1(n_173), .A2(n_146), .B1(n_161), .B2(n_145), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_171), .B(n_130), .Y(n_228) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_177), .A2(n_146), .B1(n_132), .B2(n_130), .Y(n_229) );
AO21x1_ASAP7_75t_L g230 ( .A1(n_195), .A2(n_142), .B(n_145), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_197), .A2(n_209), .B1(n_194), .B2(n_193), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_196), .B(n_165), .Y(n_232) );
OAI21x1_ASAP7_75t_L g233 ( .A1(n_227), .A2(n_190), .B(n_169), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_198), .B(n_165), .Y(n_234) );
OAI22x1_ASAP7_75t_L g235 ( .A1(n_224), .A2(n_190), .B1(n_169), .B2(n_145), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_206), .B(n_171), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_206), .B(n_180), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_199), .A2(n_188), .B(n_185), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_205), .B(n_185), .Y(n_239) );
INVx3_ASAP7_75t_L g240 ( .A(n_212), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_215), .B(n_188), .Y(n_241) );
OAI22xp5_ASAP7_75t_L g242 ( .A1(n_194), .A2(n_136), .B1(n_161), .B2(n_115), .Y(n_242) );
INVx5_ASAP7_75t_L g243 ( .A(n_194), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_199), .A2(n_187), .B(n_164), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_192), .B(n_161), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_225), .B(n_103), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_217), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_193), .A2(n_123), .B1(n_114), .B2(n_119), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_226), .A2(n_135), .B(n_122), .C(n_126), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_220), .Y(n_250) );
INVxp67_ASAP7_75t_SL g251 ( .A(n_212), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_201), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_201), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_214), .Y(n_254) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_229), .A2(n_129), .B1(n_134), .B2(n_104), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_192), .B(n_3), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_203), .Y(n_257) );
INVx2_ASAP7_75t_SL g258 ( .A(n_208), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_208), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_204), .B(n_4), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_191), .B(n_5), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_213), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_243), .B(n_208), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_244), .A2(n_222), .B(n_202), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_231), .A2(n_210), .B1(n_200), .B2(n_223), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_250), .B(n_223), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_233), .A2(n_211), .B(n_207), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_230), .A2(n_227), .B(n_204), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_254), .Y(n_269) );
BUFx4f_ASAP7_75t_SL g270 ( .A(n_259), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_254), .Y(n_271) );
AO21x2_ASAP7_75t_L g272 ( .A1(n_230), .A2(n_216), .B(n_222), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_218), .B(n_228), .Y(n_273) );
CKINVDCx11_ASAP7_75t_R g274 ( .A(n_259), .Y(n_274) );
BUFx6f_ASAP7_75t_L g275 ( .A(n_258), .Y(n_275) );
AOI21x1_ASAP7_75t_L g276 ( .A1(n_235), .A2(n_164), .B(n_166), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_262), .Y(n_277) );
NOR4xp25_ASAP7_75t_L g278 ( .A(n_255), .B(n_216), .C(n_221), .D(n_200), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_234), .A2(n_219), .B1(n_221), .B2(n_208), .Y(n_279) );
A2O1A1Ixp33_ASAP7_75t_L g280 ( .A1(n_260), .A2(n_142), .B(n_187), .C(n_174), .Y(n_280) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_233), .A2(n_166), .B(n_174), .Y(n_281) );
O2A1O1Ixp5_ASAP7_75t_L g282 ( .A1(n_256), .A2(n_155), .B(n_142), .C(n_186), .Y(n_282) );
AO32x2_ASAP7_75t_L g283 ( .A1(n_242), .A2(n_143), .A3(n_157), .B1(n_142), .B2(n_155), .Y(n_283) );
CKINVDCx5p33_ASAP7_75t_R g284 ( .A(n_243), .Y(n_284) );
O2A1O1Ixp5_ASAP7_75t_SL g285 ( .A1(n_245), .A2(n_155), .B(n_157), .C(n_143), .Y(n_285) );
INVx1_ASAP7_75t_SL g286 ( .A(n_243), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_269), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_273), .A2(n_261), .B(n_247), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g289 ( .A1(n_265), .A2(n_249), .B(n_260), .C(n_241), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_266), .B(n_232), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_276), .A2(n_248), .B(n_239), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_271), .Y(n_293) );
CKINVDCx11_ASAP7_75t_R g294 ( .A(n_274), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_267), .A2(n_247), .B(n_253), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g296 ( .A(n_274), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_264), .A2(n_235), .B(n_253), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_285), .A2(n_240), .B(n_257), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_281), .A2(n_240), .B(n_257), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_278), .B(n_237), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_270), .B(n_243), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_281), .A2(n_240), .B(n_262), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_280), .A2(n_252), .B(n_236), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_270), .Y(n_305) );
BUFx8_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_284), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_272), .Y(n_308) );
OAI33xp33_ASAP7_75t_L g309 ( .A1(n_301), .A2(n_279), .A3(n_284), .B1(n_7), .B2(n_8), .B3(n_9), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_294), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_299), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_299), .B(n_268), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_287), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_306), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_290), .B(n_286), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_306), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_289), .A2(n_243), .B1(n_272), .B2(n_263), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_295), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_293), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_295), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_295), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_291), .B(n_246), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_295), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_308), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_300), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_290), .B(n_268), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_306), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_308), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_290), .B(n_275), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_303), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_305), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_303), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_304), .B(n_275), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_304), .B(n_275), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_305), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_296), .Y(n_336) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_300), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_307), .B(n_280), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_324), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_312), .B(n_304), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_312), .B(n_281), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_326), .B(n_297), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_313), .B(n_296), .Y(n_343) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_315), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_318), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
BUFx3_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
OR2x6_ASAP7_75t_L g350 ( .A(n_327), .B(n_288), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_326), .B(n_292), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_311), .B(n_292), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_333), .B(n_298), .Y(n_353) );
INVx2_ASAP7_75t_SL g354 ( .A(n_327), .Y(n_354) );
INVx4_ASAP7_75t_L g355 ( .A(n_314), .Y(n_355) );
AND2x2_ASAP7_75t_SL g356 ( .A(n_314), .B(n_302), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_337), .Y(n_357) );
NOR2x1_ASAP7_75t_SL g358 ( .A(n_327), .B(n_275), .Y(n_358) );
INVx4_ASAP7_75t_L g359 ( .A(n_314), .Y(n_359) );
OR2x2_ASAP7_75t_L g360 ( .A(n_324), .B(n_292), .Y(n_360) );
BUFx3_ASAP7_75t_L g361 ( .A(n_316), .Y(n_361) );
NAND2x1_ASAP7_75t_L g362 ( .A(n_330), .B(n_258), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_328), .B(n_311), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_320), .Y(n_364) );
NAND2x1_ASAP7_75t_L g365 ( .A(n_330), .B(n_143), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_313), .B(n_5), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_316), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_321), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_319), .B(n_283), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_323), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_323), .Y(n_374) );
AND2x4_ASAP7_75t_L g375 ( .A(n_333), .B(n_334), .Y(n_375) );
INVxp67_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_322), .B(n_338), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_334), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_329), .B(n_283), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_332), .B(n_298), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_325), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_332), .B(n_6), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_329), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_317), .B(n_6), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_317), .B(n_283), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_325), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_331), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_335), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_337), .B(n_283), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_356), .A2(n_309), .B1(n_310), .B2(n_337), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_378), .B(n_337), .Y(n_391) );
AND2x4_ASAP7_75t_SL g392 ( .A(n_355), .B(n_337), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_339), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_377), .B(n_9), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_339), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_375), .B(n_143), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_367), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_367), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_378), .B(n_143), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_363), .B(n_10), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_371), .B(n_11), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_345), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_375), .B(n_143), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_375), .B(n_157), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_375), .B(n_157), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_373), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_340), .B(n_157), .Y(n_407) );
AND2x4_ASAP7_75t_L g408 ( .A(n_353), .B(n_157), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_340), .B(n_157), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_345), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g411 ( .A1(n_356), .A2(n_310), .B1(n_251), .B2(n_155), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_351), .B(n_157), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_355), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_344), .B(n_11), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_346), .B(n_12), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_383), .B(n_388), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_374), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_363), .B(n_12), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_374), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_353), .B(n_155), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_351), .B(n_13), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_347), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_347), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_348), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_342), .B(n_14), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_342), .B(n_14), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_352), .B(n_15), .Y(n_429) );
OR2x2_ASAP7_75t_L g430 ( .A(n_348), .B(n_15), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_365), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_352), .B(n_16), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_348), .B(n_16), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_364), .B(n_17), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_364), .Y(n_435) );
INVx4_ASAP7_75t_L g436 ( .A(n_355), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_364), .B(n_17), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_366), .B(n_20), .Y(n_438) );
AND2x4_ASAP7_75t_L g439 ( .A(n_353), .B(n_22), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_347), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_366), .B(n_24), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_366), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_361), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_370), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_370), .B(n_26), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_370), .B(n_27), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_381), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_361), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_365), .Y(n_449) );
HB1xp67_ASAP7_75t_SL g450 ( .A(n_361), .Y(n_450) );
INVx5_ASAP7_75t_L g451 ( .A(n_355), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_381), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_360), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_360), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_341), .B(n_28), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_353), .B(n_29), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_341), .B(n_31), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_382), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_372), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_387), .B(n_32), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_385), .B(n_35), .Y(n_461) );
OR2x6_ASAP7_75t_L g462 ( .A(n_359), .B(n_282), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_381), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_382), .B(n_37), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_451), .B(n_359), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_393), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_444), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_395), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_423), .B(n_372), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_395), .Y(n_470) );
NOR2xp67_ASAP7_75t_L g471 ( .A(n_451), .B(n_359), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_423), .B(n_376), .Y(n_472) );
AND3x1_ASAP7_75t_L g473 ( .A(n_450), .B(n_354), .C(n_343), .Y(n_473) );
INVxp33_ASAP7_75t_L g474 ( .A(n_413), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_418), .B(n_403), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_414), .B(n_369), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_397), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_459), .B(n_354), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_397), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_403), .B(n_369), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_398), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_429), .B(n_384), .Y(n_482) );
NAND2xp33_ASAP7_75t_SL g483 ( .A(n_436), .B(n_359), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_429), .B(n_384), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_398), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_407), .B(n_385), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_459), .B(n_369), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_407), .B(n_389), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_453), .B(n_349), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_409), .B(n_389), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_432), .B(n_379), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_404), .B(n_379), .Y(n_493) );
NOR2xp67_ASAP7_75t_R g494 ( .A(n_451), .B(n_349), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_444), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_402), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_404), .B(n_349), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_413), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_412), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_405), .B(n_356), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_405), .B(n_350), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_443), .B(n_350), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_448), .B(n_350), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_432), .B(n_350), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_406), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_453), .B(n_386), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_409), .B(n_350), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_391), .B(n_380), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_406), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_402), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_417), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_412), .B(n_358), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_410), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_427), .B(n_428), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_410), .Y(n_515) );
NAND2x1_ASAP7_75t_L g516 ( .A(n_436), .B(n_357), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_417), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_427), .B(n_358), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_454), .B(n_386), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_419), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_451), .B(n_380), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_419), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_421), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_421), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_428), .B(n_368), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_426), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_416), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_426), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_435), .Y(n_529) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_416), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_458), .B(n_386), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_442), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_391), .B(n_454), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_424), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_400), .B(n_380), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_400), .B(n_380), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_442), .B(n_362), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_433), .B(n_357), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_430), .B(n_362), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_424), .B(n_357), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_430), .B(n_357), .Y(n_541) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_431), .Y(n_542) );
INVxp67_ASAP7_75t_L g543 ( .A(n_396), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_425), .B(n_440), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_437), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_437), .B(n_38), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_425), .B(n_40), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_433), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_440), .B(n_41), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_447), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_408), .B(n_42), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_533), .B(n_434), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_499), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_483), .B(n_390), .C(n_394), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_472), .B(n_415), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_533), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_475), .B(n_508), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_476), .B(n_401), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_528), .B(n_422), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_528), .B(n_422), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_466), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_499), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_508), .B(n_396), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_468), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_470), .Y(n_565) );
O2A1O1Ixp33_ASAP7_75t_L g566 ( .A1(n_525), .A2(n_411), .B(n_420), .C(n_460), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_527), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_477), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_535), .B(n_536), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_465), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_514), .B(n_434), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_469), .B(n_463), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_483), .Y(n_573) );
OR2x2_ASAP7_75t_L g574 ( .A(n_478), .B(n_463), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_479), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_504), .A2(n_461), .B1(n_422), .B2(n_439), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_545), .B(n_399), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_481), .Y(n_578) );
INVxp33_ASAP7_75t_L g579 ( .A(n_494), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_492), .B(n_399), .Y(n_580) );
NAND2x1p5_ASAP7_75t_L g581 ( .A(n_471), .B(n_451), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_486), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_487), .B(n_396), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_487), .B(n_408), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_530), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_489), .B(n_408), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_505), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_465), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_531), .B(n_447), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_509), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_511), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_489), .B(n_439), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_498), .B(n_452), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_491), .B(n_452), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_526), .B(n_461), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_517), .Y(n_596) );
AND2x4_ASAP7_75t_L g597 ( .A(n_465), .B(n_392), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_491), .B(n_439), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_530), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_520), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_522), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_488), .B(n_457), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_523), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_506), .B(n_457), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_519), .B(n_455), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_524), .Y(n_606) );
NOR2x1_ASAP7_75t_L g607 ( .A(n_485), .B(n_431), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_529), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_501), .B(n_456), .Y(n_609) );
OR2x2_ASAP7_75t_L g610 ( .A(n_493), .B(n_455), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_532), .B(n_431), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_544), .B(n_449), .Y(n_612) );
INVxp67_ASAP7_75t_L g613 ( .A(n_473), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_490), .Y(n_614) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_474), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_544), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_485), .B(n_449), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_476), .Y(n_618) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_474), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_507), .B(n_456), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_467), .B(n_449), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_467), .B(n_456), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_500), .A2(n_462), .B1(n_464), .B2(n_441), .Y(n_623) );
OAI221xp5_ASAP7_75t_SL g624 ( .A1(n_543), .A2(n_464), .B1(n_462), .B2(n_446), .C(n_445), .Y(n_624) );
OAI221xp5_ASAP7_75t_SL g625 ( .A1(n_613), .A2(n_482), .B1(n_484), .B2(n_543), .C(n_502), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_608), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_615), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g628 ( .A(n_569), .B(n_518), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_561), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_556), .B(n_548), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_567), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g632 ( .A(n_618), .B(n_485), .Y(n_632) );
INVxp67_ASAP7_75t_L g633 ( .A(n_619), .Y(n_633) );
OAI211xp5_ASAP7_75t_SL g634 ( .A1(n_566), .A2(n_542), .B(n_539), .C(n_538), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_562), .A2(n_503), .B1(n_542), .B2(n_540), .C(n_480), .Y(n_635) );
INVx1_ASAP7_75t_SL g636 ( .A(n_597), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
INVxp67_ASAP7_75t_SL g638 ( .A(n_581), .Y(n_638) );
OAI21xp33_ASAP7_75t_SL g639 ( .A1(n_579), .A2(n_512), .B(n_497), .Y(n_639) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_554), .A2(n_555), .B(n_573), .C(n_624), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g641 ( .A1(n_554), .A2(n_516), .B1(n_537), .B2(n_546), .C(n_541), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_559), .A2(n_521), .B1(n_551), .B2(n_540), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_597), .B(n_551), .Y(n_643) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_611), .B(n_495), .C(n_550), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_607), .B(n_521), .Y(n_645) );
AOI32xp33_ASAP7_75t_L g646 ( .A1(n_570), .A2(n_521), .A3(n_392), .B1(n_438), .B2(n_441), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_564), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_565), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_553), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_568), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_575), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g652 ( .A1(n_571), .A2(n_495), .A3(n_438), .B1(n_445), .B2(n_534), .C1(n_515), .C2(n_513), .Y(n_652) );
OR2x2_ASAP7_75t_L g653 ( .A(n_594), .B(n_550), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_559), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_578), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_576), .A2(n_462), .B1(n_549), .B2(n_534), .Y(n_656) );
AND2x4_ASAP7_75t_L g657 ( .A(n_588), .B(n_510), .Y(n_657) );
INVxp67_ASAP7_75t_L g658 ( .A(n_560), .Y(n_658) );
OAI21xp33_ASAP7_75t_L g659 ( .A1(n_612), .A2(n_496), .B(n_515), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_582), .Y(n_660) );
AOI21xp33_ASAP7_75t_SL g661 ( .A1(n_581), .A2(n_446), .B(n_547), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_587), .Y(n_662) );
AOI221x1_ASAP7_75t_SL g663 ( .A1(n_614), .A2(n_513), .B1(n_510), .B2(n_496), .C(n_549), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_574), .Y(n_664) );
NOR3xp33_ASAP7_75t_L g665 ( .A(n_560), .B(n_462), .C(n_50), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_557), .B(n_49), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_590), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_592), .A2(n_186), .B1(n_183), .B2(n_55), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g669 ( .A1(n_639), .A2(n_623), .B1(n_612), .B2(n_583), .C(n_584), .Y(n_669) );
AOI211xp5_ASAP7_75t_L g670 ( .A1(n_640), .A2(n_617), .B(n_595), .C(n_611), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_663), .A2(n_563), .B(n_586), .C(n_610), .Y(n_671) );
NOR3xp33_ASAP7_75t_L g672 ( .A(n_634), .B(n_621), .C(n_591), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_626), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_654), .B(n_552), .Y(n_674) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_637), .A2(n_616), .A3(n_598), .B1(n_580), .B2(n_595), .C1(n_620), .C2(n_609), .Y(n_675) );
AND2x2_ASAP7_75t_L g676 ( .A(n_636), .B(n_572), .Y(n_676) );
OAI21xp5_ASAP7_75t_SL g677 ( .A1(n_665), .A2(n_622), .B(n_602), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g678 ( .A1(n_625), .A2(n_603), .B1(n_600), .B2(n_606), .C(n_601), .Y(n_678) );
OAI21xp33_ASAP7_75t_SL g679 ( .A1(n_638), .A2(n_621), .B(n_605), .Y(n_679) );
AOI322xp5_ASAP7_75t_L g680 ( .A1(n_627), .A2(n_596), .A3(n_577), .B1(n_585), .B2(n_599), .C1(n_589), .C2(n_622), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_629), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_643), .A2(n_604), .B1(n_589), .B2(n_593), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_658), .B(n_52), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g684 ( .A1(n_641), .A2(n_186), .B(n_183), .C(n_57), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_633), .B(n_54), .Y(n_685) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_666), .A2(n_56), .B(n_58), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g687 ( .A1(n_632), .A2(n_59), .B(n_63), .C(n_64), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_645), .B(n_186), .Y(n_688) );
NOR2xp67_ASAP7_75t_L g689 ( .A(n_645), .B(n_65), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_635), .A2(n_186), .B1(n_183), .B2(n_70), .C(n_71), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_647), .A2(n_66), .B(n_67), .C(n_75), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_659), .A2(n_183), .B1(n_81), .B2(n_82), .C(n_83), .Y(n_692) );
NAND4xp25_ASAP7_75t_SL g693 ( .A(n_646), .B(n_80), .C(n_87), .D(n_88), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g694 ( .A1(n_642), .A2(n_91), .B1(n_92), .B2(n_93), .C(n_94), .Y(n_694) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_644), .B(n_95), .Y(n_695) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_649), .Y(n_696) );
NAND4xp25_ASAP7_75t_L g697 ( .A(n_656), .B(n_96), .C(n_98), .D(n_99), .Y(n_697) );
OAI21x1_ASAP7_75t_SL g698 ( .A1(n_628), .A2(n_100), .B(n_664), .Y(n_698) );
NAND3xp33_ASAP7_75t_L g699 ( .A(n_652), .B(n_667), .C(n_660), .Y(n_699) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_661), .A2(n_653), .B1(n_657), .B2(n_630), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g701 ( .A1(n_657), .A2(n_668), .B1(n_648), .B2(n_650), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_651), .A2(n_655), .B(n_662), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_631), .A2(n_640), .B1(n_625), .B2(n_663), .C(n_634), .Y(n_703) );
AOI211x1_ASAP7_75t_L g704 ( .A1(n_700), .A2(n_699), .B(n_669), .C(n_702), .Y(n_704) );
NAND4xp25_ASAP7_75t_L g705 ( .A(n_703), .B(n_684), .C(n_697), .D(n_670), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_672), .B(n_678), .Y(n_706) );
XOR2xp5_ASAP7_75t_L g707 ( .A(n_696), .B(n_693), .Y(n_707) );
NAND3x1_ASAP7_75t_L g708 ( .A(n_695), .B(n_698), .C(n_690), .Y(n_708) );
OAI211xp5_ASAP7_75t_SL g709 ( .A1(n_679), .A2(n_680), .B(n_675), .C(n_677), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g710 ( .A(n_687), .B(n_694), .C(n_685), .Y(n_710) );
NOR3xp33_ASAP7_75t_L g711 ( .A(n_705), .B(n_691), .C(n_701), .Y(n_711) );
NOR2x1_ASAP7_75t_L g712 ( .A(n_707), .B(n_689), .Y(n_712) );
NOR3x1_ASAP7_75t_L g713 ( .A(n_706), .B(n_682), .C(n_683), .Y(n_713) );
NOR3xp33_ASAP7_75t_L g714 ( .A(n_709), .B(n_692), .C(n_688), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_712), .B(n_676), .Y(n_715) );
XOR2x2_ASAP7_75t_L g716 ( .A(n_711), .B(n_704), .Y(n_716) );
AND3x4_ASAP7_75t_L g717 ( .A(n_714), .B(n_710), .C(n_708), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_715), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_717), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_719), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_720), .A2(n_716), .B(n_713), .Y(n_722) );
NOR2xp67_ASAP7_75t_L g723 ( .A(n_722), .B(n_721), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_723), .A2(n_671), .B(n_682), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_724), .A2(n_681), .B(n_673), .Y(n_725) );
AOI21xp33_ASAP7_75t_SL g726 ( .A1(n_725), .A2(n_674), .B(n_686), .Y(n_726) );
endmodule