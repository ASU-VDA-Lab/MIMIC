module real_jpeg_10067_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_334, n_335, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_334;
input n_335;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_1),
.A2(n_24),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_36),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_1),
.A2(n_36),
.B1(n_61),
.B2(n_62),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_1),
.A2(n_36),
.B1(n_44),
.B2(n_47),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_2),
.A2(n_24),
.B1(n_33),
.B2(n_55),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_2),
.A2(n_55),
.B1(n_61),
.B2(n_62),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_2),
.A2(n_44),
.B1(n_47),
.B2(n_55),
.Y(n_219)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_4),
.A2(n_61),
.B1(n_62),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_4),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_4),
.A2(n_44),
.B1(n_47),
.B2(n_115),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_115),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_4),
.A2(n_24),
.B1(n_33),
.B2(n_115),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g112 ( 
.A(n_5),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_10),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_44),
.B1(n_47),
.B2(n_110),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_110),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_10),
.A2(n_24),
.B1(n_33),
.B2(n_110),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_11),
.A2(n_44),
.B1(n_47),
.B2(n_49),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_11),
.A2(n_49),
.B1(n_61),
.B2(n_62),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_11),
.A2(n_24),
.B1(n_33),
.B2(n_49),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_13),
.A2(n_44),
.B1(n_47),
.B2(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_13),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_13),
.A2(n_61),
.B1(n_62),
.B2(n_122),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_122),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_13),
.A2(n_24),
.B1(n_33),
.B2(n_122),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_24),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_14),
.A2(n_34),
.B1(n_61),
.B2(n_62),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_14),
.A2(n_34),
.B1(n_44),
.B2(n_47),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_15),
.A2(n_47),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_15),
.B(n_47),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_15),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_15),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_15),
.B(n_92),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_15),
.A2(n_26),
.B(n_30),
.Y(n_206)
);

OAI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_15),
.A2(n_24),
.B1(n_33),
.B2(n_131),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_98),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_96),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_83),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_19),
.B(n_83),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_70),
.C(n_74),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_20),
.A2(n_21),
.B1(n_70),
.B2(n_319),
.Y(n_325)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_37),
.B1(n_38),
.B2(n_69),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_23),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_23),
.A2(n_28),
.B1(n_226),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_23),
.A2(n_28),
.B1(n_235),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_23),
.A2(n_254),
.B(n_279),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_23),
.A2(n_91),
.B(n_300),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_24),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_24),
.A2(n_25),
.B(n_131),
.C(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_28),
.A2(n_32),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_28),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g51 ( 
.A1(n_30),
.A2(n_41),
.B(n_42),
.C(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_42),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g160 ( 
.A(n_30),
.B(n_131),
.CON(n_160),
.SN(n_160)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_56),
.B1(n_67),
.B2(n_68),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_50),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_40),
.A2(n_77),
.B(n_222),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_48),
.Y(n_40)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_41),
.A2(n_48),
.B(n_51),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_41),
.A2(n_51),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_41),
.A2(n_51),
.B1(n_79),
.B2(n_305),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_42),
.B(n_47),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_44),
.A2(n_52),
.B1(n_160),
.B2(n_166),
.Y(n_165)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_47),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_58),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_48),
.A2(n_51),
.B(n_81),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_50),
.A2(n_82),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_51),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_67),
.C(n_69),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_56),
.A2(n_68),
.B1(n_75),
.B2(n_76),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_60),
.B(n_65),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_57),
.A2(n_60),
.B1(n_119),
.B2(n_121),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_57),
.A2(n_60),
.B1(n_121),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_57),
.A2(n_60),
.B1(n_148),
.B2(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_57),
.A2(n_158),
.B(n_194),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_57),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_57),
.A2(n_60),
.B1(n_241),
.B2(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_57),
.A2(n_260),
.B(n_289),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_58),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_58),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_60),
.B(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_60),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_60),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_60),
.A2(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_61),
.B(n_112),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_61),
.B(n_64),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_61),
.B(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_123)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_66),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_66),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_70),
.C(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_70),
.A2(n_319),
.B1(n_320),
.B2(n_321),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_70),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_72),
.B(n_92),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_73),
.A2(n_92),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_74),
.B(n_325),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_80),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_77),
.A2(n_82),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_77),
.A2(n_82),
.B1(n_180),
.B2(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_82),
.B(n_131),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_84),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_92),
.B(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI321xp33_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_316),
.A3(n_326),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_268),
.A3(n_292),
.B1(n_309),
.B2(n_315),
.C(n_335),
.Y(n_99)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_228),
.C(n_264),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_199),
.B(n_227),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_103),
.A2(n_173),
.B(n_198),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_153),
.B(n_172),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_142),
.B(n_152),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_128),
.B(n_141),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_116),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_107),
.B(n_116),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_108),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_109),
.A2(n_133),
.B1(n_134),
.B2(n_135),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_111),
.B(n_170),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_114),
.A2(n_134),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_123),
.B2(n_127),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_117),
.B(n_127),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_120),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_123),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_136),
.B(n_140),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_132),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_131),
.B(n_135),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_168),
.B(n_169),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_134),
.A2(n_135),
.B1(n_184),
.B2(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_134),
.A2(n_169),
.B(n_209),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_134),
.A2(n_135),
.B(n_168),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_135),
.A2(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_143),
.B(n_144),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_154),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_147),
.CI(n_149),
.CON(n_145),
.SN(n_145)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_150),
.B(n_185),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_164),
.B2(n_171),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_157),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_163),
.C(n_171),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_161),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_167),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_175),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_190),
.B2(n_191),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_193),
.C(n_196),
.Y(n_200)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_181),
.B1(n_182),
.B2(n_189),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_178),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_186),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_186),
.B(n_187),
.C(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_193),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_194),
.B(n_242),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_200),
.B(n_201),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_213),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_203),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_203),
.B(n_212),
.C(n_213),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_207),
.B2(n_208),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_208),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_223),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_221),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_216),
.B(n_220),
.C(n_223),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_243),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_218),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_247),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_229),
.B(n_247),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.C(n_245),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_233),
.C(n_237),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_236),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_238),
.A2(n_239),
.B1(n_245),
.B2(n_246),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_244),
.Y(n_250)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_247)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_257),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_249),
.B(n_257),
.C(n_261),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_252),
.C(n_256),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_259),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_265),
.B(n_266),
.Y(n_312)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_269),
.A2(n_310),
.B(n_314),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_270),
.B(n_271),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_291),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_284),
.B2(n_285),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_285),
.C(n_291),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_275),
.B(n_277),
.C(n_283),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_281),
.B2(n_283),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_280),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_281),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_282),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_290),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_287),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_286),
.A2(n_299),
.B(n_302),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_288),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_288),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_293),
.B(n_294),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_294),
.Y(n_327)
);

FAx1_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.CI(n_308),
.CON(n_294),
.SN(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_301),
.B2(n_302),
.Y(n_295)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_306),
.B(n_307),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_306),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_307),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_307),
.A2(n_318),
.B1(n_322),
.B2(n_330),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_324),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_324),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_322),
.C(n_323),
.Y(n_317)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_329),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);


endmodule