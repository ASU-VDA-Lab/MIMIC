module fake_netlist_1_10987_n_35 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_35);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_35;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
HB1xp67_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_3), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_9), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_13), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_15), .B(n_0), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_17), .A2(n_14), .B1(n_16), .B2(n_13), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_17), .A2(n_13), .B1(n_1), .B2(n_2), .Y(n_22) );
CKINVDCx8_ASAP7_75t_R g23 ( .A(n_21), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVx3_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_23), .B(n_20), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_25), .B(n_18), .Y(n_27) );
OAI21xp33_ASAP7_75t_SL g28 ( .A1(n_25), .A2(n_19), .B(n_1), .Y(n_28) );
XNOR2xp5_ASAP7_75t_L g29 ( .A(n_27), .B(n_26), .Y(n_29) );
NAND4xp75_ASAP7_75t_L g30 ( .A(n_28), .B(n_0), .C(n_2), .D(n_3), .Y(n_30) );
NAND2xp33_ASAP7_75t_L g31 ( .A(n_27), .B(n_13), .Y(n_31) );
NAND4xp25_ASAP7_75t_SL g32 ( .A(n_30), .B(n_7), .C(n_10), .D(n_31), .Y(n_32) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_29), .Y(n_33) );
HB1xp67_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
XNOR2xp5_ASAP7_75t_L g35 ( .A(n_34), .B(n_32), .Y(n_35) );
endmodule