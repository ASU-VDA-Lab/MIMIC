module real_jpeg_12221_n_16 (n_5, n_4, n_8, n_0, n_12, n_409, n_408, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_409;
input n_408;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_2),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_43),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_3),
.B(n_48),
.Y(n_154)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_3),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_3),
.B(n_33),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_3),
.B(n_28),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_3),
.B(n_135),
.Y(n_340)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_5),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_5),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_5),
.B(n_33),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_5),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_5),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_6),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_6),
.B(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_6),
.B(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_6),
.B(n_135),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_6),
.B(n_178),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_7),
.B(n_43),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_7),
.B(n_48),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_7),
.B(n_31),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_7),
.B(n_33),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_7),
.B(n_28),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_7),
.B(n_61),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_7),
.B(n_135),
.Y(n_262)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_7),
.Y(n_300)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_10),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_10),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_10),
.B(n_28),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_61),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_10),
.B(n_135),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_11),
.B(n_43),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_11),
.B(n_48),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_11),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_11),
.B(n_33),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_11),
.B(n_28),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_11),
.B(n_61),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_11),
.B(n_135),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_12),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_13),
.B(n_28),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_13),
.B(n_48),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_13),
.B(n_31),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_13),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_13),
.B(n_61),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_13),
.B(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_13),
.B(n_178),
.Y(n_208)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_14),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_14),
.B(n_48),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_14),
.B(n_31),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_14),
.B(n_33),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_14),
.B(n_61),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_14),
.B(n_178),
.Y(n_389)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_392),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_376),
.B(n_391),
.Y(n_17)
);

OAI321xp33_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_327),
.A3(n_351),
.B1(n_374),
.B2(n_375),
.C(n_408),
.Y(n_18)
);

AOI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_249),
.A3(n_285),
.B1(n_321),
.B2(n_326),
.C(n_409),
.Y(n_19)
);

NOR3xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_182),
.C(n_244),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_143),
.B(n_181),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_108),
.B(n_142),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_76),
.B(n_107),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_51),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_25),
.B(n_51),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_35),
.C(n_45),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_26),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_53)
);

CKINVDCx5p33_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_26),
.B(n_104),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_30),
.CI(n_32),
.CON(n_26),
.SN(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_29),
.B(n_167),
.Y(n_310)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_35),
.A2(n_36),
.B1(n_45),
.B2(n_105),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_41),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_37),
.B(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_38),
.B(n_92),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_40),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_42),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_42),
.B(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_44),
.B(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_44),
.B(n_177),
.Y(n_264)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_50),
.Y(n_67)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_49),
.A2(n_50),
.B1(n_123),
.B2(n_124),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_49),
.A2(n_50),
.B1(n_171),
.B2(n_174),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_50),
.B(n_124),
.C(n_241),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_50),
.B(n_174),
.C(n_271),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_66),
.B2(n_75),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_65),
.C(n_75),
.Y(n_109)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_58),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_59),
.C(n_64),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_61),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g66 ( 
.A(n_67),
.B(n_68),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_67),
.B(n_69),
.C(n_70),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_71),
.A2(n_72),
.B1(n_282),
.B2(n_283),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_71),
.A2(n_72),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_71),
.A2(n_72),
.B1(n_118),
.B2(n_119),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_71),
.B(n_299),
.C(n_301),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_71),
.B(n_119),
.C(n_195),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_72),
.B(n_73),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_72),
.B(n_280),
.C(n_282),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_73),
.A2(n_74),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_73),
.B(n_208),
.C(n_211),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_101),
.B(n_106),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_89),
.B(n_100),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_84),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_87),
.C(n_88),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_95),
.B(n_99),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_92),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_93),
.B(n_172),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_93),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_98),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_102),
.B(n_103),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_109),
.B(n_110),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_127),
.B2(n_128),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_111),
.B(n_129),
.C(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_121),
.C(n_122),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_114),
.B(n_116),
.C(n_119),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_118),
.A2(n_119),
.B1(n_173),
.B2(n_175),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_119),
.B(n_173),
.C(n_225),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_125),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_140),
.B2(n_141),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_139),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_136),
.C(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_133),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g138 ( 
.A(n_134),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_135),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_144),
.B(n_145),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_161),
.B2(n_180),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_160),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_148),
.B(n_160),
.C(n_180),
.Y(n_245)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_150),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_156),
.B2(n_157),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_158),
.C(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g407 ( 
.A(n_152),
.Y(n_407)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_154),
.CI(n_155),
.CON(n_152),
.SN(n_152)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_153),
.B(n_154),
.C(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_161),
.Y(n_180)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_161),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.CI(n_169),
.CON(n_161),
.SN(n_161)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_163),
.C(n_169),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_166),
.B(n_168),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_166),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_165),
.B(n_200),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_167),
.B(n_361),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_168),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_173),
.B1(n_174),
.B2(n_175),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_172),
.B(n_177),
.Y(n_338)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_174),
.C(n_176),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_173),
.A2(n_175),
.B1(n_191),
.B2(n_193),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_173),
.B(n_191),
.C(n_270),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_177),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_177),
.B(n_200),
.Y(n_363)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_183),
.A2(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_217),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_184),
.B(n_217),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_205),
.C(n_216),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_204),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_196),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_187),
.B(n_196),
.C(n_204),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_194),
.B2(n_195),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_191),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_190),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_191),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_192),
.C(n_195),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_191),
.A2(n_193),
.B1(n_236),
.B2(n_237),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_193),
.B(n_236),
.C(n_306),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_194),
.A2(n_195),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_205),
.A2(n_206),
.B1(n_216),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_213),
.C(n_215),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_210),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g214 ( 
.A(n_213),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_216),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_243),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_230),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_230),
.C(n_243),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_227),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_228),
.C(n_229),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_225),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_225),
.A2(n_226),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_232),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_231),
.B(n_233),
.C(n_234),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_236),
.A2(n_237),
.B1(n_262),
.B2(n_265),
.Y(n_402)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_238),
.C(n_240),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_238),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_245),
.B(n_246),
.Y(n_323)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_250),
.A2(n_322),
.B(n_325),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_251),
.B(n_252),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_284),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_255),
.C(n_284),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_276),
.B2(n_277),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_256),
.B(n_278),
.C(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_266),
.B2(n_267),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_268),
.C(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_260),
.B(n_262),
.C(n_264),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_265),
.Y(n_261)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_274),
.B2(n_275),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_270),
.A2(n_271),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_272),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_282),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_287),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_320),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_303),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_289),
.B(n_303),
.C(n_320),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_294),
.C(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_302),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_301),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_295),
.Y(n_301)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_312),
.B2(n_313),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_304),
.B(n_314),
.C(n_319),
.Y(n_330)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_308),
.B2(n_311),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_306),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_306),
.B(n_309),
.C(n_310),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_306),
.A2(n_311),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_318),
.B2(n_319),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_328),
.B(n_329),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_352),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_331),
.CI(n_350),
.CON(n_329),
.SN(n_329)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_343),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_336),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_336),
.C(n_343),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_338),
.B1(n_339),
.B2(n_342),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_337),
.A2(n_338),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_338),
.B(n_340),
.C(n_341),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_347),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_348),
.C(n_349),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_346),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_373),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_355),
.B1(n_371),
.B2(n_372),
.Y(n_353)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_372),
.C(n_373),
.Y(n_377)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_SL g355 ( 
.A(n_356),
.B(n_364),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_365),
.C(n_370),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_360),
.C(n_362),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_362),
.B2(n_363),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_360),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_369),
.B2(n_370),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_377),
.B(n_378),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_379),
.B(n_380),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_381),
.C(n_390),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_390),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_385),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_387),
.C(n_388),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_383),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_386),
.A2(n_387),
.B1(n_388),
.B2(n_389),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_387),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_404),
.Y(n_392)
);

OR2x2_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_394),
.B(n_395),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_403),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_397),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_398),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_400),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_402),
.Y(n_401)
);


endmodule