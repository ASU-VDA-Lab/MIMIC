module fake_jpeg_26177_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_5),
.B(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_16),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_39),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_31),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_43),
.B(n_44),
.Y(n_82)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_48),
.Y(n_80)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_21),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_51),
.B(n_53),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_21),
.Y(n_53)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_62),
.B(n_73),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_33),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_65),
.A2(n_47),
.B1(n_55),
.B2(n_84),
.Y(n_99)
);

OAI32xp33_ASAP7_75t_L g66 ( 
.A1(n_46),
.A2(n_19),
.A3(n_33),
.B1(n_39),
.B2(n_32),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_66),
.B(n_41),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_69),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_58),
.A2(n_19),
.B1(n_25),
.B2(n_32),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_70),
.A2(n_22),
.B1(n_27),
.B2(n_24),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_25),
.B1(n_19),
.B2(n_29),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_74),
.A2(n_77),
.B1(n_22),
.B2(n_24),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_45),
.A2(n_25),
.B1(n_29),
.B2(n_18),
.Y(n_77)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_84),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_38),
.C(n_37),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_85),
.B(n_35),
.C(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_93),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_112),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_91),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_66),
.A2(n_22),
.B(n_24),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_92),
.A2(n_99),
.B(n_27),
.Y(n_117)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_60),
.B1(n_59),
.B2(n_38),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_94),
.A2(n_96),
.B1(n_103),
.B2(n_108),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_86),
.A2(n_59),
.B1(n_38),
.B2(n_45),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_68),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_104),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_86),
.A2(n_55),
.B1(n_41),
.B2(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_105),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_18),
.Y(n_107)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_107),
.B(n_20),
.Y(n_124)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_28),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_110),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_114),
.B(n_121),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_67),
.B1(n_83),
.B2(n_73),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_120),
.B1(n_132),
.B2(n_89),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_117),
.A2(n_20),
.B(n_23),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_95),
.A2(n_83),
.B1(n_76),
.B2(n_64),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_125),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_124),
.B(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_104),
.B1(n_108),
.B2(n_112),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_128),
.A2(n_80),
.B1(n_34),
.B2(n_35),
.Y(n_151)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_27),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_76),
.B1(n_64),
.B2(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_135),
.Y(n_158)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_35),
.Y(n_166)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_143),
.Y(n_168)
);

OA21x2_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_87),
.B(n_88),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_140),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_141),
.A2(n_147),
.B1(n_165),
.B2(n_26),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_88),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_142),
.B(n_167),
.Y(n_190)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_93),
.B1(n_87),
.B2(n_106),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_149),
.B1(n_150),
.B2(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_151),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_148),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_122),
.A2(n_106),
.B1(n_109),
.B2(n_62),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_138),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_79),
.B1(n_63),
.B2(n_101),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_79),
.B1(n_63),
.B2(n_111),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_159),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_34),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_117),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_154),
.A2(n_26),
.B(n_28),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_68),
.B1(n_17),
.B2(n_34),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_123),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_0),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_17),
.B1(n_23),
.B2(n_28),
.Y(n_165)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_166),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_35),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_140),
.Y(n_196)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_119),
.B(n_131),
.C(n_121),
.D(n_114),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_150),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_163),
.A2(n_133),
.B1(n_113),
.B2(n_135),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_180),
.B1(n_193),
.B2(n_26),
.Y(n_210)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_134),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_191),
.B(n_10),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_160),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_164),
.A2(n_113),
.B1(n_17),
.B2(n_35),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_17),
.C(n_23),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_181),
.B(n_187),
.C(n_162),
.Y(n_204)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_160),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_184),
.B(n_188),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_2),
.B(n_3),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_23),
.C(n_26),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_164),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_23),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_149),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_143),
.A2(n_26),
.B1(n_1),
.B2(n_2),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_182),
.A2(n_141),
.B1(n_145),
.B2(n_144),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_214),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_196),
.B(n_197),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_170),
.B(n_140),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_199),
.B(n_202),
.Y(n_222)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_201),
.Y(n_219)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_211),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_139),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_212),
.Y(n_227)
);

NOR2x1_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_148),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_178),
.A2(n_146),
.B1(n_157),
.B2(n_156),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_210),
.B1(n_189),
.B2(n_3),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_157),
.Y(n_209)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_209),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_175),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_8),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_213),
.A2(n_193),
.B1(n_172),
.B2(n_180),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_216),
.B(n_185),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_181),
.C(n_176),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_220),
.B(n_228),
.C(n_203),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_205),
.B1(n_210),
.B2(n_200),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_187),
.C(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_201),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_2),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_10),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_205),
.A2(n_172),
.B1(n_183),
.B2(n_191),
.Y(n_232)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_233),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_197),
.B(n_196),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_249),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_223),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_243),
.B1(n_232),
.B2(n_230),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_224),
.A2(n_225),
.B(n_229),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_240),
.A2(n_247),
.B(n_222),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_221),
.A2(n_207),
.B1(n_194),
.B2(n_213),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_212),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_246),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_220),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_244),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_218),
.B(n_216),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_10),
.B(n_14),
.Y(n_247)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_248),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_252),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_256),
.B1(n_242),
.B2(n_237),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_228),
.Y(n_252)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_259),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_241),
.A2(n_226),
.B1(n_219),
.B2(n_227),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_236),
.B(n_227),
.C(n_11),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_247),
.C(n_235),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_8),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_8),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_248),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_264),
.C(n_265),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_263),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_258),
.C(n_253),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_259),
.C(n_11),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_243),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_11),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_270),
.Y(n_275)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_261),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_3),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_242),
.B(n_238),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_5),
.B(n_6),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_274),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_262),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_278),
.B(n_280),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_279),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_267),
.B(n_12),
.C(n_13),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_275),
.B(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_285),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_273),
.Y(n_287)
);

NAND3xp33_ASAP7_75t_SL g290 ( 
.A(n_287),
.B(n_289),
.C(n_285),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_282),
.B(n_274),
.Y(n_289)
);

AO21x2_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_288),
.B(n_286),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_291),
.A2(n_283),
.B(n_266),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_292),
.B(n_267),
.C(n_265),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_293),
.B(n_12),
.C(n_3),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_294),
.B(n_4),
.Y(n_295)
);


endmodule