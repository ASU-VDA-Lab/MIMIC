module real_jpeg_25129_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_244;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_1),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_2),
.A2(n_28),
.B1(n_53),
.B2(n_54),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_21),
.B1(n_23),
.B2(n_54),
.Y(n_117)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_54),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_2),
.A2(n_54),
.B1(n_67),
.B2(n_68),
.Y(n_189)
);

BUFx8_ASAP7_75t_L g67 ( 
.A(n_3),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_6),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_21),
.B1(n_23),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_6),
.A2(n_30),
.B1(n_46),
.B2(n_48),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_6),
.A2(n_30),
.B1(n_67),
.B2(n_68),
.Y(n_131)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_7),
.A2(n_20),
.B1(n_24),
.B2(n_28),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_21),
.B1(n_23),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_8),
.A2(n_38),
.B1(n_46),
.B2(n_48),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_38),
.B1(n_67),
.B2(n_68),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_9),
.A2(n_21),
.B1(n_23),
.B2(n_33),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_33),
.B1(n_46),
.B2(n_48),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_9),
.A2(n_33),
.B1(n_67),
.B2(n_68),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_20),
.C(n_23),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_9),
.B(n_19),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_9),
.B(n_43),
.C(n_46),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_64),
.C(n_67),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_9),
.B(n_96),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_9),
.B(n_113),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_9),
.B(n_57),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_11),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_11),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_86),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_85),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_70),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_16),
.B(n_70),
.Y(n_85)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_16),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g16 ( 
.A(n_17),
.B(n_36),
.CI(n_49),
.CON(n_16),
.SN(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_25),
.B(n_31),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_18),
.A2(n_31),
.B(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_19),
.A2(n_32),
.B1(n_34),
.B2(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_34),
.Y(n_106)
);

AO22x1_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_21),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_21),
.A2(n_23),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_23),
.B(n_218),
.Y(n_217)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_41),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_40),
.A2(n_45),
.B(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_41),
.B(n_84),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_41),
.A2(n_57),
.B1(n_84),
.B2(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_45),
.Y(n_41)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_43),
.Y(n_44)
);

OA22x2_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_44),
.B1(n_46),
.B2(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_45),
.A2(n_82),
.B(n_83),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_45),
.A2(n_83),
.B(n_117),
.Y(n_138)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_46),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_48),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_46),
.B(n_231),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_55),
.C(n_58),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_72),
.B1(n_75),
.B2(n_76),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g128 ( 
.A(n_50),
.B(n_129),
.C(n_137),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_50),
.A2(n_76),
.B1(n_137),
.B2(n_138),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_50),
.A2(n_76),
.B1(n_115),
.B2(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_50),
.B(n_115),
.C(n_182),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_53),
.B(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_55),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_80),
.C(n_81),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_58),
.A2(n_74),
.B1(n_81),
.B2(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_69),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_60),
.B(n_103),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_66),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_62),
.A2(n_103),
.B1(n_113),
.B2(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_64),
.Y(n_65)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_65),
.B1(n_67),
.B2(n_68),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_66),
.A2(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_66),
.A2(n_102),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_67),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_67),
.B(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_77),
.C(n_78),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_71),
.A2(n_77),
.B1(n_80),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_77),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_77),
.A2(n_80),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_77),
.B(n_156),
.C(n_164),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_77),
.A2(n_80),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_77),
.A2(n_80),
.B1(n_164),
.B2(n_272),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_79),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_80),
.B(n_137),
.C(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_81),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_84),
.Y(n_165)
);

OAI211xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_139),
.B(n_146),
.C(n_284),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_123),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_123),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_108),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_89),
.B(n_110),
.C(n_118),
.Y(n_141)
);

AOI21xp33_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_99),
.B(n_104),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_100),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_104),
.B1(n_105),
.B2(n_126),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_90),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_90),
.A2(n_100),
.B1(n_126),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_91),
.B(n_98),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_92),
.B(n_190),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_95),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_93),
.A2(n_98),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_93),
.B(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_93),
.Y(n_188)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_97),
.A2(n_131),
.B(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g203 ( 
.A(n_97),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_99),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_100),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_118),
.B2(n_119),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_110),
.A2(n_111),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.Y(n_110)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_115),
.B(n_202),
.C(n_204),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_115),
.A2(n_192),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_127),
.C(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_127),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_152),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_130),
.Y(n_275)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_134),
.A2(n_135),
.B1(n_246),
.B2(n_247),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_134),
.A2(n_135),
.B1(n_215),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_135),
.B(n_209),
.C(n_215),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_135),
.B(n_187),
.C(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_137),
.A2(n_138),
.B1(n_178),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_137),
.A2(n_138),
.B1(n_162),
.B2(n_175),
.Y(n_252)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_138),
.B(n_162),
.C(n_253),
.Y(n_256)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

NAND3xp33_ASAP7_75t_SL g146 ( 
.A(n_140),
.B(n_147),
.C(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_141),
.B(n_142),
.Y(n_284)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_168),
.B(n_283),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_166),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_150),
.B(n_166),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.C(n_155),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_151),
.B(n_153),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_155),
.B(n_281),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_156),
.A2(n_157),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_162),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_189),
.B(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_161),
.Y(n_190)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_162),
.A2(n_175),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_162),
.B(n_232),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_164),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_278),
.B(n_282),
.Y(n_168)
);

A2O1A1Ixp33_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_205),
.B(n_264),
.C(n_277),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_194),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_171),
.B(n_194),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_181),
.B2(n_193),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_177),
.B1(n_179),
.B2(n_180),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_174),
.B(n_180),
.C(n_193),
.Y(n_265)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_191),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_183),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_186),
.A2(n_187),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_238),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_200),
.C(n_201),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_196),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_201),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_202),
.A2(n_204),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_202),
.B(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_204),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_263),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_224),
.B(n_262),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_221),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_208),
.B(n_221),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_209),
.A2(n_210),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_214),
.B(n_229),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_215),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_219),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_216),
.A2(n_217),
.B1(n_219),
.B2(n_220),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_255),
.B(n_261),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_249),
.B(n_254),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_241),
.B(n_248),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_240),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_230),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_237),
.B(n_239),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_243),
.Y(n_248)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_246),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_250),
.B(n_251),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_256),
.B(n_257),
.Y(n_261)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_266),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_273),
.B2(n_274),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_274),
.C(n_276),
.Y(n_279)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);


endmodule