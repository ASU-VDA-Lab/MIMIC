module fake_jpeg_16501_n_265 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_265);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_265;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx24_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

CKINVDCx6p67_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_18),
.B(n_13),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_41),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx2_ASAP7_75t_SL g82 ( 
.A(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_21),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_17),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_51),
.B1(n_59),
.B2(n_15),
.Y(n_67)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_53),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_41),
.A2(n_22),
.B1(n_29),
.B2(n_18),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_54),
.B(n_57),
.Y(n_66)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_33),
.A2(n_22),
.B1(n_21),
.B2(n_24),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_24),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_36),
.A2(n_22),
.B1(n_29),
.B2(n_19),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_29),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_60),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_28),
.B1(n_26),
.B2(n_31),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_23),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_23),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_74),
.B1(n_44),
.B2(n_48),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_17),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_68),
.B(n_73),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_26),
.B1(n_31),
.B2(n_20),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_77),
.Y(n_95)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_52),
.B(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_86),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_83),
.Y(n_102)
);

AND2x4_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_15),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_60),
.C(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_50),
.A2(n_20),
.B1(n_31),
.B2(n_23),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_59),
.B1(n_44),
.B2(n_48),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_57),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_65),
.B1(n_15),
.B2(n_31),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_17),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_87),
.A2(n_97),
.B1(n_99),
.B2(n_103),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_98),
.C(n_104),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_106),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_92),
.A2(n_93),
.B1(n_81),
.B2(n_74),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_76),
.A2(n_54),
.B1(n_64),
.B2(n_62),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_69),
.B(n_56),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_79),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_77),
.A2(n_64),
.B1(n_63),
.B2(n_62),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_35),
.C(n_42),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_83),
.A2(n_67),
.B1(n_66),
.B2(n_85),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_64),
.B1(n_45),
.B2(n_65),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_46),
.Y(n_104)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_72),
.A2(n_65),
.A3(n_61),
.B1(n_42),
.B2(n_35),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_58),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_58),
.C(n_25),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_80),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_110),
.B(n_113),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_118),
.C(n_98),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_116),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_104),
.B(n_72),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_85),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_117),
.B(n_131),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_80),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_124),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_101),
.A2(n_66),
.B1(n_80),
.B2(n_69),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_125),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_101),
.A2(n_80),
.B1(n_78),
.B2(n_70),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_80),
.B1(n_70),
.B2(n_82),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_91),
.B(n_75),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_127),
.B(n_128),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_96),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_87),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_8),
.B(n_13),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_96),
.B(n_25),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_133),
.A2(n_106),
.B(n_45),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_120),
.A2(n_102),
.B(n_95),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_139),
.A2(n_156),
.B(n_124),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_129),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_140),
.B(n_146),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_117),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_123),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_145),
.B(n_150),
.C(n_153),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_112),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_147),
.B(n_0),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_103),
.B1(n_93),
.B2(n_97),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_111),
.B1(n_142),
.B2(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_108),
.C(n_84),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_84),
.C(n_25),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_107),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_0),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_84),
.C(n_25),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_155),
.B(n_27),
.C(n_25),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_110),
.A2(n_15),
.B(n_1),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_159),
.A2(n_137),
.B1(n_147),
.B2(n_156),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_141),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_165),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_162),
.B(n_166),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_114),
.B(n_122),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_167),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_136),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_114),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_125),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_115),
.B1(n_100),
.B2(n_45),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_168),
.A2(n_140),
.B1(n_146),
.B2(n_141),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_171),
.B(n_174),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_25),
.C(n_27),
.Y(n_174)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_45),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g191 ( 
.A(n_176),
.B(n_138),
.CI(n_134),
.CON(n_191),
.SN(n_191)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_30),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_180),
.B(n_151),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_187),
.B1(n_199),
.B2(n_171),
.Y(n_206)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_137),
.A3(n_148),
.B1(n_138),
.B2(n_152),
.C1(n_134),
.C2(n_157),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_167),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_197),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_154),
.Y(n_189)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_189),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_178),
.B(n_151),
.Y(n_192)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_160),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_200),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_135),
.B1(n_45),
.B2(n_3),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_170),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_2),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_30),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_169),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_159),
.A2(n_172),
.B1(n_168),
.B2(n_162),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_161),
.A2(n_166),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_205),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_192),
.A2(n_176),
.B(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_188),
.B(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_206),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_158),
.C(n_163),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_209),
.B(n_213),
.C(n_214),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_215),
.Y(n_222)
);

AOI31xp67_ASAP7_75t_L g212 ( 
.A1(n_185),
.A2(n_8),
.A3(n_11),
.B(n_10),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_216),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_30),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_30),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_30),
.Y(n_215)
);

AOI31xp67_ASAP7_75t_L g216 ( 
.A1(n_185),
.A2(n_11),
.A3(n_9),
.B(n_16),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_188),
.B(n_9),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_181),
.C(n_191),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g218 ( 
.A(n_208),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_211),
.Y(n_235)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_2),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_186),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_229),
.Y(n_234)
);

OAI31xp33_ASAP7_75t_L g228 ( 
.A1(n_207),
.A2(n_200),
.A3(n_189),
.B(n_197),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_16),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_184),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_230),
.B(n_209),
.Y(n_233)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_205),
.A2(n_195),
.B(n_182),
.C(n_196),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_214),
.B(n_217),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_241),
.B(n_228),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_236),
.C(n_240),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_235),
.B(n_239),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_220),
.C(n_222),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_194),
.B1(n_181),
.B2(n_213),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_222),
.B(n_221),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_238),
.B(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_16),
.C(n_3),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_9),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_2),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_243),
.B(n_4),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_246),
.A2(n_247),
.B(n_4),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_251),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_221),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_250),
.A2(n_252),
.B(n_4),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_230),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_16),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_246),
.A2(n_244),
.B(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_253),
.B(n_254),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_5),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_256),
.B(n_6),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_258),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_257),
.C(n_7),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_7),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_259),
.Y(n_264)
);


endmodule