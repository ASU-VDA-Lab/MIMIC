module fake_jpeg_26240_n_130 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_130);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_130;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_7),
.B(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_29),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp67_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_0),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_37),
.C(n_24),
.Y(n_51)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_24),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_48),
.Y(n_61)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_18),
.B1(n_20),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_52),
.B1(n_38),
.B2(n_21),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_38),
.B1(n_18),
.B2(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_54),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_51),
.B(n_37),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_37),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_63),
.C(n_64),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_45),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_58),
.A2(n_42),
.B1(n_30),
.B2(n_43),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_66),
.B1(n_69),
.B2(n_71),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_33),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_31),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_47),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_67),
.B(n_23),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_40),
.A2(n_31),
.B1(n_17),
.B2(n_16),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_46),
.A2(n_26),
.B(n_31),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_56),
.C(n_61),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_50),
.A2(n_31),
.B1(n_34),
.B2(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_14),
.B1(n_23),
.B2(n_34),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_85),
.Y(n_93)
);

A2O1A1O1Ixp25_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_20),
.B(n_30),
.C(n_28),
.D(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_83),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_77),
.B1(n_82),
.B2(n_67),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_42),
.B1(n_44),
.B2(n_30),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_59),
.B1(n_62),
.B2(n_70),
.Y(n_90)
);

AND2x6_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_8),
.Y(n_83)
);

OAI21xp33_ASAP7_75t_SL g95 ( 
.A1(n_84),
.A2(n_65),
.B(n_60),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_63),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_28),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_65),
.C(n_67),
.Y(n_89)
);

AOI221xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_89),
.B1(n_80),
.B2(n_88),
.C(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_91),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_92),
.B(n_96),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_61),
.B1(n_71),
.B2(n_53),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_97),
.Y(n_100)
);

AO22x1_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_84),
.B1(n_94),
.B2(n_97),
.Y(n_107)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_54),
.B1(n_66),
.B2(n_69),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_91),
.C(n_57),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_102),
.A2(n_103),
.B(n_104),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_93),
.Y(n_104)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_106),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_107),
.A2(n_86),
.B(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_90),
.B1(n_74),
.B2(n_77),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_108),
.A2(n_111),
.B1(n_100),
.B2(n_107),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_114),
.B(n_106),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_83),
.C(n_57),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_105),
.A2(n_1),
.B(n_2),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_3),
.C(n_5),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_110),
.B(n_100),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_3),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_2),
.B(n_3),
.Y(n_119)
);

AOI322xp5_ASAP7_75t_L g120 ( 
.A1(n_117),
.A2(n_111),
.A3(n_114),
.B1(n_10),
.B2(n_11),
.C1(n_12),
.C2(n_7),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_120),
.A2(n_12),
.B(n_6),
.Y(n_126)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_121),
.B(n_123),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_122),
.B(n_5),
.C(n_6),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_126),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_124),
.Y(n_127)
);

OAI31xp33_ASAP7_75t_L g129 ( 
.A1(n_127),
.A2(n_122),
.A3(n_6),
.B(n_7),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_129),
.B(n_128),
.Y(n_130)
);


endmodule