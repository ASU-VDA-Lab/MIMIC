module fake_jpeg_6731_n_71 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_71);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_71;

wire n_57;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_51;
wire n_47;
wire n_22;
wire n_40;
wire n_19;
wire n_18;
wire n_59;
wire n_20;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_36;
wire n_62;
wire n_31;
wire n_25;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_50;
wire n_29;
wire n_32;
wire n_70;
wire n_66;

INVx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_39),
.Y(n_48)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_35),
.Y(n_49)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_31),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_0),
.Y(n_40)
);

BUFx24_ASAP7_75t_SL g51 ( 
.A(n_40),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_4),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_4),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.C(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_7),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_59),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_48),
.A2(n_46),
.B(n_35),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_57),
.C(n_58),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_53),
.A2(n_46),
.B(n_39),
.Y(n_57)
);

XNOR2x1_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_21),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_47),
.B(n_7),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_47),
.B1(n_54),
.B2(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_59),
.A2(n_20),
.B1(n_50),
.B2(n_29),
.Y(n_61)
);

XNOR2x1_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_52),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.C(n_20),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_65),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_62),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_22),
.B(n_14),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_67),
.C(n_16),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_8),
.Y(n_71)
);


endmodule