module fake_jpeg_484_n_438 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_438);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_0),
.B(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

NAND2xp33_ASAP7_75t_SL g106 ( 
.A(n_46),
.B(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

CKINVDCx9p33_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_61),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_52),
.Y(n_104)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_16),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_69),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g66 ( 
.A(n_31),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

BUFx12f_ASAP7_75t_SL g67 ( 
.A(n_31),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_68),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_15),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_19),
.Y(n_72)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_73),
.B(n_81),
.Y(n_135)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_74),
.B(n_76),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_78),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_79),
.Y(n_132)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_82),
.B(n_83),
.Y(n_114)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_15),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_84),
.B(n_42),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_85),
.B(n_86),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_26),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_87),
.B(n_29),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_29),
.B1(n_26),
.B2(n_27),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_93),
.B1(n_107),
.B2(n_109),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_44),
.B(n_29),
.C(n_26),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_92),
.B(n_55),
.C(n_82),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_72),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_78),
.A2(n_18),
.B1(n_42),
.B2(n_20),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_101),
.A2(n_113),
.B1(n_118),
.B2(n_127),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_27),
.B1(n_36),
.B2(n_20),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_134),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_63),
.A2(n_27),
.B1(n_36),
.B2(n_22),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_L g113 ( 
.A1(n_53),
.A2(n_36),
.B1(n_40),
.B2(n_43),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_43),
.B1(n_40),
.B2(n_25),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_58),
.B1(n_2),
.B2(n_3),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_71),
.A2(n_32),
.B1(n_24),
.B2(n_22),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_32),
.B1(n_24),
.B2(n_43),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_62),
.B(n_30),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_23),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_85),
.B(n_40),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_79),
.A2(n_23),
.B1(n_30),
.B2(n_2),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_136),
.A2(n_46),
.B1(n_30),
.B2(n_87),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g185 ( 
.A(n_137),
.B(n_142),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_129),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_88),
.B1(n_131),
.B2(n_121),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_104),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_133),
.B(n_70),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_148),
.Y(n_187)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_124),
.Y(n_147)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_0),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_90),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_150),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_90),
.B(n_1),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_92),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_151),
.B(n_176),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_60),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_152),
.Y(n_196)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_153),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_60),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_155),
.B(n_166),
.C(n_91),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_99),
.B(n_1),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_158),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_111),
.B(n_1),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_106),
.B(n_2),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_159),
.B(n_167),
.Y(n_194)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_106),
.A2(n_3),
.B(n_4),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_174),
.B(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_164),
.A2(n_125),
.B1(n_121),
.B2(n_102),
.Y(n_203)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_4),
.C(n_5),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_6),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_168),
.Y(n_208)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_170),
.Y(n_189)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_172),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_91),
.B(n_6),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_107),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_89),
.B1(n_104),
.B2(n_125),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_114),
.A2(n_7),
.B(n_8),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_89),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_175),
.B(n_178),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_123),
.B(n_7),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_114),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_8),
.Y(n_215)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_113),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_127),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_179),
.B(n_180),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_116),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_182),
.A2(n_199),
.B1(n_203),
.B2(n_140),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

NAND3xp33_ASAP7_75t_L g246 ( 
.A(n_184),
.B(n_186),
.C(n_197),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_141),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_178),
.A2(n_89),
.B1(n_103),
.B2(n_120),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_192),
.A2(n_180),
.B(n_174),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_215),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_179),
.A2(n_123),
.B1(n_116),
.B2(n_131),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_205),
.B(n_142),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_103),
.B1(n_105),
.B2(n_117),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_207),
.Y(n_221)
);

AO22x1_ASAP7_75t_SL g211 ( 
.A1(n_154),
.A2(n_112),
.B1(n_119),
.B2(n_105),
.Y(n_211)
);

OA21x2_ASAP7_75t_L g238 ( 
.A1(n_211),
.A2(n_143),
.B(n_177),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_138),
.B(n_119),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_216),
.B(n_171),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_151),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_217),
.B(n_236),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_239),
.Y(n_258)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_210),
.Y(n_219)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_200),
.B(n_148),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_220),
.B(n_222),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_144),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_159),
.B(n_161),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_229),
.B(n_241),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_143),
.B1(n_137),
.B2(n_142),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_238),
.B1(n_217),
.B2(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_181),
.Y(n_225)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_243),
.Y(n_264)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_227),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_228),
.B(n_185),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_213),
.A2(n_211),
.B1(n_184),
.B2(n_198),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_196),
.B1(n_207),
.B2(n_191),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_193),
.B(n_195),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_232),
.B(n_235),
.Y(n_267)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_191),
.C(n_196),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_165),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_187),
.B(n_149),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_176),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_240),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_189),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_150),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_213),
.A2(n_159),
.B(n_152),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_188),
.B(n_145),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_245),
.Y(n_274)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_201),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_247),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_162),
.Y(n_245)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_201),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_248),
.B(n_167),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_259),
.B1(n_246),
.B2(n_241),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g285 ( 
.A(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_252),
.B(n_255),
.C(n_265),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_254),
.A2(n_211),
.B(n_182),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_234),
.C(n_205),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_242),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_257),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_218),
.B(n_232),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_239),
.A2(n_207),
.B1(n_212),
.B2(n_189),
.Y(n_259)
);

AND2x2_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_205),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_212),
.B1(n_199),
.B2(n_211),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_261),
.A2(n_231),
.B1(n_221),
.B2(n_226),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_228),
.B(n_185),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_269),
.B(n_225),
.Y(n_299)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_230),
.A2(n_215),
.A3(n_194),
.B1(n_195),
.B2(n_185),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_276),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_193),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_271),
.B(n_240),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_234),
.B(n_185),
.C(n_152),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_273),
.B(n_155),
.C(n_152),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_SL g275 ( 
.A1(n_223),
.A2(n_194),
.B(n_214),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_275),
.A2(n_192),
.B(n_186),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_220),
.B(n_211),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_279),
.B(n_291),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_280),
.B(n_282),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_238),
.B1(n_221),
.B2(n_246),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_281),
.A2(n_289),
.B1(n_292),
.B2(n_262),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_245),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_277),
.Y(n_284)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_251),
.Y(n_287)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_287),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_224),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_288),
.B(n_293),
.Y(n_317)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_290),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_258),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_238),
.B1(n_229),
.B2(n_230),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_237),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_260),
.B(n_155),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_304),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_236),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_295),
.B(n_303),
.C(n_305),
.Y(n_307)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_298),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_299),
.B(n_302),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_265),
.B(n_227),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_258),
.B(n_204),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_252),
.B(n_247),
.C(n_243),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_306),
.A2(n_264),
.B(n_250),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_309),
.A2(n_330),
.B1(n_306),
.B2(n_270),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_286),
.A2(n_254),
.B1(n_276),
.B2(n_274),
.Y(n_310)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_269),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_322),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_260),
.C(n_273),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_325),
.C(n_331),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_286),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_318),
.B(n_321),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_285),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_260),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_292),
.A2(n_262),
.B(n_264),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_323),
.A2(n_326),
.B(n_313),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_305),
.B(n_249),
.C(n_263),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_291),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_283),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_263),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_300),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_300),
.A2(n_268),
.B1(n_274),
.B2(n_253),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_294),
.B(n_268),
.C(n_278),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_297),
.C(n_299),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_334),
.B(n_343),
.C(n_344),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_318),
.B(n_266),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_335),
.B(n_340),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_336),
.B(n_345),
.Y(n_362)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_330),
.B(n_266),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_313),
.A2(n_289),
.B1(n_284),
.B2(n_281),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_342),
.A2(n_324),
.B1(n_316),
.B2(n_327),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_307),
.B(n_297),
.C(n_303),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_279),
.C(n_296),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_325),
.B(n_298),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_346),
.A2(n_308),
.B1(n_332),
.B2(n_329),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_315),
.B(n_204),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_347),
.B(n_348),
.Y(n_360)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_311),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_328),
.B(n_219),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_353),
.Y(n_361)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_350),
.A2(n_323),
.B(n_326),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_317),
.B(n_278),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_352),
.B(n_338),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_314),
.B(n_298),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_321),
.B(n_287),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_354),
.B(n_332),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_366),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_356),
.B(n_155),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_324),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_358),
.B(n_368),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_359),
.A2(n_363),
.B1(n_367),
.B2(n_342),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_337),
.A2(n_311),
.B1(n_327),
.B2(n_308),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_350),
.Y(n_364)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_365),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_333),
.B(n_322),
.C(n_331),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_354),
.B(n_272),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_336),
.B(n_344),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_369),
.B(n_343),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_319),
.C(n_272),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_371),
.B(n_351),
.Y(n_379)
);

AND2x6_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_319),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_373),
.A2(n_233),
.B(n_244),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_376),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_364),
.A2(n_341),
.B1(n_346),
.B2(n_334),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_375),
.A2(n_359),
.B1(n_361),
.B2(n_370),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_366),
.B(n_345),
.C(n_351),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_386),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_380),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_372),
.B(n_219),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_381),
.A2(n_363),
.B1(n_358),
.B2(n_190),
.Y(n_396)
);

XOR2x2_ASAP7_75t_SL g382 ( 
.A(n_362),
.B(n_320),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_383),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_360),
.B(n_208),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_388),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_190),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_357),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_357),
.C(n_371),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_396),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_397),
.Y(n_404)
);

OAI321xp33_ASAP7_75t_L g394 ( 
.A1(n_387),
.A2(n_358),
.A3(n_378),
.B1(n_385),
.B2(n_368),
.C(n_377),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_394),
.B(n_399),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_374),
.A2(n_373),
.B1(n_182),
.B2(n_203),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_398),
.A2(n_403),
.B1(n_146),
.B2(n_210),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_382),
.C(n_375),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_190),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_400),
.B(n_160),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_169),
.B1(n_170),
.B2(n_146),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_389),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_406),
.B(n_407),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_390),
.B(n_163),
.C(n_208),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_410),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_402),
.A2(n_175),
.B(n_210),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_409),
.A2(n_167),
.B(n_160),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_395),
.B(n_166),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_411),
.B(n_414),
.Y(n_421)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_391),
.B(n_209),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_415),
.C(n_397),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_393),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_401),
.B(n_399),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_416),
.A2(n_404),
.B1(n_408),
.B2(n_147),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_412),
.B(n_209),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_424),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_405),
.A2(n_209),
.B(n_168),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_419),
.A2(n_423),
.B(n_100),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_404),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_413),
.B(n_160),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_406),
.B(n_153),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_425),
.A2(n_426),
.B(n_428),
.Y(n_432)
);

AOI221xp5_ASAP7_75t_L g431 ( 
.A1(n_427),
.A2(n_429),
.B1(n_423),
.B2(n_430),
.C(n_420),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_100),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_431),
.A2(n_433),
.B(n_11),
.Y(n_435)
);

O2A1O1Ixp33_ASAP7_75t_SL g433 ( 
.A1(n_429),
.A2(n_102),
.B(n_122),
.C(n_117),
.Y(n_433)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_432),
.B(n_122),
.C(n_12),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_434),
.B(n_435),
.C(n_11),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_436),
.A2(n_13),
.B(n_14),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_14),
.B(n_95),
.Y(n_438)
);


endmodule