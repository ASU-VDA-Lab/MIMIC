module fake_jpeg_16782_n_92 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_92);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_92;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_4),
.B(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_0),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_18),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_24),
.A2(n_29),
.B1(n_33),
.B2(n_22),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g26 ( 
.A1(n_16),
.A2(n_1),
.B(n_2),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_13),
.C(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_32),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_21),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_19),
.A2(n_20),
.B1(n_22),
.B2(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_42),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_37),
.A2(n_51),
.B1(n_49),
.B2(n_45),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_24),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_41),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_27),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_35),
.B(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_33),
.A2(n_17),
.B1(n_14),
.B2(n_5),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_47),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_31),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.C(n_50),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_29),
.A2(n_6),
.B1(n_14),
.B2(n_10),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_14),
.C(n_32),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_23),
.A2(n_10),
.B1(n_24),
.B2(n_33),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_54),
.B1(n_47),
.B2(n_48),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_51),
.B1(n_36),
.B2(n_34),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_38),
.B1(n_40),
.B2(n_52),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_50),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_39),
.C(n_41),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_68),
.C(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_67),
.B(n_71),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_38),
.B1(n_56),
.B2(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_59),
.Y(n_71)
);

OAI31xp33_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_59),
.A3(n_62),
.B(n_64),
.Y(n_72)
);

OAI21x1_ASAP7_75t_SL g75 ( 
.A1(n_72),
.A2(n_70),
.B(n_73),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_53),
.B1(n_56),
.B2(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_77),
.B(n_79),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_66),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_65),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_71),
.C(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_81),
.A2(n_74),
.B(n_68),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_72),
.B(n_69),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_83),
.A2(n_86),
.B(n_85),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_76),
.C(n_82),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_80),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_82),
.C(n_78),
.Y(n_92)
);


endmodule