module fake_jpeg_4522_n_242 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx8_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_37),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_21),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_39),
.B(n_27),
.Y(n_49)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_45),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_46),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_84),
.Y(n_101)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_52),
.Y(n_91)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_14),
.B1(n_30),
.B2(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_53),
.A2(n_77),
.B1(n_25),
.B2(n_19),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_14),
.B1(n_16),
.B2(n_31),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_86),
.B1(n_25),
.B2(n_19),
.Y(n_90)
);

BUFx8_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_55),
.Y(n_111)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_57),
.B(n_60),
.Y(n_96)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_64),
.Y(n_112)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_66),
.A2(n_76),
.B1(n_80),
.B2(n_81),
.Y(n_106)
);

CKINVDCx6p67_ASAP7_75t_R g68 ( 
.A(n_34),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_68),
.B(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_32),
.B(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_35),
.A2(n_14),
.B1(n_30),
.B2(n_24),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_72),
.A2(n_22),
.B1(n_15),
.B2(n_4),
.Y(n_99)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_35),
.A2(n_24),
.B1(n_19),
.B2(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_38),
.B(n_23),
.Y(n_79)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g84 ( 
.A(n_33),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_22),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_40),
.A2(n_16),
.B1(n_31),
.B2(n_23),
.Y(n_86)
);

INVx3_ASAP7_75t_SL g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_15),
.B1(n_27),
.B2(n_22),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_88),
.A2(n_110),
.B1(n_50),
.B2(n_71),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_89),
.B(n_104),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_97),
.B1(n_99),
.B2(n_62),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_85),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_58),
.B(n_29),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_66),
.B(n_76),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_25),
.B1(n_15),
.B2(n_28),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_81),
.B(n_29),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_98),
.B(n_2),
.Y(n_122)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_2),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_13),
.B1(n_3),
.B2(n_4),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_59),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_87),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_116),
.A2(n_121),
.B1(n_130),
.B2(n_104),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_94),
.B(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_120),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_118),
.B(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_48),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_122),
.A2(n_131),
.B(n_132),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_110),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_125),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_56),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_126),
.Y(n_157)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_128),
.B(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_114),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_106),
.A2(n_82),
.B(n_67),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_88),
.A2(n_68),
.B(n_80),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_140),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_101),
.B(n_62),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_139),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_136),
.A2(n_127),
.B1(n_135),
.B2(n_124),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_103),
.B(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_67),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_101),
.A2(n_55),
.B(n_75),
.C(n_8),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_141),
.B(n_104),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g142 ( 
.A1(n_88),
.A2(n_110),
.A3(n_99),
.B1(n_112),
.B2(n_90),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_108),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_95),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_144),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_88),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_149),
.A2(n_155),
.B(n_167),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_132),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_88),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_115),
.C(n_109),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_166),
.C(n_125),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_161),
.B(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_128),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_165),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_109),
.C(n_107),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_97),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_143),
.A2(n_107),
.B1(n_100),
.B2(n_61),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_169),
.A2(n_165),
.B1(n_148),
.B2(n_147),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_170),
.B(n_176),
.C(n_178),
.Y(n_196)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_181),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_146),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_173),
.A2(n_175),
.B1(n_178),
.B2(n_183),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_136),
.Y(n_174)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_174),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_127),
.B1(n_136),
.B2(n_139),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_167),
.A2(n_154),
.B1(n_169),
.B2(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_119),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_184),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_119),
.B1(n_92),
.B2(n_133),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_168),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_149),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g197 ( 
.A(n_185),
.B(n_187),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_149),
.B(n_118),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_179),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_190),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g193 ( 
.A1(n_187),
.A2(n_146),
.B(n_155),
.C(n_166),
.D(n_160),
.Y(n_193)
);

NOR3xp33_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_173),
.C(n_180),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_196),
.C(n_199),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_151),
.B1(n_145),
.B2(n_164),
.Y(n_198)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_164),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_150),
.C(n_145),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_203),
.C(n_157),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_157),
.C(n_158),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_195),
.A2(n_184),
.B1(n_186),
.B2(n_174),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_206),
.B1(n_212),
.B2(n_214),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_186),
.B1(n_177),
.B2(n_170),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_208),
.A2(n_210),
.B(n_201),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_209),
.A2(n_211),
.B(n_192),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_193),
.B(n_158),
.C(n_100),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_200),
.A2(n_111),
.B(n_6),
.Y(n_211)
);

NOR2xp67_ASAP7_75t_R g212 ( 
.A(n_197),
.B(n_55),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_212),
.B(n_197),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_206),
.C(n_204),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_216),
.A2(n_218),
.B(n_220),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_199),
.Y(n_229)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_219),
.B(n_221),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_213),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_202),
.B1(n_203),
.B2(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_222),
.B(n_209),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_204),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_111),
.C(n_75),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_226),
.A2(n_227),
.B(n_92),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_220),
.A2(n_208),
.B1(n_210),
.B2(n_194),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_223),
.A2(n_5),
.B(n_6),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_144),
.B1(n_140),
.B2(n_10),
.Y(n_235)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_6),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_232),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_229),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_235),
.A2(n_238),
.B(n_236),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_234),
.B(n_224),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_237),
.A2(n_227),
.B(n_9),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g241 ( 
.A1(n_239),
.A2(n_240),
.B(n_8),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_9),
.Y(n_242)
);


endmodule