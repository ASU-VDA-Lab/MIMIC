module real_aes_7581_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_555;
wire n_319;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_754;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_753;
wire n_741;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g273 ( .A1(n_0), .A2(n_274), .B(n_275), .C(n_278), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_1), .B(n_262), .Y(n_279) );
NAND3xp33_ASAP7_75t_SL g110 ( .A(n_2), .B(n_111), .C(n_112), .Y(n_110) );
INVx1_ASAP7_75t_L g125 ( .A(n_2), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_3), .B(n_190), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g533 ( .A1(n_4), .A2(n_151), .B(n_154), .C(n_534), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_5), .A2(n_146), .B(n_558), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_6), .A2(n_146), .B(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_7), .B(n_262), .Y(n_564) );
AO21x2_ASAP7_75t_L g217 ( .A1(n_8), .A2(n_181), .B(n_218), .Y(n_217) );
AND2x6_ASAP7_75t_L g151 ( .A(n_9), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g234 ( .A1(n_10), .A2(n_151), .B(n_154), .C(n_235), .Y(n_234) );
INVx1_ASAP7_75t_L g502 ( .A(n_11), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_12), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_12), .B(n_40), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g536 ( .A(n_13), .B(n_238), .Y(n_536) );
INVx1_ASAP7_75t_L g172 ( .A(n_14), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_15), .B(n_190), .Y(n_224) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_16), .A2(n_191), .B(n_520), .C(n_522), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_17), .B(n_262), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_18), .B(n_166), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_19), .A2(n_154), .B(n_157), .C(n_165), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_20), .A2(n_226), .B(n_277), .C(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_21), .B(n_238), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_22), .A2(n_54), .B1(n_756), .B2(n_757), .Y(n_755) );
CKINVDCx20_ASAP7_75t_R g756 ( .A(n_22), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_23), .B(n_238), .Y(n_475) );
CKINVDCx16_ASAP7_75t_R g549 ( .A(n_24), .Y(n_549) );
INVx1_ASAP7_75t_L g474 ( .A(n_25), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g220 ( .A1(n_26), .A2(n_154), .B(n_165), .C(n_221), .Y(n_220) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_27), .Y(n_150) );
CKINVDCx20_ASAP7_75t_R g532 ( .A(n_28), .Y(n_532) );
INVx1_ASAP7_75t_L g490 ( .A(n_29), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_30), .A2(n_146), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g149 ( .A(n_31), .Y(n_149) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_32), .A2(n_194), .B(n_203), .C(n_205), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_33), .Y(n_539) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_34), .A2(n_277), .B(n_561), .C(n_563), .Y(n_560) );
INVxp67_ASAP7_75t_L g491 ( .A(n_35), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_36), .B(n_223), .Y(n_222) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_37), .A2(n_154), .B(n_165), .C(n_473), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g559 ( .A(n_38), .Y(n_559) );
AOI222xp33_ASAP7_75t_SL g128 ( .A1(n_39), .A2(n_129), .B1(n_135), .B2(n_740), .C1(n_741), .C2(n_745), .Y(n_128) );
INVx1_ASAP7_75t_L g109 ( .A(n_40), .Y(n_109) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_41), .A2(n_278), .B(n_500), .C(n_501), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_42), .B(n_145), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g240 ( .A(n_43), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_44), .B(n_190), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_45), .B(n_146), .Y(n_219) );
CKINVDCx20_ASAP7_75t_R g477 ( .A(n_46), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_47), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_48), .A2(n_194), .B(n_203), .C(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g276 ( .A(n_49), .Y(n_276) );
OAI22xp5_ASAP7_75t_SL g753 ( .A1(n_50), .A2(n_754), .B1(n_755), .B2(n_758), .Y(n_753) );
CKINVDCx16_ASAP7_75t_R g758 ( .A(n_50), .Y(n_758) );
INVx1_ASAP7_75t_L g248 ( .A(n_51), .Y(n_248) );
INVx1_ASAP7_75t_L g508 ( .A(n_52), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_53), .B(n_146), .Y(n_245) );
CKINVDCx20_ASAP7_75t_R g757 ( .A(n_54), .Y(n_757) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_55), .Y(n_174) );
CKINVDCx14_ASAP7_75t_R g498 ( .A(n_56), .Y(n_498) );
INVx1_ASAP7_75t_L g152 ( .A(n_57), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_58), .B(n_146), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_59), .B(n_262), .Y(n_261) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_60), .A2(n_164), .B(n_187), .C(n_259), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_61), .Y(n_127) );
INVx1_ASAP7_75t_L g171 ( .A(n_62), .Y(n_171) );
OAI22xp5_ASAP7_75t_L g130 ( .A1(n_63), .A2(n_102), .B1(n_131), .B2(n_132), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g132 ( .A(n_63), .Y(n_132) );
INVx1_ASAP7_75t_SL g562 ( .A(n_64), .Y(n_562) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_65), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_66), .B(n_190), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_67), .B(n_262), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_68), .B(n_191), .Y(n_236) );
INVx1_ASAP7_75t_L g552 ( .A(n_69), .Y(n_552) );
CKINVDCx16_ASAP7_75t_R g272 ( .A(n_70), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_71), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g184 ( .A1(n_72), .A2(n_154), .B(n_185), .C(n_194), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g257 ( .A(n_73), .Y(n_257) );
INVx1_ASAP7_75t_L g114 ( .A(n_74), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_75), .A2(n_146), .B(n_497), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_76), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_77), .A2(n_146), .B(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_78), .A2(n_145), .B(n_486), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g471 ( .A(n_79), .Y(n_471) );
INVx1_ASAP7_75t_L g518 ( .A(n_80), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_81), .B(n_162), .Y(n_161) );
CKINVDCx20_ASAP7_75t_R g211 ( .A(n_82), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_83), .A2(n_146), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g521 ( .A(n_84), .Y(n_521) );
INVx2_ASAP7_75t_L g169 ( .A(n_85), .Y(n_169) );
INVx1_ASAP7_75t_L g535 ( .A(n_86), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g198 ( .A(n_87), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_88), .B(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g111 ( .A(n_89), .Y(n_111) );
OR2x2_ASAP7_75t_L g122 ( .A(n_89), .B(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g463 ( .A(n_89), .B(n_124), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g129 ( .A1(n_90), .A2(n_130), .B1(n_133), .B2(n_134), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_90), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_91), .A2(n_154), .B(n_194), .C(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_92), .B(n_146), .Y(n_201) );
INVx1_ASAP7_75t_L g206 ( .A(n_93), .Y(n_206) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_94), .A2(n_104), .B1(n_115), .B2(n_760), .Y(n_103) );
INVxp67_ASAP7_75t_L g260 ( .A(n_95), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_96), .B(n_181), .Y(n_503) );
INVx2_ASAP7_75t_L g511 ( .A(n_97), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_98), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g186 ( .A(n_99), .Y(n_186) );
INVx1_ASAP7_75t_L g232 ( .A(n_100), .Y(n_232) );
AND2x2_ASAP7_75t_L g250 ( .A(n_101), .B(n_168), .Y(n_250) );
CKINVDCx20_ASAP7_75t_R g131 ( .A(n_102), .Y(n_131) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx12_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g761 ( .A(n_107), .Y(n_761) );
OR2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
OR2x2_ASAP7_75t_L g739 ( .A(n_111), .B(n_124), .Y(n_739) );
NOR2x2_ASAP7_75t_L g747 ( .A(n_111), .B(n_123), .Y(n_747) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AOI22x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_128), .B1(n_748), .B2(n_750), .Y(n_115) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_120), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g749 ( .A(n_119), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_120), .A2(n_751), .B(n_759), .Y(n_750) );
NOR2xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_127), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
BUFx2_ASAP7_75t_L g759 ( .A(n_122), .Y(n_759) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_126), .Y(n_124) );
INVx1_ASAP7_75t_L g740 ( .A(n_129), .Y(n_740) );
INVx1_ASAP7_75t_L g133 ( .A(n_130), .Y(n_133) );
OAI22xp5_ASAP7_75t_SL g135 ( .A1(n_136), .A2(n_461), .B1(n_464), .B2(n_737), .Y(n_135) );
OAI22xp5_ASAP7_75t_SL g751 ( .A1(n_136), .A2(n_743), .B1(n_752), .B2(n_753), .Y(n_751) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx2_ASAP7_75t_L g743 ( .A(n_137), .Y(n_743) );
AND3x1_ASAP7_75t_L g137 ( .A(n_138), .B(n_365), .C(n_422), .Y(n_137) );
NOR3xp33_ASAP7_75t_L g138 ( .A(n_139), .B(n_310), .C(n_346), .Y(n_138) );
OAI211xp5_ASAP7_75t_L g139 ( .A1(n_140), .A2(n_212), .B(n_264), .C(n_297), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_176), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g267 ( .A(n_142), .B(n_268), .Y(n_267) );
INVx5_ASAP7_75t_L g296 ( .A(n_142), .Y(n_296) );
AND2x2_ASAP7_75t_L g369 ( .A(n_142), .B(n_285), .Y(n_369) );
AND2x2_ASAP7_75t_L g407 ( .A(n_142), .B(n_313), .Y(n_407) );
AND2x2_ASAP7_75t_L g427 ( .A(n_142), .B(n_269), .Y(n_427) );
OR2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_173), .Y(n_142) );
AOI21xp5_ASAP7_75t_SL g143 ( .A1(n_144), .A2(n_153), .B(n_166), .Y(n_143) );
BUFx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_147), .B(n_151), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_147), .B(n_151), .Y(n_233) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
INVx1_ASAP7_75t_L g164 ( .A(n_148), .Y(n_164) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g155 ( .A(n_149), .Y(n_155) );
INVx1_ASAP7_75t_L g227 ( .A(n_149), .Y(n_227) );
INVx1_ASAP7_75t_L g156 ( .A(n_150), .Y(n_156) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_150), .Y(n_160) );
INVx3_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
INVx1_ASAP7_75t_L g223 ( .A(n_150), .Y(n_223) );
BUFx6f_ASAP7_75t_L g238 ( .A(n_150), .Y(n_238) );
BUFx3_ASAP7_75t_L g165 ( .A(n_151), .Y(n_165) );
INVx4_ASAP7_75t_SL g195 ( .A(n_151), .Y(n_195) );
INVx5_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_155), .Y(n_193) );
BUFx3_ASAP7_75t_L g209 ( .A(n_155), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_161), .B(n_163), .Y(n_157) );
INVx2_ASAP7_75t_L g162 ( .A(n_159), .Y(n_162) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx4_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g205 ( .A1(n_162), .A2(n_206), .B(n_207), .C(n_208), .Y(n_205) );
O2A1O1Ixp33_ASAP7_75t_L g247 ( .A1(n_162), .A2(n_208), .B(n_248), .C(n_249), .Y(n_247) );
O2A1O1Ixp5_ASAP7_75t_L g534 ( .A1(n_162), .A2(n_535), .B(n_536), .C(n_537), .Y(n_534) );
O2A1O1Ixp33_ASAP7_75t_L g551 ( .A1(n_162), .A2(n_537), .B(n_552), .C(n_553), .Y(n_551) );
O2A1O1Ixp33_ASAP7_75t_L g473 ( .A1(n_163), .A2(n_190), .B(n_474), .C(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g488 ( .A(n_164), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_167), .B(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g175 ( .A(n_168), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_168), .A2(n_201), .B(n_202), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_168), .A2(n_245), .B(n_246), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g470 ( .A1(n_168), .A2(n_233), .B(n_471), .C(n_472), .Y(n_470) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_168), .A2(n_496), .B(n_503), .Y(n_495) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_169), .B(n_170), .Y(n_168) );
AND2x2_ASAP7_75t_L g182 ( .A(n_169), .B(n_170), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_172), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g173 ( .A(n_174), .B(n_175), .Y(n_173) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_175), .A2(n_531), .B(n_538), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_176), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g176 ( .A(n_177), .B(n_199), .Y(n_176) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_177), .Y(n_308) );
AND2x2_ASAP7_75t_L g322 ( .A(n_177), .B(n_268), .Y(n_322) );
INVx1_ASAP7_75t_L g345 ( .A(n_177), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_177), .B(n_296), .Y(n_384) );
OR2x2_ASAP7_75t_L g421 ( .A(n_177), .B(n_266), .Y(n_421) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_178), .Y(n_357) );
AND2x2_ASAP7_75t_L g364 ( .A(n_178), .B(n_269), .Y(n_364) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g285 ( .A(n_179), .B(n_269), .Y(n_285) );
BUFx2_ASAP7_75t_L g313 ( .A(n_179), .Y(n_313) );
AO21x2_ASAP7_75t_L g179 ( .A1(n_180), .A2(n_183), .B(n_197), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_180), .B(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_180), .B(n_211), .Y(n_210) );
AO21x2_ASAP7_75t_L g230 ( .A1(n_180), .A2(n_231), .B(n_239), .Y(n_230) );
INVx3_ASAP7_75t_L g262 ( .A(n_180), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_180), .B(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_180), .B(n_539), .Y(n_538) );
AO21x2_ASAP7_75t_L g547 ( .A1(n_180), .A2(n_548), .B(n_554), .Y(n_547) );
INVx4_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g218 ( .A1(n_181), .A2(n_219), .B(n_220), .Y(n_218) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_181), .Y(n_254) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g241 ( .A(n_182), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_196), .Y(n_183) );
O2A1O1Ixp33_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_189), .C(n_192), .Y(n_185) );
INVx1_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_188), .A2(n_190), .B1(n_490), .B2(n_491), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_188), .B(n_511), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_188), .B(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_190), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g274 ( .A(n_190), .Y(n_274) );
INVx5_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_191), .B(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx3_ASAP7_75t_L g563 ( .A(n_193), .Y(n_563) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
O2A1O1Ixp33_ASAP7_75t_L g256 ( .A1(n_195), .A2(n_204), .B(n_257), .C(n_258), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g271 ( .A1(n_195), .A2(n_204), .B(n_272), .C(n_273), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_SL g486 ( .A1(n_195), .A2(n_204), .B(n_487), .C(n_488), .Y(n_486) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_195), .A2(n_204), .B(n_498), .C(n_499), .Y(n_497) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_195), .A2(n_204), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g517 ( .A1(n_195), .A2(n_204), .B(n_518), .C(n_519), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g558 ( .A1(n_195), .A2(n_204), .B(n_559), .C(n_560), .Y(n_558) );
INVx5_ASAP7_75t_L g266 ( .A(n_199), .Y(n_266) );
BUFx2_ASAP7_75t_L g289 ( .A(n_199), .Y(n_289) );
AND2x2_ASAP7_75t_L g446 ( .A(n_199), .B(n_300), .Y(n_446) );
OR2x6_ASAP7_75t_L g199 ( .A(n_200), .B(n_210), .Y(n_199) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx2_ASAP7_75t_L g278 ( .A(n_209), .Y(n_278) );
INVx1_ASAP7_75t_L g522 ( .A(n_209), .Y(n_522) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NAND2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_251), .Y(n_213) );
OAI221xp5_ASAP7_75t_L g346 ( .A1(n_214), .A2(n_347), .B1(n_354), .B2(n_355), .C(n_358), .Y(n_346) );
OR2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_228), .Y(n_214) );
AND2x2_ASAP7_75t_L g252 ( .A(n_215), .B(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_215), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g281 ( .A(n_216), .B(n_229), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_216), .B(n_230), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_216), .B(n_253), .Y(n_302) );
AND2x2_ASAP7_75t_L g305 ( .A(n_216), .B(n_293), .Y(n_305) );
AND2x2_ASAP7_75t_L g321 ( .A(n_216), .B(n_242), .Y(n_321) );
OR2x2_ASAP7_75t_L g337 ( .A(n_216), .B(n_230), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_216), .B(n_253), .Y(n_399) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_217), .B(n_242), .Y(n_391) );
AND2x2_ASAP7_75t_L g394 ( .A(n_217), .B(n_230), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B(n_225), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_225), .A2(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
OR2x2_ASAP7_75t_L g315 ( .A(n_228), .B(n_302), .Y(n_315) );
INVx2_ASAP7_75t_L g341 ( .A(n_228), .Y(n_341) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_242), .Y(n_228) );
AND2x2_ASAP7_75t_L g263 ( .A(n_229), .B(n_243), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_229), .B(n_253), .Y(n_320) );
OR2x2_ASAP7_75t_L g331 ( .A(n_229), .B(n_243), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_229), .B(n_293), .Y(n_390) );
OAI221xp5_ASAP7_75t_L g423 ( .A1(n_229), .A2(n_424), .B1(n_426), .B2(n_428), .C(n_431), .Y(n_423) );
INVx5_ASAP7_75t_SL g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_230), .B(n_253), .Y(n_362) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
OAI21xp5_ASAP7_75t_L g531 ( .A1(n_233), .A2(n_532), .B(n_533), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g548 ( .A1(n_233), .A2(n_549), .B(n_550), .Y(n_548) );
INVx4_ASAP7_75t_L g277 ( .A(n_238), .Y(n_277) );
INVx2_ASAP7_75t_L g500 ( .A(n_238), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_L g483 ( .A(n_241), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_242), .B(n_293), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_242), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_242), .B(n_281), .Y(n_309) );
OR2x2_ASAP7_75t_L g353 ( .A(n_242), .B(n_253), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_242), .B(n_305), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_242), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g418 ( .A(n_242), .B(n_419), .Y(n_418) );
INVx5_ASAP7_75t_SL g242 ( .A(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_SL g282 ( .A(n_243), .B(n_252), .Y(n_282) );
O2A1O1Ixp33_ASAP7_75t_SL g286 ( .A1(n_243), .A2(n_287), .B(n_290), .C(n_294), .Y(n_286) );
OR2x2_ASAP7_75t_L g324 ( .A(n_243), .B(n_320), .Y(n_324) );
OR2x2_ASAP7_75t_L g360 ( .A(n_243), .B(n_302), .Y(n_360) );
OAI311xp33_ASAP7_75t_L g366 ( .A1(n_243), .A2(n_305), .A3(n_367), .B1(n_370), .C1(n_377), .Y(n_366) );
AND2x2_ASAP7_75t_L g417 ( .A(n_243), .B(n_253), .Y(n_417) );
AND2x2_ASAP7_75t_L g425 ( .A(n_243), .B(n_280), .Y(n_425) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_243), .Y(n_443) );
AND2x2_ASAP7_75t_L g460 ( .A(n_243), .B(n_281), .Y(n_460) );
OR2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_250), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_263), .Y(n_251) );
AND2x2_ASAP7_75t_L g288 ( .A(n_252), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g444 ( .A(n_252), .Y(n_444) );
AND2x2_ASAP7_75t_L g280 ( .A(n_253), .B(n_281), .Y(n_280) );
INVx3_ASAP7_75t_L g293 ( .A(n_253), .Y(n_293) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_253), .Y(n_336) );
INVxp67_ASAP7_75t_L g375 ( .A(n_253), .Y(n_375) );
OA21x2_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_255), .B(n_261), .Y(n_253) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_254), .A2(n_506), .B(n_512), .Y(n_505) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_254), .A2(n_516), .B(n_523), .Y(n_515) );
OA21x2_ASAP7_75t_L g556 ( .A1(n_254), .A2(n_557), .B(n_564), .Y(n_556) );
OA21x2_ASAP7_75t_L g269 ( .A1(n_262), .A2(n_270), .B(n_279), .Y(n_269) );
AND2x2_ASAP7_75t_L g453 ( .A(n_263), .B(n_301), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_280), .B1(n_282), .B2(n_283), .C(n_286), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_266), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g306 ( .A(n_266), .B(n_296), .Y(n_306) );
AND2x2_ASAP7_75t_L g314 ( .A(n_266), .B(n_268), .Y(n_314) );
OR2x2_ASAP7_75t_L g326 ( .A(n_266), .B(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g344 ( .A(n_266), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g368 ( .A(n_266), .B(n_369), .Y(n_368) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_266), .Y(n_388) );
AND2x2_ASAP7_75t_L g440 ( .A(n_266), .B(n_364), .Y(n_440) );
OAI31xp33_ASAP7_75t_L g448 ( .A1(n_266), .A2(n_317), .A3(n_416), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_267), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g412 ( .A(n_267), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_267), .B(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g300 ( .A(n_268), .B(n_296), .Y(n_300) );
INVx1_ASAP7_75t_L g387 ( .A(n_268), .Y(n_387) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g437 ( .A(n_269), .B(n_296), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_277), .B(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g537 ( .A(n_278), .Y(n_537) );
INVx1_ASAP7_75t_SL g447 ( .A(n_280), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_281), .B(n_352), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_282), .A2(n_394), .B1(n_432), .B2(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g295 ( .A(n_285), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g354 ( .A(n_285), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_285), .B(n_306), .Y(n_459) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g429 ( .A(n_288), .B(n_430), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_289), .A2(n_348), .B(n_350), .Y(n_347) );
OR2x2_ASAP7_75t_L g355 ( .A(n_289), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g376 ( .A(n_289), .B(n_364), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_289), .B(n_387), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_289), .B(n_427), .Y(n_426) );
OAI221xp5_ASAP7_75t_SL g403 ( .A1(n_290), .A2(n_404), .B1(n_409), .B2(n_412), .C(n_413), .Y(n_403) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
OR2x2_ASAP7_75t_L g380 ( .A(n_291), .B(n_353), .Y(n_380) );
INVx1_ASAP7_75t_L g419 ( .A(n_291), .Y(n_419) );
INVx2_ASAP7_75t_L g395 ( .A(n_292), .Y(n_395) );
INVx1_ASAP7_75t_L g329 ( .A(n_293), .Y(n_329) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
INVx2_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_296), .B(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g363 ( .A(n_296), .B(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g451 ( .A(n_296), .B(n_421), .Y(n_451) );
AOI222xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_301), .B1(n_303), .B2(n_306), .C1(n_307), .C2(n_309), .Y(n_297) );
INVxp67_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g307 ( .A(n_300), .B(n_308), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_300), .A2(n_350), .B1(n_378), .B2(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_300), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
OAI21xp33_ASAP7_75t_SL g338 ( .A1(n_309), .A2(n_339), .B(n_342), .Y(n_338) );
OAI211xp5_ASAP7_75t_SL g310 ( .A1(n_311), .A2(n_315), .B(n_316), .C(n_338), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_314), .A2(n_317), .B1(n_322), .B2(n_323), .C(n_325), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_314), .B(n_402), .Y(n_401) );
INVxp67_ASAP7_75t_L g408 ( .A(n_314), .Y(n_408) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
AND2x2_ASAP7_75t_L g410 ( .A(n_319), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g327 ( .A(n_322), .Y(n_327) );
AND2x2_ASAP7_75t_L g333 ( .A(n_322), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_328), .B1(n_332), .B2(n_335), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_329), .B(n_341), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_330), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g430 ( .A(n_334), .Y(n_430) );
AND2x2_ASAP7_75t_L g449 ( .A(n_334), .B(n_364), .Y(n_449) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_341), .B(n_398), .Y(n_457) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_344), .B(n_412), .Y(n_455) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g378 ( .A(n_356), .Y(n_378) );
BUFx2_ASAP7_75t_L g402 ( .A(n_357), .Y(n_402) );
OAI21xp5_ASAP7_75t_SL g358 ( .A1(n_359), .A2(n_361), .B(n_363), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
NOR3xp33_ASAP7_75t_L g365 ( .A(n_366), .B(n_381), .C(n_403), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B(n_376), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_SL g381 ( .A1(n_382), .A2(n_385), .B(n_389), .C(n_392), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g414 ( .A(n_382), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp67_ASAP7_75t_SL g386 ( .A(n_387), .B(n_388), .Y(n_386) );
OR2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
INVx1_ASAP7_75t_SL g411 ( .A(n_391), .Y(n_411) );
OAI21xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B(n_400), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
AND2x2_ASAP7_75t_L g416 ( .A(n_394), .B(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_408), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_418), .B2(n_420), .Y(n_413) );
INVx2_ASAP7_75t_SL g434 ( .A(n_421), .Y(n_434) );
NOR3xp33_ASAP7_75t_L g422 ( .A(n_423), .B(n_438), .C(n_450), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_434), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI221xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_441), .B1(n_445), .B2(n_447), .C(n_448), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_439), .A2(n_451), .B(n_452), .C(n_454), .Y(n_450) );
INVx1_ASAP7_75t_SL g439 ( .A(n_440), .Y(n_439) );
INVxp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_456), .B1(n_458), .B2(n_460), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g742 ( .A(n_462), .Y(n_742) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g744 ( .A(n_464), .Y(n_744) );
OR5x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_631), .C(n_695), .D(n_711), .E(n_726), .Y(n_464) );
NAND4xp25_ASAP7_75t_L g465 ( .A(n_466), .B(n_565), .C(n_592), .D(n_615), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_513), .B(n_524), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_478), .Y(n_467) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx3_ASAP7_75t_SL g544 ( .A(n_469), .Y(n_544) );
AND2x4_ASAP7_75t_L g578 ( .A(n_469), .B(n_567), .Y(n_578) );
OR2x2_ASAP7_75t_L g588 ( .A(n_469), .B(n_546), .Y(n_588) );
OR2x2_ASAP7_75t_L g634 ( .A(n_469), .B(n_481), .Y(n_634) );
AND2x2_ASAP7_75t_L g648 ( .A(n_469), .B(n_545), .Y(n_648) );
AND2x2_ASAP7_75t_L g691 ( .A(n_469), .B(n_581), .Y(n_691) );
AND2x2_ASAP7_75t_L g698 ( .A(n_469), .B(n_556), .Y(n_698) );
AND2x2_ASAP7_75t_L g717 ( .A(n_469), .B(n_607), .Y(n_717) );
AND2x2_ASAP7_75t_L g735 ( .A(n_469), .B(n_577), .Y(n_735) );
OR2x6_ASAP7_75t_L g469 ( .A(n_470), .B(n_476), .Y(n_469) );
INVx1_ASAP7_75t_L g700 ( .A(n_478), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_494), .Y(n_478) );
AND2x2_ASAP7_75t_L g610 ( .A(n_479), .B(n_545), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_479), .B(n_630), .Y(n_629) );
AOI32xp33_ASAP7_75t_L g643 ( .A1(n_479), .A2(n_644), .A3(n_647), .B1(n_649), .B2(n_653), .Y(n_643) );
AND2x2_ASAP7_75t_L g713 ( .A(n_479), .B(n_607), .Y(n_713) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g577 ( .A(n_481), .B(n_546), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_481), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g619 ( .A(n_481), .B(n_566), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_481), .B(n_698), .Y(n_697) );
AO21x2_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_484), .B(n_492), .Y(n_481) );
INVx1_ASAP7_75t_L g582 ( .A(n_482), .Y(n_582) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OA21x2_ASAP7_75t_L g581 ( .A1(n_485), .A2(n_493), .B(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g584 ( .A(n_494), .B(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g660 ( .A(n_494), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g732 ( .A(n_494), .Y(n_732) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
OR2x2_ASAP7_75t_L g527 ( .A(n_495), .B(n_505), .Y(n_527) );
AND2x2_ASAP7_75t_L g541 ( .A(n_495), .B(n_542), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_495), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g591 ( .A(n_495), .Y(n_591) );
AND2x2_ASAP7_75t_L g618 ( .A(n_495), .B(n_505), .Y(n_618) );
BUFx3_ASAP7_75t_L g621 ( .A(n_495), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_495), .B(n_596), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_495), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
AND2x2_ASAP7_75t_L g590 ( .A(n_504), .B(n_570), .Y(n_590) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x2_ASAP7_75t_L g601 ( .A(n_505), .B(n_515), .Y(n_601) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_505), .Y(n_614) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_514), .B(n_621), .Y(n_671) );
HB1xp67_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_SL g542 ( .A(n_515), .Y(n_542) );
NAND3xp33_ASAP7_75t_L g589 ( .A(n_515), .B(n_590), .C(n_591), .Y(n_589) );
OR2x2_ASAP7_75t_L g597 ( .A(n_515), .B(n_570), .Y(n_597) );
AND2x2_ASAP7_75t_L g617 ( .A(n_515), .B(n_570), .Y(n_617) );
AND2x2_ASAP7_75t_L g661 ( .A(n_515), .B(n_530), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_540), .B(n_543), .Y(n_524) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_526), .B(n_528), .Y(n_525) );
AND2x2_ASAP7_75t_L g736 ( .A(n_526), .B(n_661), .Y(n_736) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_527), .A2(n_634), .B1(n_676), .B2(n_678), .Y(n_675) );
OR2x2_ASAP7_75t_L g682 ( .A(n_527), .B(n_597), .Y(n_682) );
OR2x2_ASAP7_75t_L g706 ( .A(n_527), .B(n_707), .Y(n_706) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_527), .B(n_626), .Y(n_719) );
AND2x2_ASAP7_75t_L g612 ( .A(n_528), .B(n_613), .Y(n_612) );
AOI21xp5_ASAP7_75t_L g699 ( .A1(n_528), .A2(n_685), .B(n_700), .Y(n_699) );
AOI32xp33_ASAP7_75t_L g720 ( .A1(n_528), .A2(n_610), .A3(n_721), .B1(n_723), .B2(n_724), .Y(n_720) );
OR2x2_ASAP7_75t_L g731 ( .A(n_528), .B(n_732), .Y(n_731) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g599 ( .A(n_529), .B(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_529), .B(n_613), .Y(n_678) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g570 ( .A(n_530), .Y(n_570) );
AND2x2_ASAP7_75t_L g636 ( .A(n_530), .B(n_601), .Y(n_636) );
AND3x2_ASAP7_75t_L g645 ( .A(n_530), .B(n_541), .C(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g571 ( .A(n_542), .B(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_542), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_542), .B(n_570), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x2_ASAP7_75t_L g566 ( .A(n_544), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g606 ( .A(n_544), .B(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g624 ( .A(n_544), .B(n_556), .Y(n_624) );
AND2x2_ASAP7_75t_L g642 ( .A(n_544), .B(n_546), .Y(n_642) );
OR2x2_ASAP7_75t_L g656 ( .A(n_544), .B(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g702 ( .A(n_544), .B(n_630), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_545), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_556), .Y(n_545) );
AND2x2_ASAP7_75t_L g603 ( .A(n_546), .B(n_581), .Y(n_603) );
OR2x2_ASAP7_75t_L g657 ( .A(n_546), .B(n_581), .Y(n_657) );
AND2x2_ASAP7_75t_L g710 ( .A(n_546), .B(n_567), .Y(n_710) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g608 ( .A(n_547), .Y(n_608) );
AND2x2_ASAP7_75t_L g630 ( .A(n_547), .B(n_556), .Y(n_630) );
INVx2_ASAP7_75t_L g567 ( .A(n_556), .Y(n_567) );
INVx1_ASAP7_75t_L g587 ( .A(n_556), .Y(n_587) );
AOI211xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B(n_573), .C(n_585), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_566), .B(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g729 ( .A(n_566), .Y(n_729) );
AND2x2_ASAP7_75t_L g607 ( .A(n_567), .B(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_570), .B(n_571), .Y(n_579) );
INVx1_ASAP7_75t_L g664 ( .A(n_570), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_570), .B(n_591), .Y(n_688) );
AND2x2_ASAP7_75t_L g704 ( .A(n_570), .B(n_618), .Y(n_704) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_571), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g595 ( .A(n_572), .Y(n_595) );
OAI22xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_579), .B1(n_580), .B2(n_583), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_576), .B(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_577), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g602 ( .A(n_578), .B(n_603), .Y(n_602) );
AOI221xp5_ASAP7_75t_SL g667 ( .A1(n_578), .A2(n_620), .B1(n_668), .B2(n_673), .C(n_675), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_578), .B(n_641), .Y(n_674) );
INVx1_ASAP7_75t_L g734 ( .A(n_580), .Y(n_734) );
BUFx3_ASAP7_75t_L g641 ( .A(n_581), .Y(n_641) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AOI21xp33_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_588), .B(n_589), .Y(n_585) );
INVx1_ASAP7_75t_L g650 ( .A(n_587), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_587), .B(n_641), .Y(n_694) );
INVx1_ASAP7_75t_L g651 ( .A(n_588), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g652 ( .A(n_588), .B(n_641), .Y(n_652) );
INVxp67_ASAP7_75t_L g672 ( .A(n_590), .Y(n_672) );
AND2x2_ASAP7_75t_L g613 ( .A(n_591), .B(n_614), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_598), .B(n_602), .C(n_604), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVx1_ASAP7_75t_SL g627 ( .A(n_595), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_596), .B(n_627), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_596), .B(n_618), .Y(n_669) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_599), .A2(n_605), .B1(n_609), .B2(n_611), .Y(n_604) );
INVx1_ASAP7_75t_SL g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g620 ( .A(n_601), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g665 ( .A(n_601), .B(n_666), .Y(n_665) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_603), .A2(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_607), .A2(n_616), .B1(n_619), .B2(n_620), .C(n_622), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_607), .B(n_641), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_607), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g723 ( .A(n_613), .Y(n_723) );
INVxp67_ASAP7_75t_L g646 ( .A(n_614), .Y(n_646) );
INVx1_ASAP7_75t_L g653 ( .A(n_616), .Y(n_653) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g692 ( .A(n_617), .B(n_621), .Y(n_692) );
INVx1_ASAP7_75t_L g666 ( .A(n_621), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g696 ( .A(n_621), .B(n_636), .Y(n_696) );
OAI32xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_625), .A3(n_627), .B1(n_628), .B2(n_629), .Y(n_622) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_SL g635 ( .A(n_630), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_630), .B(n_662), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_630), .B(n_691), .Y(n_722) );
NAND2x1p5_ASAP7_75t_L g730 ( .A(n_630), .B(n_641), .Y(n_730) );
NAND5xp2_ASAP7_75t_L g631 ( .A(n_632), .B(n_654), .C(n_667), .D(n_679), .E(n_680), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B1(n_637), .B2(n_639), .C(n_643), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp33_ASAP7_75t_SL g658 ( .A(n_638), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_641), .B(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_642), .A2(n_655), .B1(n_658), .B2(n_662), .Y(n_654) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
OAI211xp5_ASAP7_75t_SL g649 ( .A1(n_645), .A2(n_650), .B(n_651), .C(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g677 ( .A(n_657), .Y(n_677) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_SL g662 ( .A(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_666), .B(n_715), .Y(n_725) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_683), .B1(n_685), .B2(n_689), .C1(n_692), .C2(n_693), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OAI221xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_699), .B2(n_701), .C(n_703), .Y(n_695) );
INVx1_ASAP7_75t_SL g701 ( .A(n_702), .Y(n_701) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_704), .A2(n_705), .B(n_708), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g715 ( .A(n_707), .Y(n_715) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B1(n_716), .B2(n_718), .C(n_720), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_SL g716 ( .A(n_717), .Y(n_716) );
INVxp67_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_730), .B(n_731), .C(n_733), .Y(n_726) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI21xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_736), .Y(n_733) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_739), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx2_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
endmodule