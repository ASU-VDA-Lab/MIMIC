module fake_jpeg_16539_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_26),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_30),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_37),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_21),
.B1(n_29),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_46),
.A2(n_49),
.B1(n_62),
.B2(n_68),
.Y(n_88)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_48),
.B(n_35),
.CON(n_81),
.SN(n_81)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_21),
.B1(n_29),
.B2(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_54),
.Y(n_102)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_35),
.A2(n_21),
.B1(n_31),
.B2(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_43),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_22),
.B1(n_24),
.B2(n_42),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_69),
.A2(n_98),
.B1(n_99),
.B2(n_20),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_71),
.B(n_76),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_45),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_72),
.B(n_74),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_77),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_45),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_45),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_53),
.B(n_56),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_SL g119 ( 
.A(n_81),
.B(n_82),
.C(n_87),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_65),
.A2(n_37),
.B(n_18),
.C(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_84),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_17),
.B(n_25),
.C(n_33),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_30),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_89),
.Y(n_127)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_90),
.Y(n_121)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_61),
.A2(n_17),
.B1(n_25),
.B2(n_28),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_40),
.Y(n_93)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_32),
.B1(n_41),
.B2(n_39),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_52),
.A2(n_32),
.B1(n_20),
.B2(n_30),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_55),
.A2(n_32),
.B1(n_20),
.B2(n_34),
.Y(n_99)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_107),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_104),
.A2(n_115),
.B1(n_101),
.B2(n_91),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_41),
.B(n_44),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_109),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_97),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_128),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_114),
.B(n_123),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g122 ( 
.A1(n_81),
.A2(n_40),
.B1(n_60),
.B2(n_50),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_85),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_90),
.Y(n_130)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_78),
.B1(n_80),
.B2(n_44),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_76),
.B(n_74),
.C(n_72),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_145),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_71),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_133),
.A2(n_144),
.B(n_34),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_88),
.B1(n_93),
.B2(n_95),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_134),
.A2(n_158),
.B1(n_163),
.B2(n_20),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_137),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_111),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_83),
.B1(n_100),
.B2(n_94),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_151),
.B1(n_36),
.B2(n_34),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_111),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_139),
.B(n_146),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_82),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_142),
.C(n_153),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_125),
.A2(n_83),
.B1(n_100),
.B2(n_80),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_141),
.A2(n_113),
.B1(n_104),
.B2(n_117),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_102),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_116),
.A2(n_87),
.A3(n_73),
.B1(n_79),
.B2(n_39),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_121),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_106),
.A2(n_116),
.B1(n_119),
.B2(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_40),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_155),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_40),
.C(n_36),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_106),
.B(n_19),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_121),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_130),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_78),
.B1(n_12),
.B2(n_13),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_159),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_131),
.B(n_19),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_161),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_23),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_114),
.A2(n_109),
.B1(n_129),
.B2(n_124),
.Y(n_163)
);

AO22x1_ASAP7_75t_SL g165 ( 
.A1(n_145),
.A2(n_129),
.B1(n_124),
.B2(n_126),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_167),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_168),
.B(n_169),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_113),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_172),
.A2(n_186),
.B1(n_189),
.B2(n_193),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_36),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_178),
.C(n_184),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_117),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_175),
.B(n_194),
.Y(n_218)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_147),
.Y(n_176)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_188),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_151),
.B(n_23),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_181),
.B(n_161),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_135),
.A2(n_16),
.B(n_19),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_140),
.C(n_135),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_143),
.A2(n_139),
.B1(n_137),
.B2(n_157),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_143),
.B(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_134),
.A2(n_23),
.B1(n_16),
.B2(n_3),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_133),
.B(n_23),
.Y(n_187)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_23),
.C(n_16),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_133),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_23),
.Y(n_190)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_138),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_8),
.Y(n_194)
);

OAI21x1_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_144),
.B(n_158),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_15),
.B(n_12),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_197),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_146),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_198),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_176),
.Y(n_199)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_201),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_210),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_173),
.A2(n_171),
.B1(n_165),
.B2(n_192),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_204),
.A2(n_212),
.B1(n_209),
.B2(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_179),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_170),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_191),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_215),
.Y(n_240)
);

NOR2x1_ASAP7_75t_R g212 ( 
.A(n_165),
.B(n_156),
.Y(n_212)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_180),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_164),
.Y(n_215)
);

INVxp67_ASAP7_75t_SL g216 ( 
.A(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_216),
.Y(n_226)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_190),
.B(n_166),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_0),
.Y(n_221)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_221),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_223),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_247),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_207),
.B(n_183),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_230),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_207),
.B(n_183),
.Y(n_230)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_221),
.Y(n_257)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_220),
.B1(n_200),
.B2(n_218),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_184),
.C(n_174),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_246),
.C(n_249),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_173),
.B1(n_166),
.B2(n_178),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_205),
.B1(n_225),
.B2(n_209),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_211),
.B(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_187),
.C(n_188),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_223),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_213),
.B(n_177),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_200),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_181),
.C(n_186),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_250),
.B(n_269),
.Y(n_277)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_201),
.B(n_224),
.C(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_232),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_258),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_233),
.B(n_202),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_204),
.C(n_214),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_262),
.C(n_263),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_214),
.C(n_198),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_199),
.C(n_215),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_264),
.A2(n_226),
.B1(n_235),
.B2(n_241),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_246),
.B(n_199),
.C(n_206),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_268),
.C(n_249),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_10),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_11),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_240),
.Y(n_270)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_244),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_276),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_256),
.B(n_243),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_281),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_252),
.B(n_253),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_241),
.C(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_283),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_248),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_261),
.A2(n_231),
.B(n_267),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_2),
.B(n_4),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_245),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_232),
.C(n_234),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_286),
.A2(n_287),
.B(n_294),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_262),
.B(n_260),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_277),
.A2(n_266),
.B1(n_268),
.B2(n_234),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_258),
.B1(n_257),
.B2(n_251),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_273),
.B1(n_5),
.B2(n_6),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_291),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_285),
.A2(n_9),
.B(n_3),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_295),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_299),
.Y(n_309)
);

XOR2x2_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_4),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_275),
.C(n_276),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_308),
.C(n_294),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_275),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_301),
.B(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_293),
.B(n_273),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_286),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_4),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_307),
.B(n_6),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_5),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_315),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_313),
.B(n_314),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_309),
.A2(n_298),
.B1(n_296),
.B2(n_287),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_304),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_289),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_318),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_299),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_312),
.A2(n_303),
.B(n_308),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_305),
.C(n_319),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_314),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_326),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_311),
.Y(n_328)
);

OAI221xp5_ASAP7_75t_L g329 ( 
.A1(n_328),
.A2(n_322),
.B1(n_321),
.B2(n_300),
.C(n_290),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_6),
.B(n_7),
.Y(n_330)
);


endmodule