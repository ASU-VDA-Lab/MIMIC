module real_aes_5560_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_357;
wire n_287;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_580;
wire n_577;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_547;
wire n_102;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_206;
wire n_307;
wire n_601;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g152 ( .A(n_0), .B(n_89), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_1), .Y(n_104) );
O2A1O1Ixp33_ASAP7_75t_SL g223 ( .A1(n_2), .A2(n_94), .B(n_224), .C(n_225), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g157 ( .A1(n_3), .A2(n_62), .B1(n_100), .B2(n_158), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_4), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g524 ( .A(n_5), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_6), .Y(n_147) );
OAI22xp5_ASAP7_75t_L g202 ( .A1(n_7), .A2(n_54), .B1(n_121), .B2(n_158), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g187 ( .A(n_8), .Y(n_187) );
INVx1_ASAP7_75t_L g479 ( .A(n_9), .Y(n_479) );
INVxp67_ASAP7_75t_L g507 ( .A(n_9), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_9), .B(n_56), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_10), .A2(n_42), .B1(n_552), .B2(n_554), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_11), .A2(n_27), .B1(n_539), .B2(n_547), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_12), .A2(n_47), .B1(n_100), .B2(n_105), .Y(n_201) );
OA21x2_ASAP7_75t_L g91 ( .A1(n_13), .A2(n_53), .B(n_92), .Y(n_91) );
OA21x2_ASAP7_75t_L g136 ( .A1(n_13), .A2(n_53), .B(n_92), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_14), .B(n_464), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g140 ( .A(n_15), .Y(n_140) );
BUFx3_ASAP7_75t_L g587 ( .A(n_16), .Y(n_587) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_17), .A2(n_102), .B(n_230), .C(n_231), .Y(n_229) );
OAI22xp33_ASAP7_75t_SL g155 ( .A1(n_18), .A2(n_33), .B1(n_97), .B2(n_100), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g116 ( .A1(n_19), .A2(n_24), .B1(n_97), .B2(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_20), .Y(n_464) );
O2A1O1Ixp5_ASAP7_75t_L g166 ( .A1(n_21), .A2(n_94), .B(n_167), .C(n_168), .Y(n_166) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_22), .Y(n_442) );
INVx1_ASAP7_75t_L g468 ( .A(n_23), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_23), .B(n_55), .Y(n_504) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_24), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_25), .A2(n_71), .B1(n_498), .B2(n_509), .Y(n_497) );
INVx1_ASAP7_75t_L g489 ( .A(n_26), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_28), .B(n_128), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_29), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_30), .Y(n_227) );
INVx1_ASAP7_75t_L g529 ( .A(n_31), .Y(n_529) );
HB1xp67_ASAP7_75t_L g450 ( .A(n_32), .Y(n_450) );
INVx1_ASAP7_75t_L g92 ( .A(n_34), .Y(n_92) );
AND2x4_ASAP7_75t_L g107 ( .A(n_35), .B(n_108), .Y(n_107) );
AND2x4_ASAP7_75t_L g134 ( .A(n_35), .B(n_108), .Y(n_134) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_35), .Y(n_597) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_36), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_37), .Y(n_101) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_38), .A2(n_94), .B(n_144), .C(n_146), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_39), .Y(n_175) );
INVx2_ASAP7_75t_L g192 ( .A(n_40), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_41), .Y(n_99) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_43), .A2(n_58), .B1(n_571), .B2(n_575), .Y(n_570) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_44), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_45), .B(n_110), .Y(n_109) );
AOI22xp5_ASAP7_75t_L g119 ( .A1(n_46), .A2(n_60), .B1(n_120), .B2(n_122), .Y(n_119) );
HB1xp67_ASAP7_75t_L g445 ( .A(n_48), .Y(n_445) );
OA22x2_ASAP7_75t_L g462 ( .A1(n_49), .A2(n_56), .B1(n_463), .B2(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g522 ( .A(n_49), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_50), .A2(n_67), .B1(n_561), .B2(n_565), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_51), .Y(n_106) );
NAND2xp33_ASAP7_75t_R g205 ( .A(n_52), .B(n_136), .Y(n_205) );
AOI22xp33_ASAP7_75t_L g249 ( .A1(n_52), .A2(n_76), .B1(n_128), .B2(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g481 ( .A(n_55), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_55), .B(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_55), .Y(n_590) );
OAI21xp33_ASAP7_75t_L g535 ( .A1(n_56), .A2(n_61), .B(n_508), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_57), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_59), .Y(n_188) );
INVx1_ASAP7_75t_L g470 ( .A(n_61), .Y(n_470) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_61), .B(n_70), .Y(n_516) );
BUFx6f_ASAP7_75t_L g98 ( .A(n_63), .Y(n_98) );
BUFx5_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g118 ( .A(n_63), .Y(n_118) );
INVx2_ASAP7_75t_L g235 ( .A(n_64), .Y(n_235) );
INVx2_ASAP7_75t_L g149 ( .A(n_65), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_66), .Y(n_232) );
INVx2_ASAP7_75t_SL g108 ( .A(n_68), .Y(n_108) );
INVx1_ASAP7_75t_L g173 ( .A(n_69), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_70), .B(n_474), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_72), .A2(n_452), .B1(n_453), .B2(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_72), .Y(n_607) );
INVx2_ASAP7_75t_L g179 ( .A(n_73), .Y(n_179) );
OAI21xp33_ASAP7_75t_SL g138 ( .A1(n_74), .A2(n_100), .B(n_139), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_75), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_76), .B(n_128), .Y(n_182) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_76), .Y(n_305) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_431), .B1(n_437), .B2(n_582), .C(n_598), .Y(n_77) );
INVxp33_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND3x4_ASAP7_75t_L g79 ( .A(n_80), .B(n_334), .C(n_385), .Y(n_79) );
NOR2x1_ASAP7_75t_L g80 ( .A(n_81), .B(n_279), .Y(n_80) );
NAND3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_252), .C(n_264), .Y(n_81) );
AOI221xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_160), .B1(n_194), .B2(n_219), .C(n_236), .Y(n_82) );
AND2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_129), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_84), .B(n_212), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_84), .B(n_293), .Y(n_329) );
AND2x2_ASAP7_75t_L g388 ( .A(n_84), .B(n_268), .Y(n_388) );
INVx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g253 ( .A(n_85), .Y(n_253) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_112), .Y(n_85) );
AND2x2_ASAP7_75t_L g213 ( .A(n_86), .B(n_214), .Y(n_213) );
AND2x4_ASAP7_75t_L g283 ( .A(n_86), .B(n_269), .Y(n_283) );
AND2x2_ASAP7_75t_L g318 ( .A(n_86), .B(n_151), .Y(n_318) );
AND2x2_ASAP7_75t_L g346 ( .A(n_86), .B(n_347), .Y(n_346) );
OA21x2_ASAP7_75t_L g86 ( .A1(n_87), .A2(n_93), .B(n_109), .Y(n_86) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_87), .A2(n_93), .B(n_109), .Y(n_210) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
OR2x2_ASAP7_75t_L g304 ( .A(n_88), .B(n_305), .Y(n_304) );
INVx2_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
NOR2xp33_ASAP7_75t_SL g233 ( .A(n_89), .B(n_176), .Y(n_233) );
INVx2_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g128 ( .A(n_90), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_90), .B(n_107), .Y(n_159) );
NOR2xp33_ASAP7_75t_SL g234 ( .A(n_90), .B(n_235), .Y(n_234) );
INVx4_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
BUFx3_ASAP7_75t_L g125 ( .A(n_91), .Y(n_125) );
OAI221xp5_ASAP7_75t_L g93 ( .A1(n_94), .A2(n_96), .B1(n_102), .B2(n_103), .C(n_107), .Y(n_93) );
INVx1_ASAP7_75t_L g193 ( .A(n_94), .Y(n_193) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_94), .A2(n_142), .B1(n_201), .B2(n_202), .Y(n_200) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_94), .A2(n_142), .B1(n_186), .B2(n_190), .Y(n_303) );
BUFx6f_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx3_ASAP7_75t_L g102 ( .A(n_95), .Y(n_102) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_95), .Y(n_115) );
INVx1_ASAP7_75t_L g123 ( .A(n_95), .Y(n_123) );
INVx4_ASAP7_75t_L g142 ( .A(n_95), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_95), .B(n_155), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_95), .B(n_173), .Y(n_172) );
AOI22xp33_ASAP7_75t_SL g96 ( .A1(n_97), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_96) );
INVx2_ASAP7_75t_SL g122 ( .A(n_97), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_97), .A2(n_100), .B1(n_187), .B2(n_188), .Y(n_186) );
INVx2_ASAP7_75t_L g226 ( .A(n_97), .Y(n_226) );
INVx6_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
INVx2_ASAP7_75t_L g105 ( .A(n_98), .Y(n_105) );
INVx3_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
INVx2_ASAP7_75t_L g158 ( .A(n_98), .Y(n_158) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_100), .A2(n_104), .B1(n_105), .B2(n_106), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_100), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_100), .B(n_169), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_100), .B(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g600 ( .A(n_101), .Y(n_600) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_102), .A2(n_157), .B(n_159), .Y(n_156) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_104), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g190 ( .A1(n_105), .A2(n_117), .B1(n_191), .B2(n_192), .Y(n_190) );
INVx1_ASAP7_75t_L g230 ( .A(n_105), .Y(n_230) );
INVx1_ASAP7_75t_L g204 ( .A(n_107), .Y(n_204) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_107), .Y(n_302) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_108), .Y(n_595) );
NOR2xp67_ASAP7_75t_L g203 ( .A(n_110), .B(n_204), .Y(n_203) );
INVx3_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_111), .B(n_149), .Y(n_148) );
BUFx3_ASAP7_75t_L g177 ( .A(n_111), .Y(n_177) );
AND2x4_ASAP7_75t_L g313 ( .A(n_112), .B(n_209), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_124), .B(n_126), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_114), .A2(n_127), .B(n_216), .Y(n_215) );
OA22x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_116), .B1(n_119), .B2(n_123), .Y(n_114) );
INVx4_ASAP7_75t_L g435 ( .A(n_115), .Y(n_435) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_117), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_117), .B(n_232), .Y(n_231) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g121 ( .A(n_118), .Y(n_121) );
INVx1_ASAP7_75t_L g224 ( .A(n_120), .Y(n_224) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_150), .Y(n_130) );
BUFx2_ASAP7_75t_L g207 ( .A(n_131), .Y(n_207) );
AND2x2_ASAP7_75t_L g212 ( .A(n_131), .B(n_151), .Y(n_212) );
INVx2_ASAP7_75t_L g240 ( .A(n_131), .Y(n_240) );
AND2x2_ASAP7_75t_L g257 ( .A(n_131), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g273 ( .A(n_131), .B(n_269), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_131), .B(n_210), .Y(n_333) );
INVx1_ASAP7_75t_L g339 ( .A(n_131), .Y(n_339) );
INVx2_ASAP7_75t_L g358 ( .A(n_131), .Y(n_358) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AOI21x1_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_137), .B(n_148), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_135), .Y(n_133) );
INVx4_ASAP7_75t_L g176 ( .A(n_134), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_134), .B(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
BUFx3_ASAP7_75t_L g218 ( .A(n_136), .Y(n_218) );
INVx2_ASAP7_75t_L g251 ( .A(n_136), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_141), .B(n_143), .Y(n_137) );
AOI221xp5_ASAP7_75t_L g184 ( .A1(n_141), .A2(n_176), .B1(n_185), .B2(n_189), .C(n_193), .Y(n_184) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g170 ( .A1(n_142), .A2(n_171), .B1(n_172), .B2(n_174), .Y(n_170) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g167 ( .A(n_145), .Y(n_167) );
INVx1_ASAP7_75t_L g171 ( .A(n_145), .Y(n_171) );
AND2x4_ASAP7_75t_L g208 ( .A(n_150), .B(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g409 ( .A(n_150), .B(n_214), .Y(n_409) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g256 ( .A(n_151), .Y(n_256) );
INVx3_ASAP7_75t_L g269 ( .A(n_151), .Y(n_269) );
AND2x4_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_154), .B(n_156), .Y(n_153) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_181), .Y(n_162) );
AND2x4_ASAP7_75t_L g196 ( .A(n_163), .B(n_197), .Y(n_196) );
OR2x2_ASAP7_75t_L g425 ( .A(n_163), .B(n_358), .Y(n_425) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g246 ( .A(n_164), .Y(n_246) );
AND2x2_ASAP7_75t_L g260 ( .A(n_164), .B(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_164), .B(n_221), .Y(n_298) );
BUFx2_ASAP7_75t_R g308 ( .A(n_164), .Y(n_308) );
AND2x2_ASAP7_75t_L g384 ( .A(n_164), .B(n_364), .Y(n_384) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_164), .Y(n_392) );
AO21x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_177), .B(n_178), .Y(n_164) );
NOR3xp33_ASAP7_75t_L g165 ( .A(n_166), .B(n_170), .C(n_176), .Y(n_165) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_177), .B(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
AND2x2_ASAP7_75t_L g220 ( .A(n_181), .B(n_221), .Y(n_220) );
OR2x2_ASAP7_75t_L g263 ( .A(n_181), .B(n_221), .Y(n_263) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_181), .Y(n_271) );
AND2x2_ASAP7_75t_L g394 ( .A(n_181), .B(n_290), .Y(n_394) );
AND2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
AND2x2_ASAP7_75t_L g247 ( .A(n_183), .B(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
OAI21xp33_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_206), .B(n_211), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g337 ( .A(n_196), .B(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g373 ( .A(n_196), .B(n_243), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_196), .B(n_340), .Y(n_375) );
NAND4xp25_ASAP7_75t_L g395 ( .A(n_196), .B(n_282), .C(n_338), .D(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g404 ( .A(n_196), .B(n_327), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_196), .B(n_309), .Y(n_417) );
INVx1_ASAP7_75t_L g278 ( .A(n_197), .Y(n_278) );
AND2x2_ASAP7_75t_L g402 ( .A(n_197), .B(n_364), .Y(n_402) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g261 ( .A(n_198), .Y(n_261) );
AND2x2_ASAP7_75t_L g299 ( .A(n_198), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g352 ( .A(n_198), .B(n_246), .Y(n_352) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_198), .Y(n_370) );
AND2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_205), .Y(n_198) );
AND2x2_ASAP7_75t_L g248 ( .A(n_199), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_203), .Y(n_199) );
OAI221xp5_ASAP7_75t_L g386 ( .A1(n_206), .A2(n_387), .B1(n_389), .B2(n_393), .C(n_395), .Y(n_386) );
NAND2x1p5_ASAP7_75t_L g206 ( .A(n_207), .B(n_208), .Y(n_206) );
NAND2x1p5_ASAP7_75t_L g292 ( .A(n_208), .B(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_208), .B(n_239), .Y(n_316) );
AND2x4_ASAP7_75t_L g342 ( .A(n_208), .B(n_331), .Y(n_342) );
AND2x2_ASAP7_75t_L g353 ( .A(n_208), .B(n_282), .Y(n_353) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g258 ( .A(n_210), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_213), .Y(n_211) );
INVx1_ASAP7_75t_L g237 ( .A(n_213), .Y(n_237) );
AOI322xp5_ASAP7_75t_L g336 ( .A1(n_213), .A2(n_245), .A3(n_326), .B1(n_337), .B2(n_340), .C1(n_342), .C2(n_343), .Y(n_336) );
INVx3_ASAP7_75t_L g267 ( .A(n_214), .Y(n_267) );
INVx1_ASAP7_75t_L g347 ( .A(n_214), .Y(n_347) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
INVx1_ASAP7_75t_L g241 ( .A(n_215), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_217), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
AOI32xp33_ASAP7_75t_L g407 ( .A1(n_219), .A2(n_408), .A3(n_410), .B1(n_411), .B2(n_412), .Y(n_407) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_220), .B(n_308), .Y(n_350) );
AND2x2_ASAP7_75t_L g354 ( .A(n_220), .B(n_260), .Y(n_354) );
INVx1_ASAP7_75t_L g244 ( .A(n_221), .Y(n_244) );
INVx1_ASAP7_75t_L g290 ( .A(n_221), .Y(n_290) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_221), .Y(n_310) );
HB1xp67_ASAP7_75t_L g320 ( .A(n_221), .Y(n_320) );
AND2x4_ASAP7_75t_L g327 ( .A(n_221), .B(n_300), .Y(n_327) );
INVx2_ASAP7_75t_L g364 ( .A(n_221), .Y(n_364) );
AO31x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_228), .A3(n_233), .B(n_234), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_227), .Y(n_225) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_230), .Y(n_436) );
AOI21xp33_ASAP7_75t_SL g236 ( .A1(n_237), .A2(n_238), .B(n_242), .Y(n_236) );
NOR2xp67_ASAP7_75t_L g366 ( .A(n_238), .B(n_283), .Y(n_366) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g365 ( .A(n_239), .B(n_283), .Y(n_365) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
INVx1_ASAP7_75t_L g294 ( .A(n_240), .Y(n_294) );
INVx1_ASAP7_75t_L g312 ( .A(n_240), .Y(n_312) );
AND2x2_ASAP7_75t_L g408 ( .A(n_240), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_241), .B(n_273), .Y(n_272) );
INVx2_ASAP7_75t_L g331 ( .A(n_241), .Y(n_331) );
OR2x2_ASAP7_75t_L g356 ( .A(n_241), .B(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g421 ( .A(n_242), .Y(n_421) );
NAND2x1p5_ASAP7_75t_SL g242 ( .A(n_243), .B(n_245), .Y(n_242) );
INVx2_ASAP7_75t_SL g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g397 ( .A(n_244), .Y(n_397) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g277 ( .A(n_246), .Y(n_277) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_246), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_247), .Y(n_287) );
INVx1_ASAP7_75t_L g291 ( .A(n_247), .Y(n_291) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_254), .B(n_259), .Y(n_252) );
AOI321xp33_ASAP7_75t_L g422 ( .A1(n_253), .A2(n_324), .A3(n_423), .B1(n_424), .B2(n_426), .C(n_427), .Y(n_422) );
AND2x4_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g332 ( .A(n_256), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_258), .B(n_339), .Y(n_413) );
INVx2_ASAP7_75t_L g429 ( .A(n_258), .Y(n_429) );
AOI22x1_ASAP7_75t_L g264 ( .A1(n_259), .A2(n_265), .B1(n_270), .B2(n_274), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_259), .A2(n_281), .B(n_284), .Y(n_280) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_262), .Y(n_259) );
AND2x4_ASAP7_75t_L g326 ( .A(n_260), .B(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g351 ( .A1(n_260), .A2(n_263), .B1(n_340), .B2(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_260), .B(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g410 ( .A(n_260), .Y(n_410) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g379 ( .A(n_263), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NOR3xp33_ASAP7_75t_L g427 ( .A(n_266), .B(n_425), .C(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx3_ASAP7_75t_L g282 ( .A(n_267), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_267), .B(n_318), .Y(n_317) );
AND2x4_ASAP7_75t_L g324 ( .A(n_267), .B(n_283), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_267), .B(n_273), .Y(n_325) );
BUFx3_ASAP7_75t_L g406 ( .A(n_268), .Y(n_406) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_269), .B(n_358), .Y(n_357) );
NOR2xp33_ASAP7_75t_SL g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp33_ASAP7_75t_L g355 ( .A(n_272), .B(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g315 ( .A(n_276), .B(n_310), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g279 ( .A(n_280), .B(n_295), .C(n_321), .Y(n_279) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
AND2x2_ASAP7_75t_L g372 ( .A(n_282), .B(n_318), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_282), .B(n_283), .Y(n_381) );
OAI22xp33_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_288), .B1(n_289), .B2(n_292), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g423 ( .A(n_289), .Y(n_423) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
AND2x2_ASAP7_75t_L g411 ( .A(n_290), .B(n_299), .Y(n_411) );
OR2x2_ASAP7_75t_L g319 ( .A(n_291), .B(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
O2A1O1Ixp5_ASAP7_75t_SL g295 ( .A1(n_296), .A2(n_306), .B(n_311), .C(n_314), .Y(n_295) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_296), .A2(n_342), .B1(n_346), .B2(n_383), .Y(n_382) );
AND2x4_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_299), .A2(n_322), .B1(n_326), .B2(n_328), .Y(n_321) );
AND2x2_ASAP7_75t_L g383 ( .A(n_299), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g341 ( .A(n_300), .Y(n_341) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B(n_304), .Y(n_300) );
AND2x2_ASAP7_75t_L g432 ( .A(n_302), .B(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g400 ( .A(n_312), .Y(n_400) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_316), .B1(n_317), .B2(n_319), .Y(n_314) );
NOR2x1_ASAP7_75t_L g426 ( .A(n_319), .B(n_425), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_324), .B(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_324), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_327), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g390 ( .A(n_327), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
BUFx2_ASAP7_75t_SL g419 ( .A(n_332), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g334 ( .A(n_335), .B(n_359), .C(n_378), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_336), .B(n_348), .Y(n_335) );
INVx1_ASAP7_75t_L g344 ( .A(n_338), .Y(n_344) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2x1_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
INVx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g376 ( .A(n_346), .B(n_377), .Y(n_376) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_353), .B1(n_354), .B2(n_355), .Y(n_348) );
NAND2xp33_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_L g361 ( .A(n_352), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g380 ( .A(n_352), .Y(n_380) );
INVx1_ASAP7_75t_L g420 ( .A(n_357), .Y(n_420) );
BUFx2_ASAP7_75t_L g377 ( .A(n_358), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_371), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_365), .B1(n_366), .B2(n_367), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_364), .Y(n_430) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_373), .B1(n_374), .B2(n_376), .Y(n_371) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g378 ( .A1(n_379), .A2(n_381), .B(n_382), .Y(n_378) );
NOR3xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_398), .C(n_414), .Y(n_385) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_401), .B1(n_403), .B2(n_405), .C(n_407), .Y(n_398) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_418), .C(n_422), .Y(n_414) );
INVxp67_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_420), .B(n_421), .Y(n_418) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
BUFx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OA21x2_ASAP7_75t_L g609 ( .A1(n_433), .A2(n_610), .B(n_611), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
XNOR2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_451), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_440), .B1(n_449), .B2(n_450), .Y(n_438) );
CKINVDCx20_ASAP7_75t_R g439 ( .A(n_440), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_442), .B1(n_443), .B2(n_444), .Y(n_440) );
CKINVDCx16_ASAP7_75t_R g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_447), .B2(n_448), .Y(n_444) );
CKINVDCx14_ASAP7_75t_R g448 ( .A(n_445), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g447 ( .A(n_446), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B1(n_580), .B2(n_581), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_452), .A2(n_453), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_536), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_488), .C(n_523), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_482), .B2(n_483), .Y(n_456) );
INVx4_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_471), .Y(n_460) );
AND2x4_ASAP7_75t_L g528 ( .A(n_461), .B(n_495), .Y(n_528) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_465), .Y(n_461) );
AND2x2_ASAP7_75t_L g487 ( .A(n_462), .B(n_466), .Y(n_487) );
AND2x2_ASAP7_75t_L g505 ( .A(n_462), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g543 ( .A(n_462), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_463), .B(n_470), .Y(n_469) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
NAND2xp33_ASAP7_75t_L g467 ( .A(n_464), .B(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g474 ( .A(n_464), .Y(n_474) );
NAND2xp33_ASAP7_75t_L g480 ( .A(n_464), .B(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
INVx1_ASAP7_75t_L g508 ( .A(n_464), .Y(n_508) );
AND2x4_ASAP7_75t_L g542 ( .A(n_465), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_468), .B(n_522), .Y(n_521) );
INVxp67_ASAP7_75t_L g591 ( .A(n_468), .Y(n_591) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_470), .A2(n_507), .B(n_508), .Y(n_506) );
AND2x2_ASAP7_75t_L g486 ( .A(n_471), .B(n_487), .Y(n_486) );
AND2x4_ASAP7_75t_L g564 ( .A(n_471), .B(n_542), .Y(n_564) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_476), .Y(n_471) );
INVx2_ASAP7_75t_L g496 ( .A(n_472), .Y(n_496) );
AND2x2_ASAP7_75t_L g501 ( .A(n_472), .B(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g544 ( .A(n_472), .B(n_545), .Y(n_544) );
OR2x2_ASAP7_75t_L g558 ( .A(n_472), .B(n_546), .Y(n_558) );
AND2x4_ASAP7_75t_L g472 ( .A(n_473), .B(n_475), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_474), .B(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_L g519 ( .A(n_474), .Y(n_519) );
NAND3xp33_ASAP7_75t_L g517 ( .A(n_475), .B(n_518), .C(n_520), .Y(n_517) );
AND2x4_ASAP7_75t_L g495 ( .A(n_476), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g546 ( .A(n_477), .Y(n_546) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_480), .Y(n_477) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g494 ( .A(n_487), .B(n_495), .Y(n_494) );
AND2x2_ASAP7_75t_L g553 ( .A(n_487), .B(n_544), .Y(n_553) );
AND2x4_ASAP7_75t_L g556 ( .A(n_487), .B(n_557), .Y(n_556) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_490), .B(n_497), .Y(n_488) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g533 ( .A(n_495), .B(n_534), .Y(n_533) );
AND2x2_ASAP7_75t_L g569 ( .A(n_495), .B(n_542), .Y(n_569) );
INVx4_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx5_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_501), .B(n_505), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g513 ( .A(n_503), .Y(n_513) );
HB1xp67_ASAP7_75t_L g588 ( .A(n_504), .Y(n_588) );
INVx4_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx3_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_517), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_519), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g534 ( .A(n_520), .B(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_522), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B1(n_529), .B2(n_530), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx6f_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g550 ( .A(n_534), .B(n_544), .Y(n_550) );
AND2x4_ASAP7_75t_L g579 ( .A(n_534), .B(n_574), .Y(n_579) );
NOR2xp67_ASAP7_75t_L g536 ( .A(n_537), .B(n_559), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_551), .Y(n_537) );
BUFx12f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
BUFx12f_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
AND2x4_ASAP7_75t_L g573 ( .A(n_542), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx4_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx8_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
BUFx8_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx3_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx12f_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g574 ( .A(n_558), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_570), .Y(n_559) );
BUFx4f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx3_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx6_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_580), .Y(n_581) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_593), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g603 ( .A(n_586), .B(n_593), .Y(n_603) );
AOI211xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_588), .B(n_589), .C(n_592), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
OR2x2_ASAP7_75t_L g605 ( .A(n_594), .B(n_597), .Y(n_605) );
INVx1_ASAP7_75t_L g610 ( .A(n_594), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_594), .B(n_596), .Y(n_611) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI222xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_602), .B1(n_604), .B2(n_606), .C1(n_608), .C2(n_612), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_600), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
endmodule