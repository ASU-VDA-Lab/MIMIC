module fake_ariane_813_n_5221 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_636, n_427, n_108, n_587, n_497, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_5221);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_5221;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_4824;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_3482;
wire n_823;
wire n_1900;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_3359;
wire n_3841;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_1032;
wire n_1592;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_688;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_986;
wire n_1104;
wire n_2802;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1044;
wire n_1714;
wire n_4429;
wire n_3340;
wire n_5053;
wire n_1243;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_1256;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_1048;
wire n_2343;
wire n_775;
wire n_3380;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_1056;
wire n_3168;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_3645;
wire n_793;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_1141;
wire n_3457;
wire n_840;
wire n_2324;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_3941;
wire n_1915;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_1091;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_998;
wire n_3592;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_1001;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_1169;
wire n_789;
wire n_3181;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_721;
wire n_1084;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_3391;
wire n_912;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_3508;
wire n_4129;
wire n_1105;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1614;
wire n_1377;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_1747;
wire n_3990;
wire n_1171;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_4097;
wire n_4162;
wire n_779;
wire n_4790;
wire n_4173;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_3738;
wire n_894;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_918;
wire n_1968;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_4333;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_994;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_856;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_831;
wire n_3681;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_684;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2085;
wire n_2432;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_1410;
wire n_939;
wire n_2297;
wire n_4203;
wire n_1325;
wire n_1223;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_3763;
wire n_933;
wire n_3499;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_1421;
wire n_2423;
wire n_2208;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_1069;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_2407;
wire n_690;
wire n_2243;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_2731;
wire n_3703;
wire n_1246;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5050;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1468;
wire n_1253;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_2072;
wire n_3852;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_686;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_1864;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_2133;
wire n_2497;
wire n_879;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_2749;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_1022;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_4435;
wire n_3248;
wire n_2387;
wire n_4318;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_4673;
wire n_2793;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2597;
wire n_1077;
wire n_2321;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_2039;
wire n_1285;
wire n_761;
wire n_733;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1982;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_938;
wire n_1891;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_1314;
wire n_1512;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_693;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_2727;
wire n_942;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_3562;
wire n_2281;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2499;
wire n_2549;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_4794;
wire n_4843;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_824;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5112;
wire n_1627;
wire n_2903;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_4836;
wire n_3889;
wire n_3262;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_3682;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_861;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_3648;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_876;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_790;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_1426;
wire n_4969;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_3470;
wire n_1407;
wire n_2865;
wire n_973;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_5133;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;

INVx1_ASAP7_75t_SL g684 ( 
.A(n_661),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_282),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_156),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_405),
.Y(n_687)
);

CKINVDCx20_ASAP7_75t_R g688 ( 
.A(n_635),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_46),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_414),
.Y(n_690)
);

BUFx10_ASAP7_75t_L g691 ( 
.A(n_314),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_637),
.Y(n_692)
);

BUFx2_ASAP7_75t_L g693 ( 
.A(n_238),
.Y(n_693)
);

BUFx5_ASAP7_75t_L g694 ( 
.A(n_660),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_533),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_664),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_578),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_235),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_513),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_531),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_493),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_342),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_624),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_218),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_418),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_424),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_258),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_470),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_537),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_36),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_163),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_434),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_77),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_268),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_256),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_611),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_421),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_437),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_585),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_44),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_673),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_345),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_627),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_282),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_312),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_267),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_537),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_331),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_555),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_357),
.Y(n_730)
);

CKINVDCx16_ASAP7_75t_R g731 ( 
.A(n_68),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_432),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_543),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_326),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_295),
.Y(n_735)
);

CKINVDCx16_ASAP7_75t_R g736 ( 
.A(n_267),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_351),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_578),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_429),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_462),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_168),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_257),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_285),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_573),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_232),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_318),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_675),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_525),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_298),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_403),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_13),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_649),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_392),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_557),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_541),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_306),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_430),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_62),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_679),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_622),
.Y(n_760)
);

CKINVDCx20_ASAP7_75t_R g761 ( 
.A(n_587),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_397),
.Y(n_762)
);

BUFx5_ASAP7_75t_L g763 ( 
.A(n_565),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_590),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_417),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_218),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_672),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_490),
.Y(n_768)
);

INVx1_ASAP7_75t_SL g769 ( 
.A(n_377),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_432),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_133),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_413),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_401),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_454),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_46),
.Y(n_775)
);

HB1xp67_ASAP7_75t_L g776 ( 
.A(n_573),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_117),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_22),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_332),
.Y(n_779)
);

BUFx10_ASAP7_75t_L g780 ( 
.A(n_122),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_98),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_374),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_470),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_562),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_70),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_586),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_671),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_580),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_84),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_307),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_144),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_647),
.Y(n_792)
);

BUFx6f_ASAP7_75t_L g793 ( 
.A(n_136),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_598),
.Y(n_794)
);

BUFx3_ASAP7_75t_L g795 ( 
.A(n_541),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_25),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_407),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_405),
.Y(n_798)
);

CKINVDCx16_ASAP7_75t_R g799 ( 
.A(n_487),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_116),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_47),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_146),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_180),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_127),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_37),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_623),
.Y(n_806)
);

CKINVDCx14_ASAP7_75t_R g807 ( 
.A(n_565),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_159),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_535),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_480),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_643),
.Y(n_811)
);

CKINVDCx16_ASAP7_75t_R g812 ( 
.A(n_510),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_663),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_39),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_289),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_656),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_447),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_404),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_618),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_525),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_533),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_677),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_231),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_229),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_638),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_25),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_596),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_651),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_420),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_474),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_209),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_268),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_428),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_269),
.Y(n_834)
);

BUFx8_ASAP7_75t_SL g835 ( 
.A(n_445),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_118),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_435),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_655),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_676),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_119),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_579),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_95),
.Y(n_842)
);

BUFx10_ASAP7_75t_L g843 ( 
.A(n_597),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_442),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_667),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_236),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_659),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_127),
.Y(n_848)
);

INVxp67_ASAP7_75t_L g849 ( 
.A(n_207),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_645),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_119),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_518),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_135),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_491),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_156),
.Y(n_855)
);

BUFx3_ASAP7_75t_L g856 ( 
.A(n_95),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_614),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_325),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_448),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_670),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_254),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_45),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_199),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_641),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_341),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_215),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_630),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_604),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_225),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_549),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_148),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_640),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_359),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_658),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_580),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_250),
.Y(n_876)
);

CKINVDCx5p33_ASAP7_75t_R g877 ( 
.A(n_487),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_152),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_532),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_224),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_250),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_154),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_301),
.Y(n_883)
);

BUFx10_ASAP7_75t_L g884 ( 
.A(n_491),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_357),
.Y(n_885)
);

BUFx8_ASAP7_75t_SL g886 ( 
.A(n_666),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_180),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_94),
.Y(n_888)
);

CKINVDCx20_ASAP7_75t_R g889 ( 
.A(n_258),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_548),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_612),
.Y(n_891)
);

CKINVDCx16_ASAP7_75t_R g892 ( 
.A(n_518),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_527),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_344),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_123),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_589),
.Y(n_896)
);

CKINVDCx16_ASAP7_75t_R g897 ( 
.A(n_452),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_49),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_646),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_648),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_540),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_40),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_228),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_493),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_338),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_147),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_530),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_37),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_581),
.Y(n_909)
);

CKINVDCx20_ASAP7_75t_R g910 ( 
.A(n_334),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_225),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_373),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_100),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_181),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_639),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_680),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_668),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_615),
.Y(n_918)
);

INVx2_ASAP7_75t_SL g919 ( 
.A(n_582),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_62),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_184),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_188),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_204),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_184),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_3),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_40),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_59),
.Y(n_927)
);

BUFx10_ASAP7_75t_L g928 ( 
.A(n_488),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_277),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_30),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_135),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_365),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_466),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_316),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_519),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_188),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_304),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_23),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_125),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_6),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_528),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_136),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_299),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_389),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_1),
.Y(n_945)
);

BUFx2_ASAP7_75t_SL g946 ( 
.A(n_217),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_208),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_130),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_41),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_391),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_205),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_481),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_257),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_559),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_519),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_463),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_220),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_446),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_665),
.Y(n_959)
);

CKINVDCx16_ASAP7_75t_R g960 ( 
.A(n_176),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_132),
.Y(n_961)
);

INVx2_ASAP7_75t_SL g962 ( 
.A(n_416),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_431),
.Y(n_963)
);

CKINVDCx14_ASAP7_75t_R g964 ( 
.A(n_193),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_1),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_654),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_118),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_521),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_246),
.Y(n_969)
);

CKINVDCx20_ASAP7_75t_R g970 ( 
.A(n_547),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_181),
.Y(n_971)
);

INVx2_ASAP7_75t_SL g972 ( 
.A(n_593),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_449),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_185),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_404),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_253),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_261),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_355),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_411),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_237),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_344),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_396),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_682),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_130),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_242),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_476),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_78),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_595),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_305),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_387),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_549),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_314),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_463),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_227),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_616),
.Y(n_995)
);

BUFx3_ASAP7_75t_L g996 ( 
.A(n_26),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_293),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_550),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_2),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_650),
.Y(n_1000)
);

BUFx3_ASAP7_75t_L g1001 ( 
.A(n_662),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_302),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_468),
.Y(n_1003)
);

CKINVDCx20_ASAP7_75t_R g1004 ( 
.A(n_553),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_419),
.Y(n_1005)
);

INVxp67_ASAP7_75t_L g1006 ( 
.A(n_204),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_21),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_528),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_397),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_385),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_108),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_145),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_292),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_251),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_9),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_56),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_452),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_657),
.Y(n_1018)
);

INVx2_ASAP7_75t_SL g1019 ( 
.A(n_17),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_695),
.Y(n_1020)
);

CKINVDCx16_ASAP7_75t_R g1021 ( 
.A(n_807),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_835),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_886),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_695),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_731),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_718),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_736),
.Y(n_1027)
);

BUFx10_ASAP7_75t_L g1028 ( 
.A(n_723),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_799),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_705),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_812),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_763),
.Y(n_1032)
);

INVx1_ASAP7_75t_SL g1033 ( 
.A(n_705),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_718),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_892),
.Y(n_1035)
);

CKINVDCx20_ASAP7_75t_R g1036 ( 
.A(n_713),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_713),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_897),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_864),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_960),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_964),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_744),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_685),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_744),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_714),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_763),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_757),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_786),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_891),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_757),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_763),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_688),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_795),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_688),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_795),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_830),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_761),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_830),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_856),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_761),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_856),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_899),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_942),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_942),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_899),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_714),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_949),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_983),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_754),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_983),
.Y(n_1070)
);

CKINVDCx16_ASAP7_75t_R g1071 ( 
.A(n_691),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_843),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_843),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_864),
.Y(n_1074)
);

BUFx10_ASAP7_75t_L g1075 ( 
.A(n_732),
.Y(n_1075)
);

CKINVDCx16_ASAP7_75t_R g1076 ( 
.A(n_691),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_949),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_693),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_954),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_754),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_954),
.Y(n_1081)
);

NOR2xp67_ASAP7_75t_L g1082 ( 
.A(n_1019),
.B(n_0),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_687),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_996),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_996),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_763),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_690),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_763),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_763),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_691),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_741),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_762),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_697),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_763),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_699),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_701),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_700),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_706),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_702),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_707),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_881),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_709),
.Y(n_1102)
);

INVx2_ASAP7_75t_SL g1103 ( 
.A(n_741),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_956),
.Y(n_1104)
);

HB1xp67_ASAP7_75t_L g1105 ( 
.A(n_708),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_710),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_843),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_733),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_734),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_732),
.Y(n_1110)
);

CKINVDCx20_ASAP7_75t_R g1111 ( 
.A(n_762),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_735),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_732),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_984),
.Y(n_1114)
);

CKINVDCx20_ASAP7_75t_R g1115 ( 
.A(n_774),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_711),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_991),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_732),
.Y(n_1118)
);

INVx1_ASAP7_75t_SL g1119 ( 
.A(n_774),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_732),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_726),
.Y(n_1121)
);

CKINVDCx16_ASAP7_75t_R g1122 ( 
.A(n_741),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_737),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_738),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_739),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_L g1126 ( 
.A(n_1019),
.B(n_0),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_740),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_729),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_793),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_730),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_742),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_753),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_766),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_770),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_745),
.Y(n_1135)
);

CKINVDCx16_ASAP7_75t_R g1136 ( 
.A(n_780),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_746),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_748),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_749),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_772),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_797),
.Y(n_1141)
);

CKINVDCx16_ASAP7_75t_R g1142 ( 
.A(n_780),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_750),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_751),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_797),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_773),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_782),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_788),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_791),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_808),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_918),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_834),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_776),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_918),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_756),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_765),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_768),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_840),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_851),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_853),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_858),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_878),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_771),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_885),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_775),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_801),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_898),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_777),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_904),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_778),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_909),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_779),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_911),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_781),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_913),
.Y(n_1175)
);

CKINVDCx16_ASAP7_75t_R g1176 ( 
.A(n_780),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1001),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_801),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_793),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_784),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_785),
.Y(n_1181)
);

INVx2_ASAP7_75t_SL g1182 ( 
.A(n_809),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_922),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_809),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_923),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_927),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_930),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_809),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_937),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_938),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_939),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_716),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_716),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_940),
.Y(n_1194)
);

CKINVDCx16_ASAP7_75t_R g1195 ( 
.A(n_884),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_719),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_865),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_719),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_837),
.B(n_2),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_941),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_789),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_951),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_968),
.Y(n_1203)
);

BUFx3_ASAP7_75t_L g1204 ( 
.A(n_1001),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_971),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_793),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_790),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_976),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_796),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_798),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_800),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_981),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_883),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_985),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_986),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_989),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_802),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_994),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_804),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_805),
.Y(n_1220)
);

INVxp33_ASAP7_75t_L g1221 ( 
.A(n_689),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1012),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_793),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_689),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_725),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_725),
.Y(n_1226)
);

CKINVDCx14_ASAP7_75t_R g1227 ( 
.A(n_721),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_743),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_743),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_755),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_793),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_755),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_810),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_814),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_758),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_815),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_884),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_817),
.Y(n_1238)
);

INVx4_ASAP7_75t_R g1239 ( 
.A(n_1018),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_758),
.Y(n_1240)
);

CKINVDCx5p33_ASAP7_75t_R g1241 ( 
.A(n_818),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_686),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_820),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1018),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_821),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_823),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_803),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_824),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_865),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_826),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_829),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1011),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_831),
.Y(n_1253)
);

BUFx5_ASAP7_75t_L g1254 ( 
.A(n_692),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_803),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1011),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1011),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_696),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_888),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_888),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_686),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_907),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_833),
.Y(n_1263)
);

BUFx2_ASAP7_75t_SL g1264 ( 
.A(n_972),
.Y(n_1264)
);

INVx2_ASAP7_75t_L g1265 ( 
.A(n_1011),
.Y(n_1265)
);

OR2x2_ASAP7_75t_L g1266 ( 
.A(n_837),
.B(n_3),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_836),
.Y(n_1267)
);

NOR2xp67_ASAP7_75t_L g1268 ( 
.A(n_919),
.B(n_4),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_841),
.Y(n_1269)
);

CKINVDCx20_ASAP7_75t_R g1270 ( 
.A(n_889),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_842),
.Y(n_1271)
);

NOR2xp33_ASAP7_75t_L g1272 ( 
.A(n_919),
.B(n_5),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_844),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1011),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_846),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_848),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_852),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_854),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_907),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_855),
.Y(n_1280)
);

BUFx2_ASAP7_75t_L g1281 ( 
.A(n_712),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_859),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_908),
.Y(n_1283)
);

CKINVDCx14_ASAP7_75t_R g1284 ( 
.A(n_721),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_703),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_889),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_908),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_861),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_912),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_862),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_816),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_890),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_912),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_921),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_921),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_935),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_935),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_747),
.Y(n_1298)
);

BUFx10_ASAP7_75t_L g1299 ( 
.A(n_972),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_957),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_890),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_957),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_910),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_792),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_863),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_967),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_794),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_967),
.Y(n_1308)
);

INVx2_ASAP7_75t_SL g1309 ( 
.A(n_884),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_980),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_828),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_980),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_L g1313 ( 
.A(n_816),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_998),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_998),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_866),
.Y(n_1316)
);

HB1xp67_ASAP7_75t_L g1317 ( 
.A(n_712),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_869),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_850),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_870),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_962),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_871),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_962),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_928),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_715),
.Y(n_1325)
);

CKINVDCx14_ASAP7_75t_R g1326 ( 
.A(n_959),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_873),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_715),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_928),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_928),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_910),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_959),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_946),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_896),
.Y(n_1334)
);

CKINVDCx14_ASAP7_75t_R g1335 ( 
.A(n_752),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_915),
.Y(n_1336)
);

CKINVDCx16_ASAP7_75t_R g1337 ( 
.A(n_944),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_917),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_875),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_876),
.Y(n_1340)
);

BUFx3_ASAP7_75t_L g1341 ( 
.A(n_966),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_944),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_877),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_717),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_995),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_783),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_879),
.Y(n_1347)
);

INVxp67_ASAP7_75t_L g1348 ( 
.A(n_717),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_849),
.B(n_4),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_838),
.Y(n_1350)
);

BUFx2_ASAP7_75t_L g1351 ( 
.A(n_720),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_694),
.Y(n_1352)
);

CKINVDCx20_ASAP7_75t_R g1353 ( 
.A(n_970),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1006),
.Y(n_1354)
);

BUFx2_ASAP7_75t_L g1355 ( 
.A(n_720),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_722),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_880),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_882),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_887),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_893),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_894),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_722),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_694),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_724),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_724),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_694),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_727),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_727),
.Y(n_1368)
);

CKINVDCx5p33_ASAP7_75t_R g1369 ( 
.A(n_895),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_901),
.Y(n_1370)
);

CKINVDCx16_ASAP7_75t_R g1371 ( 
.A(n_970),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_950),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_902),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_903),
.Y(n_1374)
);

CKINVDCx20_ASAP7_75t_R g1375 ( 
.A(n_973),
.Y(n_1375)
);

CKINVDCx20_ASAP7_75t_R g1376 ( 
.A(n_973),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_950),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_952),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_952),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_905),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_953),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_698),
.B(n_5),
.Y(n_1382)
);

INVx3_ASAP7_75t_L g1383 ( 
.A(n_838),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1023),
.Y(n_1384)
);

CKINVDCx20_ASAP7_75t_R g1385 ( 
.A(n_1030),
.Y(n_1385)
);

NOR2xp33_ASAP7_75t_L g1386 ( 
.A(n_1227),
.B(n_684),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1086),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1088),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1052),
.Y(n_1389)
);

NOR2xp33_ASAP7_75t_L g1390 ( 
.A(n_1227),
.B(n_1284),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1025),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1052),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1252),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1264),
.B(n_806),
.Y(n_1394)
);

NOR2xp67_ASAP7_75t_L g1395 ( 
.A(n_1072),
.B(n_759),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_1054),
.Y(n_1396)
);

NOR2xp67_ASAP7_75t_L g1397 ( 
.A(n_1072),
.B(n_760),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1089),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1284),
.B(n_764),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1094),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1095),
.Y(n_1401)
);

CKINVDCx20_ASAP7_75t_R g1402 ( 
.A(n_1030),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1054),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1057),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1036),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1073),
.B(n_767),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1097),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1099),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1057),
.Y(n_1409)
);

HB1xp67_ASAP7_75t_L g1410 ( 
.A(n_1027),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1060),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1100),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1102),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_1060),
.Y(n_1414)
);

INVxp67_ASAP7_75t_L g1415 ( 
.A(n_1261),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1106),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1116),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1252),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1036),
.Y(n_1419)
);

INVxp67_ASAP7_75t_SL g1420 ( 
.A(n_1074),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1121),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1062),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1062),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1128),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1130),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1065),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1045),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1131),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1065),
.Y(n_1429)
);

INVxp67_ASAP7_75t_SL g1430 ( 
.A(n_1074),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1132),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1133),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1281),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1134),
.Y(n_1434)
);

INVxp67_ASAP7_75t_L g1435 ( 
.A(n_1325),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1140),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1326),
.B(n_787),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1146),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1068),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1147),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1029),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_1045),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1326),
.B(n_811),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1068),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1148),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1149),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1070),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1150),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1070),
.Y(n_1449)
);

INVxp67_ASAP7_75t_L g1450 ( 
.A(n_1328),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1152),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_1022),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1066),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1158),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1031),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_1192),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1066),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1159),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1160),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1161),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1192),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1162),
.Y(n_1462)
);

CKINVDCx20_ASAP7_75t_R g1463 ( 
.A(n_1080),
.Y(n_1463)
);

INVxp67_ASAP7_75t_L g1464 ( 
.A(n_1351),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1252),
.Y(n_1465)
);

INVxp67_ASAP7_75t_SL g1466 ( 
.A(n_1154),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1335),
.B(n_813),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1164),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1335),
.B(n_819),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1167),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1169),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1171),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1021),
.B(n_953),
.Y(n_1473)
);

HB1xp67_ASAP7_75t_L g1474 ( 
.A(n_1035),
.Y(n_1474)
);

INVxp67_ASAP7_75t_L g1475 ( 
.A(n_1355),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1193),
.Y(n_1476)
);

CKINVDCx16_ASAP7_75t_R g1477 ( 
.A(n_1071),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1080),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_1193),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1092),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_1196),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1173),
.Y(n_1482)
);

CKINVDCx20_ASAP7_75t_R g1483 ( 
.A(n_1092),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1175),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1183),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1196),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1185),
.Y(n_1487)
);

NOR2xp67_ASAP7_75t_L g1488 ( 
.A(n_1073),
.B(n_822),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1186),
.Y(n_1489)
);

NOR2xp33_ASAP7_75t_L g1490 ( 
.A(n_1198),
.B(n_1332),
.Y(n_1490)
);

INVxp67_ASAP7_75t_SL g1491 ( 
.A(n_1154),
.Y(n_1491)
);

CKINVDCx20_ASAP7_75t_R g1492 ( 
.A(n_1111),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1111),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1115),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1198),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_1115),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1204),
.B(n_825),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1332),
.Y(n_1498)
);

INVxp67_ASAP7_75t_SL g1499 ( 
.A(n_1204),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1043),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1187),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1189),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1190),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_1141),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1191),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1083),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1194),
.Y(n_1507)
);

HB1xp67_ASAP7_75t_L g1508 ( 
.A(n_1038),
.Y(n_1508)
);

INVxp33_ASAP7_75t_L g1509 ( 
.A(n_1242),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1141),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1200),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_1087),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1145),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1040),
.Y(n_1514)
);

CKINVDCx20_ASAP7_75t_R g1515 ( 
.A(n_1145),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1202),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1203),
.Y(n_1517)
);

NOR2xp67_ASAP7_75t_L g1518 ( 
.A(n_1107),
.B(n_827),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1166),
.Y(n_1519)
);

HB1xp67_ASAP7_75t_L g1520 ( 
.A(n_1033),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1205),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1208),
.Y(n_1522)
);

NOR2xp67_ASAP7_75t_L g1523 ( 
.A(n_1107),
.B(n_839),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1212),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_1093),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1214),
.Y(n_1526)
);

BUFx6f_ASAP7_75t_L g1527 ( 
.A(n_1252),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1215),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1037),
.Y(n_1529)
);

INVxp67_ASAP7_75t_L g1530 ( 
.A(n_1317),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1166),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1096),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1216),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1257),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1218),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1257),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1257),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1178),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1178),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1069),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1098),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1222),
.Y(n_1542)
);

CKINVDCx20_ASAP7_75t_R g1543 ( 
.A(n_1197),
.Y(n_1543)
);

INVxp67_ASAP7_75t_SL g1544 ( 
.A(n_1244),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1039),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1039),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_1108),
.Y(n_1547)
);

CKINVDCx20_ASAP7_75t_R g1548 ( 
.A(n_1197),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1109),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1112),
.Y(n_1550)
);

INVxp67_ASAP7_75t_SL g1551 ( 
.A(n_1244),
.Y(n_1551)
);

INVxp67_ASAP7_75t_SL g1552 ( 
.A(n_1039),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1039),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1123),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1299),
.B(n_845),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1151),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1151),
.Y(n_1557)
);

CKINVDCx20_ASAP7_75t_R g1558 ( 
.A(n_1270),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_1124),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1151),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1125),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_1257),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1299),
.B(n_847),
.Y(n_1563)
);

CKINVDCx20_ASAP7_75t_R g1564 ( 
.A(n_1270),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_1127),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_1135),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1137),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_1138),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1151),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1177),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_1139),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1177),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1286),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1177),
.Y(n_1574)
);

INVxp67_ASAP7_75t_SL g1575 ( 
.A(n_1177),
.Y(n_1575)
);

NOR2xp67_ASAP7_75t_L g1576 ( 
.A(n_1048),
.B(n_1344),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_1143),
.Y(n_1577)
);

XOR2xp5_ASAP7_75t_L g1578 ( 
.A(n_1286),
.B(n_1292),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1231),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1333),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1291),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1144),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1155),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1291),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1291),
.Y(n_1585)
);

NOR2xp67_ASAP7_75t_L g1586 ( 
.A(n_1048),
.B(n_857),
.Y(n_1586)
);

INVxp67_ASAP7_75t_SL g1587 ( 
.A(n_1231),
.Y(n_1587)
);

CKINVDCx16_ASAP7_75t_R g1588 ( 
.A(n_1076),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1291),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1156),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1292),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1231),
.Y(n_1592)
);

INVxp33_ASAP7_75t_SL g1593 ( 
.A(n_1157),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1313),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1119),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1163),
.Y(n_1596)
);

INVxp33_ASAP7_75t_SL g1597 ( 
.A(n_1165),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1313),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1168),
.Y(n_1599)
);

CKINVDCx20_ASAP7_75t_R g1600 ( 
.A(n_1301),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1301),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1170),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1299),
.B(n_860),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1313),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1313),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_1303),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1249),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1350),
.Y(n_1608)
);

CKINVDCx5p33_ASAP7_75t_R g1609 ( 
.A(n_1172),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1350),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1350),
.Y(n_1611)
);

INVxp67_ASAP7_75t_L g1612 ( 
.A(n_1078),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1174),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1101),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1350),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1020),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1180),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_1303),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1024),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1026),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1110),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1034),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1041),
.B(n_867),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1110),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1042),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1044),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1221),
.B(n_955),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_1181),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1201),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1047),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1050),
.Y(n_1631)
);

INVxp67_ASAP7_75t_SL g1632 ( 
.A(n_1221),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1053),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1055),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1207),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1209),
.Y(n_1636)
);

HB1xp67_ASAP7_75t_L g1637 ( 
.A(n_1342),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1056),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1210),
.Y(n_1639)
);

CKINVDCx20_ASAP7_75t_R g1640 ( 
.A(n_1331),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1075),
.Y(n_1641)
);

NOR2xp67_ASAP7_75t_L g1642 ( 
.A(n_1348),
.B(n_868),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1331),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_1211),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1058),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1217),
.Y(n_1646)
);

CKINVDCx20_ASAP7_75t_R g1647 ( 
.A(n_1353),
.Y(n_1647)
);

INVxp33_ASAP7_75t_L g1648 ( 
.A(n_1105),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1219),
.Y(n_1649)
);

CKINVDCx16_ASAP7_75t_R g1650 ( 
.A(n_1090),
.Y(n_1650)
);

CKINVDCx20_ASAP7_75t_R g1651 ( 
.A(n_1353),
.Y(n_1651)
);

CKINVDCx20_ASAP7_75t_R g1652 ( 
.A(n_1375),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1362),
.B(n_872),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1059),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1220),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1113),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1061),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1356),
.B(n_874),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_1233),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1063),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1064),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1234),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1067),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1364),
.B(n_900),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_1375),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1077),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1236),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1367),
.B(n_916),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1122),
.B(n_955),
.Y(n_1669)
);

INVxp67_ASAP7_75t_SL g1670 ( 
.A(n_1383),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1079),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1238),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1081),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1241),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1075),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_1243),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1084),
.Y(n_1677)
);

INVxp33_ASAP7_75t_L g1678 ( 
.A(n_1153),
.Y(n_1678)
);

NAND2xp33_ASAP7_75t_R g1679 ( 
.A(n_1339),
.B(n_958),
.Y(n_1679)
);

INVxp67_ASAP7_75t_SL g1680 ( 
.A(n_1383),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1085),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1376),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1376),
.Y(n_1683)
);

CKINVDCx5p33_ASAP7_75t_R g1684 ( 
.A(n_1245),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1298),
.Y(n_1685)
);

CKINVDCx20_ASAP7_75t_R g1686 ( 
.A(n_1337),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1298),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1304),
.Y(n_1688)
);

CKINVDCx20_ASAP7_75t_R g1689 ( 
.A(n_1371),
.Y(n_1689)
);

BUFx3_ASAP7_75t_L g1690 ( 
.A(n_1384),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1386),
.B(n_1254),
.Y(n_1691)
);

INVxp67_ASAP7_75t_L g1692 ( 
.A(n_1520),
.Y(n_1692)
);

INVx5_ASAP7_75t_L g1693 ( 
.A(n_1465),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1632),
.B(n_1136),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1616),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1619),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_SL g1697 ( 
.A(n_1390),
.B(n_1254),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1627),
.B(n_1142),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1620),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1465),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1545),
.Y(n_1701)
);

INVx2_ASAP7_75t_SL g1702 ( 
.A(n_1529),
.Y(n_1702)
);

BUFx6f_ASAP7_75t_L g1703 ( 
.A(n_1465),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1546),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1387),
.A2(n_1398),
.B(n_1388),
.Y(n_1705)
);

INVx2_ASAP7_75t_L g1706 ( 
.A(n_1553),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1622),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1556),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1625),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1469),
.B(n_1258),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1626),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1420),
.B(n_1324),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1540),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1630),
.Y(n_1714)
);

OAI22xp5_ASAP7_75t_L g1715 ( 
.A1(n_1490),
.A2(n_978),
.B1(n_1003),
.B2(n_997),
.Y(n_1715)
);

AND2x2_ASAP7_75t_SL g1716 ( 
.A(n_1590),
.B(n_1266),
.Y(n_1716)
);

AND2x4_ASAP7_75t_L g1717 ( 
.A(n_1430),
.B(n_1329),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1400),
.B(n_1254),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1631),
.Y(n_1719)
);

NAND2xp33_ASAP7_75t_L g1720 ( 
.A(n_1672),
.B(n_1456),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1466),
.B(n_1330),
.Y(n_1721)
);

BUFx2_ASAP7_75t_L g1722 ( 
.A(n_1612),
.Y(n_1722)
);

OA21x2_ASAP7_75t_L g1723 ( 
.A1(n_1581),
.A2(n_1046),
.B(n_1032),
.Y(n_1723)
);

OAI22x1_ASAP7_75t_SL g1724 ( 
.A1(n_1385),
.A2(n_978),
.B1(n_1003),
.B2(n_997),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1579),
.B(n_1254),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1633),
.Y(n_1726)
);

BUFx8_ASAP7_75t_L g1727 ( 
.A(n_1655),
.Y(n_1727)
);

BUFx6f_ASAP7_75t_L g1728 ( 
.A(n_1465),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1587),
.B(n_1254),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1527),
.Y(n_1730)
);

HB1xp67_ASAP7_75t_L g1731 ( 
.A(n_1614),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1557),
.Y(n_1732)
);

INVx6_ASAP7_75t_L g1733 ( 
.A(n_1641),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1527),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1634),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1638),
.Y(n_1736)
);

INVx5_ASAP7_75t_L g1737 ( 
.A(n_1527),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1461),
.A2(n_1004),
.B1(n_1014),
.B2(n_1005),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1645),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1560),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1569),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1595),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1607),
.Y(n_1743)
);

CKINVDCx20_ASAP7_75t_R g1744 ( 
.A(n_1385),
.Y(n_1744)
);

CKINVDCx11_ASAP7_75t_R g1745 ( 
.A(n_1686),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1491),
.B(n_1091),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1654),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1657),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1570),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1499),
.B(n_1368),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1592),
.B(n_1254),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1544),
.B(n_1372),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1660),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1661),
.Y(n_1754)
);

BUFx3_ASAP7_75t_L g1755 ( 
.A(n_1452),
.Y(n_1755)
);

BUFx6f_ASAP7_75t_L g1756 ( 
.A(n_1527),
.Y(n_1756)
);

CKINVDCx20_ASAP7_75t_R g1757 ( 
.A(n_1402),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1663),
.Y(n_1758)
);

HB1xp67_ASAP7_75t_L g1759 ( 
.A(n_1637),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1572),
.Y(n_1760)
);

NOR2x1_ASAP7_75t_L g1761 ( 
.A(n_1437),
.B(n_1258),
.Y(n_1761)
);

AND2x4_ASAP7_75t_L g1762 ( 
.A(n_1551),
.B(n_1103),
.Y(n_1762)
);

OA21x2_ASAP7_75t_L g1763 ( 
.A1(n_1584),
.A2(n_1046),
.B(n_1032),
.Y(n_1763)
);

INVx2_ASAP7_75t_SL g1764 ( 
.A(n_1473),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1666),
.Y(n_1765)
);

CKINVDCx11_ASAP7_75t_R g1766 ( 
.A(n_1686),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1670),
.B(n_1254),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1680),
.B(n_1182),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_SL g1769 ( 
.A1(n_1402),
.A2(n_1004),
.B1(n_1014),
.B2(n_1005),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1500),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1405),
.A2(n_1049),
.B1(n_1195),
.B2(n_1176),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1675),
.B(n_1051),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1574),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1675),
.B(n_1051),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1580),
.B(n_1184),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1671),
.Y(n_1776)
);

OAI21x1_ASAP7_75t_L g1777 ( 
.A1(n_1675),
.A2(n_1497),
.B(n_1363),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1673),
.Y(n_1778)
);

BUFx6f_ASAP7_75t_L g1779 ( 
.A(n_1562),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1677),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1681),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1648),
.B(n_1339),
.Y(n_1782)
);

INVx2_ASAP7_75t_SL g1783 ( 
.A(n_1506),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1512),
.Y(n_1784)
);

BUFx2_ASAP7_75t_L g1785 ( 
.A(n_1525),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1648),
.B(n_1340),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1585),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1589),
.Y(n_1788)
);

BUFx6f_ASAP7_75t_L g1789 ( 
.A(n_1562),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1401),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1678),
.B(n_1509),
.Y(n_1791)
);

AND2x2_ASAP7_75t_L g1792 ( 
.A(n_1678),
.B(n_1340),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1641),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1407),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1532),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1685),
.Y(n_1796)
);

INVx6_ASAP7_75t_L g1797 ( 
.A(n_1562),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1594),
.Y(n_1798)
);

BUFx8_ASAP7_75t_SL g1799 ( 
.A(n_1689),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1552),
.B(n_1352),
.Y(n_1800)
);

AND2x4_ASAP7_75t_L g1801 ( 
.A(n_1576),
.B(n_1188),
.Y(n_1801)
);

INVx2_ASAP7_75t_L g1802 ( 
.A(n_1598),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1408),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_L g1804 ( 
.A(n_1562),
.Y(n_1804)
);

OR2x6_ASAP7_75t_L g1805 ( 
.A(n_1391),
.B(n_1237),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1604),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1509),
.B(n_1343),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1412),
.B(n_1309),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1413),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1605),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1608),
.Y(n_1811)
);

OAI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1555),
.A2(n_1363),
.B(n_1352),
.Y(n_1812)
);

OAI22xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1405),
.A2(n_1049),
.B1(n_1114),
.B2(n_1104),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1541),
.Y(n_1814)
);

AND2x6_ASAP7_75t_L g1815 ( 
.A(n_1669),
.B(n_1687),
.Y(n_1815)
);

AND2x4_ASAP7_75t_L g1816 ( 
.A(n_1416),
.B(n_1377),
.Y(n_1816)
);

OA21x2_ASAP7_75t_L g1817 ( 
.A1(n_1610),
.A2(n_1366),
.B(n_1611),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1547),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1415),
.B(n_1343),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1417),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1615),
.Y(n_1821)
);

INVx5_ASAP7_75t_L g1822 ( 
.A(n_1393),
.Y(n_1822)
);

INVx2_ASAP7_75t_L g1823 ( 
.A(n_1621),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1433),
.B(n_1347),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1421),
.Y(n_1825)
);

BUFx8_ASAP7_75t_L g1826 ( 
.A(n_1477),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1435),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1424),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1679),
.A2(n_1272),
.B1(n_1126),
.B2(n_1199),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1653),
.B(n_1378),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1425),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1621),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1450),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1624),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1549),
.Y(n_1835)
);

INVx3_ASAP7_75t_L g1836 ( 
.A(n_1688),
.Y(n_1836)
);

INVx2_ASAP7_75t_L g1837 ( 
.A(n_1624),
.Y(n_1837)
);

INVx4_ASAP7_75t_L g1838 ( 
.A(n_1550),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1464),
.B(n_1475),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1575),
.B(n_1366),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_SL g1841 ( 
.A1(n_1419),
.A2(n_1117),
.B1(n_1213),
.B2(n_1357),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1428),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1431),
.Y(n_1843)
);

OA21x2_ASAP7_75t_L g1844 ( 
.A1(n_1393),
.A2(n_1338),
.B(n_1336),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1530),
.B(n_1347),
.Y(n_1845)
);

BUFx2_ASAP7_75t_L g1846 ( 
.A(n_1554),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1656),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1656),
.Y(n_1848)
);

NOR2x1_ASAP7_75t_L g1849 ( 
.A(n_1467),
.B(n_1399),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1432),
.B(n_1434),
.Y(n_1850)
);

BUFx6f_ASAP7_75t_L g1851 ( 
.A(n_1418),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1418),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1436),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_SL g1854 ( 
.A(n_1593),
.B(n_1246),
.Y(n_1854)
);

INVx5_ASAP7_75t_L g1855 ( 
.A(n_1534),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1438),
.B(n_1345),
.Y(n_1856)
);

INVx3_ASAP7_75t_L g1857 ( 
.A(n_1534),
.Y(n_1857)
);

AND2x4_ASAP7_75t_L g1858 ( 
.A(n_1440),
.B(n_1379),
.Y(n_1858)
);

BUFx2_ASAP7_75t_L g1859 ( 
.A(n_1559),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_SL g1860 ( 
.A(n_1597),
.B(n_1359),
.Y(n_1860)
);

BUFx6f_ASAP7_75t_L g1861 ( 
.A(n_1536),
.Y(n_1861)
);

AND2x6_ASAP7_75t_L g1862 ( 
.A(n_1445),
.B(n_1446),
.Y(n_1862)
);

OAI22x1_ASAP7_75t_L g1863 ( 
.A1(n_1578),
.A2(n_1382),
.B1(n_1358),
.B2(n_1357),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1588),
.B(n_1365),
.Y(n_1864)
);

OA21x2_ASAP7_75t_L g1865 ( 
.A1(n_1536),
.A2(n_1537),
.B(n_1451),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1537),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1448),
.B(n_1304),
.Y(n_1867)
);

OA21x2_ASAP7_75t_L g1868 ( 
.A1(n_1454),
.A2(n_1319),
.B(n_1311),
.Y(n_1868)
);

BUFx6f_ASAP7_75t_L g1869 ( 
.A(n_1458),
.Y(n_1869)
);

INVx3_ASAP7_75t_L g1870 ( 
.A(n_1459),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1460),
.Y(n_1871)
);

INVx5_ASAP7_75t_L g1872 ( 
.A(n_1650),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1462),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1468),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1470),
.Y(n_1875)
);

BUFx6f_ASAP7_75t_L g1876 ( 
.A(n_1471),
.Y(n_1876)
);

AOI22xp5_ASAP7_75t_L g1877 ( 
.A1(n_1476),
.A2(n_1268),
.B1(n_1082),
.B2(n_1349),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1472),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1482),
.B(n_1311),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1484),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1485),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1410),
.B(n_1358),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1487),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1489),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1501),
.B(n_1381),
.Y(n_1885)
);

AND2x4_ASAP7_75t_L g1886 ( 
.A(n_1502),
.B(n_1285),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1503),
.B(n_1285),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1505),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1561),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1507),
.Y(n_1890)
);

INVx6_ASAP7_75t_L g1891 ( 
.A(n_1511),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1516),
.Y(n_1892)
);

NOR2xp33_ASAP7_75t_L g1893 ( 
.A(n_1664),
.B(n_1248),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1517),
.Y(n_1894)
);

BUFx6f_ASAP7_75t_L g1895 ( 
.A(n_1521),
.Y(n_1895)
);

BUFx6f_ASAP7_75t_L g1896 ( 
.A(n_1522),
.Y(n_1896)
);

OAI22xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1419),
.A2(n_1442),
.B1(n_1483),
.B2(n_1453),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_SL g1898 ( 
.A1(n_1442),
.A2(n_1008),
.B1(n_1009),
.B2(n_958),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1524),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1441),
.B(n_1250),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1526),
.Y(n_1901)
);

BUFx2_ASAP7_75t_L g1902 ( 
.A(n_1565),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1528),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1533),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1535),
.Y(n_1905)
);

OA21x2_ASAP7_75t_L g1906 ( 
.A1(n_1542),
.A2(n_1334),
.B(n_1319),
.Y(n_1906)
);

BUFx6f_ASAP7_75t_L g1907 ( 
.A(n_1394),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1455),
.B(n_1251),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1668),
.Y(n_1909)
);

AND2x4_ASAP7_75t_L g1910 ( 
.A(n_1586),
.B(n_1341),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1642),
.Y(n_1911)
);

BUFx2_ASAP7_75t_L g1912 ( 
.A(n_1566),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1603),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1658),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1443),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1563),
.B(n_1334),
.Y(n_1916)
);

BUFx2_ASAP7_75t_L g1917 ( 
.A(n_1567),
.Y(n_1917)
);

AND2x4_ASAP7_75t_L g1918 ( 
.A(n_1395),
.B(n_1341),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1568),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1571),
.Y(n_1920)
);

INVx2_ASAP7_75t_SL g1921 ( 
.A(n_1577),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1623),
.Y(n_1922)
);

INVx3_ASAP7_75t_L g1923 ( 
.A(n_1582),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1649),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1397),
.B(n_1383),
.Y(n_1925)
);

AOI22xp5_ASAP7_75t_L g1926 ( 
.A1(n_1479),
.A2(n_704),
.B1(n_769),
.B2(n_728),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1667),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1474),
.B(n_1253),
.Y(n_1928)
);

BUFx6f_ASAP7_75t_L g1929 ( 
.A(n_1583),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1406),
.Y(n_1930)
);

BUFx3_ASAP7_75t_L g1931 ( 
.A(n_1596),
.Y(n_1931)
);

INVxp67_ASAP7_75t_L g1932 ( 
.A(n_1508),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1488),
.B(n_1307),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1518),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1523),
.B(n_1307),
.Y(n_1935)
);

AND2x6_ASAP7_75t_L g1936 ( 
.A(n_1599),
.B(n_1113),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1602),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1389),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1609),
.Y(n_1939)
);

BUFx6f_ASAP7_75t_L g1940 ( 
.A(n_1613),
.Y(n_1940)
);

INVx2_ASAP7_75t_L g1941 ( 
.A(n_1617),
.Y(n_1941)
);

HB1xp67_ASAP7_75t_L g1942 ( 
.A(n_1392),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1514),
.B(n_1263),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1481),
.A2(n_832),
.B1(n_1009),
.B2(n_1008),
.Y(n_1944)
);

BUFx6f_ASAP7_75t_L g1945 ( 
.A(n_1628),
.Y(n_1945)
);

AND2x4_ASAP7_75t_L g1946 ( 
.A(n_1629),
.B(n_1346),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1486),
.Y(n_1947)
);

NOR2x1_ASAP7_75t_L g1948 ( 
.A(n_1689),
.B(n_1354),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1635),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1495),
.Y(n_1950)
);

NOR2x1_ASAP7_75t_L g1951 ( 
.A(n_1684),
.B(n_1321),
.Y(n_1951)
);

BUFx6f_ASAP7_75t_L g1952 ( 
.A(n_1636),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1639),
.B(n_1267),
.Y(n_1953)
);

OA21x2_ASAP7_75t_L g1954 ( 
.A1(n_1498),
.A2(n_1120),
.B(n_1118),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1644),
.B(n_1269),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1646),
.B(n_1118),
.Y(n_1956)
);

NOR2x1_ASAP7_75t_L g1957 ( 
.A(n_1659),
.B(n_1323),
.Y(n_1957)
);

INVx5_ASAP7_75t_L g1958 ( 
.A(n_1662),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1674),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1676),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1396),
.A2(n_1010),
.B1(n_906),
.B2(n_920),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1403),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1404),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1409),
.B(n_1327),
.Y(n_1964)
);

BUFx6f_ASAP7_75t_L g1965 ( 
.A(n_1411),
.Y(n_1965)
);

OA21x2_ASAP7_75t_L g1966 ( 
.A1(n_1414),
.A2(n_1129),
.B(n_1120),
.Y(n_1966)
);

INVx3_ASAP7_75t_L g1967 ( 
.A(n_1422),
.Y(n_1967)
);

AOI22xp5_ASAP7_75t_L g1968 ( 
.A1(n_1423),
.A2(n_1010),
.B1(n_914),
.B2(n_925),
.Y(n_1968)
);

NOR2x1_ASAP7_75t_L g1969 ( 
.A(n_1427),
.B(n_1283),
.Y(n_1969)
);

INVx4_ASAP7_75t_L g1970 ( 
.A(n_1426),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1429),
.Y(n_1971)
);

BUFx6f_ASAP7_75t_L g1972 ( 
.A(n_1439),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1444),
.Y(n_1973)
);

OAI22xp5_ASAP7_75t_L g1974 ( 
.A1(n_1447),
.A2(n_926),
.B1(n_929),
.B2(n_924),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1449),
.Y(n_1975)
);

AND2x4_ASAP7_75t_L g1976 ( 
.A(n_1457),
.B(n_1283),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1463),
.B(n_1271),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1478),
.B(n_1273),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1695),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1922),
.B(n_1275),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1868),
.Y(n_1981)
);

OAI21x1_ASAP7_75t_L g1982 ( 
.A1(n_1812),
.A2(n_1179),
.B(n_1129),
.Y(n_1982)
);

BUFx6f_ASAP7_75t_L g1983 ( 
.A(n_1700),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1696),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1723),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1699),
.Y(n_1986)
);

INVx2_ASAP7_75t_L g1987 ( 
.A(n_1723),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_1700),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1713),
.B(n_1276),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1713),
.B(n_1277),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1909),
.B(n_1278),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1707),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1716),
.B(n_1280),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1763),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1709),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1763),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_L g1997 ( 
.A(n_1830),
.B(n_1282),
.Y(n_1997)
);

CKINVDCx16_ASAP7_75t_R g1998 ( 
.A(n_1744),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1711),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1714),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1830),
.B(n_1288),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1719),
.Y(n_2002)
);

BUFx8_ASAP7_75t_L g2003 ( 
.A(n_1785),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1916),
.B(n_1290),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1722),
.Y(n_2005)
);

BUFx6f_ASAP7_75t_L g2006 ( 
.A(n_1700),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1726),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1735),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1736),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1916),
.B(n_1305),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1703),
.Y(n_2011)
);

BUFx6f_ASAP7_75t_L g2012 ( 
.A(n_1703),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1739),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1893),
.B(n_1316),
.Y(n_2014)
);

HB1xp67_ASAP7_75t_L g2015 ( 
.A(n_1791),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1747),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1748),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1865),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1753),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1754),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1758),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1765),
.Y(n_2022)
);

BUFx6f_ASAP7_75t_L g2023 ( 
.A(n_1703),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1694),
.B(n_1028),
.Y(n_2024)
);

BUFx3_ASAP7_75t_L g2025 ( 
.A(n_1690),
.Y(n_2025)
);

CKINVDCx8_ASAP7_75t_R g2026 ( 
.A(n_1872),
.Y(n_2026)
);

INVx1_ASAP7_75t_SL g2027 ( 
.A(n_1742),
.Y(n_2027)
);

AND2x2_ASAP7_75t_L g2028 ( 
.A(n_1782),
.B(n_1028),
.Y(n_2028)
);

CKINVDCx16_ASAP7_75t_R g2029 ( 
.A(n_1744),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1776),
.Y(n_2030)
);

BUFx2_ASAP7_75t_L g2031 ( 
.A(n_1759),
.Y(n_2031)
);

BUFx6f_ASAP7_75t_L g2032 ( 
.A(n_1728),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1778),
.Y(n_2033)
);

INVxp67_ASAP7_75t_L g2034 ( 
.A(n_1759),
.Y(n_2034)
);

BUFx6f_ASAP7_75t_L g2035 ( 
.A(n_1728),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1780),
.Y(n_2036)
);

INVx1_ASAP7_75t_L g2037 ( 
.A(n_1781),
.Y(n_2037)
);

HB1xp67_ASAP7_75t_L g2038 ( 
.A(n_1976),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1865),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1692),
.B(n_1318),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1790),
.Y(n_2041)
);

BUFx6f_ASAP7_75t_L g2042 ( 
.A(n_1728),
.Y(n_2042)
);

BUFx3_ASAP7_75t_L g2043 ( 
.A(n_1755),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1817),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_1794),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1817),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1803),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1823),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1809),
.Y(n_2049)
);

BUFx2_ASAP7_75t_L g2050 ( 
.A(n_1692),
.Y(n_2050)
);

OAI22xp5_ASAP7_75t_SL g2051 ( 
.A1(n_1769),
.A2(n_1483),
.B1(n_1492),
.B2(n_1453),
.Y(n_2051)
);

OA21x2_ASAP7_75t_L g2052 ( 
.A1(n_1705),
.A2(n_1206),
.B(n_1179),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1820),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1832),
.Y(n_2054)
);

HB1xp67_ASAP7_75t_L g2055 ( 
.A(n_1976),
.Y(n_2055)
);

BUFx6f_ASAP7_75t_L g2056 ( 
.A(n_1730),
.Y(n_2056)
);

INVx3_ASAP7_75t_L g2057 ( 
.A(n_1868),
.Y(n_2057)
);

OAI22xp5_ASAP7_75t_L g2058 ( 
.A1(n_1893),
.A2(n_932),
.B1(n_933),
.B2(n_931),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1834),
.Y(n_2059)
);

INVx3_ASAP7_75t_L g2060 ( 
.A(n_1906),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_1730),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1837),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1825),
.Y(n_2063)
);

AND2x6_ASAP7_75t_L g2064 ( 
.A(n_1849),
.B(n_1224),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1743),
.B(n_1320),
.Y(n_2065)
);

INVx2_ASAP7_75t_L g2066 ( 
.A(n_1847),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1915),
.B(n_1322),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1828),
.Y(n_2068)
);

INVx4_ASAP7_75t_L g2069 ( 
.A(n_1862),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1848),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1906),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1730),
.Y(n_2072)
);

BUFx6f_ASAP7_75t_L g2073 ( 
.A(n_1734),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1844),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1831),
.Y(n_2075)
);

OA21x2_ASAP7_75t_L g2076 ( 
.A1(n_1777),
.A2(n_1223),
.B(n_1206),
.Y(n_2076)
);

BUFx6f_ASAP7_75t_L g2077 ( 
.A(n_1734),
.Y(n_2077)
);

INVx1_ASAP7_75t_SL g2078 ( 
.A(n_1702),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1842),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1843),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1853),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_1874),
.Y(n_2082)
);

INVx4_ASAP7_75t_L g2083 ( 
.A(n_1862),
.Y(n_2083)
);

AND2x4_ASAP7_75t_L g2084 ( 
.A(n_1815),
.B(n_1283),
.Y(n_2084)
);

BUFx2_ASAP7_75t_L g2085 ( 
.A(n_1743),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1878),
.Y(n_2086)
);

OAI21x1_ASAP7_75t_L g2087 ( 
.A1(n_1718),
.A2(n_1256),
.B(n_1223),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1880),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1913),
.B(n_1360),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_1881),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1844),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_1796),
.Y(n_2092)
);

INVx2_ASAP7_75t_L g2093 ( 
.A(n_1796),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_1836),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1884),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1888),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_1890),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_1836),
.Y(n_2098)
);

BUFx3_ASAP7_75t_L g2099 ( 
.A(n_1770),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_1786),
.B(n_1028),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1892),
.Y(n_2101)
);

CKINVDCx5p33_ASAP7_75t_R g2102 ( 
.A(n_1784),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1907),
.B(n_1361),
.Y(n_2103)
);

CKINVDCx5p33_ASAP7_75t_R g2104 ( 
.A(n_1784),
.Y(n_2104)
);

INVx3_ASAP7_75t_L g2105 ( 
.A(n_1851),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1894),
.Y(n_2106)
);

BUFx2_ASAP7_75t_L g2107 ( 
.A(n_1757),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1852),
.Y(n_2108)
);

INVx1_ASAP7_75t_SL g2109 ( 
.A(n_1757),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1899),
.Y(n_2110)
);

OAI21x1_ASAP7_75t_L g2111 ( 
.A1(n_1718),
.A2(n_1265),
.B(n_1256),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1901),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1904),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_1870),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_1731),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1954),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_1954),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1857),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1870),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1857),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1787),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1873),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1792),
.B(n_1369),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1788),
.Y(n_2124)
);

BUFx6f_ASAP7_75t_L g2125 ( 
.A(n_1734),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_1697),
.A2(n_1274),
.B(n_1265),
.Y(n_2126)
);

INVx2_ASAP7_75t_L g2127 ( 
.A(n_1798),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1802),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1806),
.Y(n_2129)
);

INVx3_ASAP7_75t_L g2130 ( 
.A(n_1851),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1883),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1756),
.Y(n_2132)
);

INVx2_ASAP7_75t_L g2133 ( 
.A(n_1810),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1811),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_1756),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_1716),
.B(n_1370),
.Y(n_2136)
);

INVx3_ASAP7_75t_L g2137 ( 
.A(n_1851),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1821),
.Y(n_2138)
);

BUFx6f_ASAP7_75t_L g2139 ( 
.A(n_1756),
.Y(n_2139)
);

BUFx6f_ASAP7_75t_L g2140 ( 
.A(n_1779),
.Y(n_2140)
);

AND2x2_ASAP7_75t_L g2141 ( 
.A(n_1807),
.B(n_1373),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1701),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1704),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_1946),
.B(n_1374),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_1861),
.Y(n_2145)
);

BUFx6f_ASAP7_75t_L g2146 ( 
.A(n_1779),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1903),
.Y(n_2147)
);

NAND2xp33_ASAP7_75t_SL g2148 ( 
.A(n_1838),
.B(n_1380),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1706),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1907),
.B(n_934),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1907),
.B(n_936),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1905),
.Y(n_2152)
);

INVx2_ASAP7_75t_L g2153 ( 
.A(n_1708),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_1839),
.B(n_1480),
.Y(n_2154)
);

BUFx6f_ASAP7_75t_L g2155 ( 
.A(n_1779),
.Y(n_2155)
);

BUFx2_ASAP7_75t_L g2156 ( 
.A(n_1731),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1867),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1867),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1879),
.Y(n_2159)
);

HB1xp67_ASAP7_75t_L g2160 ( 
.A(n_1827),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1879),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1750),
.B(n_943),
.Y(n_2162)
);

BUFx2_ASAP7_75t_L g2163 ( 
.A(n_1827),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1850),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1850),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_1732),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_1833),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1740),
.Y(n_2168)
);

AND2x4_ASAP7_75t_L g2169 ( 
.A(n_1815),
.B(n_1225),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1869),
.Y(n_2170)
);

NAND2xp5_ASAP7_75t_L g2171 ( 
.A(n_1750),
.B(n_945),
.Y(n_2171)
);

INVx3_ASAP7_75t_L g2172 ( 
.A(n_1861),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1741),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1869),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1869),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1871),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1871),
.Y(n_2177)
);

INVx2_ASAP7_75t_L g2178 ( 
.A(n_1749),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_1871),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_1977),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1752),
.B(n_947),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_1760),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1875),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_1789),
.Y(n_2184)
);

AND2x6_ASAP7_75t_L g2185 ( 
.A(n_1698),
.B(n_1226),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1875),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_1789),
.Y(n_2187)
);

BUFx2_ASAP7_75t_L g2188 ( 
.A(n_1833),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_1773),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1752),
.B(n_948),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1861),
.Y(n_2191)
);

CKINVDCx8_ASAP7_75t_R g2192 ( 
.A(n_1872),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1866),
.Y(n_2193)
);

BUFx2_ASAP7_75t_L g2194 ( 
.A(n_1978),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1866),
.Y(n_2195)
);

INVx4_ASAP7_75t_L g2196 ( 
.A(n_1862),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1875),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1866),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_1845),
.B(n_1228),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_1876),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_1966),
.Y(n_2201)
);

OA21x2_ASAP7_75t_L g2202 ( 
.A1(n_1725),
.A2(n_1274),
.B(n_1230),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_1876),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_1876),
.B(n_961),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1895),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1966),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_1895),
.Y(n_2207)
);

BUFx6f_ASAP7_75t_L g2208 ( 
.A(n_1789),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_1800),
.Y(n_2209)
);

AOI22xp5_ASAP7_75t_L g2210 ( 
.A1(n_1815),
.A2(n_1829),
.B1(n_1877),
.B2(n_1862),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_SL g2211 ( 
.A(n_1946),
.B(n_694),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1895),
.B(n_963),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1804),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1896),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1896),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1896),
.Y(n_2216)
);

INVx3_ASAP7_75t_L g2217 ( 
.A(n_1862),
.Y(n_2217)
);

HB1xp67_ASAP7_75t_L g2218 ( 
.A(n_1872),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1891),
.Y(n_2219)
);

BUFx6f_ASAP7_75t_L g2220 ( 
.A(n_1804),
.Y(n_2220)
);

INVx3_ASAP7_75t_L g2221 ( 
.A(n_1804),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1891),
.Y(n_2222)
);

OAI21x1_ASAP7_75t_L g2223 ( 
.A1(n_1697),
.A2(n_1232),
.B(n_1229),
.Y(n_2223)
);

NAND2x1p5_ASAP7_75t_L g2224 ( 
.A(n_1958),
.B(n_1235),
.Y(n_2224)
);

AND2x4_ASAP7_75t_L g2225 ( 
.A(n_1815),
.B(n_1240),
.Y(n_2225)
);

INVx1_ASAP7_75t_SL g2226 ( 
.A(n_1819),
.Y(n_2226)
);

NAND2x1p5_ASAP7_75t_L g2227 ( 
.A(n_1958),
.B(n_1247),
.Y(n_2227)
);

INVx3_ASAP7_75t_L g2228 ( 
.A(n_1797),
.Y(n_2228)
);

XOR2xp5_ASAP7_75t_L g2229 ( 
.A(n_1818),
.B(n_1492),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1800),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1797),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_SL g2232 ( 
.A(n_1958),
.B(n_694),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1891),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1725),
.A2(n_1259),
.B(n_1255),
.Y(n_2234)
);

NOR2x1_ASAP7_75t_L g2235 ( 
.A(n_1838),
.B(n_1260),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1793),
.B(n_965),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1840),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_1797),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1856),
.Y(n_2239)
);

INVx3_ASAP7_75t_L g2240 ( 
.A(n_1822),
.Y(n_2240)
);

HB1xp67_ASAP7_75t_L g2241 ( 
.A(n_1872),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1856),
.Y(n_2242)
);

INVx3_ASAP7_75t_L g2243 ( 
.A(n_1822),
.Y(n_2243)
);

INVx2_ASAP7_75t_L g2244 ( 
.A(n_1840),
.Y(n_2244)
);

BUFx3_ASAP7_75t_L g2245 ( 
.A(n_1931),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_1824),
.B(n_1262),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_1795),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_1772),
.Y(n_2248)
);

NAND2xp33_ASAP7_75t_SL g2249 ( 
.A(n_1919),
.B(n_969),
.Y(n_2249)
);

CKINVDCx16_ASAP7_75t_R g2250 ( 
.A(n_1814),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_1886),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_1886),
.Y(n_2252)
);

AND2x2_ASAP7_75t_L g2253 ( 
.A(n_1953),
.B(n_1882),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1887),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1793),
.B(n_974),
.Y(n_2255)
);

NAND2xp5_ASAP7_75t_L g2256 ( 
.A(n_1918),
.B(n_1933),
.Y(n_2256)
);

NAND2x1_ASAP7_75t_L g2257 ( 
.A(n_1733),
.B(n_1239),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1772),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1887),
.Y(n_2259)
);

INVx1_ASAP7_75t_SL g2260 ( 
.A(n_1846),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1816),
.Y(n_2261)
);

BUFx2_ASAP7_75t_L g2262 ( 
.A(n_1814),
.Y(n_2262)
);

INVx3_ASAP7_75t_L g2263 ( 
.A(n_1822),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1816),
.Y(n_2264)
);

OA21x2_ASAP7_75t_L g2265 ( 
.A1(n_1729),
.A2(n_1751),
.B(n_1774),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1858),
.Y(n_2266)
);

INVx3_ASAP7_75t_L g2267 ( 
.A(n_1822),
.Y(n_2267)
);

BUFx8_ASAP7_75t_L g2268 ( 
.A(n_1859),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1858),
.Y(n_2269)
);

INVx2_ASAP7_75t_L g2270 ( 
.A(n_1774),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_1918),
.B(n_975),
.Y(n_2271)
);

INVx2_ASAP7_75t_L g2272 ( 
.A(n_1729),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_1900),
.B(n_1279),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1885),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1885),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_1751),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_1767),
.Y(n_2277)
);

INVx2_ASAP7_75t_L g2278 ( 
.A(n_1767),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1855),
.Y(n_2279)
);

BUFx6f_ASAP7_75t_L g2280 ( 
.A(n_1693),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1712),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1712),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_1717),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_SL g2284 ( 
.A(n_1958),
.B(n_694),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_1908),
.B(n_1287),
.Y(n_2285)
);

AND2x2_ASAP7_75t_L g2286 ( 
.A(n_1928),
.B(n_1289),
.Y(n_2286)
);

AOI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_1815),
.A2(n_1000),
.B1(n_988),
.B2(n_977),
.Y(n_2287)
);

BUFx6f_ASAP7_75t_L g2288 ( 
.A(n_1693),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_1717),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1933),
.B(n_979),
.Y(n_2290)
);

INVx1_ASAP7_75t_SL g2291 ( 
.A(n_1889),
.Y(n_2291)
);

AND2x2_ASAP7_75t_SL g2292 ( 
.A(n_1829),
.B(n_1293),
.Y(n_2292)
);

BUFx2_ASAP7_75t_L g2293 ( 
.A(n_1727),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_1721),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1855),
.Y(n_2295)
);

INVx1_ASAP7_75t_SL g2296 ( 
.A(n_1902),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_1955),
.B(n_1294),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_1721),
.Y(n_2298)
);

INVx2_ASAP7_75t_L g2299 ( 
.A(n_1855),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_2092),
.Y(n_2300)
);

BUFx4f_ASAP7_75t_L g2301 ( 
.A(n_2005),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2272),
.B(n_1955),
.Y(n_2302)
);

BUFx4f_ASAP7_75t_L g2303 ( 
.A(n_2262),
.Y(n_2303)
);

INVxp67_ASAP7_75t_SL g2304 ( 
.A(n_2074),
.Y(n_2304)
);

INVx2_ASAP7_75t_L g2305 ( 
.A(n_2092),
.Y(n_2305)
);

INVx2_ASAP7_75t_SL g2306 ( 
.A(n_2027),
.Y(n_2306)
);

BUFx10_ASAP7_75t_L g2307 ( 
.A(n_2102),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2272),
.B(n_1691),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2093),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2276),
.B(n_1691),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_1979),
.Y(n_2311)
);

INVx2_ASAP7_75t_L g2312 ( 
.A(n_2093),
.Y(n_2312)
);

NOR2xp33_ASAP7_75t_L g2313 ( 
.A(n_1997),
.B(n_1764),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1984),
.Y(n_2314)
);

INVxp33_ASAP7_75t_L g2315 ( 
.A(n_1989),
.Y(n_2315)
);

BUFx8_ASAP7_75t_SL g2316 ( 
.A(n_2102),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1986),
.Y(n_2317)
);

BUFx3_ASAP7_75t_L g2318 ( 
.A(n_2025),
.Y(n_2318)
);

INVx3_ASAP7_75t_L g2319 ( 
.A(n_2069),
.Y(n_2319)
);

NOR2xp33_ASAP7_75t_L g2320 ( 
.A(n_2001),
.B(n_1923),
.Y(n_2320)
);

INVx2_ASAP7_75t_L g2321 ( 
.A(n_2094),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2239),
.A2(n_1715),
.B1(n_1769),
.B2(n_1898),
.Y(n_2322)
);

INVx4_ASAP7_75t_L g2323 ( 
.A(n_2025),
.Y(n_2323)
);

BUFx3_ASAP7_75t_L g2324 ( 
.A(n_2043),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_2094),
.Y(n_2325)
);

AOI22xp5_ASAP7_75t_L g2326 ( 
.A1(n_2067),
.A2(n_2014),
.B1(n_2253),
.B2(n_2185),
.Y(n_2326)
);

INVx2_ASAP7_75t_L g2327 ( 
.A(n_2098),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_1983),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_1992),
.Y(n_2329)
);

INVx1_ASAP7_75t_SL g2330 ( 
.A(n_2078),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_2098),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_2276),
.B(n_1768),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_1995),
.Y(n_2333)
);

HB1xp67_ASAP7_75t_L g2334 ( 
.A(n_2031),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1999),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_2118),
.Y(n_2336)
);

AOI22xp33_ASAP7_75t_L g2337 ( 
.A1(n_2242),
.A2(n_1715),
.B1(n_1898),
.B2(n_1738),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2118),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2120),
.Y(n_2339)
);

INVx3_ASAP7_75t_L g2340 ( 
.A(n_2069),
.Y(n_2340)
);

INVx2_ASAP7_75t_SL g2341 ( 
.A(n_2260),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_SL g2342 ( 
.A(n_1990),
.B(n_1919),
.Y(n_2342)
);

INVx1_ASAP7_75t_L g2343 ( 
.A(n_2000),
.Y(n_2343)
);

NOR2xp33_ASAP7_75t_SL g2344 ( 
.A(n_2069),
.B(n_2083),
.Y(n_2344)
);

NOR2xp33_ASAP7_75t_L g2345 ( 
.A(n_2004),
.B(n_1923),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2002),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2007),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2008),
.Y(n_2348)
);

OAI22xp33_ASAP7_75t_L g2349 ( 
.A1(n_2210),
.A2(n_1877),
.B1(n_1926),
.B2(n_1944),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_2278),
.B(n_1768),
.Y(n_2350)
);

INVx3_ASAP7_75t_L g2351 ( 
.A(n_2083),
.Y(n_2351)
);

INVx5_ASAP7_75t_L g2352 ( 
.A(n_2083),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2009),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2043),
.B(n_1919),
.Y(n_2354)
);

BUFx6f_ASAP7_75t_L g2355 ( 
.A(n_1983),
.Y(n_2355)
);

OAI22xp5_ASAP7_75t_L g2356 ( 
.A1(n_2277),
.A2(n_1944),
.B1(n_1968),
.B2(n_1961),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2010),
.B(n_2226),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_1983),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2067),
.B(n_1937),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_2013),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_2120),
.Y(n_2361)
);

OR2x2_ASAP7_75t_L g2362 ( 
.A(n_2109),
.B(n_1897),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2016),
.Y(n_2363)
);

INVx3_ASAP7_75t_L g2364 ( 
.A(n_2196),
.Y(n_2364)
);

INVx2_ASAP7_75t_L g2365 ( 
.A(n_2108),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2099),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2278),
.B(n_1746),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2108),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2017),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_2048),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2019),
.Y(n_2371)
);

OAI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2162),
.A2(n_1968),
.B1(n_1961),
.B2(n_1818),
.Y(n_2372)
);

NOR2x1p5_ASAP7_75t_L g2373 ( 
.A(n_2104),
.B(n_1835),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2050),
.B(n_1945),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2020),
.Y(n_2375)
);

INVx3_ASAP7_75t_L g2376 ( 
.A(n_2196),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2048),
.Y(n_2377)
);

OAI22xp5_ASAP7_75t_L g2378 ( 
.A1(n_2171),
.A2(n_1835),
.B1(n_1941),
.B2(n_1939),
.Y(n_2378)
);

BUFx4f_ASAP7_75t_L g2379 ( 
.A(n_2185),
.Y(n_2379)
);

XNOR2x1_ASAP7_75t_L g2380 ( 
.A(n_2229),
.B(n_1738),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_1983),
.Y(n_2381)
);

INVx2_ASAP7_75t_L g2382 ( 
.A(n_2054),
.Y(n_2382)
);

OR2x2_ASAP7_75t_L g2383 ( 
.A(n_2156),
.B(n_2163),
.Y(n_2383)
);

INVx3_ASAP7_75t_L g2384 ( 
.A(n_2196),
.Y(n_2384)
);

INVx4_ASAP7_75t_L g2385 ( 
.A(n_2099),
.Y(n_2385)
);

OR2x2_ASAP7_75t_L g2386 ( 
.A(n_2188),
.B(n_1897),
.Y(n_2386)
);

INVxp67_ASAP7_75t_SL g2387 ( 
.A(n_2074),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2280),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2021),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2024),
.B(n_1912),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2022),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_2054),
.Y(n_2392)
);

NOR2xp33_ASAP7_75t_L g2393 ( 
.A(n_2089),
.B(n_1949),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_SL g2394 ( 
.A(n_2085),
.B(n_1929),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2059),
.Y(n_2395)
);

INVx3_ASAP7_75t_L g2396 ( 
.A(n_2280),
.Y(n_2396)
);

INVx2_ASAP7_75t_L g2397 ( 
.A(n_2059),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2030),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2062),
.Y(n_2399)
);

INVxp67_ASAP7_75t_SL g2400 ( 
.A(n_2091),
.Y(n_2400)
);

AOI22xp5_ASAP7_75t_L g2401 ( 
.A1(n_2185),
.A2(n_2136),
.B1(n_2297),
.B2(n_1993),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2033),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2157),
.B(n_1746),
.Y(n_2403)
);

NAND3xp33_ASAP7_75t_L g2404 ( 
.A(n_2034),
.B(n_1720),
.C(n_1917),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_SL g2405 ( 
.A(n_2291),
.B(n_1929),
.Y(n_2405)
);

INVx2_ASAP7_75t_SL g2406 ( 
.A(n_2296),
.Y(n_2406)
);

NOR3xp33_ASAP7_75t_L g2407 ( 
.A(n_1993),
.B(n_1720),
.C(n_1967),
.Y(n_2407)
);

INVx1_ASAP7_75t_SL g2408 ( 
.A(n_2180),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2036),
.Y(n_2409)
);

AOI22xp5_ASAP7_75t_L g2410 ( 
.A1(n_2185),
.A2(n_1920),
.B1(n_1921),
.B2(n_1783),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2037),
.Y(n_2411)
);

BUFx3_ASAP7_75t_L g2412 ( 
.A(n_2245),
.Y(n_2412)
);

OAI22xp33_ASAP7_75t_L g2413 ( 
.A1(n_2181),
.A2(n_1926),
.B1(n_1940),
.B2(n_1929),
.Y(n_2413)
);

INVx2_ASAP7_75t_L g2414 ( 
.A(n_2062),
.Y(n_2414)
);

XOR2xp5_ASAP7_75t_L g2415 ( 
.A(n_2104),
.B(n_1493),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2041),
.Y(n_2416)
);

BUFx6f_ASAP7_75t_L g2417 ( 
.A(n_1988),
.Y(n_2417)
);

INVx1_ASAP7_75t_SL g2418 ( 
.A(n_2154),
.Y(n_2418)
);

INVx4_ASAP7_75t_L g2419 ( 
.A(n_2245),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2045),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2158),
.B(n_1762),
.Y(n_2421)
);

CKINVDCx5p33_ASAP7_75t_R g2422 ( 
.A(n_2250),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_L g2423 ( 
.A(n_2058),
.B(n_1950),
.C(n_1947),
.Y(n_2423)
);

NAND2xp33_ASAP7_75t_L g2424 ( 
.A(n_2148),
.B(n_1940),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2159),
.B(n_1762),
.Y(n_2425)
);

NAND2xp33_ASAP7_75t_R g2426 ( 
.A(n_2293),
.B(n_1967),
.Y(n_2426)
);

INVxp67_ASAP7_75t_L g2427 ( 
.A(n_2115),
.Y(n_2427)
);

AND2x6_ASAP7_75t_L g2428 ( 
.A(n_2217),
.B(n_1952),
.Y(n_2428)
);

NAND2xp33_ASAP7_75t_L g2429 ( 
.A(n_2148),
.B(n_1940),
.Y(n_2429)
);

BUFx3_ASAP7_75t_L g2430 ( 
.A(n_2003),
.Y(n_2430)
);

BUFx2_ASAP7_75t_L g2431 ( 
.A(n_2107),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2066),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_SL g2433 ( 
.A(n_2123),
.B(n_1945),
.Y(n_2433)
);

OR2x6_ASAP7_75t_L g2434 ( 
.A(n_2194),
.B(n_1945),
.Y(n_2434)
);

AND2x6_ASAP7_75t_L g2435 ( 
.A(n_2217),
.B(n_1952),
.Y(n_2435)
);

BUFx3_ASAP7_75t_L g2436 ( 
.A(n_2003),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_SL g2437 ( 
.A(n_2141),
.B(n_1952),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2161),
.B(n_2248),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2047),
.Y(n_2439)
);

INVx2_ASAP7_75t_SL g2440 ( 
.A(n_2003),
.Y(n_2440)
);

AOI22xp33_ASAP7_75t_L g2441 ( 
.A1(n_2292),
.A2(n_1813),
.B1(n_1863),
.B2(n_1771),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2049),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2053),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2063),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_2248),
.B(n_2258),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_L g2446 ( 
.A(n_2015),
.B(n_1959),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2068),
.Y(n_2447)
);

INVx4_ASAP7_75t_L g2448 ( 
.A(n_2217),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2015),
.B(n_1960),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_SL g2450 ( 
.A(n_2040),
.B(n_1965),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2075),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2079),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2066),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2080),
.Y(n_2454)
);

AND2x2_ASAP7_75t_L g2455 ( 
.A(n_2024),
.B(n_1943),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_2280),
.Y(n_2456)
);

BUFx8_ASAP7_75t_SL g2457 ( 
.A(n_2065),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2081),
.Y(n_2458)
);

AOI22xp33_ASAP7_75t_L g2459 ( 
.A1(n_2292),
.A2(n_1813),
.B1(n_1771),
.B2(n_1775),
.Y(n_2459)
);

INVx1_ASAP7_75t_L g2460 ( 
.A(n_2082),
.Y(n_2460)
);

INVxp67_ASAP7_75t_L g2461 ( 
.A(n_2115),
.Y(n_2461)
);

AOI22xp33_ASAP7_75t_L g2462 ( 
.A1(n_2209),
.A2(n_2230),
.B1(n_2244),
.B2(n_2237),
.Y(n_2462)
);

AOI22xp33_ASAP7_75t_SL g2463 ( 
.A1(n_2051),
.A2(n_1841),
.B1(n_1493),
.B2(n_1496),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2070),
.Y(n_2464)
);

INVx2_ASAP7_75t_L g2465 ( 
.A(n_2070),
.Y(n_2465)
);

INVx2_ASAP7_75t_L g2466 ( 
.A(n_2121),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2086),
.Y(n_2467)
);

CKINVDCx16_ASAP7_75t_R g2468 ( 
.A(n_1998),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2121),
.Y(n_2469)
);

INVx2_ASAP7_75t_L g2470 ( 
.A(n_2124),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2258),
.B(n_1910),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_2088),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_L g2473 ( 
.A(n_2160),
.B(n_1932),
.C(n_1860),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2090),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_L g2475 ( 
.A(n_2270),
.B(n_1910),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2095),
.Y(n_2476)
);

INVx2_ASAP7_75t_L g2477 ( 
.A(n_2124),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2028),
.B(n_1938),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2268),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_SL g2480 ( 
.A(n_2103),
.B(n_1965),
.Y(n_2480)
);

BUFx6f_ASAP7_75t_L g2481 ( 
.A(n_1988),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2028),
.B(n_1938),
.Y(n_2482)
);

INVx4_ASAP7_75t_L g2483 ( 
.A(n_2231),
.Y(n_2483)
);

INVx4_ASAP7_75t_L g2484 ( 
.A(n_2231),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2029),
.B(n_1864),
.Y(n_2485)
);

INVx2_ASAP7_75t_L g2486 ( 
.A(n_2127),
.Y(n_2486)
);

AOI22xp5_ASAP7_75t_L g2487 ( 
.A1(n_2185),
.A2(n_1860),
.B1(n_1854),
.B2(n_1932),
.Y(n_2487)
);

INVx4_ASAP7_75t_L g2488 ( 
.A(n_2231),
.Y(n_2488)
);

AOI22xp33_ASAP7_75t_L g2489 ( 
.A1(n_2209),
.A2(n_1775),
.B1(n_1974),
.B2(n_1808),
.Y(n_2489)
);

AOI22xp5_ASAP7_75t_L g2490 ( 
.A1(n_2136),
.A2(n_1854),
.B1(n_1971),
.B2(n_1963),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2127),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_SL g2492 ( 
.A(n_2297),
.B(n_1965),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_1991),
.B(n_1956),
.Y(n_2493)
);

INVx4_ASAP7_75t_L g2494 ( 
.A(n_2231),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2128),
.Y(n_2495)
);

OR2x6_ASAP7_75t_L g2496 ( 
.A(n_2256),
.B(n_1972),
.Y(n_2496)
);

INVx1_ASAP7_75t_SL g2497 ( 
.A(n_2160),
.Y(n_2497)
);

BUFx3_ASAP7_75t_L g2498 ( 
.A(n_2268),
.Y(n_2498)
);

BUFx2_ASAP7_75t_L g2499 ( 
.A(n_2167),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2096),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2097),
.Y(n_2501)
);

OR2x6_ASAP7_75t_L g2502 ( 
.A(n_2261),
.B(n_1972),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2101),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_2026),
.B(n_1972),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2106),
.Y(n_2505)
);

OAI22xp33_ASAP7_75t_L g2506 ( 
.A1(n_2190),
.A2(n_2165),
.B1(n_2164),
.B2(n_2264),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2110),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_2268),
.Y(n_2508)
);

AOI22xp33_ASAP7_75t_L g2509 ( 
.A1(n_2230),
.A2(n_1974),
.B1(n_1808),
.B2(n_1936),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_SL g2510 ( 
.A(n_2026),
.B(n_1970),
.Y(n_2510)
);

INVx2_ASAP7_75t_L g2511 ( 
.A(n_2128),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_SL g2512 ( 
.A(n_2192),
.B(n_1970),
.Y(n_2512)
);

CKINVDCx20_ASAP7_75t_R g2513 ( 
.A(n_2247),
.Y(n_2513)
);

NOR2xp33_ASAP7_75t_L g2514 ( 
.A(n_1991),
.B(n_1956),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2112),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2113),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_2192),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2270),
.B(n_1761),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2122),
.Y(n_2519)
);

NOR2xp33_ASAP7_75t_L g2520 ( 
.A(n_1980),
.B(n_1942),
.Y(n_2520)
);

INVx2_ASAP7_75t_L g2521 ( 
.A(n_2129),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2129),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2280),
.Y(n_2523)
);

OR2x6_ASAP7_75t_L g2524 ( 
.A(n_2266),
.B(n_1805),
.Y(n_2524)
);

INVx1_ASAP7_75t_L g2525 ( 
.A(n_2131),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2100),
.B(n_1942),
.Y(n_2526)
);

OR2x6_ASAP7_75t_L g2527 ( 
.A(n_2269),
.B(n_1805),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_1988),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2237),
.B(n_1710),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2147),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_L g2531 ( 
.A(n_1980),
.B(n_1924),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_2100),
.A2(n_1973),
.B1(n_1975),
.B2(n_1962),
.Y(n_2532)
);

AND2x2_ASAP7_75t_L g2533 ( 
.A(n_2167),
.B(n_1841),
.Y(n_2533)
);

BUFx6f_ASAP7_75t_L g2534 ( 
.A(n_1988),
.Y(n_2534)
);

NOR2xp33_ASAP7_75t_L g2535 ( 
.A(n_2281),
.B(n_1927),
.Y(n_2535)
);

INVx3_ASAP7_75t_L g2536 ( 
.A(n_2288),
.Y(n_2536)
);

CKINVDCx16_ASAP7_75t_R g2537 ( 
.A(n_2249),
.Y(n_2537)
);

OR2x6_ASAP7_75t_L g2538 ( 
.A(n_2274),
.B(n_1805),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2244),
.A2(n_2282),
.B1(n_2289),
.B2(n_2283),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2133),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2152),
.Y(n_2541)
);

BUFx2_ASAP7_75t_L g2542 ( 
.A(n_2038),
.Y(n_2542)
);

AOI22xp33_ASAP7_75t_L g2543 ( 
.A1(n_2294),
.A2(n_1936),
.B1(n_1948),
.B2(n_1801),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2133),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2134),
.Y(n_2545)
);

NAND2xp5_ASAP7_75t_L g2546 ( 
.A(n_2265),
.B(n_1911),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2134),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2265),
.B(n_1914),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_2084),
.B(n_1801),
.Y(n_2549)
);

INVx5_ASAP7_75t_L g2550 ( 
.A(n_2288),
.Y(n_2550)
);

INVx2_ASAP7_75t_SL g2551 ( 
.A(n_2273),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2138),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2138),
.Y(n_2553)
);

INVx2_ASAP7_75t_L g2554 ( 
.A(n_2142),
.Y(n_2554)
);

INVx3_ASAP7_75t_L g2555 ( 
.A(n_2288),
.Y(n_2555)
);

BUFx3_ASAP7_75t_L g2556 ( 
.A(n_2285),
.Y(n_2556)
);

OR2x2_ASAP7_75t_L g2557 ( 
.A(n_2286),
.B(n_1964),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2142),
.Y(n_2558)
);

INVx1_ASAP7_75t_SL g2559 ( 
.A(n_2084),
.Y(n_2559)
);

INVx2_ASAP7_75t_SL g2560 ( 
.A(n_2199),
.Y(n_2560)
);

CKINVDCx5p33_ASAP7_75t_R g2561 ( 
.A(n_2218),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2143),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2143),
.Y(n_2563)
);

OR2x6_ASAP7_75t_L g2564 ( 
.A(n_2275),
.B(n_1969),
.Y(n_2564)
);

BUFx6f_ASAP7_75t_L g2565 ( 
.A(n_2006),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2246),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2149),
.Y(n_2567)
);

INVx3_ASAP7_75t_L g2568 ( 
.A(n_2288),
.Y(n_2568)
);

AO21x2_ASAP7_75t_L g2569 ( 
.A1(n_2116),
.A2(n_1925),
.B(n_1935),
.Y(n_2569)
);

OAI22xp33_ASAP7_75t_SL g2570 ( 
.A1(n_2144),
.A2(n_1964),
.B1(n_1925),
.B2(n_1935),
.Y(n_2570)
);

INVx4_ASAP7_75t_L g2571 ( 
.A(n_2084),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_L g2572 ( 
.A1(n_2298),
.A2(n_1936),
.B1(n_1934),
.B2(n_1930),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2149),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2265),
.B(n_1936),
.Y(n_2574)
);

BUFx10_ASAP7_75t_L g2575 ( 
.A(n_2169),
.Y(n_2575)
);

AND2x6_ASAP7_75t_L g2576 ( 
.A(n_2091),
.B(n_1951),
.Y(n_2576)
);

XNOR2xp5_ASAP7_75t_L g2577 ( 
.A(n_2218),
.B(n_1494),
.Y(n_2577)
);

INVx4_ASAP7_75t_L g2578 ( 
.A(n_2006),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2153),
.Y(n_2579)
);

INVxp67_ASAP7_75t_SL g2580 ( 
.A(n_2071),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2153),
.Y(n_2581)
);

NAND3xp33_ASAP7_75t_L g2582 ( 
.A(n_2150),
.B(n_1727),
.C(n_1826),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2166),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_SL g2584 ( 
.A(n_2287),
.B(n_1957),
.Y(n_2584)
);

BUFx4f_ASAP7_75t_L g2585 ( 
.A(n_2064),
.Y(n_2585)
);

BUFx2_ASAP7_75t_L g2586 ( 
.A(n_2038),
.Y(n_2586)
);

NOR3xp33_ASAP7_75t_L g2587 ( 
.A(n_2144),
.B(n_1766),
.C(n_1745),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2166),
.Y(n_2588)
);

BUFx2_ASAP7_75t_L g2589 ( 
.A(n_2055),
.Y(n_2589)
);

INVx2_ASAP7_75t_L g2590 ( 
.A(n_2168),
.Y(n_2590)
);

AND2x6_ASAP7_75t_L g2591 ( 
.A(n_2169),
.B(n_1936),
.Y(n_2591)
);

NAND2xp33_ASAP7_75t_L g2592 ( 
.A(n_2224),
.B(n_982),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2055),
.B(n_1494),
.Y(n_2593)
);

INVx5_ASAP7_75t_L g2594 ( 
.A(n_2006),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2168),
.Y(n_2595)
);

NAND2xp5_ASAP7_75t_L g2596 ( 
.A(n_2114),
.B(n_1733),
.Y(n_2596)
);

NAND3xp33_ASAP7_75t_L g2597 ( 
.A(n_2151),
.B(n_1826),
.C(n_1766),
.Y(n_2597)
);

HB1xp67_ASAP7_75t_L g2598 ( 
.A(n_2169),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2241),
.Y(n_2599)
);

AOI21x1_ASAP7_75t_L g2600 ( 
.A1(n_2232),
.A2(n_1296),
.B(n_1295),
.Y(n_2600)
);

INVx3_ASAP7_75t_L g2601 ( 
.A(n_2006),
.Y(n_2601)
);

NOR2xp33_ASAP7_75t_L g2602 ( 
.A(n_2119),
.B(n_1733),
.Y(n_2602)
);

INVx5_ASAP7_75t_L g2603 ( 
.A(n_2011),
.Y(n_2603)
);

AND2x2_ASAP7_75t_SL g2604 ( 
.A(n_2241),
.B(n_1724),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2011),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2173),
.Y(n_2606)
);

INVx1_ASAP7_75t_SL g2607 ( 
.A(n_2225),
.Y(n_2607)
);

INVx3_ASAP7_75t_L g2608 ( 
.A(n_2011),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2011),
.Y(n_2609)
);

NAND2xp33_ASAP7_75t_L g2610 ( 
.A(n_2224),
.B(n_987),
.Y(n_2610)
);

BUFx6f_ASAP7_75t_L g2611 ( 
.A(n_2012),
.Y(n_2611)
);

CKINVDCx20_ASAP7_75t_R g2612 ( 
.A(n_2249),
.Y(n_2612)
);

INVxp33_ASAP7_75t_L g2613 ( 
.A(n_2271),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2173),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2178),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_L g2616 ( 
.A(n_2064),
.B(n_2225),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2211),
.B(n_990),
.Y(n_2617)
);

AND2x4_ASAP7_75t_L g2618 ( 
.A(n_2251),
.B(n_2252),
.Y(n_2618)
);

NAND2xp33_ASAP7_75t_L g2619 ( 
.A(n_2227),
.B(n_992),
.Y(n_2619)
);

INVx4_ASAP7_75t_L g2620 ( 
.A(n_2012),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2254),
.B(n_1496),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_SL g2622 ( 
.A(n_2225),
.B(n_1693),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2178),
.Y(n_2623)
);

INVx3_ASAP7_75t_L g2624 ( 
.A(n_2012),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2182),
.Y(n_2625)
);

INVx2_ASAP7_75t_SL g2626 ( 
.A(n_2235),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_L g2627 ( 
.A(n_2211),
.B(n_993),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2182),
.Y(n_2628)
);

BUFx3_ASAP7_75t_L g2629 ( 
.A(n_2259),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2189),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2219),
.B(n_2222),
.Y(n_2631)
);

INVx5_ASAP7_75t_L g2632 ( 
.A(n_2012),
.Y(n_2632)
);

BUFx6f_ASAP7_75t_L g2633 ( 
.A(n_2023),
.Y(n_2633)
);

INVx3_ASAP7_75t_L g2634 ( 
.A(n_2023),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_SL g2635 ( 
.A(n_2233),
.B(n_2236),
.Y(n_2635)
);

BUFx2_ASAP7_75t_L g2636 ( 
.A(n_2064),
.Y(n_2636)
);

NOR2xp33_ASAP7_75t_L g2637 ( 
.A(n_2290),
.B(n_999),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2189),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2044),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_2255),
.B(n_1693),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2170),
.Y(n_2641)
);

BUFx2_ASAP7_75t_L g2642 ( 
.A(n_2064),
.Y(n_2642)
);

INVx5_ASAP7_75t_L g2643 ( 
.A(n_2023),
.Y(n_2643)
);

INVx8_ASAP7_75t_L g2644 ( 
.A(n_2064),
.Y(n_2644)
);

NOR2xp33_ASAP7_75t_L g2645 ( 
.A(n_2204),
.B(n_1504),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2174),
.Y(n_2646)
);

CKINVDCx5p33_ASAP7_75t_R g2647 ( 
.A(n_2212),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2044),
.Y(n_2648)
);

INVx2_ASAP7_75t_SL g2649 ( 
.A(n_2257),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2175),
.A2(n_1002),
.B1(n_1013),
.B2(n_1007),
.Y(n_2650)
);

INVx4_ASAP7_75t_L g2651 ( 
.A(n_2023),
.Y(n_2651)
);

NOR2xp33_ASAP7_75t_L g2652 ( 
.A(n_2176),
.B(n_1015),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2177),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2179),
.Y(n_2654)
);

BUFx6f_ASAP7_75t_L g2655 ( 
.A(n_2594),
.Y(n_2655)
);

INVx3_ASAP7_75t_L g2656 ( 
.A(n_2448),
.Y(n_2656)
);

NAND2xp5_ASAP7_75t_L g2657 ( 
.A(n_2359),
.B(n_2205),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2359),
.B(n_2183),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2311),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_L g2660 ( 
.A(n_2315),
.B(n_1504),
.Y(n_2660)
);

NOR2xp33_ASAP7_75t_L g2661 ( 
.A(n_2320),
.B(n_1510),
.Y(n_2661)
);

NAND3xp33_ASAP7_75t_L g2662 ( 
.A(n_2372),
.B(n_1745),
.C(n_2186),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2357),
.B(n_2200),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2314),
.Y(n_2664)
);

NOR3xp33_ASAP7_75t_L g2665 ( 
.A(n_2372),
.B(n_2284),
.C(n_2232),
.Y(n_2665)
);

BUFx6f_ASAP7_75t_L g2666 ( 
.A(n_2594),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2317),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2329),
.Y(n_2668)
);

NAND2x1p5_ASAP7_75t_L g2669 ( 
.A(n_2323),
.B(n_2197),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2594),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2333),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_SL g2672 ( 
.A(n_2301),
.B(n_2203),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_L g2673 ( 
.A(n_2357),
.B(n_2207),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2335),
.Y(n_2674)
);

INVxp67_ASAP7_75t_SL g2675 ( 
.A(n_2304),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2466),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2302),
.B(n_2214),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_2302),
.B(n_2215),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2343),
.Y(n_2679)
);

INVx4_ASAP7_75t_L g2680 ( 
.A(n_2422),
.Y(n_2680)
);

NOR3xp33_ASAP7_75t_L g2681 ( 
.A(n_2356),
.B(n_2284),
.C(n_1017),
.Y(n_2681)
);

CKINVDCx5p33_ASAP7_75t_R g2682 ( 
.A(n_2316),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2320),
.B(n_2216),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2390),
.B(n_1510),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_SL g2685 ( 
.A(n_2301),
.B(n_2227),
.Y(n_2685)
);

NAND2xp5_ASAP7_75t_L g2686 ( 
.A(n_2313),
.B(n_2345),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2346),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2469),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2470),
.Y(n_2689)
);

XOR2xp5_ASAP7_75t_L g2690 ( 
.A(n_2415),
.B(n_1513),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2347),
.Y(n_2691)
);

NAND3xp33_ASAP7_75t_L g2692 ( 
.A(n_2326),
.B(n_1515),
.C(n_1513),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_SL g2693 ( 
.A(n_2413),
.B(n_2032),
.Y(n_2693)
);

NAND2xp33_ASAP7_75t_SL g2694 ( 
.A(n_2378),
.B(n_2032),
.Y(n_2694)
);

NOR2xp33_ASAP7_75t_R g2695 ( 
.A(n_2517),
.B(n_1515),
.Y(n_2695)
);

HB1xp67_ASAP7_75t_L g2696 ( 
.A(n_2334),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2348),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2533),
.B(n_1519),
.Y(n_2698)
);

NOR3xp33_ASAP7_75t_L g2699 ( 
.A(n_2356),
.B(n_1016),
.C(n_2228),
.Y(n_2699)
);

INVx8_ASAP7_75t_L g2700 ( 
.A(n_2434),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2313),
.B(n_2105),
.Y(n_2701)
);

NAND2xp5_ASAP7_75t_L g2702 ( 
.A(n_2345),
.B(n_2105),
.Y(n_2702)
);

NOR3xp33_ASAP7_75t_L g2703 ( 
.A(n_2413),
.B(n_2238),
.C(n_2228),
.Y(n_2703)
);

NOR2xp33_ASAP7_75t_L g2704 ( 
.A(n_2393),
.B(n_1519),
.Y(n_2704)
);

NAND3xp33_ASAP7_75t_L g2705 ( 
.A(n_2393),
.B(n_1538),
.C(n_1531),
.Y(n_2705)
);

INVxp67_ASAP7_75t_SL g2706 ( 
.A(n_2304),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2353),
.Y(n_2707)
);

AND2x4_ASAP7_75t_L g2708 ( 
.A(n_2354),
.B(n_2228),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2455),
.B(n_1531),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2360),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2363),
.Y(n_2711)
);

XOR2x2_ASAP7_75t_L g2712 ( 
.A(n_2380),
.B(n_1538),
.Y(n_2712)
);

BUFx6f_ASAP7_75t_L g2713 ( 
.A(n_2594),
.Y(n_2713)
);

NOR3xp33_ASAP7_75t_L g2714 ( 
.A(n_2378),
.B(n_2238),
.C(n_2221),
.Y(n_2714)
);

NAND2x1_ASAP7_75t_L g2715 ( 
.A(n_2448),
.B(n_2221),
.Y(n_2715)
);

NAND2xp5_ASAP7_75t_L g2716 ( 
.A(n_2367),
.B(n_2105),
.Y(n_2716)
);

INVxp67_ASAP7_75t_L g2717 ( 
.A(n_2306),
.Y(n_2717)
);

NAND3xp33_ASAP7_75t_L g2718 ( 
.A(n_2337),
.B(n_1543),
.C(n_1539),
.Y(n_2718)
);

AND2x6_ASAP7_75t_SL g2719 ( 
.A(n_2434),
.B(n_1799),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2367),
.B(n_2130),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2369),
.Y(n_2721)
);

BUFx6f_ASAP7_75t_L g2722 ( 
.A(n_2603),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_L g2723 ( 
.A(n_2332),
.B(n_2130),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2445),
.Y(n_2724)
);

NAND3xp33_ASAP7_75t_L g2725 ( 
.A(n_2337),
.B(n_2322),
.C(n_2637),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2332),
.B(n_2350),
.Y(n_2726)
);

INVx8_ASAP7_75t_L g2727 ( 
.A(n_2434),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2350),
.B(n_2130),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2403),
.B(n_2137),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2477),
.Y(n_2730)
);

INVx2_ASAP7_75t_SL g2731 ( 
.A(n_2303),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2403),
.B(n_2137),
.Y(n_2732)
);

NAND2xp5_ASAP7_75t_L g2733 ( 
.A(n_2421),
.B(n_2425),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2421),
.B(n_2137),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2425),
.B(n_2145),
.Y(n_2735)
);

INVx2_ASAP7_75t_SL g2736 ( 
.A(n_2303),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2371),
.Y(n_2737)
);

INVx2_ASAP7_75t_L g2738 ( 
.A(n_2486),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2375),
.Y(n_2739)
);

NOR2xp33_ASAP7_75t_L g2740 ( 
.A(n_2349),
.B(n_1539),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2349),
.B(n_2145),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2389),
.Y(n_2742)
);

AND2x2_ASAP7_75t_L g2743 ( 
.A(n_2478),
.B(n_1543),
.Y(n_2743)
);

BUFx6f_ASAP7_75t_L g2744 ( 
.A(n_2603),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2489),
.B(n_2145),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2391),
.Y(n_2746)
);

INVxp33_ASAP7_75t_L g2747 ( 
.A(n_2577),
.Y(n_2747)
);

NOR3xp33_ASAP7_75t_L g2748 ( 
.A(n_2433),
.B(n_2238),
.C(n_2221),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2487),
.B(n_2032),
.Y(n_2749)
);

INVx2_ASAP7_75t_SL g2750 ( 
.A(n_2341),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2489),
.B(n_2172),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2398),
.Y(n_2752)
);

BUFx6f_ASAP7_75t_L g2753 ( 
.A(n_2603),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_L g2754 ( 
.A(n_2482),
.B(n_1548),
.Y(n_2754)
);

OR2x6_ASAP7_75t_L g2755 ( 
.A(n_2524),
.B(n_1799),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2526),
.B(n_1548),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2491),
.Y(n_2757)
);

NAND2xp5_ASAP7_75t_SL g2758 ( 
.A(n_2330),
.B(n_2032),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_SL g2759 ( 
.A(n_2330),
.B(n_2035),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2402),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2493),
.B(n_2172),
.Y(n_2761)
);

AOI22xp5_ASAP7_75t_L g2762 ( 
.A1(n_2459),
.A2(n_1652),
.B1(n_1600),
.B2(n_1564),
.Y(n_2762)
);

AND2x2_ASAP7_75t_L g2763 ( 
.A(n_2497),
.B(n_1558),
.Y(n_2763)
);

NAND2xp5_ASAP7_75t_L g2764 ( 
.A(n_2493),
.B(n_2514),
.Y(n_2764)
);

BUFx6f_ASAP7_75t_L g2765 ( 
.A(n_2603),
.Y(n_2765)
);

AOI22xp5_ASAP7_75t_L g2766 ( 
.A1(n_2459),
.A2(n_1652),
.B1(n_1600),
.B2(n_1564),
.Y(n_2766)
);

AND2x2_ASAP7_75t_L g2767 ( 
.A(n_2497),
.B(n_1558),
.Y(n_2767)
);

NOR3xp33_ASAP7_75t_L g2768 ( 
.A(n_2437),
.B(n_1300),
.C(n_1297),
.Y(n_2768)
);

AOI22xp33_ASAP7_75t_L g2769 ( 
.A1(n_2322),
.A2(n_1591),
.B1(n_1601),
.B2(n_1573),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_SL g2770 ( 
.A(n_2406),
.B(n_2035),
.Y(n_2770)
);

INVx3_ASAP7_75t_L g2771 ( 
.A(n_2571),
.Y(n_2771)
);

AOI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2645),
.A2(n_1643),
.B1(n_1591),
.B2(n_1601),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2514),
.B(n_2172),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2383),
.B(n_1573),
.Y(n_2774)
);

INVx2_ASAP7_75t_L g2775 ( 
.A(n_2495),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_2520),
.B(n_2490),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2560),
.B(n_2191),
.Y(n_2777)
);

INVx2_ASAP7_75t_L g2778 ( 
.A(n_2511),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2418),
.B(n_1606),
.Y(n_2779)
);

INVx1_ASAP7_75t_L g2780 ( 
.A(n_2409),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2411),
.Y(n_2781)
);

NOR2xp33_ASAP7_75t_L g2782 ( 
.A(n_2418),
.B(n_1606),
.Y(n_2782)
);

NOR2xp33_ASAP7_75t_L g2783 ( 
.A(n_2401),
.B(n_1618),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2521),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2416),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2420),
.Y(n_2786)
);

NAND3xp33_ASAP7_75t_L g2787 ( 
.A(n_2637),
.B(n_1640),
.C(n_1618),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2566),
.B(n_2195),
.Y(n_2788)
);

AND2x2_ASAP7_75t_L g2789 ( 
.A(n_2499),
.B(n_1640),
.Y(n_2789)
);

NAND2xp5_ASAP7_75t_SL g2790 ( 
.A(n_2410),
.B(n_2537),
.Y(n_2790)
);

NAND2xp33_ASAP7_75t_SL g2791 ( 
.A(n_2373),
.B(n_2035),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2439),
.Y(n_2792)
);

INVx2_ASAP7_75t_SL g2793 ( 
.A(n_2318),
.Y(n_2793)
);

INVx2_ASAP7_75t_L g2794 ( 
.A(n_2522),
.Y(n_2794)
);

INVx1_ASAP7_75t_L g2795 ( 
.A(n_2442),
.Y(n_2795)
);

NAND3xp33_ASAP7_75t_L g2796 ( 
.A(n_2423),
.B(n_1647),
.C(n_1643),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2540),
.Y(n_2797)
);

NAND3xp33_ASAP7_75t_L g2798 ( 
.A(n_2407),
.B(n_1651),
.C(n_1647),
.Y(n_2798)
);

NOR3xp33_ASAP7_75t_L g2799 ( 
.A(n_2404),
.B(n_1306),
.C(n_1302),
.Y(n_2799)
);

INVx2_ASAP7_75t_SL g2800 ( 
.A(n_2324),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_SL g2801 ( 
.A(n_2532),
.B(n_2035),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2334),
.B(n_1651),
.Y(n_2802)
);

AO221x1_ASAP7_75t_L g2803 ( 
.A1(n_2506),
.A2(n_2056),
.B1(n_2072),
.B2(n_2061),
.C(n_2042),
.Y(n_2803)
);

INVx1_ASAP7_75t_L g2804 ( 
.A(n_2443),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2544),
.Y(n_2805)
);

BUFx6f_ASAP7_75t_L g2806 ( 
.A(n_2632),
.Y(n_2806)
);

INVx2_ASAP7_75t_L g2807 ( 
.A(n_2545),
.Y(n_2807)
);

OR2x2_ASAP7_75t_L g2808 ( 
.A(n_2386),
.B(n_1665),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2427),
.B(n_1665),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2444),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2551),
.B(n_2195),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2446),
.B(n_2198),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2632),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2556),
.B(n_1682),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2447),
.Y(n_2815)
);

BUFx6f_ASAP7_75t_SL g2816 ( 
.A(n_2430),
.Y(n_2816)
);

NAND2xp5_ASAP7_75t_SL g2817 ( 
.A(n_2354),
.B(n_2042),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2446),
.B(n_2198),
.Y(n_2818)
);

NOR2xp67_ASAP7_75t_SL g2819 ( 
.A(n_2479),
.B(n_2508),
.Y(n_2819)
);

OR2x6_ASAP7_75t_L g2820 ( 
.A(n_2524),
.B(n_2191),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2451),
.Y(n_2821)
);

NOR2xp33_ASAP7_75t_L g2822 ( 
.A(n_2427),
.B(n_1682),
.Y(n_2822)
);

INVx1_ASAP7_75t_L g2823 ( 
.A(n_2445),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2449),
.B(n_2193),
.Y(n_2824)
);

NAND2xp5_ASAP7_75t_L g2825 ( 
.A(n_2449),
.B(n_2462),
.Y(n_2825)
);

BUFx6f_ASAP7_75t_L g2826 ( 
.A(n_2632),
.Y(n_2826)
);

NAND2xp5_ASAP7_75t_L g2827 ( 
.A(n_2462),
.B(n_2193),
.Y(n_2827)
);

NOR2xp33_ASAP7_75t_L g2828 ( 
.A(n_2461),
.B(n_1683),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2438),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_L g2830 ( 
.A(n_2531),
.B(n_2018),
.Y(n_2830)
);

NOR2xp33_ASAP7_75t_SL g2831 ( 
.A(n_2436),
.B(n_1683),
.Y(n_2831)
);

INVxp67_ASAP7_75t_L g2832 ( 
.A(n_2593),
.Y(n_2832)
);

NOR2xp33_ASAP7_75t_L g2833 ( 
.A(n_2461),
.B(n_2042),
.Y(n_2833)
);

NAND2xp5_ASAP7_75t_L g2834 ( 
.A(n_2531),
.B(n_2039),
.Y(n_2834)
);

INVxp67_ASAP7_75t_L g2835 ( 
.A(n_2408),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2438),
.B(n_2039),
.Y(n_2836)
);

AO221x1_ASAP7_75t_L g2837 ( 
.A1(n_2506),
.A2(n_2056),
.B1(n_2072),
.B2(n_2061),
.C(n_2042),
.Y(n_2837)
);

NAND2xp5_ASAP7_75t_SL g2838 ( 
.A(n_2352),
.B(n_2056),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_SL g2839 ( 
.A(n_2352),
.B(n_2056),
.Y(n_2839)
);

AND2x2_ASAP7_75t_L g2840 ( 
.A(n_2408),
.B(n_1308),
.Y(n_2840)
);

INVx2_ASAP7_75t_SL g2841 ( 
.A(n_2366),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_SL g2842 ( 
.A(n_2352),
.B(n_2061),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2452),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2632),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2547),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2471),
.B(n_2018),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2454),
.Y(n_2847)
);

AND2x6_ASAP7_75t_L g2848 ( 
.A(n_2319),
.B(n_2071),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2458),
.Y(n_2849)
);

NOR2xp33_ASAP7_75t_L g2850 ( 
.A(n_2362),
.B(n_2061),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_SL g2851 ( 
.A(n_2352),
.B(n_2647),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_L g2852 ( 
.A(n_2557),
.B(n_2513),
.Y(n_2852)
);

BUFx6f_ASAP7_75t_L g2853 ( 
.A(n_2643),
.Y(n_2853)
);

AND2x2_ASAP7_75t_L g2854 ( 
.A(n_2542),
.B(n_1310),
.Y(n_2854)
);

BUFx6f_ASAP7_75t_SL g2855 ( 
.A(n_2498),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2471),
.B(n_2060),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_SL g2857 ( 
.A(n_2473),
.B(n_2072),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_SL g2858 ( 
.A(n_2379),
.B(n_2072),
.Y(n_2858)
);

AO221x1_ASAP7_75t_L g2859 ( 
.A1(n_2441),
.A2(n_2125),
.B1(n_2132),
.B2(n_2077),
.C(n_2073),
.Y(n_2859)
);

INVx1_ASAP7_75t_L g2860 ( 
.A(n_2460),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2475),
.B(n_2060),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_SL g2862 ( 
.A(n_2379),
.B(n_2073),
.Y(n_2862)
);

BUFx6f_ASAP7_75t_L g2863 ( 
.A(n_2643),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2467),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2472),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2553),
.Y(n_2866)
);

NOR2xp33_ASAP7_75t_L g2867 ( 
.A(n_2613),
.B(n_2073),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2554),
.Y(n_2868)
);

INVx2_ASAP7_75t_SL g2869 ( 
.A(n_2412),
.Y(n_2869)
);

OR2x6_ASAP7_75t_L g2870 ( 
.A(n_2524),
.B(n_2295),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2474),
.Y(n_2871)
);

NAND2xp5_ASAP7_75t_L g2872 ( 
.A(n_2475),
.B(n_2060),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2476),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_SL g2874 ( 
.A(n_2509),
.B(n_2570),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2539),
.B(n_1981),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2539),
.B(n_1981),
.Y(n_2876)
);

BUFx5_ASAP7_75t_L g2877 ( 
.A(n_2591),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2500),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2535),
.B(n_1981),
.Y(n_2879)
);

INVx2_ASAP7_75t_L g2880 ( 
.A(n_2558),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2562),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2501),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2573),
.Y(n_2883)
);

INVx2_ASAP7_75t_SL g2884 ( 
.A(n_2307),
.Y(n_2884)
);

INVx2_ASAP7_75t_L g2885 ( 
.A(n_2581),
.Y(n_2885)
);

BUFx6f_ASAP7_75t_L g2886 ( 
.A(n_2643),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_SL g2887 ( 
.A(n_2509),
.B(n_2073),
.Y(n_2887)
);

NOR2xp33_ASAP7_75t_L g2888 ( 
.A(n_2549),
.B(n_2077),
.Y(n_2888)
);

INVxp33_ASAP7_75t_L g2889 ( 
.A(n_2457),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_L g2890 ( 
.A(n_2485),
.B(n_2077),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2503),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2505),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2507),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2492),
.B(n_2077),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_SL g2895 ( 
.A(n_2323),
.B(n_2125),
.Y(n_2895)
);

AOI221xp5_ASAP7_75t_L g2896 ( 
.A1(n_2441),
.A2(n_1315),
.B1(n_1314),
.B2(n_1312),
.C(n_2240),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_2431),
.B(n_2125),
.Y(n_2897)
);

INVxp33_ASAP7_75t_L g2898 ( 
.A(n_2621),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2535),
.B(n_2057),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2515),
.B(n_2057),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2516),
.B(n_2607),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_SL g2902 ( 
.A(n_2385),
.B(n_2125),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2519),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2607),
.B(n_2057),
.Y(n_2904)
);

AND2x2_ASAP7_75t_L g2905 ( 
.A(n_2586),
.B(n_2202),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_SL g2906 ( 
.A(n_2385),
.B(n_2132),
.Y(n_2906)
);

NAND2xp5_ASAP7_75t_SL g2907 ( 
.A(n_2419),
.B(n_2132),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_SL g2908 ( 
.A(n_2419),
.B(n_2132),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2525),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2307),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2589),
.B(n_2135),
.Y(n_2911)
);

INVx1_ASAP7_75t_L g2912 ( 
.A(n_2530),
.Y(n_2912)
);

NOR2xp33_ASAP7_75t_L g2913 ( 
.A(n_2561),
.B(n_2135),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2541),
.Y(n_2914)
);

INVx8_ASAP7_75t_L g2915 ( 
.A(n_2502),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2590),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2407),
.B(n_2135),
.Y(n_2917)
);

BUFx6f_ASAP7_75t_L g2918 ( 
.A(n_2643),
.Y(n_2918)
);

INVx2_ASAP7_75t_L g2919 ( 
.A(n_2595),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2552),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_SL g2921 ( 
.A(n_2599),
.B(n_2571),
.Y(n_2921)
);

NOR2xp33_ASAP7_75t_L g2922 ( 
.A(n_2342),
.B(n_2135),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2563),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2559),
.B(n_2046),
.Y(n_2924)
);

INVx8_ASAP7_75t_L g2925 ( 
.A(n_2502),
.Y(n_2925)
);

NAND2xp5_ASAP7_75t_L g2926 ( 
.A(n_2559),
.B(n_2046),
.Y(n_2926)
);

NOR2xp33_ASAP7_75t_SL g2927 ( 
.A(n_2468),
.B(n_2279),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2598),
.B(n_1985),
.Y(n_2928)
);

NAND2xp5_ASAP7_75t_SL g2929 ( 
.A(n_2344),
.B(n_2139),
.Y(n_2929)
);

NOR3xp33_ASAP7_75t_L g2930 ( 
.A(n_2450),
.B(n_2243),
.C(n_2240),
.Y(n_2930)
);

HB1xp67_ASAP7_75t_L g2931 ( 
.A(n_2527),
.Y(n_2931)
);

INVx2_ASAP7_75t_L g2932 ( 
.A(n_2625),
.Y(n_2932)
);

NOR2xp33_ASAP7_75t_L g2933 ( 
.A(n_2527),
.B(n_2139),
.Y(n_2933)
);

NAND2xp5_ASAP7_75t_SL g2934 ( 
.A(n_2344),
.B(n_2139),
.Y(n_2934)
);

NOR3xp33_ASAP7_75t_L g2935 ( 
.A(n_2424),
.B(n_2243),
.C(n_2240),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2598),
.B(n_1985),
.Y(n_2936)
);

INVx2_ASAP7_75t_SL g2937 ( 
.A(n_2440),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_SL g2938 ( 
.A(n_2575),
.B(n_2139),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2543),
.B(n_1987),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2567),
.Y(n_2940)
);

BUFx6f_ASAP7_75t_SL g2941 ( 
.A(n_2527),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2543),
.B(n_1987),
.Y(n_2942)
);

BUFx6f_ASAP7_75t_L g2943 ( 
.A(n_2328),
.Y(n_2943)
);

AND2x4_ASAP7_75t_L g2944 ( 
.A(n_2496),
.B(n_2140),
.Y(n_2944)
);

NAND2x1p5_ASAP7_75t_L g2945 ( 
.A(n_2550),
.B(n_2146),
.Y(n_2945)
);

NAND3xp33_ASAP7_75t_L g2946 ( 
.A(n_2429),
.B(n_2295),
.C(n_2279),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_SL g2947 ( 
.A(n_2538),
.Y(n_2947)
);

AOI22xp33_ASAP7_75t_L g2948 ( 
.A1(n_2725),
.A2(n_2463),
.B1(n_2612),
.B2(n_2604),
.Y(n_2948)
);

INVx1_ASAP7_75t_L g2949 ( 
.A(n_2659),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2664),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2764),
.B(n_2463),
.Y(n_2951)
);

NAND2xp5_ASAP7_75t_L g2952 ( 
.A(n_2686),
.B(n_2618),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_SL g2953 ( 
.A(n_2661),
.B(n_2585),
.Y(n_2953)
);

INVx1_ASAP7_75t_SL g2954 ( 
.A(n_2696),
.Y(n_2954)
);

OAI22xp5_ASAP7_75t_L g2955 ( 
.A1(n_2776),
.A2(n_2617),
.B1(n_2627),
.B2(n_2496),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_SL g2956 ( 
.A(n_2733),
.B(n_2585),
.Y(n_2956)
);

INVx8_ASAP7_75t_L g2957 ( 
.A(n_2700),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2667),
.Y(n_2958)
);

NAND2xp5_ASAP7_75t_L g2959 ( 
.A(n_2704),
.B(n_2618),
.Y(n_2959)
);

NAND2xp33_ASAP7_75t_SL g2960 ( 
.A(n_2884),
.B(n_2910),
.Y(n_2960)
);

AOI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2740),
.A2(n_2617),
.B1(n_2627),
.B2(n_2587),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2668),
.Y(n_2962)
);

AOI22xp33_ASAP7_75t_L g2963 ( 
.A1(n_2718),
.A2(n_2587),
.B1(n_2629),
.B2(n_2564),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2676),
.Y(n_2964)
);

INVx2_ASAP7_75t_SL g2965 ( 
.A(n_2700),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2829),
.B(n_2538),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2829),
.B(n_2538),
.Y(n_2967)
);

NOR2xp33_ASAP7_75t_L g2968 ( 
.A(n_2809),
.B(n_2405),
.Y(n_2968)
);

BUFx3_ASAP7_75t_L g2969 ( 
.A(n_2793),
.Y(n_2969)
);

AOI22xp5_ASAP7_75t_L g2970 ( 
.A1(n_2699),
.A2(n_2426),
.B1(n_2502),
.B2(n_2435),
.Y(n_2970)
);

BUFx8_ASAP7_75t_L g2971 ( 
.A(n_2816),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2663),
.B(n_2652),
.Y(n_2972)
);

INVx5_ASAP7_75t_L g2973 ( 
.A(n_2655),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2671),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2673),
.B(n_2850),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2674),
.Y(n_2976)
);

AND2x6_ASAP7_75t_L g2977 ( 
.A(n_2655),
.B(n_2616),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2679),
.Y(n_2978)
);

OR2x6_ASAP7_75t_L g2979 ( 
.A(n_2727),
.B(n_2644),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2657),
.B(n_2652),
.Y(n_2980)
);

A2O1A1Ixp33_ASAP7_75t_L g2981 ( 
.A1(n_2681),
.A2(n_2584),
.B(n_2518),
.C(n_2529),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2658),
.B(n_2496),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2835),
.B(n_2529),
.Y(n_2983)
);

A2O1A1Ixp33_ASAP7_75t_L g2984 ( 
.A1(n_2874),
.A2(n_2518),
.B(n_2602),
.C(n_2480),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_SL g2985 ( 
.A(n_2913),
.B(n_2616),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2687),
.Y(n_2986)
);

AOI22xp5_ASAP7_75t_L g2987 ( 
.A1(n_2783),
.A2(n_2435),
.B1(n_2428),
.B2(n_2597),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_2655),
.Y(n_2988)
);

AO22x1_ASAP7_75t_L g2989 ( 
.A1(n_2747),
.A2(n_2435),
.B1(n_2428),
.B2(n_2591),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2840),
.B(n_2825),
.Y(n_2990)
);

INVx1_ASAP7_75t_L g2991 ( 
.A(n_2691),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2697),
.Y(n_2992)
);

INVx2_ASAP7_75t_SL g2993 ( 
.A(n_2727),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2726),
.B(n_2374),
.Y(n_2994)
);

BUFx3_ASAP7_75t_L g2995 ( 
.A(n_2800),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2854),
.B(n_2394),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_L g2997 ( 
.A(n_2901),
.B(n_2504),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_L g2998 ( 
.A(n_2852),
.B(n_2754),
.Y(n_2998)
);

NOR2x1p5_ASAP7_75t_L g2999 ( 
.A(n_2662),
.B(n_2582),
.Y(n_2999)
);

INVxp67_ASAP7_75t_L g3000 ( 
.A(n_2779),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2707),
.Y(n_3001)
);

NAND2x1_ASAP7_75t_L g3002 ( 
.A(n_2656),
.B(n_2578),
.Y(n_3002)
);

AND2x2_ASAP7_75t_L g3003 ( 
.A(n_2743),
.B(n_2564),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2688),
.Y(n_3004)
);

AOI22xp5_ASAP7_75t_L g3005 ( 
.A1(n_2756),
.A2(n_2435),
.B1(n_2428),
.B2(n_2592),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_SL g3006 ( 
.A(n_2927),
.B(n_2636),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2724),
.B(n_2428),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2822),
.B(n_2510),
.Y(n_3008)
);

OAI21xp5_ASAP7_75t_L g3009 ( 
.A1(n_2761),
.A2(n_2548),
.B(n_2546),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2897),
.B(n_2787),
.Y(n_3010)
);

NOR2xp33_ASAP7_75t_L g3011 ( 
.A(n_2828),
.B(n_2512),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2724),
.B(n_2823),
.Y(n_3012)
);

AOI22xp5_ASAP7_75t_L g3013 ( 
.A1(n_2802),
.A2(n_2435),
.B1(n_2428),
.B2(n_2610),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2823),
.B(n_2641),
.Y(n_3014)
);

INVx2_ASAP7_75t_L g3015 ( 
.A(n_2689),
.Y(n_3015)
);

AOI21xp5_ASAP7_75t_L g3016 ( 
.A1(n_2675),
.A2(n_2574),
.B(n_2310),
.Y(n_3016)
);

NOR2xp33_ASAP7_75t_L g3017 ( 
.A(n_2690),
.B(n_2626),
.Y(n_3017)
);

NOR2xp33_ASAP7_75t_L g3018 ( 
.A(n_2772),
.B(n_2631),
.Y(n_3018)
);

INVx2_ASAP7_75t_SL g3019 ( 
.A(n_2695),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2782),
.B(n_2646),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2710),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2763),
.B(n_2653),
.Y(n_3022)
);

OAI22xp5_ASAP7_75t_L g3023 ( 
.A1(n_2701),
.A2(n_2602),
.B1(n_2596),
.B2(n_2572),
.Y(n_3023)
);

AOI22xp5_ASAP7_75t_L g3024 ( 
.A1(n_2705),
.A2(n_2619),
.B1(n_2572),
.B2(n_2591),
.Y(n_3024)
);

INVx1_ASAP7_75t_L g3025 ( 
.A(n_2711),
.Y(n_3025)
);

INVx8_ASAP7_75t_L g3026 ( 
.A(n_2915),
.Y(n_3026)
);

INVxp67_ASAP7_75t_L g3027 ( 
.A(n_2767),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2730),
.Y(n_3028)
);

AO22x1_ASAP7_75t_L g3029 ( 
.A1(n_2898),
.A2(n_2591),
.B1(n_2576),
.B2(n_2642),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2721),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2737),
.Y(n_3031)
);

O2A1O1Ixp33_ASAP7_75t_L g3032 ( 
.A1(n_2774),
.A2(n_2635),
.B(n_2596),
.C(n_2640),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2684),
.B(n_2654),
.Y(n_3033)
);

NAND2xp5_ASAP7_75t_L g3034 ( 
.A(n_2709),
.B(n_2890),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2677),
.B(n_2678),
.Y(n_3035)
);

BUFx3_ASAP7_75t_L g3036 ( 
.A(n_2841),
.Y(n_3036)
);

AOI22xp33_ASAP7_75t_L g3037 ( 
.A1(n_2769),
.A2(n_2564),
.B1(n_2576),
.B2(n_2579),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2832),
.B(n_2583),
.Y(n_3038)
);

AOI21x1_ASAP7_75t_L g3039 ( 
.A1(n_2917),
.A2(n_2548),
.B(n_2546),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2812),
.B(n_2588),
.Y(n_3040)
);

AOI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2712),
.A2(n_2762),
.B1(n_2766),
.B2(n_2698),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2738),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2739),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2789),
.B(n_2650),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2666),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2814),
.B(n_2483),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2757),
.Y(n_3047)
);

BUFx6f_ASAP7_75t_L g3048 ( 
.A(n_2666),
.Y(n_3048)
);

BUFx3_ASAP7_75t_L g3049 ( 
.A(n_2869),
.Y(n_3049)
);

OAI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2692),
.A2(n_2644),
.B1(n_2340),
.B2(n_2351),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2775),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_2798),
.B(n_2483),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_2660),
.A2(n_2576),
.B1(n_2614),
.B2(n_2606),
.Y(n_3053)
);

NOR2xp33_ASAP7_75t_L g3054 ( 
.A(n_2808),
.B(n_2484),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2755),
.B(n_2575),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2742),
.Y(n_3056)
);

AOI22xp33_ASAP7_75t_L g3057 ( 
.A1(n_2796),
.A2(n_2576),
.B1(n_2623),
.B2(n_2615),
.Y(n_3057)
);

OR2x2_ASAP7_75t_L g3058 ( 
.A(n_2755),
.B(n_2628),
.Y(n_3058)
);

NAND2x1p5_ASAP7_75t_L g3059 ( 
.A(n_2666),
.B(n_2550),
.Y(n_3059)
);

HB1xp67_ASAP7_75t_SL g3060 ( 
.A(n_2682),
.Y(n_3060)
);

BUFx3_ASAP7_75t_L g3061 ( 
.A(n_2750),
.Y(n_3061)
);

NAND2xp33_ASAP7_75t_SL g3062 ( 
.A(n_2819),
.B(n_2319),
.Y(n_3062)
);

NAND2xp5_ASAP7_75t_SL g3063 ( 
.A(n_2911),
.B(n_2550),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2818),
.B(n_2630),
.Y(n_3064)
);

AOI21xp5_ASAP7_75t_L g3065 ( 
.A1(n_2706),
.A2(n_2574),
.B(n_2310),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2746),
.Y(n_3066)
);

AOI22xp33_ASAP7_75t_L g3067 ( 
.A1(n_2859),
.A2(n_2576),
.B1(n_2638),
.B2(n_2368),
.Y(n_3067)
);

OR2x6_ASAP7_75t_L g3068 ( 
.A(n_2915),
.B(n_2644),
.Y(n_3068)
);

INVx3_ASAP7_75t_L g3069 ( 
.A(n_2670),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_L g3070 ( 
.A(n_2824),
.B(n_2300),
.Y(n_3070)
);

NOR3xp33_ASAP7_75t_L g3071 ( 
.A(n_2791),
.B(n_2488),
.C(n_2484),
.Y(n_3071)
);

INVx2_ASAP7_75t_SL g3072 ( 
.A(n_2731),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2717),
.B(n_2305),
.Y(n_3073)
);

AND2x6_ASAP7_75t_SL g3074 ( 
.A(n_2867),
.B(n_2308),
.Y(n_3074)
);

AND2x2_ASAP7_75t_SL g3075 ( 
.A(n_2831),
.B(n_2578),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_2752),
.B(n_2309),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2760),
.B(n_2312),
.Y(n_3077)
);

INVx2_ASAP7_75t_L g3078 ( 
.A(n_2778),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2780),
.B(n_2321),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2784),
.Y(n_3080)
);

CKINVDCx5p33_ASAP7_75t_R g3081 ( 
.A(n_2816),
.Y(n_3081)
);

NOR2xp33_ASAP7_75t_L g3082 ( 
.A(n_2790),
.B(n_2488),
.Y(n_3082)
);

AOI22xp33_ASAP7_75t_L g3083 ( 
.A1(n_2794),
.A2(n_2370),
.B1(n_2377),
.B2(n_2365),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_SL g3084 ( 
.A(n_2833),
.B(n_2550),
.Y(n_3084)
);

NOR2xp33_ASAP7_75t_L g3085 ( 
.A(n_2680),
.B(n_2494),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2797),
.Y(n_3086)
);

INVx2_ASAP7_75t_L g3087 ( 
.A(n_2805),
.Y(n_3087)
);

INVx4_ASAP7_75t_L g3088 ( 
.A(n_2670),
.Y(n_3088)
);

NAND2xp5_ASAP7_75t_SL g3089 ( 
.A(n_2670),
.B(n_2328),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_SL g3090 ( 
.A(n_2713),
.B(n_2328),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_2680),
.B(n_2736),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2781),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2785),
.Y(n_3093)
);

NAND2xp5_ASAP7_75t_L g3094 ( 
.A(n_2786),
.B(n_2325),
.Y(n_3094)
);

AOI22xp33_ASAP7_75t_L g3095 ( 
.A1(n_2807),
.A2(n_2866),
.B1(n_2868),
.B2(n_2845),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2792),
.B(n_2327),
.Y(n_3096)
);

A2O1A1Ixp33_ASAP7_75t_L g3097 ( 
.A1(n_2694),
.A2(n_2308),
.B(n_2351),
.C(n_2340),
.Y(n_3097)
);

AOI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2741),
.A2(n_2591),
.B1(n_2622),
.B2(n_2331),
.Y(n_3098)
);

AOI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_2745),
.A2(n_2376),
.B1(n_2384),
.B2(n_2364),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_SL g3100 ( 
.A(n_2713),
.B(n_2355),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2880),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_SL g3102 ( 
.A(n_2713),
.B(n_2355),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2795),
.B(n_2336),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_SL g3104 ( 
.A(n_2722),
.B(n_2355),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_SL g3105 ( 
.A(n_2722),
.B(n_2744),
.Y(n_3105)
);

NOR2xp33_ASAP7_75t_L g3106 ( 
.A(n_2708),
.B(n_2494),
.Y(n_3106)
);

OR2x2_ASAP7_75t_L g3107 ( 
.A(n_2804),
.B(n_2338),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2881),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2810),
.B(n_2339),
.Y(n_3109)
);

OR2x2_ASAP7_75t_L g3110 ( 
.A(n_2815),
.B(n_2361),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2821),
.B(n_2382),
.Y(n_3111)
);

AOI22xp33_ASAP7_75t_L g3112 ( 
.A1(n_2883),
.A2(n_2395),
.B1(n_2397),
.B2(n_2392),
.Y(n_3112)
);

NOR2xp33_ASAP7_75t_L g3113 ( 
.A(n_2708),
.B(n_2388),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2843),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2722),
.B(n_2358),
.Y(n_3115)
);

NAND2xp5_ASAP7_75t_L g3116 ( 
.A(n_2847),
.B(n_2399),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2849),
.Y(n_3117)
);

NAND2xp5_ASAP7_75t_L g3118 ( 
.A(n_2860),
.B(n_2414),
.Y(n_3118)
);

BUFx2_ASAP7_75t_L g3119 ( 
.A(n_2870),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_L g3120 ( 
.A(n_2864),
.B(n_2432),
.Y(n_3120)
);

NAND2xp5_ASAP7_75t_L g3121 ( 
.A(n_2865),
.B(n_2453),
.Y(n_3121)
);

AOI22xp33_ASAP7_75t_L g3122 ( 
.A1(n_2885),
.A2(n_2465),
.B1(n_2464),
.B2(n_2569),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2871),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2873),
.B(n_2387),
.Y(n_3124)
);

NAND2xp5_ASAP7_75t_L g3125 ( 
.A(n_2878),
.B(n_2387),
.Y(n_3125)
);

NOR2xp33_ASAP7_75t_L g3126 ( 
.A(n_2685),
.B(n_2388),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2882),
.B(n_2400),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_2931),
.B(n_2601),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2891),
.B(n_2400),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_SL g3130 ( 
.A(n_2744),
.B(n_2358),
.Y(n_3130)
);

NOR2xp33_ASAP7_75t_L g3131 ( 
.A(n_2672),
.B(n_2396),
.Y(n_3131)
);

AND2x2_ASAP7_75t_L g3132 ( 
.A(n_2892),
.B(n_2601),
.Y(n_3132)
);

OR2x2_ASAP7_75t_L g3133 ( 
.A(n_2893),
.B(n_2605),
.Y(n_3133)
);

AO22x1_ASAP7_75t_L g3134 ( 
.A1(n_2889),
.A2(n_2649),
.B1(n_2396),
.B2(n_2523),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2916),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2919),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2830),
.B(n_2580),
.Y(n_3137)
);

INVx2_ASAP7_75t_L g3138 ( 
.A(n_2932),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2903),
.Y(n_3139)
);

AOI22xp33_ASAP7_75t_L g3140 ( 
.A1(n_2941),
.A2(n_2569),
.B1(n_2201),
.B2(n_2580),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2909),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_2912),
.B(n_2605),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2834),
.B(n_2639),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2914),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2920),
.Y(n_3145)
);

INVxp67_ASAP7_75t_SL g3146 ( 
.A(n_2928),
.Y(n_3146)
);

NAND2xp5_ASAP7_75t_L g3147 ( 
.A(n_2925),
.B(n_2648),
.Y(n_3147)
);

INVx4_ASAP7_75t_L g3148 ( 
.A(n_2744),
.Y(n_3148)
);

INVx4_ASAP7_75t_L g3149 ( 
.A(n_2753),
.Y(n_3149)
);

OAI22xp5_ASAP7_75t_L g3150 ( 
.A1(n_2683),
.A2(n_2364),
.B1(n_2384),
.B2(n_2376),
.Y(n_3150)
);

NOR2xp67_ASAP7_75t_L g3151 ( 
.A(n_2937),
.B(n_2456),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2925),
.B(n_2608),
.Y(n_3152)
);

NOR3xp33_ASAP7_75t_SL g3153 ( 
.A(n_2921),
.B(n_6),
.C(n_7),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2923),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2940),
.Y(n_3155)
);

BUFx6f_ASAP7_75t_L g3156 ( 
.A(n_2753),
.Y(n_3156)
);

AOI22xp5_ASAP7_75t_L g3157 ( 
.A1(n_2751),
.A2(n_2609),
.B1(n_2624),
.B2(n_2608),
.Y(n_3157)
);

NAND2xp5_ASAP7_75t_SL g3158 ( 
.A(n_2753),
.B(n_2358),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2933),
.B(n_2609),
.Y(n_3159)
);

OAI22xp33_ASAP7_75t_L g3160 ( 
.A1(n_2729),
.A2(n_2651),
.B1(n_2620),
.B2(n_2523),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2777),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2773),
.B(n_2624),
.Y(n_3162)
);

A2O1A1Ixp33_ASAP7_75t_L g3163 ( 
.A1(n_2665),
.A2(n_2223),
.B(n_2536),
.C(n_2456),
.Y(n_3163)
);

AOI22xp33_ASAP7_75t_L g3164 ( 
.A1(n_2941),
.A2(n_2201),
.B1(n_2117),
.B2(n_2116),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_SL g3165 ( 
.A(n_2765),
.B(n_2381),
.Y(n_3165)
);

NOR2xp33_ASAP7_75t_L g3166 ( 
.A(n_2851),
.B(n_2536),
.Y(n_3166)
);

NOR2xp33_ASAP7_75t_SL g3167 ( 
.A(n_2877),
.B(n_2855),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2788),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2944),
.B(n_2634),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2811),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2944),
.B(n_2634),
.Y(n_3171)
);

AOI22xp5_ASAP7_75t_L g3172 ( 
.A1(n_2961),
.A2(n_2855),
.B1(n_2801),
.B2(n_2947),
.Y(n_3172)
);

OAI21x1_ASAP7_75t_L g3173 ( 
.A1(n_3016),
.A2(n_1982),
.B(n_2087),
.Y(n_3173)
);

AOI21xp5_ASAP7_75t_L g3174 ( 
.A1(n_3035),
.A2(n_2702),
.B(n_2929),
.Y(n_3174)
);

AOI21xp5_ASAP7_75t_L g3175 ( 
.A1(n_3097),
.A2(n_2934),
.B(n_2837),
.Y(n_3175)
);

NOR2xp67_ASAP7_75t_L g3176 ( 
.A(n_3019),
.B(n_2946),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2952),
.B(n_2896),
.Y(n_3177)
);

AOI21xp5_ASAP7_75t_L g3178 ( 
.A1(n_3163),
.A2(n_2803),
.B(n_2879),
.Y(n_3178)
);

NAND2xp5_ASAP7_75t_L g3179 ( 
.A(n_2972),
.B(n_2905),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_3141),
.Y(n_3180)
);

INVx3_ASAP7_75t_L g3181 ( 
.A(n_3059),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2949),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2990),
.B(n_2899),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_L g3184 ( 
.A(n_2980),
.B(n_2799),
.Y(n_3184)
);

NAND2x1p5_ASAP7_75t_L g3185 ( 
.A(n_2973),
.B(n_2765),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2950),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_3107),
.Y(n_3187)
);

HB1xp67_ASAP7_75t_L g3188 ( 
.A(n_2954),
.Y(n_3188)
);

HB1xp67_ASAP7_75t_L g3189 ( 
.A(n_2954),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_3110),
.Y(n_3190)
);

AOI22xp5_ASAP7_75t_L g3191 ( 
.A1(n_2955),
.A2(n_2947),
.B1(n_2888),
.B2(n_2870),
.Y(n_3191)
);

NAND2xp5_ASAP7_75t_L g3192 ( 
.A(n_2975),
.B(n_2820),
.Y(n_3192)
);

INVx1_ASAP7_75t_SL g3193 ( 
.A(n_3128),
.Y(n_3193)
);

BUFx2_ASAP7_75t_L g3194 ( 
.A(n_3055),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_L g3195 ( 
.A(n_2951),
.B(n_2959),
.Y(n_3195)
);

NOR2xp33_ASAP7_75t_L g3196 ( 
.A(n_2998),
.B(n_2719),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_3034),
.B(n_2820),
.Y(n_3197)
);

NOR2xp33_ASAP7_75t_SL g3198 ( 
.A(n_2955),
.B(n_2877),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2958),
.Y(n_3199)
);

AOI21xp33_ASAP7_75t_L g3200 ( 
.A1(n_3032),
.A2(n_2922),
.B(n_2894),
.Y(n_3200)
);

O2A1O1Ixp33_ASAP7_75t_L g3201 ( 
.A1(n_3010),
.A2(n_2693),
.B(n_2714),
.C(n_2857),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_3020),
.B(n_2732),
.Y(n_3202)
);

OAI22xp5_ASAP7_75t_L g3203 ( 
.A1(n_2968),
.A2(n_3044),
.B1(n_3008),
.B2(n_3011),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_2983),
.B(n_2734),
.Y(n_3204)
);

NOR2xp33_ASAP7_75t_SL g3205 ( 
.A(n_3075),
.B(n_2877),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_3033),
.B(n_2735),
.Y(n_3206)
);

INVx1_ASAP7_75t_L g3207 ( 
.A(n_2962),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_3003),
.B(n_2768),
.Y(n_3208)
);

AOI33xp33_ASAP7_75t_L g3209 ( 
.A1(n_3041),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_8),
.B3(n_10),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_3000),
.B(n_2936),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_2970),
.B(n_2703),
.Y(n_3211)
);

NOR2xp33_ASAP7_75t_L g3212 ( 
.A(n_3046),
.B(n_2771),
.Y(n_3212)
);

NAND2xp5_ASAP7_75t_L g3213 ( 
.A(n_3022),
.B(n_2836),
.Y(n_3213)
);

INVx2_ASAP7_75t_SL g3214 ( 
.A(n_2957),
.Y(n_3214)
);

AOI22xp5_ASAP7_75t_L g3215 ( 
.A1(n_3018),
.A2(n_2749),
.B1(n_2817),
.B2(n_2887),
.Y(n_3215)
);

OAI22xp5_ASAP7_75t_L g3216 ( 
.A1(n_3005),
.A2(n_2771),
.B1(n_2656),
.B2(n_2720),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3161),
.B(n_2716),
.Y(n_3217)
);

BUFx2_ASAP7_75t_SL g3218 ( 
.A(n_2965),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_3154),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_3168),
.B(n_2723),
.Y(n_3220)
);

A2O1A1Ixp33_ASAP7_75t_L g3221 ( 
.A1(n_3024),
.A2(n_2728),
.B(n_2748),
.C(n_2930),
.Y(n_3221)
);

NOR2xp33_ASAP7_75t_L g3222 ( 
.A(n_3054),
.B(n_2943),
.Y(n_3222)
);

A2O1A1Ixp33_ASAP7_75t_L g3223 ( 
.A1(n_3024),
.A2(n_2935),
.B(n_2770),
.C(n_2758),
.Y(n_3223)
);

OR2x2_ASAP7_75t_L g3224 ( 
.A(n_3155),
.B(n_2875),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2974),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2964),
.Y(n_3226)
);

AOI21xp5_ASAP7_75t_L g3227 ( 
.A1(n_3137),
.A2(n_2900),
.B(n_2861),
.Y(n_3227)
);

AOI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_3150),
.A2(n_2872),
.B(n_2856),
.Y(n_3228)
);

AO22x1_ASAP7_75t_L g3229 ( 
.A1(n_2971),
.A2(n_2806),
.B1(n_2813),
.B2(n_2765),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_2976),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2978),
.Y(n_3231)
);

BUFx2_ASAP7_75t_L g3232 ( 
.A(n_2960),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3004),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_2970),
.B(n_2918),
.Y(n_3234)
);

AOI21xp5_ASAP7_75t_L g3235 ( 
.A1(n_3009),
.A2(n_2839),
.B(n_2838),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3170),
.B(n_2846),
.Y(n_3236)
);

O2A1O1Ixp5_ASAP7_75t_L g3237 ( 
.A1(n_2953),
.A2(n_2902),
.B(n_2906),
.C(n_2895),
.Y(n_3237)
);

BUFx6f_ASAP7_75t_L g3238 ( 
.A(n_2957),
.Y(n_3238)
);

AOI21xp5_ASAP7_75t_L g3239 ( 
.A1(n_3009),
.A2(n_2842),
.B(n_2715),
.Y(n_3239)
);

AND2x2_ASAP7_75t_SL g3240 ( 
.A(n_3167),
.B(n_2844),
.Y(n_3240)
);

AOI21xp5_ASAP7_75t_L g3241 ( 
.A1(n_3065),
.A2(n_2876),
.B(n_2904),
.Y(n_3241)
);

AOI21xp5_ASAP7_75t_L g3242 ( 
.A1(n_3012),
.A2(n_2862),
.B(n_2858),
.Y(n_3242)
);

NAND2xp5_ASAP7_75t_L g3243 ( 
.A(n_2994),
.B(n_2943),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3023),
.A2(n_2981),
.B(n_2956),
.Y(n_3244)
);

AOI21xp5_ASAP7_75t_L g3245 ( 
.A1(n_3124),
.A2(n_2827),
.B(n_2907),
.Y(n_3245)
);

O2A1O1Ixp33_ASAP7_75t_L g3246 ( 
.A1(n_3153),
.A2(n_2908),
.B(n_2759),
.C(n_2938),
.Y(n_3246)
);

INVxp33_ASAP7_75t_SL g3247 ( 
.A(n_3081),
.Y(n_3247)
);

AOI21xp5_ASAP7_75t_L g3248 ( 
.A1(n_3125),
.A2(n_2942),
.B(n_2939),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2986),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_3027),
.B(n_7),
.Y(n_3250)
);

AOI21xp5_ASAP7_75t_L g3251 ( 
.A1(n_3127),
.A2(n_2234),
.B(n_2924),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3015),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_3073),
.B(n_2943),
.Y(n_3253)
);

AOI21xp5_ASAP7_75t_L g3254 ( 
.A1(n_3129),
.A2(n_3007),
.B(n_3162),
.Y(n_3254)
);

AOI221x1_ASAP7_75t_L g3255 ( 
.A1(n_2984),
.A2(n_2926),
.B1(n_2201),
.B2(n_2568),
.C(n_2555),
.Y(n_3255)
);

OAI22xp5_ASAP7_75t_L g3256 ( 
.A1(n_3005),
.A2(n_2669),
.B1(n_2568),
.B2(n_2555),
.Y(n_3256)
);

INVx3_ASAP7_75t_L g3257 ( 
.A(n_3059),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_2997),
.B(n_2996),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3146),
.B(n_2806),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_3061),
.B(n_2620),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_3013),
.B(n_2806),
.Y(n_3261)
);

INVx2_ASAP7_75t_L g3262 ( 
.A(n_3028),
.Y(n_3262)
);

OAI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_3099),
.A2(n_2223),
.B(n_2234),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_L g3264 ( 
.A(n_2991),
.B(n_2813),
.Y(n_3264)
);

OAI21xp5_ASAP7_75t_L g3265 ( 
.A1(n_3099),
.A2(n_2126),
.B(n_2111),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_SL g3266 ( 
.A(n_3013),
.B(n_2813),
.Y(n_3266)
);

NOR2xp67_ASAP7_75t_L g3267 ( 
.A(n_3085),
.B(n_3091),
.Y(n_3267)
);

O2A1O1Ixp33_ASAP7_75t_L g3268 ( 
.A1(n_2982),
.A2(n_2945),
.B(n_2243),
.C(n_2267),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_2992),
.B(n_2826),
.Y(n_3269)
);

AND2x4_ASAP7_75t_L g3270 ( 
.A(n_3068),
.B(n_2979),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_SL g3271 ( 
.A(n_2987),
.B(n_2826),
.Y(n_3271)
);

O2A1O1Ixp33_ASAP7_75t_L g3272 ( 
.A1(n_2985),
.A2(n_2263),
.B(n_2267),
.C(n_2299),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_3014),
.A2(n_2111),
.B(n_2087),
.Y(n_3273)
);

O2A1O1Ixp33_ASAP7_75t_L g3274 ( 
.A1(n_2966),
.A2(n_2967),
.B(n_3052),
.C(n_3050),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_SL g3275 ( 
.A(n_2987),
.B(n_2844),
.Y(n_3275)
);

HB1xp67_ASAP7_75t_L g3276 ( 
.A(n_3132),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_3082),
.B(n_2844),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3001),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_SL g3279 ( 
.A(n_3167),
.B(n_2877),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3021),
.B(n_2826),
.Y(n_3280)
);

NAND2xp5_ASAP7_75t_L g3281 ( 
.A(n_3025),
.B(n_2853),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_L g3282 ( 
.A(n_3030),
.B(n_2853),
.Y(n_3282)
);

O2A1O1Ixp33_ASAP7_75t_L g3283 ( 
.A1(n_2999),
.A2(n_2263),
.B(n_2267),
.C(n_2299),
.Y(n_3283)
);

NOR2xp33_ASAP7_75t_L g3284 ( 
.A(n_3017),
.B(n_2651),
.Y(n_3284)
);

AOI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_3160),
.A2(n_2052),
.B(n_2076),
.Y(n_3285)
);

NAND2xp5_ASAP7_75t_L g3286 ( 
.A(n_3031),
.B(n_3043),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3056),
.B(n_2853),
.Y(n_3287)
);

AOI21x1_ASAP7_75t_L g3288 ( 
.A1(n_3134),
.A2(n_1982),
.B(n_2076),
.Y(n_3288)
);

A2O1A1Ixp33_ASAP7_75t_L g3289 ( 
.A1(n_2948),
.A2(n_3053),
.B(n_3126),
.C(n_3057),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3042),
.Y(n_3290)
);

O2A1O1Ixp5_ASAP7_75t_L g3291 ( 
.A1(n_3084),
.A2(n_2600),
.B(n_2263),
.C(n_1994),
.Y(n_3291)
);

OAI21xp5_ASAP7_75t_L g3292 ( 
.A1(n_3157),
.A2(n_2126),
.B(n_2848),
.Y(n_3292)
);

AO21x1_ASAP7_75t_L g3293 ( 
.A1(n_3157),
.A2(n_2206),
.B(n_2117),
.Y(n_3293)
);

O2A1O1Ixp5_ASAP7_75t_L g3294 ( 
.A1(n_3062),
.A2(n_1994),
.B(n_1996),
.C(n_2206),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_SL g3295 ( 
.A(n_3068),
.B(n_2877),
.Y(n_3295)
);

A2O1A1Ixp33_ASAP7_75t_L g3296 ( 
.A1(n_3098),
.A2(n_2886),
.B(n_2918),
.C(n_2863),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3066),
.B(n_2863),
.Y(n_3297)
);

NAND2xp5_ASAP7_75t_L g3298 ( 
.A(n_3092),
.B(n_2863),
.Y(n_3298)
);

INVx2_ASAP7_75t_L g3299 ( 
.A(n_3047),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_3051),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_L g3301 ( 
.A(n_3093),
.B(n_3114),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3117),
.B(n_2886),
.Y(n_3302)
);

AO21x1_ASAP7_75t_L g3303 ( 
.A1(n_3040),
.A2(n_2848),
.B(n_1996),
.Y(n_3303)
);

BUFx6f_ASAP7_75t_L g3304 ( 
.A(n_2957),
.Y(n_3304)
);

AO21x2_ASAP7_75t_L g3305 ( 
.A1(n_3039),
.A2(n_2848),
.B(n_2202),
.Y(n_3305)
);

NAND2xp5_ASAP7_75t_L g3306 ( 
.A(n_3123),
.B(n_2886),
.Y(n_3306)
);

INVx3_ASAP7_75t_L g3307 ( 
.A(n_2988),
.Y(n_3307)
);

O2A1O1Ixp33_ASAP7_75t_L g3308 ( 
.A1(n_3038),
.A2(n_2052),
.B(n_2076),
.C(n_2202),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_3078),
.Y(n_3309)
);

BUFx6f_ASAP7_75t_L g3310 ( 
.A(n_3026),
.Y(n_3310)
);

AOI21xp5_ASAP7_75t_L g3311 ( 
.A1(n_2989),
.A2(n_2052),
.B(n_2381),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_SL g3312 ( 
.A(n_2973),
.B(n_2918),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_L g3313 ( 
.A(n_3139),
.B(n_2381),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_3144),
.B(n_2417),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_SL g3315 ( 
.A(n_2973),
.B(n_2417),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3142),
.B(n_3113),
.Y(n_3316)
);

NAND2xp5_ASAP7_75t_L g3317 ( 
.A(n_3145),
.B(n_2417),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_R g3318 ( 
.A(n_3060),
.B(n_2481),
.Y(n_3318)
);

AOI21xp5_ASAP7_75t_L g3319 ( 
.A1(n_3064),
.A2(n_2528),
.B(n_2481),
.Y(n_3319)
);

NOR3xp33_ASAP7_75t_L g3320 ( 
.A(n_3166),
.B(n_8),
.C(n_10),
.Y(n_3320)
);

HB1xp67_ASAP7_75t_L g3321 ( 
.A(n_3133),
.Y(n_3321)
);

NOR2xp33_ASAP7_75t_SL g3322 ( 
.A(n_3068),
.B(n_2848),
.Y(n_3322)
);

AOI21xp5_ASAP7_75t_L g3323 ( 
.A1(n_3143),
.A2(n_2528),
.B(n_2481),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2988),
.B(n_2528),
.Y(n_3324)
);

AOI21xp5_ASAP7_75t_L g3325 ( 
.A1(n_3029),
.A2(n_2565),
.B(n_2534),
.Y(n_3325)
);

AOI21xp5_ASAP7_75t_L g3326 ( 
.A1(n_3070),
.A2(n_2565),
.B(n_2534),
.Y(n_3326)
);

AOI21xp5_ASAP7_75t_L g3327 ( 
.A1(n_3002),
.A2(n_2565),
.B(n_2534),
.Y(n_3327)
);

AOI21xp5_ASAP7_75t_L g3328 ( 
.A1(n_3098),
.A2(n_2633),
.B(n_2611),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_3080),
.Y(n_3329)
);

OAI22xp5_ASAP7_75t_L g3330 ( 
.A1(n_2963),
.A2(n_2611),
.B1(n_2633),
.B2(n_2140),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_3106),
.B(n_2611),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_3086),
.Y(n_3332)
);

O2A1O1Ixp33_ASAP7_75t_SL g3333 ( 
.A1(n_3063),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_3333)
);

INVx2_ASAP7_75t_L g3334 ( 
.A(n_3087),
.Y(n_3334)
);

OAI21xp5_ASAP7_75t_L g3335 ( 
.A1(n_3067),
.A2(n_1737),
.B(n_1855),
.Y(n_3335)
);

OAI21xp5_ASAP7_75t_L g3336 ( 
.A1(n_3131),
.A2(n_1737),
.B(n_2633),
.Y(n_3336)
);

AOI21xp5_ASAP7_75t_L g3337 ( 
.A1(n_3089),
.A2(n_2146),
.B(n_2140),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_2969),
.B(n_14),
.Y(n_3338)
);

NOR2x2_ASAP7_75t_L g3339 ( 
.A(n_2979),
.B(n_14),
.Y(n_3339)
);

OAI21xp5_ASAP7_75t_L g3340 ( 
.A1(n_3071),
.A2(n_1737),
.B(n_2140),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3090),
.A2(n_2155),
.B(n_2146),
.Y(n_3341)
);

INVx3_ASAP7_75t_L g3342 ( 
.A(n_2988),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3111),
.B(n_2146),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3101),
.Y(n_3344)
);

BUFx3_ASAP7_75t_L g3345 ( 
.A(n_2995),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3116),
.B(n_2155),
.Y(n_3346)
);

AND2x2_ASAP7_75t_L g3347 ( 
.A(n_2993),
.B(n_15),
.Y(n_3347)
);

NAND2xp5_ASAP7_75t_SL g3348 ( 
.A(n_3048),
.B(n_2220),
.Y(n_3348)
);

AND2x2_ASAP7_75t_L g3349 ( 
.A(n_3036),
.B(n_15),
.Y(n_3349)
);

AOI21xp5_ASAP7_75t_L g3350 ( 
.A1(n_3100),
.A2(n_2184),
.B(n_2155),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_3108),
.Y(n_3351)
);

AOI21xp5_ASAP7_75t_L g3352 ( 
.A1(n_3102),
.A2(n_2184),
.B(n_2155),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3135),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_3136),
.Y(n_3354)
);

NOR2xp33_ASAP7_75t_L g3355 ( 
.A(n_3049),
.B(n_16),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_3048),
.B(n_2184),
.Y(n_3356)
);

AOI211xp5_ASAP7_75t_L g3357 ( 
.A1(n_3058),
.A2(n_2187),
.B(n_2208),
.C(n_2184),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_L g3358 ( 
.A(n_3118),
.B(n_2187),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3138),
.Y(n_3359)
);

AND2x2_ASAP7_75t_L g3360 ( 
.A(n_3072),
.B(n_16),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_3120),
.B(n_2187),
.Y(n_3361)
);

AOI21x1_ASAP7_75t_L g3362 ( 
.A1(n_3104),
.A2(n_2208),
.B(n_2187),
.Y(n_3362)
);

AOI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3115),
.A2(n_2213),
.B(n_2208),
.Y(n_3363)
);

BUFx6f_ASAP7_75t_L g3364 ( 
.A(n_3026),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3121),
.B(n_2208),
.Y(n_3365)
);

AOI21xp5_ASAP7_75t_L g3366 ( 
.A1(n_3130),
.A2(n_2220),
.B(n_2213),
.Y(n_3366)
);

O2A1O1Ixp5_ASAP7_75t_L g3367 ( 
.A1(n_3158),
.A2(n_2213),
.B(n_2220),
.C(n_1737),
.Y(n_3367)
);

O2A1O1Ixp33_ASAP7_75t_L g3368 ( 
.A1(n_3159),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_SL g3369 ( 
.A(n_3048),
.B(n_2213),
.Y(n_3369)
);

OAI21xp5_ASAP7_75t_L g3370 ( 
.A1(n_3140),
.A2(n_2220),
.B(n_1075),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3076),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_SL g3372 ( 
.A(n_3156),
.B(n_694),
.Y(n_3372)
);

AOI21xp5_ASAP7_75t_L g3373 ( 
.A1(n_3165),
.A2(n_18),
.B(n_19),
.Y(n_3373)
);

NOR2xp33_ASAP7_75t_L g3374 ( 
.A(n_3152),
.B(n_20),
.Y(n_3374)
);

AOI21xp5_ASAP7_75t_L g3375 ( 
.A1(n_3006),
.A2(n_20),
.B(n_21),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3077),
.B(n_22),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3079),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_3094),
.Y(n_3378)
);

NOR2x1p5_ASAP7_75t_L g3379 ( 
.A(n_3045),
.B(n_23),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3096),
.Y(n_3380)
);

CKINVDCx20_ASAP7_75t_R g3381 ( 
.A(n_2971),
.Y(n_3381)
);

BUFx2_ASAP7_75t_L g3382 ( 
.A(n_3276),
.Y(n_3382)
);

INVx1_ASAP7_75t_SL g3383 ( 
.A(n_3345),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_3203),
.A2(n_3037),
.B1(n_2977),
.B2(n_2979),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3182),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_3219),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3258),
.B(n_3074),
.Y(n_3387)
);

BUFx6f_ASAP7_75t_L g3388 ( 
.A(n_3238),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3193),
.B(n_3119),
.Y(n_3389)
);

INVx3_ASAP7_75t_L g3390 ( 
.A(n_3270),
.Y(n_3390)
);

INVx1_ASAP7_75t_L g3391 ( 
.A(n_3186),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3199),
.Y(n_3392)
);

BUFx4f_ASAP7_75t_L g3393 ( 
.A(n_3238),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_3179),
.B(n_3074),
.Y(n_3394)
);

AND2x2_ASAP7_75t_L g3395 ( 
.A(n_3193),
.B(n_3045),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3180),
.Y(n_3396)
);

INVx1_ASAP7_75t_L g3397 ( 
.A(n_3207),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_3225),
.Y(n_3398)
);

INVx5_ASAP7_75t_L g3399 ( 
.A(n_3270),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3230),
.Y(n_3400)
);

INVx2_ASAP7_75t_L g3401 ( 
.A(n_3226),
.Y(n_3401)
);

AND2x2_ASAP7_75t_L g3402 ( 
.A(n_3194),
.B(n_3069),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3210),
.B(n_3188),
.Y(n_3403)
);

INVx2_ASAP7_75t_L g3404 ( 
.A(n_3233),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_3231),
.Y(n_3405)
);

NOR2xp67_ASAP7_75t_L g3406 ( 
.A(n_3267),
.B(n_3088),
.Y(n_3406)
);

AND2x4_ASAP7_75t_L g3407 ( 
.A(n_3321),
.B(n_3088),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3189),
.B(n_3103),
.Y(n_3408)
);

INVx2_ASAP7_75t_L g3409 ( 
.A(n_3252),
.Y(n_3409)
);

OR2x6_ASAP7_75t_L g3410 ( 
.A(n_3229),
.B(n_3026),
.Y(n_3410)
);

OR2x6_ASAP7_75t_L g3411 ( 
.A(n_3234),
.B(n_3151),
.Y(n_3411)
);

OAI22xp5_ASAP7_75t_L g3412 ( 
.A1(n_3184),
.A2(n_3169),
.B1(n_3171),
.B2(n_3164),
.Y(n_3412)
);

BUFx12f_ASAP7_75t_L g3413 ( 
.A(n_3238),
.Y(n_3413)
);

INVxp67_ASAP7_75t_L g3414 ( 
.A(n_3253),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3202),
.B(n_3109),
.Y(n_3415)
);

INVx3_ASAP7_75t_L g3416 ( 
.A(n_3307),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3249),
.Y(n_3417)
);

INVx3_ASAP7_75t_L g3418 ( 
.A(n_3304),
.Y(n_3418)
);

BUFx2_ASAP7_75t_L g3419 ( 
.A(n_3318),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3204),
.B(n_3069),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3262),
.Y(n_3421)
);

AND2x2_ASAP7_75t_L g3422 ( 
.A(n_3316),
.B(n_3156),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3278),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_3290),
.Y(n_3424)
);

AND2x4_ASAP7_75t_L g3425 ( 
.A(n_3259),
.B(n_3148),
.Y(n_3425)
);

INVx1_ASAP7_75t_L g3426 ( 
.A(n_3286),
.Y(n_3426)
);

INVx2_ASAP7_75t_L g3427 ( 
.A(n_3299),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3206),
.B(n_3195),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3301),
.Y(n_3429)
);

NAND2xp5_ASAP7_75t_L g3430 ( 
.A(n_3183),
.B(n_2977),
.Y(n_3430)
);

INVx3_ASAP7_75t_L g3431 ( 
.A(n_3307),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3213),
.B(n_2977),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3224),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3300),
.Y(n_3434)
);

BUFx3_ASAP7_75t_L g3435 ( 
.A(n_3381),
.Y(n_3435)
);

INVx1_ASAP7_75t_SL g3436 ( 
.A(n_3218),
.Y(n_3436)
);

INVx4_ASAP7_75t_L g3437 ( 
.A(n_3304),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_3187),
.B(n_2977),
.Y(n_3438)
);

AOI22xp5_ASAP7_75t_L g3439 ( 
.A1(n_3196),
.A2(n_3147),
.B1(n_3105),
.B2(n_3148),
.Y(n_3439)
);

O2A1O1Ixp33_ASAP7_75t_L g3440 ( 
.A1(n_3320),
.A2(n_3095),
.B(n_3112),
.C(n_3083),
.Y(n_3440)
);

OR2x6_ASAP7_75t_L g3441 ( 
.A(n_3379),
.B(n_3156),
.Y(n_3441)
);

AND2x4_ASAP7_75t_L g3442 ( 
.A(n_3222),
.B(n_3149),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_SL g3443 ( 
.A(n_3232),
.B(n_3149),
.Y(n_3443)
);

OR2x6_ASAP7_75t_L g3444 ( 
.A(n_3271),
.B(n_3122),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3309),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3378),
.Y(n_3446)
);

BUFx8_ASAP7_75t_L g3447 ( 
.A(n_3304),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3329),
.Y(n_3448)
);

INVx3_ASAP7_75t_L g3449 ( 
.A(n_3342),
.Y(n_3449)
);

BUFx6f_ASAP7_75t_L g3450 ( 
.A(n_3310),
.Y(n_3450)
);

INVx5_ASAP7_75t_L g3451 ( 
.A(n_3310),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3190),
.B(n_24),
.Y(n_3452)
);

INVx2_ASAP7_75t_L g3453 ( 
.A(n_3334),
.Y(n_3453)
);

NOR2xp33_ASAP7_75t_L g3454 ( 
.A(n_3247),
.B(n_24),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3332),
.Y(n_3455)
);

AND2x4_ASAP7_75t_L g3456 ( 
.A(n_3275),
.B(n_669),
.Y(n_3456)
);

OR2x6_ASAP7_75t_L g3457 ( 
.A(n_3192),
.B(n_588),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_3310),
.Y(n_3458)
);

INVx5_ASAP7_75t_L g3459 ( 
.A(n_3364),
.Y(n_3459)
);

NAND2xp5_ASAP7_75t_L g3460 ( 
.A(n_3217),
.B(n_26),
.Y(n_3460)
);

HB1xp67_ASAP7_75t_L g3461 ( 
.A(n_3243),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3220),
.B(n_27),
.Y(n_3462)
);

INVx2_ASAP7_75t_L g3463 ( 
.A(n_3351),
.Y(n_3463)
);

NAND2xp5_ASAP7_75t_L g3464 ( 
.A(n_3371),
.B(n_27),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3359),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3344),
.Y(n_3466)
);

BUFx12f_ASAP7_75t_L g3467 ( 
.A(n_3364),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3353),
.Y(n_3468)
);

BUFx6f_ASAP7_75t_L g3469 ( 
.A(n_3364),
.Y(n_3469)
);

INVx2_ASAP7_75t_L g3470 ( 
.A(n_3354),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_3377),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3380),
.B(n_28),
.Y(n_3472)
);

NOR2xp67_ASAP7_75t_L g3473 ( 
.A(n_3214),
.B(n_28),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3313),
.Y(n_3474)
);

INVx5_ASAP7_75t_L g3475 ( 
.A(n_3181),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_3314),
.Y(n_3476)
);

AND2x4_ASAP7_75t_L g3477 ( 
.A(n_3342),
.B(n_681),
.Y(n_3477)
);

OR2x2_ASAP7_75t_L g3478 ( 
.A(n_3197),
.B(n_29),
.Y(n_3478)
);

NAND2xp33_ASAP7_75t_SL g3479 ( 
.A(n_3209),
.B(n_29),
.Y(n_3479)
);

OR2x6_ASAP7_75t_L g3480 ( 
.A(n_3274),
.B(n_591),
.Y(n_3480)
);

AOI21xp5_ASAP7_75t_L g3481 ( 
.A1(n_3178),
.A2(n_32),
.B(n_31),
.Y(n_3481)
);

INVx1_ASAP7_75t_L g3482 ( 
.A(n_3317),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_L g3483 ( 
.A(n_3236),
.B(n_30),
.Y(n_3483)
);

NAND2xp5_ASAP7_75t_L g3484 ( 
.A(n_3212),
.B(n_31),
.Y(n_3484)
);

BUFx6f_ASAP7_75t_L g3485 ( 
.A(n_3240),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3264),
.B(n_32),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3269),
.B(n_33),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3280),
.Y(n_3488)
);

AOI22xp5_ASAP7_75t_L g3489 ( 
.A1(n_3211),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3281),
.B(n_34),
.Y(n_3490)
);

NAND2xp5_ASAP7_75t_SL g3491 ( 
.A(n_3172),
.B(n_592),
.Y(n_3491)
);

NAND2x1p5_ASAP7_75t_L g3492 ( 
.A(n_3312),
.B(n_594),
.Y(n_3492)
);

AND2x6_ASAP7_75t_L g3493 ( 
.A(n_3191),
.B(n_599),
.Y(n_3493)
);

INVx1_ASAP7_75t_L g3494 ( 
.A(n_3282),
.Y(n_3494)
);

NOR2xp67_ASAP7_75t_L g3495 ( 
.A(n_3284),
.B(n_3260),
.Y(n_3495)
);

BUFx2_ASAP7_75t_L g3496 ( 
.A(n_3287),
.Y(n_3496)
);

NOR2xp33_ASAP7_75t_L g3497 ( 
.A(n_3338),
.B(n_35),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_3297),
.B(n_36),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_L g3499 ( 
.A(n_3298),
.B(n_38),
.Y(n_3499)
);

AND2x4_ASAP7_75t_L g3500 ( 
.A(n_3261),
.B(n_674),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3302),
.B(n_38),
.Y(n_3501)
);

BUFx2_ASAP7_75t_L g3502 ( 
.A(n_3306),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3343),
.Y(n_3503)
);

INVx5_ASAP7_75t_L g3504 ( 
.A(n_3181),
.Y(n_3504)
);

INVx4_ASAP7_75t_L g3505 ( 
.A(n_3185),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3346),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3358),
.Y(n_3507)
);

AOI22x1_ASAP7_75t_L g3508 ( 
.A1(n_3373),
.A2(n_42),
.B1(n_39),
.B2(n_41),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3361),
.Y(n_3509)
);

BUFx2_ASAP7_75t_L g3510 ( 
.A(n_3331),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3174),
.B(n_42),
.Y(n_3511)
);

INVxp67_ASAP7_75t_SL g3512 ( 
.A(n_3293),
.Y(n_3512)
);

INVx4_ASAP7_75t_L g3513 ( 
.A(n_3185),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3365),
.Y(n_3514)
);

INVx5_ASAP7_75t_L g3515 ( 
.A(n_3257),
.Y(n_3515)
);

CKINVDCx20_ASAP7_75t_R g3516 ( 
.A(n_3349),
.Y(n_3516)
);

OAI22xp5_ASAP7_75t_SL g3517 ( 
.A1(n_3355),
.A2(n_52),
.B1(n_60),
.B2(n_43),
.Y(n_3517)
);

AOI22xp33_ASAP7_75t_L g3518 ( 
.A1(n_3208),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3254),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3376),
.Y(n_3520)
);

BUFx6f_ASAP7_75t_L g3521 ( 
.A(n_3257),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3305),
.Y(n_3522)
);

OR2x2_ASAP7_75t_L g3523 ( 
.A(n_3250),
.B(n_47),
.Y(n_3523)
);

INVx3_ASAP7_75t_L g3524 ( 
.A(n_3362),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_SL g3525 ( 
.A(n_3205),
.B(n_600),
.Y(n_3525)
);

HB1xp67_ASAP7_75t_L g3526 ( 
.A(n_3216),
.Y(n_3526)
);

AND2x6_ASAP7_75t_L g3527 ( 
.A(n_3215),
.B(n_601),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3177),
.B(n_48),
.Y(n_3528)
);

NAND2xp5_ASAP7_75t_L g3529 ( 
.A(n_3244),
.B(n_48),
.Y(n_3529)
);

INVx2_ASAP7_75t_L g3530 ( 
.A(n_3305),
.Y(n_3530)
);

NAND2xp5_ASAP7_75t_L g3531 ( 
.A(n_3374),
.B(n_49),
.Y(n_3531)
);

A2O1A1Ixp33_ASAP7_75t_L g3532 ( 
.A1(n_3289),
.A2(n_52),
.B(n_50),
.C(n_51),
.Y(n_3532)
);

INVx3_ASAP7_75t_L g3533 ( 
.A(n_3360),
.Y(n_3533)
);

CKINVDCx5p33_ASAP7_75t_R g3534 ( 
.A(n_3347),
.Y(n_3534)
);

INVx3_ASAP7_75t_L g3535 ( 
.A(n_3288),
.Y(n_3535)
);

INVx2_ASAP7_75t_L g3536 ( 
.A(n_3294),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3303),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3266),
.Y(n_3538)
);

BUFx2_ASAP7_75t_L g3539 ( 
.A(n_3336),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3291),
.Y(n_3540)
);

HB1xp67_ASAP7_75t_L g3541 ( 
.A(n_3336),
.Y(n_3541)
);

NOR2xp33_ASAP7_75t_L g3542 ( 
.A(n_3277),
.B(n_50),
.Y(n_3542)
);

AND3x1_ASAP7_75t_L g3543 ( 
.A(n_3339),
.B(n_51),
.C(n_53),
.Y(n_3543)
);

INVx2_ASAP7_75t_L g3544 ( 
.A(n_3237),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3248),
.Y(n_3545)
);

INVx3_ASAP7_75t_L g3546 ( 
.A(n_3173),
.Y(n_3546)
);

NAND2xp5_ASAP7_75t_L g3547 ( 
.A(n_3227),
.B(n_53),
.Y(n_3547)
);

AND3x1_ASAP7_75t_SL g3548 ( 
.A(n_3368),
.B(n_54),
.C(n_55),
.Y(n_3548)
);

INVx3_ASAP7_75t_L g3549 ( 
.A(n_3322),
.Y(n_3549)
);

OR2x2_ASAP7_75t_L g3550 ( 
.A(n_3330),
.B(n_3296),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3245),
.Y(n_3551)
);

INVx4_ASAP7_75t_L g3552 ( 
.A(n_3324),
.Y(n_3552)
);

INVx1_ASAP7_75t_SL g3553 ( 
.A(n_3315),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3201),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3200),
.B(n_54),
.Y(n_3555)
);

INVx2_ASAP7_75t_SL g3556 ( 
.A(n_3348),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3241),
.Y(n_3557)
);

BUFx6f_ASAP7_75t_L g3558 ( 
.A(n_3356),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3369),
.Y(n_3559)
);

INVx3_ASAP7_75t_L g3560 ( 
.A(n_3322),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3367),
.Y(n_3561)
);

AND2x4_ASAP7_75t_L g3562 ( 
.A(n_3176),
.B(n_678),
.Y(n_3562)
);

NAND2xp5_ASAP7_75t_L g3563 ( 
.A(n_3235),
.B(n_55),
.Y(n_3563)
);

NAND2xp5_ASAP7_75t_L g3564 ( 
.A(n_3242),
.B(n_3175),
.Y(n_3564)
);

INVx3_ASAP7_75t_L g3565 ( 
.A(n_3295),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3256),
.Y(n_3566)
);

AOI22xp33_ASAP7_75t_L g3567 ( 
.A1(n_3198),
.A2(n_58),
.B1(n_56),
.B2(n_57),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_3308),
.Y(n_3568)
);

HB1xp67_ASAP7_75t_L g3569 ( 
.A(n_3292),
.Y(n_3569)
);

INVx2_ASAP7_75t_L g3570 ( 
.A(n_3372),
.Y(n_3570)
);

BUFx6f_ASAP7_75t_L g3571 ( 
.A(n_3295),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3221),
.B(n_57),
.Y(n_3572)
);

A2O1A1Ixp33_ASAP7_75t_L g3573 ( 
.A1(n_3198),
.A2(n_60),
.B(n_58),
.C(n_59),
.Y(n_3573)
);

INVx2_ASAP7_75t_L g3574 ( 
.A(n_3263),
.Y(n_3574)
);

INVx4_ASAP7_75t_SL g3575 ( 
.A(n_3205),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_SL g3576 ( 
.A(n_3357),
.B(n_602),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3251),
.Y(n_3577)
);

INVx2_ASAP7_75t_L g3578 ( 
.A(n_3263),
.Y(n_3578)
);

NAND2xp5_ASAP7_75t_L g3579 ( 
.A(n_3223),
.B(n_61),
.Y(n_3579)
);

HB1xp67_ASAP7_75t_L g3580 ( 
.A(n_3292),
.Y(n_3580)
);

INVx4_ASAP7_75t_L g3581 ( 
.A(n_3246),
.Y(n_3581)
);

INVx1_ASAP7_75t_L g3582 ( 
.A(n_3370),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3370),
.Y(n_3583)
);

CKINVDCx16_ASAP7_75t_R g3584 ( 
.A(n_3279),
.Y(n_3584)
);

AOI22xp5_ASAP7_75t_L g3585 ( 
.A1(n_3279),
.A2(n_3335),
.B1(n_3375),
.B2(n_3333),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_L g3586 ( 
.A(n_3228),
.B(n_61),
.Y(n_3586)
);

NAND2xp5_ASAP7_75t_L g3587 ( 
.A(n_3319),
.B(n_63),
.Y(n_3587)
);

INVx2_ASAP7_75t_L g3588 ( 
.A(n_3335),
.Y(n_3588)
);

CKINVDCx5p33_ASAP7_75t_R g3589 ( 
.A(n_3327),
.Y(n_3589)
);

INVx3_ASAP7_75t_L g3590 ( 
.A(n_3328),
.Y(n_3590)
);

BUFx2_ASAP7_75t_L g3591 ( 
.A(n_3382),
.Y(n_3591)
);

NOR2xp33_ASAP7_75t_L g3592 ( 
.A(n_3383),
.B(n_63),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3402),
.B(n_3340),
.Y(n_3593)
);

INVx4_ASAP7_75t_L g3594 ( 
.A(n_3413),
.Y(n_3594)
);

A2O1A1Ixp33_ASAP7_75t_L g3595 ( 
.A1(n_3532),
.A2(n_3479),
.B(n_3481),
.C(n_3572),
.Y(n_3595)
);

INVx6_ASAP7_75t_L g3596 ( 
.A(n_3447),
.Y(n_3596)
);

HB1xp67_ASAP7_75t_L g3597 ( 
.A(n_3510),
.Y(n_3597)
);

INVx3_ASAP7_75t_L g3598 ( 
.A(n_3467),
.Y(n_3598)
);

INVx2_ASAP7_75t_SL g3599 ( 
.A(n_3419),
.Y(n_3599)
);

CKINVDCx20_ASAP7_75t_R g3600 ( 
.A(n_3435),
.Y(n_3600)
);

AOI21xp5_ASAP7_75t_L g3601 ( 
.A1(n_3564),
.A2(n_3255),
.B(n_3268),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3385),
.Y(n_3602)
);

NAND2x1_ASAP7_75t_SL g3603 ( 
.A(n_3581),
.B(n_3283),
.Y(n_3603)
);

INVx3_ASAP7_75t_L g3604 ( 
.A(n_3447),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3396),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3470),
.Y(n_3606)
);

NAND2xp5_ASAP7_75t_L g3607 ( 
.A(n_3403),
.B(n_3239),
.Y(n_3607)
);

HB1xp67_ASAP7_75t_L g3608 ( 
.A(n_3526),
.Y(n_3608)
);

BUFx6f_ASAP7_75t_L g3609 ( 
.A(n_3410),
.Y(n_3609)
);

OR2x2_ASAP7_75t_L g3610 ( 
.A(n_3391),
.B(n_3323),
.Y(n_3610)
);

OAI22x1_ASAP7_75t_L g3611 ( 
.A1(n_3497),
.A2(n_3387),
.B1(n_3384),
.B2(n_3520),
.Y(n_3611)
);

INVx2_ASAP7_75t_SL g3612 ( 
.A(n_3436),
.Y(n_3612)
);

INVx1_ASAP7_75t_L g3613 ( 
.A(n_3392),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_3397),
.Y(n_3614)
);

BUFx6f_ASAP7_75t_L g3615 ( 
.A(n_3410),
.Y(n_3615)
);

OAI21x1_ASAP7_75t_L g3616 ( 
.A1(n_3535),
.A2(n_3285),
.B(n_3273),
.Y(n_3616)
);

AOI22xp33_ASAP7_75t_L g3617 ( 
.A1(n_3527),
.A2(n_3326),
.B1(n_3311),
.B2(n_3325),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_SL g3618 ( 
.A(n_3495),
.B(n_3337),
.Y(n_3618)
);

AOI22xp5_ASAP7_75t_L g3619 ( 
.A1(n_3527),
.A2(n_3341),
.B1(n_3352),
.B2(n_3350),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_3398),
.Y(n_3620)
);

AOI21xp5_ASAP7_75t_SL g3621 ( 
.A1(n_3480),
.A2(n_3272),
.B(n_3265),
.Y(n_3621)
);

INVx1_ASAP7_75t_L g3622 ( 
.A(n_3400),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_3405),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3480),
.A2(n_3265),
.B(n_3363),
.Y(n_3624)
);

INVx1_ASAP7_75t_SL g3625 ( 
.A(n_3534),
.Y(n_3625)
);

CKINVDCx5p33_ASAP7_75t_R g3626 ( 
.A(n_3516),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3471),
.Y(n_3627)
);

BUFx2_ASAP7_75t_L g3628 ( 
.A(n_3407),
.Y(n_3628)
);

AOI22xp5_ASAP7_75t_L g3629 ( 
.A1(n_3527),
.A2(n_3366),
.B1(n_66),
.B2(n_64),
.Y(n_3629)
);

NAND2xp5_ASAP7_75t_L g3630 ( 
.A(n_3428),
.B(n_64),
.Y(n_3630)
);

AOI22xp33_ASAP7_75t_L g3631 ( 
.A1(n_3493),
.A2(n_67),
.B1(n_65),
.B2(n_66),
.Y(n_3631)
);

INVx2_ASAP7_75t_L g3632 ( 
.A(n_3455),
.Y(n_3632)
);

INVx2_ASAP7_75t_L g3633 ( 
.A(n_3466),
.Y(n_3633)
);

BUFx2_ASAP7_75t_L g3634 ( 
.A(n_3407),
.Y(n_3634)
);

INVx8_ASAP7_75t_L g3635 ( 
.A(n_3441),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3417),
.Y(n_3636)
);

NAND2xp5_ASAP7_75t_SL g3637 ( 
.A(n_3589),
.B(n_65),
.Y(n_3637)
);

INVx1_ASAP7_75t_L g3638 ( 
.A(n_3423),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3468),
.Y(n_3639)
);

BUFx6f_ASAP7_75t_L g3640 ( 
.A(n_3388),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_3386),
.Y(n_3641)
);

INVx4_ASAP7_75t_L g3642 ( 
.A(n_3388),
.Y(n_3642)
);

AND2x4_ASAP7_75t_L g3643 ( 
.A(n_3399),
.B(n_3390),
.Y(n_3643)
);

INVx1_ASAP7_75t_L g3644 ( 
.A(n_3426),
.Y(n_3644)
);

NOR2xp33_ASAP7_75t_L g3645 ( 
.A(n_3454),
.B(n_67),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3394),
.B(n_68),
.Y(n_3646)
);

INVxp67_ASAP7_75t_L g3647 ( 
.A(n_3461),
.Y(n_3647)
);

NOR2xp33_ASAP7_75t_L g3648 ( 
.A(n_3531),
.B(n_69),
.Y(n_3648)
);

BUFx6f_ASAP7_75t_L g3649 ( 
.A(n_3388),
.Y(n_3649)
);

INVx1_ASAP7_75t_SL g3650 ( 
.A(n_3422),
.Y(n_3650)
);

BUFx2_ASAP7_75t_L g3651 ( 
.A(n_3395),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_3401),
.Y(n_3652)
);

AND2x4_ASAP7_75t_L g3653 ( 
.A(n_3399),
.B(n_69),
.Y(n_3653)
);

O2A1O1Ixp33_ASAP7_75t_L g3654 ( 
.A1(n_3579),
.A2(n_72),
.B(n_70),
.C(n_71),
.Y(n_3654)
);

BUFx12f_ASAP7_75t_L g3655 ( 
.A(n_3450),
.Y(n_3655)
);

INVx5_ASAP7_75t_L g3656 ( 
.A(n_3493),
.Y(n_3656)
);

INVx3_ASAP7_75t_SL g3657 ( 
.A(n_3442),
.Y(n_3657)
);

INVx2_ASAP7_75t_L g3658 ( 
.A(n_3404),
.Y(n_3658)
);

BUFx6f_ASAP7_75t_L g3659 ( 
.A(n_3450),
.Y(n_3659)
);

INVx1_ASAP7_75t_L g3660 ( 
.A(n_3429),
.Y(n_3660)
);

BUFx6f_ASAP7_75t_L g3661 ( 
.A(n_3450),
.Y(n_3661)
);

AO21x2_ASAP7_75t_L g3662 ( 
.A1(n_3537),
.A2(n_71),
.B(n_72),
.Y(n_3662)
);

INVx2_ASAP7_75t_SL g3663 ( 
.A(n_3389),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3474),
.Y(n_3664)
);

INVx4_ASAP7_75t_L g3665 ( 
.A(n_3458),
.Y(n_3665)
);

AOI22xp5_ASAP7_75t_L g3666 ( 
.A1(n_3493),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_3666)
);

AND2x4_ASAP7_75t_L g3667 ( 
.A(n_3399),
.B(n_73),
.Y(n_3667)
);

BUFx8_ASAP7_75t_L g3668 ( 
.A(n_3458),
.Y(n_3668)
);

AOI22xp33_ASAP7_75t_L g3669 ( 
.A1(n_3444),
.A2(n_76),
.B1(n_74),
.B2(n_75),
.Y(n_3669)
);

A2O1A1Ixp33_ASAP7_75t_L g3670 ( 
.A1(n_3573),
.A2(n_78),
.B(n_76),
.C(n_77),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3476),
.Y(n_3671)
);

BUFx2_ASAP7_75t_L g3672 ( 
.A(n_3442),
.Y(n_3672)
);

BUFx6f_ASAP7_75t_L g3673 ( 
.A(n_3458),
.Y(n_3673)
);

AO221x1_ASAP7_75t_L g3674 ( 
.A1(n_3517),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.C(n_82),
.Y(n_3674)
);

INVx4_ASAP7_75t_L g3675 ( 
.A(n_3469),
.Y(n_3675)
);

AOI22xp33_ASAP7_75t_L g3676 ( 
.A1(n_3444),
.A2(n_81),
.B1(n_79),
.B2(n_80),
.Y(n_3676)
);

BUFx12f_ASAP7_75t_L g3677 ( 
.A(n_3469),
.Y(n_3677)
);

BUFx2_ASAP7_75t_L g3678 ( 
.A(n_3390),
.Y(n_3678)
);

AND2x4_ASAP7_75t_L g3679 ( 
.A(n_3575),
.B(n_82),
.Y(n_3679)
);

CKINVDCx5p33_ASAP7_75t_R g3680 ( 
.A(n_3469),
.Y(n_3680)
);

INVx1_ASAP7_75t_SL g3681 ( 
.A(n_3496),
.Y(n_3681)
);

INVx2_ASAP7_75t_SL g3682 ( 
.A(n_3451),
.Y(n_3682)
);

AO22x1_ASAP7_75t_L g3683 ( 
.A1(n_3485),
.A2(n_85),
.B1(n_83),
.B2(n_84),
.Y(n_3683)
);

NOR2xp67_ASAP7_75t_L g3684 ( 
.A(n_3581),
.B(n_83),
.Y(n_3684)
);

INVx2_ASAP7_75t_SL g3685 ( 
.A(n_3451),
.Y(n_3685)
);

OR2x2_ASAP7_75t_L g3686 ( 
.A(n_3408),
.B(n_85),
.Y(n_3686)
);

INVx1_ASAP7_75t_L g3687 ( 
.A(n_3482),
.Y(n_3687)
);

CKINVDCx20_ASAP7_75t_R g3688 ( 
.A(n_3502),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3409),
.Y(n_3689)
);

AOI21xp5_ASAP7_75t_L g3690 ( 
.A1(n_3586),
.A2(n_86),
.B(n_87),
.Y(n_3690)
);

INVx4_ASAP7_75t_L g3691 ( 
.A(n_3393),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3420),
.B(n_86),
.Y(n_3692)
);

AOI21xp5_ASAP7_75t_L g3693 ( 
.A1(n_3525),
.A2(n_87),
.B(n_88),
.Y(n_3693)
);

AND2x4_ASAP7_75t_L g3694 ( 
.A(n_3575),
.B(n_88),
.Y(n_3694)
);

INVx3_ASAP7_75t_L g3695 ( 
.A(n_3437),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3421),
.Y(n_3696)
);

INVx3_ASAP7_75t_L g3697 ( 
.A(n_3437),
.Y(n_3697)
);

INVx2_ASAP7_75t_L g3698 ( 
.A(n_3424),
.Y(n_3698)
);

AOI22xp33_ASAP7_75t_L g3699 ( 
.A1(n_3508),
.A2(n_91),
.B1(n_89),
.B2(n_90),
.Y(n_3699)
);

BUFx2_ASAP7_75t_L g3700 ( 
.A(n_3425),
.Y(n_3700)
);

BUFx2_ASAP7_75t_L g3701 ( 
.A(n_3425),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3433),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3503),
.Y(n_3703)
);

BUFx6f_ASAP7_75t_L g3704 ( 
.A(n_3451),
.Y(n_3704)
);

AOI21xp5_ASAP7_75t_L g3705 ( 
.A1(n_3576),
.A2(n_89),
.B(n_90),
.Y(n_3705)
);

AOI22xp5_ASAP7_75t_L g3706 ( 
.A1(n_3548),
.A2(n_93),
.B1(n_91),
.B2(n_92),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3533),
.B(n_92),
.Y(n_3707)
);

AOI21xp5_ASAP7_75t_L g3708 ( 
.A1(n_3557),
.A2(n_93),
.B(n_94),
.Y(n_3708)
);

CKINVDCx5p33_ASAP7_75t_R g3709 ( 
.A(n_3418),
.Y(n_3709)
);

AND2x4_ASAP7_75t_L g3710 ( 
.A(n_3539),
.B(n_96),
.Y(n_3710)
);

AND2x4_ASAP7_75t_L g3711 ( 
.A(n_3565),
.B(n_96),
.Y(n_3711)
);

NAND3xp33_ASAP7_75t_SL g3712 ( 
.A(n_3528),
.B(n_97),
.C(n_98),
.Y(n_3712)
);

NOR2xp33_ASAP7_75t_L g3713 ( 
.A(n_3523),
.B(n_97),
.Y(n_3713)
);

BUFx3_ASAP7_75t_L g3714 ( 
.A(n_3485),
.Y(n_3714)
);

O2A1O1Ixp33_ASAP7_75t_L g3715 ( 
.A1(n_3529),
.A2(n_101),
.B(n_99),
.C(n_100),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3507),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3427),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3434),
.Y(n_3718)
);

INVx2_ASAP7_75t_L g3719 ( 
.A(n_3445),
.Y(n_3719)
);

CKINVDCx5p33_ASAP7_75t_R g3720 ( 
.A(n_3414),
.Y(n_3720)
);

NOR2xp33_ASAP7_75t_L g3721 ( 
.A(n_3484),
.B(n_99),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3509),
.Y(n_3722)
);

BUFx2_ASAP7_75t_L g3723 ( 
.A(n_3416),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3569),
.B(n_101),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3448),
.Y(n_3725)
);

A2O1A1Ixp33_ASAP7_75t_L g3726 ( 
.A1(n_3473),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_3726)
);

BUFx6f_ASAP7_75t_L g3727 ( 
.A(n_3459),
.Y(n_3727)
);

INVxp67_ASAP7_75t_SL g3728 ( 
.A(n_3519),
.Y(n_3728)
);

OAI22xp5_ASAP7_75t_SL g3729 ( 
.A1(n_3543),
.A2(n_104),
.B1(n_102),
.B2(n_103),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3547),
.A2(n_105),
.B(n_106),
.Y(n_3730)
);

BUFx6f_ASAP7_75t_L g3731 ( 
.A(n_3459),
.Y(n_3731)
);

BUFx12f_ASAP7_75t_L g3732 ( 
.A(n_3478),
.Y(n_3732)
);

AND2x2_ASAP7_75t_L g3733 ( 
.A(n_3580),
.B(n_105),
.Y(n_3733)
);

NAND2x1p5_ASAP7_75t_L g3734 ( 
.A(n_3459),
.B(n_603),
.Y(n_3734)
);

NOR2xp33_ASAP7_75t_L g3735 ( 
.A(n_3483),
.B(n_106),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3514),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3506),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3446),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_SL g3739 ( 
.A(n_3406),
.B(n_107),
.Y(n_3739)
);

NAND2x1p5_ASAP7_75t_L g3740 ( 
.A(n_3485),
.B(n_605),
.Y(n_3740)
);

BUFx2_ASAP7_75t_L g3741 ( 
.A(n_3416),
.Y(n_3741)
);

OAI22xp5_ASAP7_75t_L g3742 ( 
.A1(n_3567),
.A2(n_109),
.B1(n_107),
.B2(n_108),
.Y(n_3742)
);

AOI22xp33_ASAP7_75t_L g3743 ( 
.A1(n_3554),
.A2(n_111),
.B1(n_109),
.B2(n_110),
.Y(n_3743)
);

AOI22xp33_ASAP7_75t_L g3744 ( 
.A1(n_3544),
.A2(n_112),
.B1(n_110),
.B2(n_111),
.Y(n_3744)
);

AND2x4_ASAP7_75t_L g3745 ( 
.A(n_3565),
.B(n_112),
.Y(n_3745)
);

AOI21xp5_ASAP7_75t_L g3746 ( 
.A1(n_3568),
.A2(n_113),
.B(n_114),
.Y(n_3746)
);

AOI22xp5_ASAP7_75t_L g3747 ( 
.A1(n_3489),
.A2(n_115),
.B1(n_113),
.B2(n_114),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_3488),
.B(n_115),
.Y(n_3748)
);

INVx3_ASAP7_75t_L g3749 ( 
.A(n_3521),
.Y(n_3749)
);

BUFx3_ASAP7_75t_L g3750 ( 
.A(n_3521),
.Y(n_3750)
);

INVxp67_ASAP7_75t_L g3751 ( 
.A(n_3460),
.Y(n_3751)
);

INVx1_ASAP7_75t_SL g3752 ( 
.A(n_3441),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3494),
.Y(n_3753)
);

AND2x4_ASAP7_75t_L g3754 ( 
.A(n_3571),
.B(n_116),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3453),
.Y(n_3755)
);

AOI21xp5_ASAP7_75t_L g3756 ( 
.A1(n_3545),
.A2(n_117),
.B(n_120),
.Y(n_3756)
);

OAI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_3518),
.A2(n_122),
.B1(n_120),
.B2(n_121),
.Y(n_3757)
);

OAI22xp5_ASAP7_75t_L g3758 ( 
.A1(n_3555),
.A2(n_124),
.B1(n_121),
.B2(n_123),
.Y(n_3758)
);

INVx3_ASAP7_75t_SL g3759 ( 
.A(n_3457),
.Y(n_3759)
);

OAI22xp5_ASAP7_75t_L g3760 ( 
.A1(n_3585),
.A2(n_126),
.B1(n_124),
.B2(n_125),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3463),
.Y(n_3761)
);

OAI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_3563),
.A2(n_129),
.B1(n_126),
.B2(n_128),
.Y(n_3762)
);

OAI22xp5_ASAP7_75t_L g3763 ( 
.A1(n_3542),
.A2(n_131),
.B1(n_128),
.B2(n_129),
.Y(n_3763)
);

INVx2_ASAP7_75t_SL g3764 ( 
.A(n_3521),
.Y(n_3764)
);

AOI22xp5_ASAP7_75t_L g3765 ( 
.A1(n_3457),
.A2(n_3491),
.B1(n_3456),
.B2(n_3500),
.Y(n_3765)
);

OAI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3511),
.A2(n_131),
.B(n_132),
.Y(n_3766)
);

NAND2x1_ASAP7_75t_L g3767 ( 
.A(n_3551),
.B(n_133),
.Y(n_3767)
);

HB1xp67_ASAP7_75t_L g3768 ( 
.A(n_3566),
.Y(n_3768)
);

NOR2xp33_ASAP7_75t_L g3769 ( 
.A(n_3462),
.B(n_3486),
.Y(n_3769)
);

BUFx2_ASAP7_75t_L g3770 ( 
.A(n_3431),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3465),
.Y(n_3771)
);

AOI21xp5_ASAP7_75t_L g3772 ( 
.A1(n_3577),
.A2(n_134),
.B(n_137),
.Y(n_3772)
);

NAND2xp5_ASAP7_75t_L g3773 ( 
.A(n_3415),
.B(n_134),
.Y(n_3773)
);

INVx2_ASAP7_75t_L g3774 ( 
.A(n_3538),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_3432),
.B(n_3430),
.Y(n_3775)
);

INVx1_ASAP7_75t_SL g3776 ( 
.A(n_3553),
.Y(n_3776)
);

INVxp33_ASAP7_75t_SL g3777 ( 
.A(n_3439),
.Y(n_3777)
);

O2A1O1Ixp33_ASAP7_75t_SL g3778 ( 
.A1(n_3443),
.A2(n_139),
.B(n_137),
.C(n_138),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3438),
.Y(n_3779)
);

A2O1A1Ixp33_ASAP7_75t_L g3780 ( 
.A1(n_3582),
.A2(n_140),
.B(n_138),
.C(n_139),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3522),
.Y(n_3781)
);

AOI21x1_ASAP7_75t_L g3782 ( 
.A1(n_3530),
.A2(n_3540),
.B(n_3536),
.Y(n_3782)
);

INVx3_ASAP7_75t_L g3783 ( 
.A(n_3505),
.Y(n_3783)
);

O2A1O1Ixp33_ASAP7_75t_L g3784 ( 
.A1(n_3587),
.A2(n_142),
.B(n_140),
.C(n_141),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_L g3785 ( 
.A(n_3541),
.B(n_141),
.Y(n_3785)
);

OAI22xp5_ASAP7_75t_L g3786 ( 
.A1(n_3583),
.A2(n_144),
.B1(n_142),
.B2(n_143),
.Y(n_3786)
);

O2A1O1Ixp33_ASAP7_75t_L g3787 ( 
.A1(n_3464),
.A2(n_146),
.B(n_143),
.C(n_145),
.Y(n_3787)
);

HB1xp67_ASAP7_75t_L g3788 ( 
.A(n_3559),
.Y(n_3788)
);

AOI22xp5_ASAP7_75t_L g3789 ( 
.A1(n_3456),
.A2(n_149),
.B1(n_147),
.B2(n_148),
.Y(n_3789)
);

NOR2xp33_ASAP7_75t_L g3790 ( 
.A(n_3487),
.B(n_149),
.Y(n_3790)
);

O2A1O1Ixp33_ASAP7_75t_L g3791 ( 
.A1(n_3472),
.A2(n_152),
.B(n_150),
.C(n_151),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3431),
.B(n_150),
.Y(n_3792)
);

BUFx6f_ASAP7_75t_L g3793 ( 
.A(n_3505),
.Y(n_3793)
);

OAI22xp5_ASAP7_75t_L g3794 ( 
.A1(n_3584),
.A2(n_154),
.B1(n_151),
.B2(n_153),
.Y(n_3794)
);

INVx3_ASAP7_75t_L g3795 ( 
.A(n_3513),
.Y(n_3795)
);

AOI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_3561),
.A2(n_153),
.B(n_155),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3449),
.B(n_155),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3571),
.Y(n_3798)
);

OR2x6_ASAP7_75t_SL g3799 ( 
.A(n_3452),
.B(n_157),
.Y(n_3799)
);

AND2x2_ASAP7_75t_SL g3800 ( 
.A(n_3571),
.B(n_3549),
.Y(n_3800)
);

AND2x4_ASAP7_75t_L g3801 ( 
.A(n_3549),
.B(n_157),
.Y(n_3801)
);

BUFx8_ASAP7_75t_L g3802 ( 
.A(n_3562),
.Y(n_3802)
);

AOI222xp33_ASAP7_75t_L g3803 ( 
.A1(n_3412),
.A2(n_160),
.B1(n_162),
.B2(n_158),
.C1(n_159),
.C2(n_161),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3449),
.B(n_158),
.Y(n_3804)
);

A2O1A1Ixp33_ASAP7_75t_L g3805 ( 
.A1(n_3562),
.A2(n_162),
.B(n_160),
.C(n_161),
.Y(n_3805)
);

INVx5_ASAP7_75t_L g3806 ( 
.A(n_3411),
.Y(n_3806)
);

INVx2_ASAP7_75t_SL g3807 ( 
.A(n_3475),
.Y(n_3807)
);

AOI22xp33_ASAP7_75t_L g3808 ( 
.A1(n_3560),
.A2(n_165),
.B1(n_163),
.B2(n_164),
.Y(n_3808)
);

NAND2xp5_ASAP7_75t_L g3809 ( 
.A(n_3490),
.B(n_164),
.Y(n_3809)
);

AO32x1_ASAP7_75t_L g3810 ( 
.A1(n_3552),
.A2(n_3556),
.A3(n_3513),
.B1(n_3570),
.B2(n_3574),
.Y(n_3810)
);

INVx3_ASAP7_75t_L g3811 ( 
.A(n_3552),
.Y(n_3811)
);

BUFx6f_ASAP7_75t_L g3812 ( 
.A(n_3411),
.Y(n_3812)
);

OAI22xp5_ASAP7_75t_L g3813 ( 
.A1(n_3498),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_3813)
);

BUFx3_ASAP7_75t_L g3814 ( 
.A(n_3475),
.Y(n_3814)
);

OR2x6_ASAP7_75t_SL g3815 ( 
.A(n_3499),
.B(n_3501),
.Y(n_3815)
);

A2O1A1Ixp33_ASAP7_75t_L g3816 ( 
.A1(n_3440),
.A2(n_168),
.B(n_166),
.C(n_167),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_SL g3817 ( 
.A(n_3656),
.B(n_3558),
.Y(n_3817)
);

OR2x6_ASAP7_75t_L g3818 ( 
.A(n_3635),
.B(n_3560),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3664),
.Y(n_3819)
);

AOI22xp33_ASAP7_75t_L g3820 ( 
.A1(n_3674),
.A2(n_3588),
.B1(n_3500),
.B2(n_3550),
.Y(n_3820)
);

BUFx3_ASAP7_75t_L g3821 ( 
.A(n_3600),
.Y(n_3821)
);

NOR2xp33_ASAP7_75t_L g3822 ( 
.A(n_3799),
.B(n_3558),
.Y(n_3822)
);

BUFx3_ASAP7_75t_L g3823 ( 
.A(n_3688),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3608),
.B(n_3578),
.Y(n_3824)
);

INVx1_ASAP7_75t_L g3825 ( 
.A(n_3671),
.Y(n_3825)
);

OR2x6_ASAP7_75t_L g3826 ( 
.A(n_3635),
.B(n_3558),
.Y(n_3826)
);

AOI22xp5_ASAP7_75t_L g3827 ( 
.A1(n_3674),
.A2(n_3512),
.B1(n_3477),
.B2(n_3590),
.Y(n_3827)
);

OAI22xp33_ASAP7_75t_L g3828 ( 
.A1(n_3656),
.A2(n_3504),
.B1(n_3515),
.B2(n_3475),
.Y(n_3828)
);

BUFx2_ASAP7_75t_L g3829 ( 
.A(n_3728),
.Y(n_3829)
);

INVx2_ASAP7_75t_L g3830 ( 
.A(n_3774),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_L g3831 ( 
.A(n_3597),
.B(n_3590),
.Y(n_3831)
);

OAI22xp5_ASAP7_75t_L g3832 ( 
.A1(n_3666),
.A2(n_3631),
.B1(n_3629),
.B2(n_3706),
.Y(n_3832)
);

INVx1_ASAP7_75t_L g3833 ( 
.A(n_3687),
.Y(n_3833)
);

A2O1A1Ixp33_ASAP7_75t_L g3834 ( 
.A1(n_3787),
.A2(n_3477),
.B(n_3515),
.C(n_3504),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3632),
.Y(n_3835)
);

BUFx6f_ASAP7_75t_L g3836 ( 
.A(n_3655),
.Y(n_3836)
);

A2O1A1Ixp33_ASAP7_75t_L g3837 ( 
.A1(n_3791),
.A2(n_3504),
.B(n_3515),
.C(n_3524),
.Y(n_3837)
);

BUFx6f_ASAP7_75t_L g3838 ( 
.A(n_3677),
.Y(n_3838)
);

AOI22xp33_ASAP7_75t_L g3839 ( 
.A1(n_3729),
.A2(n_3524),
.B1(n_3535),
.B2(n_3492),
.Y(n_3839)
);

BUFx6f_ASAP7_75t_L g3840 ( 
.A(n_3640),
.Y(n_3840)
);

AND2x2_ASAP7_75t_L g3841 ( 
.A(n_3651),
.B(n_3546),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3607),
.B(n_3546),
.Y(n_3842)
);

A2O1A1Ixp33_ASAP7_75t_SL g3843 ( 
.A1(n_3766),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_3843)
);

OA22x2_ASAP7_75t_L g3844 ( 
.A1(n_3611),
.A2(n_171),
.B1(n_169),
.B2(n_170),
.Y(n_3844)
);

AND2x2_ASAP7_75t_L g3845 ( 
.A(n_3591),
.B(n_172),
.Y(n_3845)
);

OAI22xp5_ASAP7_75t_SL g3846 ( 
.A1(n_3596),
.A2(n_3656),
.B1(n_3759),
.B2(n_3645),
.Y(n_3846)
);

BUFx2_ASAP7_75t_L g3847 ( 
.A(n_3723),
.Y(n_3847)
);

AND2x4_ASAP7_75t_L g3848 ( 
.A(n_3628),
.B(n_172),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_L g3849 ( 
.A(n_3647),
.B(n_3681),
.Y(n_3849)
);

INVx3_ASAP7_75t_L g3850 ( 
.A(n_3596),
.Y(n_3850)
);

BUFx3_ASAP7_75t_L g3851 ( 
.A(n_3626),
.Y(n_3851)
);

INVx1_ASAP7_75t_L g3852 ( 
.A(n_3703),
.Y(n_3852)
);

AO21x2_ASAP7_75t_L g3853 ( 
.A1(n_3782),
.A2(n_173),
.B(n_174),
.Y(n_3853)
);

NOR2xp33_ASAP7_75t_L g3854 ( 
.A(n_3657),
.B(n_173),
.Y(n_3854)
);

INVx1_ASAP7_75t_L g3855 ( 
.A(n_3716),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3672),
.B(n_174),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3722),
.Y(n_3857)
);

AND2x4_ASAP7_75t_L g3858 ( 
.A(n_3634),
.B(n_175),
.Y(n_3858)
);

AND2x4_ASAP7_75t_L g3859 ( 
.A(n_3700),
.B(n_175),
.Y(n_3859)
);

BUFx3_ASAP7_75t_L g3860 ( 
.A(n_3612),
.Y(n_3860)
);

OR2x6_ASAP7_75t_L g3861 ( 
.A(n_3609),
.B(n_176),
.Y(n_3861)
);

INVx1_ASAP7_75t_L g3862 ( 
.A(n_3736),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3602),
.Y(n_3863)
);

INVx8_ASAP7_75t_L g3864 ( 
.A(n_3653),
.Y(n_3864)
);

AND2x4_ASAP7_75t_L g3865 ( 
.A(n_3701),
.B(n_3643),
.Y(n_3865)
);

OAI22xp5_ASAP7_75t_L g3866 ( 
.A1(n_3789),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3613),
.Y(n_3867)
);

INVx6_ASAP7_75t_L g3868 ( 
.A(n_3668),
.Y(n_3868)
);

NAND2xp5_ASAP7_75t_L g3869 ( 
.A(n_3776),
.B(n_177),
.Y(n_3869)
);

OAI22xp5_ASAP7_75t_L g3870 ( 
.A1(n_3669),
.A2(n_182),
.B1(n_178),
.B2(n_179),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3614),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3620),
.Y(n_3872)
);

AO21x2_ASAP7_75t_L g3873 ( 
.A1(n_3782),
.A2(n_182),
.B(n_183),
.Y(n_3873)
);

BUFx6f_ASAP7_75t_L g3874 ( 
.A(n_3640),
.Y(n_3874)
);

BUFx6f_ASAP7_75t_L g3875 ( 
.A(n_3640),
.Y(n_3875)
);

AND2x4_ASAP7_75t_L g3876 ( 
.A(n_3678),
.B(n_183),
.Y(n_3876)
);

AOI22xp33_ASAP7_75t_L g3877 ( 
.A1(n_3662),
.A2(n_3712),
.B1(n_3779),
.B2(n_3803),
.Y(n_3877)
);

BUFx12f_ASAP7_75t_L g3878 ( 
.A(n_3594),
.Y(n_3878)
);

INVx2_ASAP7_75t_L g3879 ( 
.A(n_3633),
.Y(n_3879)
);

INVx6_ASAP7_75t_L g3880 ( 
.A(n_3668),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3775),
.B(n_185),
.Y(n_3881)
);

AND2x2_ASAP7_75t_L g3882 ( 
.A(n_3663),
.B(n_186),
.Y(n_3882)
);

BUFx12f_ASAP7_75t_L g3883 ( 
.A(n_3680),
.Y(n_3883)
);

INVx6_ASAP7_75t_L g3884 ( 
.A(n_3802),
.Y(n_3884)
);

INVx3_ASAP7_75t_L g3885 ( 
.A(n_3604),
.Y(n_3885)
);

BUFx6f_ASAP7_75t_L g3886 ( 
.A(n_3649),
.Y(n_3886)
);

BUFx2_ASAP7_75t_L g3887 ( 
.A(n_3741),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_3768),
.B(n_186),
.Y(n_3888)
);

AOI22xp5_ASAP7_75t_L g3889 ( 
.A1(n_3777),
.A2(n_190),
.B1(n_187),
.B2(n_189),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3676),
.A2(n_190),
.B1(n_187),
.B2(n_189),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3639),
.Y(n_3891)
);

BUFx12f_ASAP7_75t_L g3892 ( 
.A(n_3679),
.Y(n_3892)
);

BUFx2_ASAP7_75t_L g3893 ( 
.A(n_3770),
.Y(n_3893)
);

INVx1_ASAP7_75t_L g3894 ( 
.A(n_3622),
.Y(n_3894)
);

AND2x4_ASAP7_75t_L g3895 ( 
.A(n_3643),
.B(n_191),
.Y(n_3895)
);

INVx1_ASAP7_75t_L g3896 ( 
.A(n_3623),
.Y(n_3896)
);

CKINVDCx6p67_ASAP7_75t_R g3897 ( 
.A(n_3625),
.Y(n_3897)
);

AND2x2_ASAP7_75t_L g3898 ( 
.A(n_3599),
.B(n_191),
.Y(n_3898)
);

BUFx2_ASAP7_75t_L g3899 ( 
.A(n_3811),
.Y(n_3899)
);

BUFx3_ASAP7_75t_L g3900 ( 
.A(n_3720),
.Y(n_3900)
);

AOI21xp33_ASAP7_75t_L g3901 ( 
.A1(n_3715),
.A2(n_192),
.B(n_193),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3636),
.Y(n_3902)
);

BUFx2_ASAP7_75t_L g3903 ( 
.A(n_3814),
.Y(n_3903)
);

INVx1_ASAP7_75t_SL g3904 ( 
.A(n_3732),
.Y(n_3904)
);

INVx1_ASAP7_75t_SL g3905 ( 
.A(n_3650),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3769),
.B(n_192),
.Y(n_3906)
);

NAND2x1p5_ASAP7_75t_L g3907 ( 
.A(n_3679),
.B(n_194),
.Y(n_3907)
);

INVx2_ASAP7_75t_SL g3908 ( 
.A(n_3598),
.Y(n_3908)
);

AOI21xp5_ASAP7_75t_L g3909 ( 
.A1(n_3621),
.A2(n_194),
.B(n_195),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3638),
.Y(n_3910)
);

BUFx2_ASAP7_75t_L g3911 ( 
.A(n_3750),
.Y(n_3911)
);

INVx1_ASAP7_75t_L g3912 ( 
.A(n_3753),
.Y(n_3912)
);

OR2x6_ASAP7_75t_L g3913 ( 
.A(n_3609),
.B(n_3615),
.Y(n_3913)
);

INVx2_ASAP7_75t_SL g3914 ( 
.A(n_3709),
.Y(n_3914)
);

NOR2xp33_ASAP7_75t_SL g3915 ( 
.A(n_3691),
.B(n_195),
.Y(n_3915)
);

AOI22xp33_ASAP7_75t_L g3916 ( 
.A1(n_3637),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3644),
.Y(n_3917)
);

INVx1_ASAP7_75t_L g3918 ( 
.A(n_3660),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3605),
.Y(n_3919)
);

INVx1_ASAP7_75t_L g3920 ( 
.A(n_3738),
.Y(n_3920)
);

INVx2_ASAP7_75t_SL g3921 ( 
.A(n_3802),
.Y(n_3921)
);

NOR2xp67_ASAP7_75t_L g3922 ( 
.A(n_3806),
.B(n_196),
.Y(n_3922)
);

OAI22xp5_ASAP7_75t_L g3923 ( 
.A1(n_3765),
.A2(n_3595),
.B1(n_3805),
.B2(n_3670),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_L g3924 ( 
.A(n_3751),
.B(n_197),
.Y(n_3924)
);

INVxp67_ASAP7_75t_L g3925 ( 
.A(n_3815),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_L g3926 ( 
.A(n_3788),
.B(n_3724),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3733),
.B(n_198),
.Y(n_3927)
);

AOI22xp5_ASAP7_75t_L g3928 ( 
.A1(n_3794),
.A2(n_201),
.B1(n_199),
.B2(n_200),
.Y(n_3928)
);

INVx2_ASAP7_75t_SL g3929 ( 
.A(n_3702),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3735),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3593),
.B(n_202),
.Y(n_3931)
);

O2A1O1Ixp33_ASAP7_75t_L g3932 ( 
.A1(n_3816),
.A2(n_206),
.B(n_203),
.C(n_205),
.Y(n_3932)
);

INVx2_ASAP7_75t_SL g3933 ( 
.A(n_3714),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3785),
.B(n_203),
.Y(n_3934)
);

INVx3_ASAP7_75t_L g3935 ( 
.A(n_3704),
.Y(n_3935)
);

INVx2_ASAP7_75t_L g3936 ( 
.A(n_3606),
.Y(n_3936)
);

BUFx2_ASAP7_75t_L g3937 ( 
.A(n_3807),
.Y(n_3937)
);

INVx1_ASAP7_75t_L g3938 ( 
.A(n_3627),
.Y(n_3938)
);

BUFx6f_ASAP7_75t_L g3939 ( 
.A(n_3649),
.Y(n_3939)
);

BUFx2_ASAP7_75t_L g3940 ( 
.A(n_3610),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_3686),
.B(n_206),
.Y(n_3941)
);

OAI22xp5_ASAP7_75t_L g3942 ( 
.A1(n_3699),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_3942)
);

A2O1A1Ixp33_ASAP7_75t_L g3943 ( 
.A1(n_3654),
.A2(n_212),
.B(n_210),
.C(n_211),
.Y(n_3943)
);

AOI22xp5_ASAP7_75t_L g3944 ( 
.A1(n_3694),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3641),
.Y(n_3945)
);

INVxp67_ASAP7_75t_L g3946 ( 
.A(n_3646),
.Y(n_3946)
);

BUFx3_ASAP7_75t_L g3947 ( 
.A(n_3801),
.Y(n_3947)
);

BUFx6f_ASAP7_75t_L g3948 ( 
.A(n_3649),
.Y(n_3948)
);

NOR3xp33_ASAP7_75t_L g3949 ( 
.A(n_3758),
.B(n_213),
.C(n_214),
.Y(n_3949)
);

AND2x4_ASAP7_75t_L g3950 ( 
.A(n_3609),
.B(n_213),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3737),
.Y(n_3951)
);

BUFx6f_ASAP7_75t_L g3952 ( 
.A(n_3659),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3692),
.B(n_214),
.Y(n_3953)
);

AOI221xp5_ASAP7_75t_L g3954 ( 
.A1(n_3784),
.A2(n_217),
.B1(n_215),
.B2(n_216),
.C(n_219),
.Y(n_3954)
);

OR2x6_ASAP7_75t_L g3955 ( 
.A(n_3615),
.B(n_216),
.Y(n_3955)
);

INVx3_ASAP7_75t_L g3956 ( 
.A(n_3704),
.Y(n_3956)
);

OAI22xp5_ASAP7_75t_L g3957 ( 
.A1(n_3747),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3652),
.Y(n_3958)
);

OAI22xp33_ASAP7_75t_L g3959 ( 
.A1(n_3684),
.A2(n_223),
.B1(n_221),
.B2(n_222),
.Y(n_3959)
);

INVx1_ASAP7_75t_SL g3960 ( 
.A(n_3752),
.Y(n_3960)
);

CKINVDCx5p33_ASAP7_75t_R g3961 ( 
.A(n_3659),
.Y(n_3961)
);

INVx1_ASAP7_75t_SL g3962 ( 
.A(n_3801),
.Y(n_3962)
);

NAND2xp5_ASAP7_75t_SL g3963 ( 
.A(n_3615),
.B(n_3806),
.Y(n_3963)
);

NAND3xp33_ASAP7_75t_L g3964 ( 
.A(n_3690),
.B(n_222),
.C(n_223),
.Y(n_3964)
);

INVx2_ASAP7_75t_L g3965 ( 
.A(n_3658),
.Y(n_3965)
);

AOI22xp5_ASAP7_75t_L g3966 ( 
.A1(n_3694),
.A2(n_3763),
.B1(n_3760),
.B2(n_3721),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3689),
.Y(n_3967)
);

AND2x4_ASAP7_75t_L g3968 ( 
.A(n_3806),
.B(n_224),
.Y(n_3968)
);

INVx2_ASAP7_75t_L g3969 ( 
.A(n_3696),
.Y(n_3969)
);

AOI21xp5_ASAP7_75t_L g3970 ( 
.A1(n_3624),
.A2(n_226),
.B(n_227),
.Y(n_3970)
);

INVx2_ASAP7_75t_L g3971 ( 
.A(n_3698),
.Y(n_3971)
);

BUFx4f_ASAP7_75t_SL g3972 ( 
.A(n_3710),
.Y(n_3972)
);

AOI22xp5_ASAP7_75t_L g3973 ( 
.A1(n_3757),
.A2(n_229),
.B1(n_226),
.B2(n_228),
.Y(n_3973)
);

INVx1_ASAP7_75t_L g3974 ( 
.A(n_3755),
.Y(n_3974)
);

INVx1_ASAP7_75t_L g3975 ( 
.A(n_3771),
.Y(n_3975)
);

AOI21xp5_ASAP7_75t_L g3976 ( 
.A1(n_3601),
.A2(n_230),
.B(n_231),
.Y(n_3976)
);

INVx3_ASAP7_75t_L g3977 ( 
.A(n_3704),
.Y(n_3977)
);

AOI222xp33_ASAP7_75t_L g3978 ( 
.A1(n_3762),
.A2(n_233),
.B1(n_235),
.B2(n_230),
.C1(n_232),
.C2(n_234),
.Y(n_3978)
);

CKINVDCx20_ASAP7_75t_R g3979 ( 
.A(n_3592),
.Y(n_3979)
);

INVx1_ASAP7_75t_L g3980 ( 
.A(n_3717),
.Y(n_3980)
);

BUFx8_ASAP7_75t_L g3981 ( 
.A(n_3707),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3718),
.Y(n_3982)
);

NOR2xp33_ASAP7_75t_L g3983 ( 
.A(n_3648),
.B(n_233),
.Y(n_3983)
);

HB1xp67_ASAP7_75t_L g3984 ( 
.A(n_3748),
.Y(n_3984)
);

AND2x4_ASAP7_75t_L g3985 ( 
.A(n_3798),
.B(n_234),
.Y(n_3985)
);

INVx2_ASAP7_75t_SL g3986 ( 
.A(n_3659),
.Y(n_3986)
);

BUFx12f_ASAP7_75t_L g3987 ( 
.A(n_3653),
.Y(n_3987)
);

INVx4_ASAP7_75t_L g3988 ( 
.A(n_3661),
.Y(n_3988)
);

BUFx12f_ASAP7_75t_L g3989 ( 
.A(n_3667),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3719),
.Y(n_3990)
);

CKINVDCx20_ASAP7_75t_R g3991 ( 
.A(n_3713),
.Y(n_3991)
);

NOR2xp33_ASAP7_75t_L g3992 ( 
.A(n_3630),
.B(n_236),
.Y(n_3992)
);

BUFx4f_ASAP7_75t_SL g3993 ( 
.A(n_3710),
.Y(n_3993)
);

BUFx2_ASAP7_75t_L g3994 ( 
.A(n_3764),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3773),
.B(n_237),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3790),
.B(n_238),
.Y(n_3996)
);

AOI21xp5_ASAP7_75t_L g3997 ( 
.A1(n_3618),
.A2(n_239),
.B(n_240),
.Y(n_3997)
);

INVx3_ASAP7_75t_SL g3998 ( 
.A(n_3884),
.Y(n_3998)
);

OAI21x1_ASAP7_75t_SL g3999 ( 
.A1(n_3921),
.A2(n_3797),
.B(n_3792),
.Y(n_3999)
);

AOI21x1_ASAP7_75t_L g4000 ( 
.A1(n_3888),
.A2(n_3767),
.B(n_3804),
.Y(n_4000)
);

INVx2_ASAP7_75t_SL g4001 ( 
.A(n_3884),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3830),
.Y(n_4002)
);

AND2x2_ASAP7_75t_L g4003 ( 
.A(n_3865),
.B(n_3749),
.Y(n_4003)
);

AO31x2_ASAP7_75t_L g4004 ( 
.A1(n_3837),
.A2(n_3923),
.A3(n_3832),
.B(n_3909),
.Y(n_4004)
);

INVx2_ASAP7_75t_L g4005 ( 
.A(n_3835),
.Y(n_4005)
);

OAI21x1_ASAP7_75t_L g4006 ( 
.A1(n_3963),
.A2(n_3616),
.B(n_3767),
.Y(n_4006)
);

INVx2_ASAP7_75t_SL g4007 ( 
.A(n_3868),
.Y(n_4007)
);

OA21x2_ASAP7_75t_L g4008 ( 
.A1(n_3842),
.A2(n_3781),
.B(n_3617),
.Y(n_4008)
);

INVx2_ASAP7_75t_L g4009 ( 
.A(n_3879),
.Y(n_4009)
);

OAI21x1_ASAP7_75t_L g4010 ( 
.A1(n_3831),
.A2(n_3603),
.B(n_3783),
.Y(n_4010)
);

OAI21x1_ASAP7_75t_L g4011 ( 
.A1(n_3817),
.A2(n_3795),
.B(n_3697),
.Y(n_4011)
);

BUFx3_ASAP7_75t_L g4012 ( 
.A(n_3821),
.Y(n_4012)
);

INVx2_ASAP7_75t_L g4013 ( 
.A(n_3891),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_3829),
.Y(n_4014)
);

AO21x2_ASAP7_75t_L g4015 ( 
.A1(n_3970),
.A2(n_3809),
.B(n_3730),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3940),
.B(n_3711),
.Y(n_4016)
);

AO21x1_ASAP7_75t_L g4017 ( 
.A1(n_3822),
.A2(n_3745),
.B(n_3711),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3863),
.Y(n_4018)
);

AND2x2_ASAP7_75t_L g4019 ( 
.A(n_3940),
.B(n_3695),
.Y(n_4019)
);

AOI22xp5_ASAP7_75t_L g4020 ( 
.A1(n_3844),
.A2(n_3754),
.B1(n_3745),
.B2(n_3667),
.Y(n_4020)
);

CKINVDCx20_ASAP7_75t_R g4021 ( 
.A(n_3823),
.Y(n_4021)
);

OAI21xp5_ASAP7_75t_L g4022 ( 
.A1(n_3906),
.A2(n_3780),
.B(n_3746),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3867),
.Y(n_4023)
);

OA21x2_ASAP7_75t_L g4024 ( 
.A1(n_3925),
.A2(n_3761),
.B(n_3725),
.Y(n_4024)
);

AO31x2_ASAP7_75t_L g4025 ( 
.A1(n_3834),
.A2(n_3813),
.A3(n_3786),
.B(n_3756),
.Y(n_4025)
);

AOI22xp33_ASAP7_75t_L g4026 ( 
.A1(n_3976),
.A2(n_3796),
.B1(n_3812),
.B2(n_3705),
.Y(n_4026)
);

OAI21x1_ASAP7_75t_L g4027 ( 
.A1(n_3935),
.A2(n_3619),
.B(n_3772),
.Y(n_4027)
);

OAI21x1_ASAP7_75t_L g4028 ( 
.A1(n_3956),
.A2(n_3708),
.B(n_3740),
.Y(n_4028)
);

INVx3_ASAP7_75t_L g4029 ( 
.A(n_3829),
.Y(n_4029)
);

OAI22xp5_ASAP7_75t_L g4030 ( 
.A1(n_3820),
.A2(n_3808),
.B1(n_3744),
.B2(n_3743),
.Y(n_4030)
);

AND2x2_ASAP7_75t_L g4031 ( 
.A(n_3847),
.B(n_3682),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3984),
.B(n_3661),
.Y(n_4032)
);

OAI21x1_ASAP7_75t_L g4033 ( 
.A1(n_3977),
.A2(n_3739),
.B(n_3734),
.Y(n_4033)
);

BUFx12f_ASAP7_75t_L g4034 ( 
.A(n_3878),
.Y(n_4034)
);

BUFx2_ASAP7_75t_L g4035 ( 
.A(n_3903),
.Y(n_4035)
);

INVx2_ASAP7_75t_SL g4036 ( 
.A(n_3868),
.Y(n_4036)
);

CKINVDCx6p67_ASAP7_75t_R g4037 ( 
.A(n_3851),
.Y(n_4037)
);

AND2x2_ASAP7_75t_L g4038 ( 
.A(n_3847),
.B(n_3685),
.Y(n_4038)
);

AOI221xp5_ASAP7_75t_L g4039 ( 
.A1(n_3901),
.A2(n_3683),
.B1(n_3726),
.B2(n_3742),
.C(n_3778),
.Y(n_4039)
);

OAI21x1_ASAP7_75t_L g4040 ( 
.A1(n_3824),
.A2(n_3693),
.B(n_3810),
.Y(n_4040)
);

INVx4_ASAP7_75t_L g4041 ( 
.A(n_3880),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3871),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3929),
.B(n_3661),
.Y(n_4043)
);

INVx1_ASAP7_75t_L g4044 ( 
.A(n_3872),
.Y(n_4044)
);

BUFx8_ASAP7_75t_SL g4045 ( 
.A(n_3883),
.Y(n_4045)
);

OAI221xp5_ASAP7_75t_L g4046 ( 
.A1(n_3877),
.A2(n_3812),
.B1(n_3793),
.B2(n_3675),
.C(n_3665),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_L g4047 ( 
.A(n_3887),
.B(n_3673),
.Y(n_4047)
);

AOI21xp5_ASAP7_75t_L g4048 ( 
.A1(n_3828),
.A2(n_3810),
.B(n_3800),
.Y(n_4048)
);

AND2x2_ASAP7_75t_L g4049 ( 
.A(n_3887),
.B(n_3642),
.Y(n_4049)
);

INVx1_ASAP7_75t_SL g4050 ( 
.A(n_3897),
.Y(n_4050)
);

OAI21x1_ASAP7_75t_L g4051 ( 
.A1(n_3827),
.A2(n_3812),
.B(n_3793),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3894),
.Y(n_4052)
);

BUFx6f_ASAP7_75t_L g4053 ( 
.A(n_3836),
.Y(n_4053)
);

INVx1_ASAP7_75t_L g4054 ( 
.A(n_3896),
.Y(n_4054)
);

OA21x2_ASAP7_75t_L g4055 ( 
.A1(n_3937),
.A2(n_3754),
.B(n_3793),
.Y(n_4055)
);

BUFx3_ASAP7_75t_L g4056 ( 
.A(n_3900),
.Y(n_4056)
);

OAI21x1_ASAP7_75t_L g4057 ( 
.A1(n_3839),
.A2(n_3731),
.B(n_3727),
.Y(n_4057)
);

OAI222xp33_ASAP7_75t_L g4058 ( 
.A1(n_3966),
.A2(n_3673),
.B1(n_3731),
.B2(n_3727),
.C1(n_241),
.C2(n_243),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_L g4059 ( 
.A(n_3893),
.B(n_3673),
.Y(n_4059)
);

NOR2x1_ASAP7_75t_SL g4060 ( 
.A(n_3818),
.B(n_3727),
.Y(n_4060)
);

OAI21x1_ASAP7_75t_L g4061 ( 
.A1(n_3849),
.A2(n_3731),
.B(n_239),
.Y(n_4061)
);

INVx1_ASAP7_75t_L g4062 ( 
.A(n_3902),
.Y(n_4062)
);

AOI21xp5_ASAP7_75t_L g4063 ( 
.A1(n_3932),
.A2(n_240),
.B(n_241),
.Y(n_4063)
);

AOI221xp5_ASAP7_75t_L g4064 ( 
.A1(n_3954),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.C(n_245),
.Y(n_4064)
);

INVx1_ASAP7_75t_L g4065 ( 
.A(n_3910),
.Y(n_4065)
);

OAI21x1_ASAP7_75t_L g4066 ( 
.A1(n_3885),
.A2(n_244),
.B(n_245),
.Y(n_4066)
);

OA21x2_ASAP7_75t_L g4067 ( 
.A1(n_3937),
.A2(n_246),
.B(n_247),
.Y(n_4067)
);

CKINVDCx6p67_ASAP7_75t_R g4068 ( 
.A(n_3836),
.Y(n_4068)
);

NAND3xp33_ASAP7_75t_L g4069 ( 
.A(n_3949),
.B(n_247),
.C(n_248),
.Y(n_4069)
);

AO22x2_ASAP7_75t_L g4070 ( 
.A1(n_3951),
.A2(n_251),
.B1(n_248),
.B2(n_249),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_L g4071 ( 
.A(n_3893),
.B(n_249),
.Y(n_4071)
);

INVx1_ASAP7_75t_L g4072 ( 
.A(n_3920),
.Y(n_4072)
);

OR2x6_ASAP7_75t_L g4073 ( 
.A(n_3864),
.B(n_3846),
.Y(n_4073)
);

OAI21x1_ASAP7_75t_L g4074 ( 
.A1(n_3926),
.A2(n_252),
.B(n_253),
.Y(n_4074)
);

O2A1O1Ixp33_ASAP7_75t_L g4075 ( 
.A1(n_3943),
.A2(n_255),
.B(n_252),
.C(n_254),
.Y(n_4075)
);

OAI21x1_ASAP7_75t_L g4076 ( 
.A1(n_3881),
.A2(n_255),
.B(n_256),
.Y(n_4076)
);

INVx3_ASAP7_75t_L g4077 ( 
.A(n_3860),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3819),
.Y(n_4078)
);

CKINVDCx5p33_ASAP7_75t_R g4079 ( 
.A(n_3914),
.Y(n_4079)
);

AOI21xp5_ASAP7_75t_L g4080 ( 
.A1(n_3843),
.A2(n_3964),
.B(n_3997),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3919),
.Y(n_4081)
);

INVx1_ASAP7_75t_L g4082 ( 
.A(n_3825),
.Y(n_4082)
);

BUFx2_ASAP7_75t_L g4083 ( 
.A(n_3903),
.Y(n_4083)
);

INVx1_ASAP7_75t_L g4084 ( 
.A(n_3833),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3852),
.B(n_259),
.Y(n_4085)
);

AOI22xp33_ASAP7_75t_L g4086 ( 
.A1(n_3853),
.A2(n_261),
.B1(n_259),
.B2(n_260),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3855),
.Y(n_4087)
);

OAI21x1_ASAP7_75t_L g4088 ( 
.A1(n_3841),
.A2(n_260),
.B(n_262),
.Y(n_4088)
);

BUFx6f_ASAP7_75t_L g4089 ( 
.A(n_3838),
.Y(n_4089)
);

OAI21x1_ASAP7_75t_L g4090 ( 
.A1(n_3850),
.A2(n_262),
.B(n_263),
.Y(n_4090)
);

OAI21x1_ASAP7_75t_L g4091 ( 
.A1(n_3974),
.A2(n_263),
.B(n_264),
.Y(n_4091)
);

INVx2_ASAP7_75t_L g4092 ( 
.A(n_3936),
.Y(n_4092)
);

A2O1A1Ixp33_ASAP7_75t_L g4093 ( 
.A1(n_3983),
.A2(n_266),
.B(n_264),
.C(n_265),
.Y(n_4093)
);

OR2x2_ASAP7_75t_L g4094 ( 
.A(n_3905),
.B(n_265),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_3857),
.Y(n_4095)
);

AOI22xp33_ASAP7_75t_L g4096 ( 
.A1(n_3873),
.A2(n_270),
.B1(n_266),
.B2(n_269),
.Y(n_4096)
);

NAND2xp5_ASAP7_75t_L g4097 ( 
.A(n_3862),
.B(n_270),
.Y(n_4097)
);

OAI21x1_ASAP7_75t_L g4098 ( 
.A1(n_3975),
.A2(n_271),
.B(n_272),
.Y(n_4098)
);

O2A1O1Ixp33_ASAP7_75t_SL g4099 ( 
.A1(n_3996),
.A2(n_273),
.B(n_271),
.C(n_272),
.Y(n_4099)
);

AO21x2_ASAP7_75t_L g4100 ( 
.A1(n_3922),
.A2(n_273),
.B(n_274),
.Y(n_4100)
);

OAI21x1_ASAP7_75t_L g4101 ( 
.A1(n_3912),
.A2(n_274),
.B(n_275),
.Y(n_4101)
);

CKINVDCx20_ASAP7_75t_R g4102 ( 
.A(n_3979),
.Y(n_4102)
);

OAI21x1_ASAP7_75t_L g4103 ( 
.A1(n_3917),
.A2(n_275),
.B(n_276),
.Y(n_4103)
);

NOR2x1_ASAP7_75t_R g4104 ( 
.A(n_3880),
.B(n_276),
.Y(n_4104)
);

INVx3_ASAP7_75t_L g4105 ( 
.A(n_3947),
.Y(n_4105)
);

HB1xp67_ASAP7_75t_L g4106 ( 
.A(n_3918),
.Y(n_4106)
);

OR2x2_ASAP7_75t_L g4107 ( 
.A(n_3899),
.B(n_277),
.Y(n_4107)
);

OAI21xp5_ASAP7_75t_L g4108 ( 
.A1(n_3992),
.A2(n_278),
.B(n_279),
.Y(n_4108)
);

AOI22x1_ASAP7_75t_L g4109 ( 
.A1(n_3978),
.A2(n_280),
.B1(n_278),
.B2(n_279),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_3938),
.Y(n_4110)
);

INVx2_ASAP7_75t_SL g4111 ( 
.A(n_3864),
.Y(n_4111)
);

INVx1_ASAP7_75t_L g4112 ( 
.A(n_3980),
.Y(n_4112)
);

INVx2_ASAP7_75t_L g4113 ( 
.A(n_3945),
.Y(n_4113)
);

AOI221xp5_ASAP7_75t_L g4114 ( 
.A1(n_3959),
.A2(n_283),
.B1(n_280),
.B2(n_281),
.C(n_284),
.Y(n_4114)
);

NAND2x1p5_ASAP7_75t_L g4115 ( 
.A(n_3968),
.B(n_3848),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_3982),
.Y(n_4116)
);

OAI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_3972),
.A2(n_284),
.B1(n_281),
.B2(n_283),
.Y(n_4117)
);

INVx1_ASAP7_75t_L g4118 ( 
.A(n_3990),
.Y(n_4118)
);

OAI21xp5_ASAP7_75t_L g4119 ( 
.A1(n_3889),
.A2(n_285),
.B(n_286),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3899),
.B(n_286),
.Y(n_4120)
);

HB1xp67_ASAP7_75t_L g4121 ( 
.A(n_3994),
.Y(n_4121)
);

OAI21xp5_ASAP7_75t_L g4122 ( 
.A1(n_3934),
.A2(n_287),
.B(n_288),
.Y(n_4122)
);

AOI31xp67_ASAP7_75t_L g4123 ( 
.A1(n_3876),
.A2(n_289),
.A3(n_287),
.B(n_288),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_3911),
.B(n_290),
.Y(n_4124)
);

AND2x2_ASAP7_75t_L g4125 ( 
.A(n_3911),
.B(n_3994),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_3958),
.Y(n_4126)
);

AOI22xp33_ASAP7_75t_L g4127 ( 
.A1(n_3866),
.A2(n_292),
.B1(n_290),
.B2(n_291),
.Y(n_4127)
);

OAI21x1_ASAP7_75t_L g4128 ( 
.A1(n_3931),
.A2(n_291),
.B(n_293),
.Y(n_4128)
);

OAI21x1_ASAP7_75t_L g4129 ( 
.A1(n_3907),
.A2(n_3924),
.B(n_3869),
.Y(n_4129)
);

OAI21x1_ASAP7_75t_SL g4130 ( 
.A1(n_3908),
.A2(n_294),
.B(n_295),
.Y(n_4130)
);

AOI31xp33_ASAP7_75t_L g4131 ( 
.A1(n_3848),
.A2(n_297),
.A3(n_294),
.B(n_296),
.Y(n_4131)
);

INVx2_ASAP7_75t_SL g4132 ( 
.A(n_3892),
.Y(n_4132)
);

BUFx10_ASAP7_75t_L g4133 ( 
.A(n_3968),
.Y(n_4133)
);

NOR2xp33_ASAP7_75t_L g4134 ( 
.A(n_3946),
.B(n_296),
.Y(n_4134)
);

OAI21x1_ASAP7_75t_L g4135 ( 
.A1(n_3856),
.A2(n_297),
.B(n_298),
.Y(n_4135)
);

OAI21x1_ASAP7_75t_L g4136 ( 
.A1(n_3941),
.A2(n_299),
.B(n_300),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3965),
.Y(n_4137)
);

OAI21x1_ASAP7_75t_L g4138 ( 
.A1(n_3845),
.A2(n_300),
.B(n_301),
.Y(n_4138)
);

O2A1O1Ixp33_ASAP7_75t_SL g4139 ( 
.A1(n_3854),
.A2(n_304),
.B(n_302),
.C(n_303),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3962),
.B(n_303),
.Y(n_4140)
);

HB1xp67_ASAP7_75t_L g4141 ( 
.A(n_3933),
.Y(n_4141)
);

OAI22xp5_ASAP7_75t_SL g4142 ( 
.A1(n_3991),
.A2(n_3993),
.B1(n_3989),
.B2(n_3987),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_3967),
.Y(n_4143)
);

AO21x2_ASAP7_75t_L g4144 ( 
.A1(n_3953),
.A2(n_305),
.B(n_306),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3969),
.Y(n_4145)
);

AOI22xp33_ASAP7_75t_SL g4146 ( 
.A1(n_3915),
.A2(n_309),
.B1(n_307),
.B2(n_308),
.Y(n_4146)
);

INVx1_ASAP7_75t_L g4147 ( 
.A(n_3971),
.Y(n_4147)
);

BUFx3_ASAP7_75t_L g4148 ( 
.A(n_3981),
.Y(n_4148)
);

OR2x2_ASAP7_75t_L g4149 ( 
.A(n_3960),
.B(n_308),
.Y(n_4149)
);

HB1xp67_ASAP7_75t_L g4150 ( 
.A(n_4014),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4106),
.Y(n_4151)
);

INVx2_ASAP7_75t_L g4152 ( 
.A(n_4024),
.Y(n_4152)
);

CKINVDCx5p33_ASAP7_75t_R g4153 ( 
.A(n_4045),
.Y(n_4153)
);

INVx3_ASAP7_75t_L g4154 ( 
.A(n_4073),
.Y(n_4154)
);

AOI22xp33_ASAP7_75t_L g4155 ( 
.A1(n_4015),
.A2(n_3957),
.B1(n_3870),
.B2(n_3890),
.Y(n_4155)
);

BUFx8_ASAP7_75t_L g4156 ( 
.A(n_4034),
.Y(n_4156)
);

INVx1_ASAP7_75t_L g4157 ( 
.A(n_4042),
.Y(n_4157)
);

BUFx6f_ASAP7_75t_L g4158 ( 
.A(n_3998),
.Y(n_4158)
);

INVx4_ASAP7_75t_L g4159 ( 
.A(n_4041),
.Y(n_4159)
);

AOI21x1_ASAP7_75t_L g4160 ( 
.A1(n_4073),
.A2(n_3876),
.B(n_3858),
.Y(n_4160)
);

OAI21x1_ASAP7_75t_L g4161 ( 
.A1(n_4051),
.A2(n_3927),
.B(n_3995),
.Y(n_4161)
);

INVx2_ASAP7_75t_SL g4162 ( 
.A(n_4133),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_4024),
.Y(n_4163)
);

OAI21x1_ASAP7_75t_L g4164 ( 
.A1(n_4010),
.A2(n_3882),
.B(n_3898),
.Y(n_4164)
);

OAI21x1_ASAP7_75t_L g4165 ( 
.A1(n_4011),
.A2(n_3944),
.B(n_3930),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_4055),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_4055),
.Y(n_4167)
);

AND2x4_ASAP7_75t_L g4168 ( 
.A(n_4035),
.B(n_3858),
.Y(n_4168)
);

OAI21x1_ASAP7_75t_L g4169 ( 
.A1(n_4057),
.A2(n_3916),
.B(n_3928),
.Y(n_4169)
);

OA21x2_ASAP7_75t_L g4170 ( 
.A1(n_4040),
.A2(n_3904),
.B(n_3961),
.Y(n_4170)
);

AOI22xp33_ASAP7_75t_SL g4171 ( 
.A1(n_4022),
.A2(n_3859),
.B1(n_3955),
.B2(n_3861),
.Y(n_4171)
);

INVx1_ASAP7_75t_SL g4172 ( 
.A(n_4102),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4042),
.Y(n_4173)
);

HB1xp67_ASAP7_75t_L g4174 ( 
.A(n_4014),
.Y(n_4174)
);

INVx2_ASAP7_75t_SL g4175 ( 
.A(n_4133),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4044),
.Y(n_4176)
);

INVx2_ASAP7_75t_L g4177 ( 
.A(n_4044),
.Y(n_4177)
);

BUFx12f_ASAP7_75t_L g4178 ( 
.A(n_4053),
.Y(n_4178)
);

BUFx2_ASAP7_75t_L g4179 ( 
.A(n_4083),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_4054),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4054),
.Y(n_4181)
);

BUFx6f_ASAP7_75t_L g4182 ( 
.A(n_4053),
.Y(n_4182)
);

INVx3_ASAP7_75t_L g4183 ( 
.A(n_4041),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4125),
.B(n_3986),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_L g4185 ( 
.A(n_4062),
.B(n_4065),
.Y(n_4185)
);

AOI22xp33_ASAP7_75t_L g4186 ( 
.A1(n_4015),
.A2(n_3942),
.B1(n_3955),
.B2(n_3861),
.Y(n_4186)
);

INVx1_ASAP7_75t_L g4187 ( 
.A(n_4062),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_4065),
.Y(n_4188)
);

OR2x2_ASAP7_75t_L g4189 ( 
.A(n_4016),
.B(n_3988),
.Y(n_4189)
);

AND2x2_ASAP7_75t_L g4190 ( 
.A(n_4019),
.B(n_3838),
.Y(n_4190)
);

BUFx10_ASAP7_75t_L g4191 ( 
.A(n_4053),
.Y(n_4191)
);

HB1xp67_ASAP7_75t_L g4192 ( 
.A(n_4121),
.Y(n_4192)
);

AOI22xp33_ASAP7_75t_SL g4193 ( 
.A1(n_4108),
.A2(n_3950),
.B1(n_3985),
.B2(n_3895),
.Y(n_4193)
);

AO21x1_ASAP7_75t_L g4194 ( 
.A1(n_4131),
.A2(n_3950),
.B(n_3985),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4072),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4072),
.Y(n_4196)
);

AOI22xp33_ASAP7_75t_L g4197 ( 
.A1(n_4109),
.A2(n_3973),
.B1(n_3818),
.B2(n_3826),
.Y(n_4197)
);

AOI21x1_ASAP7_75t_L g4198 ( 
.A1(n_4000),
.A2(n_3913),
.B(n_3826),
.Y(n_4198)
);

AOI21x1_ASAP7_75t_L g4199 ( 
.A1(n_4017),
.A2(n_3913),
.B(n_3874),
.Y(n_4199)
);

INVx3_ASAP7_75t_L g4200 ( 
.A(n_4029),
.Y(n_4200)
);

INVx2_ASAP7_75t_L g4201 ( 
.A(n_4078),
.Y(n_4201)
);

OAI21x1_ASAP7_75t_L g4202 ( 
.A1(n_4029),
.A2(n_4048),
.B(n_4006),
.Y(n_4202)
);

OAI22xp5_ASAP7_75t_L g4203 ( 
.A1(n_4069),
.A2(n_3874),
.B1(n_3875),
.B2(n_3840),
.Y(n_4203)
);

NAND2x1p5_ASAP7_75t_L g4204 ( 
.A(n_4077),
.B(n_3840),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4078),
.Y(n_4205)
);

INVx1_ASAP7_75t_SL g4206 ( 
.A(n_4021),
.Y(n_4206)
);

BUFx2_ASAP7_75t_L g4207 ( 
.A(n_4077),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4082),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4082),
.Y(n_4209)
);

INVx4_ASAP7_75t_L g4210 ( 
.A(n_4068),
.Y(n_4210)
);

OAI21x1_ASAP7_75t_SL g4211 ( 
.A1(n_4060),
.A2(n_3886),
.B(n_3875),
.Y(n_4211)
);

AO21x2_ASAP7_75t_L g4212 ( 
.A1(n_4085),
.A2(n_3939),
.B(n_3886),
.Y(n_4212)
);

BUFx6f_ASAP7_75t_L g4213 ( 
.A(n_4089),
.Y(n_4213)
);

INVx3_ASAP7_75t_SL g4214 ( 
.A(n_4037),
.Y(n_4214)
);

INVx1_ASAP7_75t_L g4215 ( 
.A(n_4084),
.Y(n_4215)
);

INVx2_ASAP7_75t_SL g4216 ( 
.A(n_4148),
.Y(n_4216)
);

INVx4_ASAP7_75t_L g4217 ( 
.A(n_4089),
.Y(n_4217)
);

AOI21x1_ASAP7_75t_L g4218 ( 
.A1(n_4071),
.A2(n_4120),
.B(n_3999),
.Y(n_4218)
);

AOI22xp33_ASAP7_75t_SL g4219 ( 
.A1(n_4067),
.A2(n_3948),
.B1(n_3952),
.B2(n_3939),
.Y(n_4219)
);

INVx2_ASAP7_75t_SL g4220 ( 
.A(n_4089),
.Y(n_4220)
);

OAI21x1_ASAP7_75t_L g4221 ( 
.A1(n_4047),
.A2(n_3952),
.B(n_3948),
.Y(n_4221)
);

BUFx8_ASAP7_75t_SL g4222 ( 
.A(n_4012),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_4084),
.Y(n_4223)
);

INVx2_ASAP7_75t_L g4224 ( 
.A(n_4087),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_L g4225 ( 
.A(n_4087),
.B(n_309),
.Y(n_4225)
);

AOI22xp33_ASAP7_75t_L g4226 ( 
.A1(n_4030),
.A2(n_312),
.B1(n_310),
.B2(n_311),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_4095),
.Y(n_4227)
);

INVx2_ASAP7_75t_L g4228 ( 
.A(n_4095),
.Y(n_4228)
);

AO21x1_ASAP7_75t_L g4229 ( 
.A1(n_4094),
.A2(n_4149),
.B(n_4134),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_4112),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_4112),
.Y(n_4231)
);

INVx3_ASAP7_75t_L g4232 ( 
.A(n_4067),
.Y(n_4232)
);

AO21x2_ASAP7_75t_L g4233 ( 
.A1(n_4097),
.A2(n_310),
.B(n_311),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4116),
.Y(n_4234)
);

AOI22xp33_ASAP7_75t_SL g4235 ( 
.A1(n_4119),
.A2(n_316),
.B1(n_313),
.B2(n_315),
.Y(n_4235)
);

AO21x1_ASAP7_75t_SL g4236 ( 
.A1(n_4107),
.A2(n_313),
.B(n_315),
.Y(n_4236)
);

INVx1_ASAP7_75t_L g4237 ( 
.A(n_4116),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_4118),
.Y(n_4238)
);

AO21x2_ASAP7_75t_L g4239 ( 
.A1(n_4140),
.A2(n_317),
.B(n_318),
.Y(n_4239)
);

OR2x6_ASAP7_75t_L g4240 ( 
.A(n_4115),
.B(n_317),
.Y(n_4240)
);

INVx4_ASAP7_75t_L g4241 ( 
.A(n_4124),
.Y(n_4241)
);

OAI22xp33_ASAP7_75t_L g4242 ( 
.A1(n_4020),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_4002),
.Y(n_4243)
);

INVx2_ASAP7_75t_L g4244 ( 
.A(n_4005),
.Y(n_4244)
);

INVx2_ASAP7_75t_L g4245 ( 
.A(n_4009),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_4013),
.Y(n_4246)
);

AOI22xp33_ASAP7_75t_L g4247 ( 
.A1(n_4063),
.A2(n_321),
.B1(n_319),
.B2(n_320),
.Y(n_4247)
);

NAND2xp5_ASAP7_75t_L g4248 ( 
.A(n_4018),
.B(n_322),
.Y(n_4248)
);

OAI22xp5_ASAP7_75t_L g4249 ( 
.A1(n_4093),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_4023),
.B(n_323),
.Y(n_4250)
);

INVx2_ASAP7_75t_L g4251 ( 
.A(n_4118),
.Y(n_4251)
);

INVx3_ASAP7_75t_L g4252 ( 
.A(n_4105),
.Y(n_4252)
);

NAND2x1p5_ASAP7_75t_L g4253 ( 
.A(n_4105),
.B(n_324),
.Y(n_4253)
);

HB1xp67_ASAP7_75t_L g4254 ( 
.A(n_4052),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4110),
.Y(n_4255)
);

NAND2x1p5_ASAP7_75t_L g4256 ( 
.A(n_4033),
.B(n_325),
.Y(n_4256)
);

INVx2_ASAP7_75t_L g4257 ( 
.A(n_4081),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_4092),
.Y(n_4258)
);

INVx2_ASAP7_75t_L g4259 ( 
.A(n_4113),
.Y(n_4259)
);

OA21x2_ASAP7_75t_L g4260 ( 
.A1(n_4129),
.A2(n_326),
.B(n_327),
.Y(n_4260)
);

INVx2_ASAP7_75t_L g4261 ( 
.A(n_4126),
.Y(n_4261)
);

AOI22xp33_ASAP7_75t_L g4262 ( 
.A1(n_4080),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.Y(n_4262)
);

BUFx4f_ASAP7_75t_SL g4263 ( 
.A(n_4050),
.Y(n_4263)
);

CKINVDCx20_ASAP7_75t_R g4264 ( 
.A(n_4079),
.Y(n_4264)
);

HB1xp67_ASAP7_75t_L g4265 ( 
.A(n_4144),
.Y(n_4265)
);

NOR2x1_ASAP7_75t_SL g4266 ( 
.A(n_4049),
.B(n_4031),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_4137),
.Y(n_4267)
);

INVx3_ASAP7_75t_L g4268 ( 
.A(n_4056),
.Y(n_4268)
);

OAI22xp33_ASAP7_75t_L g4269 ( 
.A1(n_4046),
.A2(n_330),
.B1(n_328),
.B2(n_329),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4137),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4143),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_4143),
.Y(n_4272)
);

OR2x2_ASAP7_75t_L g4273 ( 
.A(n_4032),
.B(n_330),
.Y(n_4273)
);

HB1xp67_ASAP7_75t_L g4274 ( 
.A(n_4008),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4145),
.Y(n_4275)
);

AOI22xp33_ASAP7_75t_SL g4276 ( 
.A1(n_4070),
.A2(n_333),
.B1(n_331),
.B2(n_332),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_4145),
.Y(n_4277)
);

INVx1_ASAP7_75t_L g4278 ( 
.A(n_4147),
.Y(n_4278)
);

BUFx4f_ASAP7_75t_L g4279 ( 
.A(n_4001),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4147),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_4141),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_4008),
.Y(n_4282)
);

INVx3_ASAP7_75t_L g4283 ( 
.A(n_4038),
.Y(n_4283)
);

BUFx6f_ASAP7_75t_L g4284 ( 
.A(n_4090),
.Y(n_4284)
);

INVxp67_ASAP7_75t_L g4285 ( 
.A(n_4144),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4003),
.B(n_333),
.Y(n_4286)
);

BUFx6f_ASAP7_75t_L g4287 ( 
.A(n_4066),
.Y(n_4287)
);

OAI21x1_ASAP7_75t_L g4288 ( 
.A1(n_4059),
.A2(n_334),
.B(n_335),
.Y(n_4288)
);

AOI22xp33_ASAP7_75t_SL g4289 ( 
.A1(n_4070),
.A2(n_337),
.B1(n_335),
.B2(n_336),
.Y(n_4289)
);

INVx1_ASAP7_75t_L g4290 ( 
.A(n_4043),
.Y(n_4290)
);

BUFx3_ASAP7_75t_L g4291 ( 
.A(n_4142),
.Y(n_4291)
);

HB1xp67_ASAP7_75t_L g4292 ( 
.A(n_4004),
.Y(n_4292)
);

INVx2_ASAP7_75t_L g4293 ( 
.A(n_4074),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_4027),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4091),
.Y(n_4295)
);

BUFx2_ASAP7_75t_L g4296 ( 
.A(n_4007),
.Y(n_4296)
);

AOI22xp5_ASAP7_75t_L g4297 ( 
.A1(n_4039),
.A2(n_338),
.B1(n_336),
.B2(n_337),
.Y(n_4297)
);

OAI21x1_ASAP7_75t_L g4298 ( 
.A1(n_4028),
.A2(n_339),
.B(n_340),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_4260),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4260),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_4292),
.B(n_4232),
.Y(n_4301)
);

INVx1_ASAP7_75t_L g4302 ( 
.A(n_4254),
.Y(n_4302)
);

INVx2_ASAP7_75t_L g4303 ( 
.A(n_4232),
.Y(n_4303)
);

BUFx2_ASAP7_75t_L g4304 ( 
.A(n_4222),
.Y(n_4304)
);

OAI221xp5_ASAP7_75t_L g4305 ( 
.A1(n_4292),
.A2(n_4122),
.B1(n_4026),
.B2(n_4096),
.C(n_4086),
.Y(n_4305)
);

BUFx2_ASAP7_75t_L g4306 ( 
.A(n_4154),
.Y(n_4306)
);

INVx2_ASAP7_75t_L g4307 ( 
.A(n_4152),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4254),
.Y(n_4308)
);

CKINVDCx5p33_ASAP7_75t_R g4309 ( 
.A(n_4153),
.Y(n_4309)
);

INVx1_ASAP7_75t_L g4310 ( 
.A(n_4255),
.Y(n_4310)
);

INVx2_ASAP7_75t_L g4311 ( 
.A(n_4163),
.Y(n_4311)
);

AND2x2_ASAP7_75t_L g4312 ( 
.A(n_4266),
.B(n_4111),
.Y(n_4312)
);

NOR2x1_ASAP7_75t_L g4313 ( 
.A(n_4159),
.B(n_4058),
.Y(n_4313)
);

AND2x4_ASAP7_75t_L g4314 ( 
.A(n_4154),
.B(n_4004),
.Y(n_4314)
);

HB1xp67_ASAP7_75t_L g4315 ( 
.A(n_4150),
.Y(n_4315)
);

INVx2_ASAP7_75t_L g4316 ( 
.A(n_4295),
.Y(n_4316)
);

OAI21xp5_ASAP7_75t_L g4317 ( 
.A1(n_4219),
.A2(n_4123),
.B(n_4075),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4157),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4173),
.Y(n_4319)
);

OAI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_4219),
.A2(n_4297),
.B(n_4285),
.Y(n_4320)
);

NAND2x1p5_ASAP7_75t_L g4321 ( 
.A(n_4199),
.B(n_4036),
.Y(n_4321)
);

INVx1_ASAP7_75t_L g4322 ( 
.A(n_4176),
.Y(n_4322)
);

BUFx12f_ASAP7_75t_L g4323 ( 
.A(n_4156),
.Y(n_4323)
);

AOI222xp33_ASAP7_75t_L g4324 ( 
.A1(n_4285),
.A2(n_4064),
.B1(n_4114),
.B2(n_4104),
.C1(n_4117),
.C2(n_4127),
.Y(n_4324)
);

OA21x2_ASAP7_75t_L g4325 ( 
.A1(n_4202),
.A2(n_4061),
.B(n_4088),
.Y(n_4325)
);

INVx1_ASAP7_75t_L g4326 ( 
.A(n_4181),
.Y(n_4326)
);

INVx1_ASAP7_75t_L g4327 ( 
.A(n_4187),
.Y(n_4327)
);

INVx1_ASAP7_75t_L g4328 ( 
.A(n_4188),
.Y(n_4328)
);

AND2x4_ASAP7_75t_L g4329 ( 
.A(n_4294),
.B(n_4004),
.Y(n_4329)
);

INVx2_ASAP7_75t_L g4330 ( 
.A(n_4293),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_4283),
.B(n_4132),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_4282),
.Y(n_4332)
);

AND2x2_ASAP7_75t_L g4333 ( 
.A(n_4283),
.B(n_4025),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_4195),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4177),
.Y(n_4335)
);

BUFx2_ASAP7_75t_L g4336 ( 
.A(n_4158),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4241),
.B(n_4025),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4180),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4201),
.Y(n_4339)
);

AOI22xp33_ASAP7_75t_L g4340 ( 
.A1(n_4229),
.A2(n_4100),
.B1(n_4146),
.B2(n_4130),
.Y(n_4340)
);

AOI22xp5_ASAP7_75t_L g4341 ( 
.A1(n_4276),
.A2(n_4100),
.B1(n_4139),
.B2(n_4099),
.Y(n_4341)
);

INVx2_ASAP7_75t_L g4342 ( 
.A(n_4224),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4196),
.Y(n_4343)
);

AND2x4_ASAP7_75t_L g4344 ( 
.A(n_4212),
.B(n_4025),
.Y(n_4344)
);

CKINVDCx16_ASAP7_75t_R g4345 ( 
.A(n_4264),
.Y(n_4345)
);

AND2x2_ASAP7_75t_L g4346 ( 
.A(n_4241),
.B(n_4207),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4228),
.Y(n_4347)
);

CKINVDCx5p33_ASAP7_75t_R g4348 ( 
.A(n_4156),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4251),
.Y(n_4349)
);

NAND2x1p5_ASAP7_75t_L g4350 ( 
.A(n_4160),
.B(n_4135),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_4205),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_4166),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4208),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_4167),
.Y(n_4354)
);

BUFx3_ASAP7_75t_L g4355 ( 
.A(n_4158),
.Y(n_4355)
);

BUFx3_ASAP7_75t_L g4356 ( 
.A(n_4158),
.Y(n_4356)
);

INVx2_ASAP7_75t_SL g4357 ( 
.A(n_4279),
.Y(n_4357)
);

INVx3_ASAP7_75t_L g4358 ( 
.A(n_4159),
.Y(n_4358)
);

INVx1_ASAP7_75t_L g4359 ( 
.A(n_4209),
.Y(n_4359)
);

INVxp33_ASAP7_75t_L g4360 ( 
.A(n_4170),
.Y(n_4360)
);

HB1xp67_ASAP7_75t_L g4361 ( 
.A(n_4150),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4215),
.Y(n_4362)
);

OAI22xp5_ASAP7_75t_L g4363 ( 
.A1(n_4155),
.A2(n_4138),
.B1(n_4076),
.B2(n_4128),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4223),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4271),
.Y(n_4365)
);

INVx2_ASAP7_75t_L g4366 ( 
.A(n_4277),
.Y(n_4366)
);

INVx1_ASAP7_75t_L g4367 ( 
.A(n_4227),
.Y(n_4367)
);

INVx3_ASAP7_75t_L g4368 ( 
.A(n_4217),
.Y(n_4368)
);

INVx1_ASAP7_75t_L g4369 ( 
.A(n_4185),
.Y(n_4369)
);

BUFx2_ASAP7_75t_SL g4370 ( 
.A(n_4206),
.Y(n_4370)
);

BUFx3_ASAP7_75t_L g4371 ( 
.A(n_4214),
.Y(n_4371)
);

AND2x2_ASAP7_75t_L g4372 ( 
.A(n_4168),
.B(n_4136),
.Y(n_4372)
);

INVx3_ASAP7_75t_L g4373 ( 
.A(n_4217),
.Y(n_4373)
);

AND2x2_ASAP7_75t_L g4374 ( 
.A(n_4168),
.B(n_4101),
.Y(n_4374)
);

NAND2x1p5_ASAP7_75t_L g4375 ( 
.A(n_4198),
.B(n_4098),
.Y(n_4375)
);

INVx1_ASAP7_75t_L g4376 ( 
.A(n_4185),
.Y(n_4376)
);

OAI21x1_ASAP7_75t_L g4377 ( 
.A1(n_4252),
.A2(n_4103),
.B(n_339),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4225),
.Y(n_4378)
);

HB1xp67_ASAP7_75t_L g4379 ( 
.A(n_4174),
.Y(n_4379)
);

INVx2_ASAP7_75t_L g4380 ( 
.A(n_4287),
.Y(n_4380)
);

INVx1_ASAP7_75t_SL g4381 ( 
.A(n_4206),
.Y(n_4381)
);

AO21x2_ASAP7_75t_L g4382 ( 
.A1(n_4274),
.A2(n_340),
.B(n_341),
.Y(n_4382)
);

HB1xp67_ASAP7_75t_L g4383 ( 
.A(n_4174),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4287),
.Y(n_4384)
);

INVx2_ASAP7_75t_L g4385 ( 
.A(n_4287),
.Y(n_4385)
);

INVx1_ASAP7_75t_L g4386 ( 
.A(n_4225),
.Y(n_4386)
);

INVx2_ASAP7_75t_L g4387 ( 
.A(n_4239),
.Y(n_4387)
);

AND2x4_ASAP7_75t_L g4388 ( 
.A(n_4183),
.B(n_342),
.Y(n_4388)
);

INVx3_ASAP7_75t_L g4389 ( 
.A(n_4210),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_4265),
.B(n_343),
.Y(n_4390)
);

BUFx3_ASAP7_75t_L g4391 ( 
.A(n_4178),
.Y(n_4391)
);

INVx1_ASAP7_75t_L g4392 ( 
.A(n_4230),
.Y(n_4392)
);

AND2x2_ASAP7_75t_L g4393 ( 
.A(n_4162),
.B(n_343),
.Y(n_4393)
);

INVx2_ASAP7_75t_L g4394 ( 
.A(n_4239),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4231),
.Y(n_4395)
);

INVx1_ASAP7_75t_L g4396 ( 
.A(n_4234),
.Y(n_4396)
);

INVx1_ASAP7_75t_SL g4397 ( 
.A(n_4172),
.Y(n_4397)
);

INVx2_ASAP7_75t_L g4398 ( 
.A(n_4237),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4238),
.Y(n_4399)
);

INVx1_ASAP7_75t_L g4400 ( 
.A(n_4151),
.Y(n_4400)
);

INVx2_ASAP7_75t_L g4401 ( 
.A(n_4284),
.Y(n_4401)
);

INVx2_ASAP7_75t_L g4402 ( 
.A(n_4284),
.Y(n_4402)
);

OAI21x1_ASAP7_75t_L g4403 ( 
.A1(n_4252),
.A2(n_345),
.B(n_346),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4248),
.Y(n_4404)
);

INVx1_ASAP7_75t_L g4405 ( 
.A(n_4248),
.Y(n_4405)
);

INVx1_ASAP7_75t_L g4406 ( 
.A(n_4250),
.Y(n_4406)
);

INVx1_ASAP7_75t_L g4407 ( 
.A(n_4250),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4284),
.Y(n_4408)
);

OAI21x1_ASAP7_75t_L g4409 ( 
.A1(n_4200),
.A2(n_346),
.B(n_347),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4267),
.Y(n_4410)
);

AND2x4_ASAP7_75t_L g4411 ( 
.A(n_4212),
.B(n_347),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4270),
.Y(n_4412)
);

INVx1_ASAP7_75t_L g4413 ( 
.A(n_4272),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4275),
.Y(n_4414)
);

INVx2_ASAP7_75t_L g4415 ( 
.A(n_4256),
.Y(n_4415)
);

INVx1_ASAP7_75t_L g4416 ( 
.A(n_4278),
.Y(n_4416)
);

AOI22xp33_ASAP7_75t_L g4417 ( 
.A1(n_4276),
.A2(n_350),
.B1(n_348),
.B2(n_349),
.Y(n_4417)
);

BUFx2_ASAP7_75t_L g4418 ( 
.A(n_4291),
.Y(n_4418)
);

INVx1_ASAP7_75t_L g4419 ( 
.A(n_4280),
.Y(n_4419)
);

INVx1_ASAP7_75t_L g4420 ( 
.A(n_4281),
.Y(n_4420)
);

O2A1O1Ixp33_ASAP7_75t_SL g4421 ( 
.A1(n_4172),
.A2(n_350),
.B(n_348),
.C(n_349),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4192),
.Y(n_4422)
);

AO21x2_ASAP7_75t_L g4423 ( 
.A1(n_4274),
.A2(n_351),
.B(n_352),
.Y(n_4423)
);

NAND2x1p5_ASAP7_75t_L g4424 ( 
.A(n_4210),
.B(n_352),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4179),
.Y(n_4425)
);

INVx1_ASAP7_75t_L g4426 ( 
.A(n_4233),
.Y(n_4426)
);

INVx1_ASAP7_75t_L g4427 ( 
.A(n_4233),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4218),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_4256),
.Y(n_4429)
);

HB1xp67_ASAP7_75t_L g4430 ( 
.A(n_4170),
.Y(n_4430)
);

BUFx2_ASAP7_75t_L g4431 ( 
.A(n_4183),
.Y(n_4431)
);

AND2x2_ASAP7_75t_L g4432 ( 
.A(n_4175),
.B(n_353),
.Y(n_4432)
);

OAI21x1_ASAP7_75t_L g4433 ( 
.A1(n_4200),
.A2(n_353),
.B(n_354),
.Y(n_4433)
);

INVx1_ASAP7_75t_L g4434 ( 
.A(n_4290),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4296),
.B(n_354),
.Y(n_4435)
);

OAI21x1_ASAP7_75t_L g4436 ( 
.A1(n_4164),
.A2(n_355),
.B(n_356),
.Y(n_4436)
);

AND2x2_ASAP7_75t_L g4437 ( 
.A(n_4190),
.B(n_356),
.Y(n_4437)
);

AO21x2_ASAP7_75t_L g4438 ( 
.A1(n_4297),
.A2(n_358),
.B(n_359),
.Y(n_4438)
);

HB1xp67_ASAP7_75t_L g4439 ( 
.A(n_4165),
.Y(n_4439)
);

INVx1_ASAP7_75t_L g4440 ( 
.A(n_4273),
.Y(n_4440)
);

INVx2_ASAP7_75t_L g4441 ( 
.A(n_4243),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_4244),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_4288),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4161),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4189),
.Y(n_4445)
);

INVx1_ASAP7_75t_L g4446 ( 
.A(n_4298),
.Y(n_4446)
);

HB1xp67_ASAP7_75t_L g4447 ( 
.A(n_4240),
.Y(n_4447)
);

INVx1_ASAP7_75t_SL g4448 ( 
.A(n_4263),
.Y(n_4448)
);

AND2x2_ASAP7_75t_L g4449 ( 
.A(n_4184),
.B(n_358),
.Y(n_4449)
);

OAI21xp5_ASAP7_75t_L g4450 ( 
.A1(n_4289),
.A2(n_360),
.B(n_361),
.Y(n_4450)
);

OR2x2_ASAP7_75t_L g4451 ( 
.A(n_4404),
.B(n_4268),
.Y(n_4451)
);

OR2x6_ASAP7_75t_L g4452 ( 
.A(n_4323),
.B(n_4240),
.Y(n_4452)
);

AOI211xp5_ASAP7_75t_L g4453 ( 
.A1(n_4317),
.A2(n_4320),
.B(n_4360),
.C(n_4337),
.Y(n_4453)
);

NAND3xp33_ASAP7_75t_L g4454 ( 
.A(n_4340),
.B(n_4289),
.C(n_4235),
.Y(n_4454)
);

OR2x4_ASAP7_75t_L g4455 ( 
.A(n_4425),
.B(n_4182),
.Y(n_4455)
);

AOI21xp33_ASAP7_75t_L g4456 ( 
.A1(n_4360),
.A2(n_4249),
.B(n_4203),
.Y(n_4456)
);

AOI221xp5_ASAP7_75t_L g4457 ( 
.A1(n_4439),
.A2(n_4249),
.B1(n_4242),
.B2(n_4226),
.C(n_4186),
.Y(n_4457)
);

AND2x2_ASAP7_75t_L g4458 ( 
.A(n_4346),
.B(n_4268),
.Y(n_4458)
);

AND2x2_ASAP7_75t_L g4459 ( 
.A(n_4418),
.B(n_4182),
.Y(n_4459)
);

AOI22xp33_ASAP7_75t_L g4460 ( 
.A1(n_4299),
.A2(n_4194),
.B1(n_4235),
.B2(n_4236),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_4397),
.B(n_4193),
.Y(n_4461)
);

AOI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_4341),
.A2(n_4171),
.B1(n_4203),
.B2(n_4193),
.Y(n_4462)
);

INVx1_ASAP7_75t_L g4463 ( 
.A(n_4315),
.Y(n_4463)
);

OAI221xp5_ASAP7_75t_L g4464 ( 
.A1(n_4340),
.A2(n_4171),
.B1(n_4262),
.B2(n_4247),
.C(n_4240),
.Y(n_4464)
);

OR2x2_ASAP7_75t_L g4465 ( 
.A(n_4405),
.B(n_4220),
.Y(n_4465)
);

BUFx2_ASAP7_75t_L g4466 ( 
.A(n_4323),
.Y(n_4466)
);

NAND4xp25_ASAP7_75t_L g4467 ( 
.A(n_4381),
.B(n_4197),
.C(n_4286),
.D(n_4279),
.Y(n_4467)
);

BUFx2_ASAP7_75t_L g4468 ( 
.A(n_4371),
.Y(n_4468)
);

OR2x2_ASAP7_75t_L g4469 ( 
.A(n_4406),
.B(n_4407),
.Y(n_4469)
);

INVx2_ASAP7_75t_SL g4470 ( 
.A(n_4345),
.Y(n_4470)
);

OAI22xp5_ASAP7_75t_L g4471 ( 
.A1(n_4313),
.A2(n_4253),
.B1(n_4182),
.B2(n_4213),
.Y(n_4471)
);

AOI22xp33_ASAP7_75t_L g4472 ( 
.A1(n_4299),
.A2(n_4169),
.B1(n_4246),
.B2(n_4245),
.Y(n_4472)
);

OAI21x1_ASAP7_75t_L g4473 ( 
.A1(n_4321),
.A2(n_4221),
.B(n_4204),
.Y(n_4473)
);

INVxp67_ASAP7_75t_SL g4474 ( 
.A(n_4447),
.Y(n_4474)
);

AOI222xp33_ASAP7_75t_L g4475 ( 
.A1(n_4450),
.A2(n_4269),
.B1(n_4261),
.B2(n_4259),
.C1(n_4258),
.C2(n_4257),
.Y(n_4475)
);

AOI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_4390),
.A2(n_4216),
.B(n_4253),
.Y(n_4476)
);

AND2x2_ASAP7_75t_L g4477 ( 
.A(n_4374),
.B(n_4213),
.Y(n_4477)
);

BUFx12f_ASAP7_75t_L g4478 ( 
.A(n_4348),
.Y(n_4478)
);

HB1xp67_ASAP7_75t_L g4479 ( 
.A(n_4306),
.Y(n_4479)
);

OAI22xp5_ASAP7_75t_L g4480 ( 
.A1(n_4430),
.A2(n_4213),
.B1(n_4204),
.B2(n_4191),
.Y(n_4480)
);

OAI22xp5_ASAP7_75t_L g4481 ( 
.A1(n_4430),
.A2(n_4191),
.B1(n_4211),
.B2(n_362),
.Y(n_4481)
);

AOI221xp5_ASAP7_75t_L g4482 ( 
.A1(n_4439),
.A2(n_360),
.B1(n_361),
.B2(n_362),
.C(n_363),
.Y(n_4482)
);

BUFx3_ASAP7_75t_L g4483 ( 
.A(n_4304),
.Y(n_4483)
);

OAI211xp5_ASAP7_75t_L g4484 ( 
.A1(n_4324),
.A2(n_365),
.B(n_363),
.C(n_364),
.Y(n_4484)
);

OAI22xp33_ASAP7_75t_L g4485 ( 
.A1(n_4300),
.A2(n_367),
.B1(n_364),
.B2(n_366),
.Y(n_4485)
);

OAI21xp33_ASAP7_75t_L g4486 ( 
.A1(n_4333),
.A2(n_366),
.B(n_367),
.Y(n_4486)
);

AOI22xp33_ASAP7_75t_L g4487 ( 
.A1(n_4300),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_4487)
);

AOI22xp33_ASAP7_75t_L g4488 ( 
.A1(n_4387),
.A2(n_370),
.B1(n_368),
.B2(n_369),
.Y(n_4488)
);

INVx2_ASAP7_75t_L g4489 ( 
.A(n_4411),
.Y(n_4489)
);

INVx1_ASAP7_75t_L g4490 ( 
.A(n_4315),
.Y(n_4490)
);

OAI22xp5_ASAP7_75t_L g4491 ( 
.A1(n_4447),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_4491)
);

NAND2x1_ASAP7_75t_L g4492 ( 
.A(n_4344),
.B(n_371),
.Y(n_4492)
);

OAI22xp5_ASAP7_75t_L g4493 ( 
.A1(n_4350),
.A2(n_375),
.B1(n_372),
.B2(n_374),
.Y(n_4493)
);

OAI22xp5_ASAP7_75t_L g4494 ( 
.A1(n_4350),
.A2(n_377),
.B1(n_375),
.B2(n_376),
.Y(n_4494)
);

INVx1_ASAP7_75t_L g4495 ( 
.A(n_4361),
.Y(n_4495)
);

AND2x2_ASAP7_75t_L g4496 ( 
.A(n_4331),
.B(n_376),
.Y(n_4496)
);

AOI22xp33_ASAP7_75t_L g4497 ( 
.A1(n_4387),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_4497)
);

OAI211xp5_ASAP7_75t_L g4498 ( 
.A1(n_4301),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_4498)
);

OAI221xp5_ASAP7_75t_L g4499 ( 
.A1(n_4426),
.A2(n_4427),
.B1(n_4305),
.B2(n_4394),
.C(n_4375),
.Y(n_4499)
);

AOI22xp33_ASAP7_75t_L g4500 ( 
.A1(n_4394),
.A2(n_383),
.B1(n_381),
.B2(n_382),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4372),
.B(n_381),
.Y(n_4501)
);

OAI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_4428),
.A2(n_384),
.B1(n_382),
.B2(n_383),
.Y(n_4502)
);

INVx2_ASAP7_75t_L g4503 ( 
.A(n_4411),
.Y(n_4503)
);

AOI22xp5_ASAP7_75t_L g4504 ( 
.A1(n_4438),
.A2(n_386),
.B1(n_384),
.B2(n_385),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4411),
.Y(n_4505)
);

INVx1_ASAP7_75t_L g4506 ( 
.A(n_4361),
.Y(n_4506)
);

INVx1_ASAP7_75t_L g4507 ( 
.A(n_4379),
.Y(n_4507)
);

AOI221xp5_ASAP7_75t_L g4508 ( 
.A1(n_4329),
.A2(n_386),
.B1(n_387),
.B2(n_388),
.C(n_389),
.Y(n_4508)
);

AND2x2_ASAP7_75t_L g4509 ( 
.A(n_4312),
.B(n_4336),
.Y(n_4509)
);

INVx1_ASAP7_75t_L g4510 ( 
.A(n_4379),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4436),
.Y(n_4511)
);

INVx3_ASAP7_75t_L g4512 ( 
.A(n_4371),
.Y(n_4512)
);

BUFx5_ASAP7_75t_L g4513 ( 
.A(n_4355),
.Y(n_4513)
);

OAI22xp33_ASAP7_75t_L g4514 ( 
.A1(n_4303),
.A2(n_391),
.B1(n_388),
.B2(n_390),
.Y(n_4514)
);

A2O1A1Ixp33_ASAP7_75t_L g4515 ( 
.A1(n_4314),
.A2(n_393),
.B(n_390),
.C(n_392),
.Y(n_4515)
);

NAND2xp5_ASAP7_75t_L g4516 ( 
.A(n_4378),
.B(n_4386),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_4382),
.B(n_393),
.Y(n_4517)
);

AOI211xp5_ASAP7_75t_L g4518 ( 
.A1(n_4421),
.A2(n_396),
.B(n_394),
.C(n_395),
.Y(n_4518)
);

NAND2xp5_ASAP7_75t_L g4519 ( 
.A(n_4382),
.B(n_394),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4355),
.Y(n_4520)
);

INVx1_ASAP7_75t_L g4521 ( 
.A(n_4383),
.Y(n_4521)
);

AOI22xp33_ASAP7_75t_L g4522 ( 
.A1(n_4332),
.A2(n_399),
.B1(n_395),
.B2(n_398),
.Y(n_4522)
);

INVx2_ASAP7_75t_SL g4523 ( 
.A(n_4448),
.Y(n_4523)
);

AOI22xp33_ASAP7_75t_L g4524 ( 
.A1(n_4332),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_4524)
);

AOI222xp33_ASAP7_75t_SL g4525 ( 
.A1(n_4302),
.A2(n_400),
.B1(n_401),
.B2(n_402),
.C1(n_403),
.C2(n_406),
.Y(n_4525)
);

AOI22xp33_ASAP7_75t_L g4526 ( 
.A1(n_4438),
.A2(n_407),
.B1(n_402),
.B2(n_406),
.Y(n_4526)
);

AO21x2_ASAP7_75t_L g4527 ( 
.A1(n_4303),
.A2(n_408),
.B(n_409),
.Y(n_4527)
);

OAI21x1_ASAP7_75t_L g4528 ( 
.A1(n_4321),
.A2(n_408),
.B(n_409),
.Y(n_4528)
);

AOI22xp33_ASAP7_75t_L g4529 ( 
.A1(n_4352),
.A2(n_412),
.B1(n_410),
.B2(n_411),
.Y(n_4529)
);

AND2x4_ASAP7_75t_L g4530 ( 
.A(n_4356),
.B(n_410),
.Y(n_4530)
);

INVx3_ASAP7_75t_L g4531 ( 
.A(n_4356),
.Y(n_4531)
);

AOI22xp33_ASAP7_75t_L g4532 ( 
.A1(n_4352),
.A2(n_414),
.B1(n_412),
.B2(n_413),
.Y(n_4532)
);

AOI21xp5_ASAP7_75t_L g4533 ( 
.A1(n_4344),
.A2(n_415),
.B(n_416),
.Y(n_4533)
);

AOI22xp33_ASAP7_75t_L g4534 ( 
.A1(n_4354),
.A2(n_418),
.B1(n_415),
.B2(n_417),
.Y(n_4534)
);

AOI22xp33_ASAP7_75t_SL g4535 ( 
.A1(n_4314),
.A2(n_421),
.B1(n_419),
.B2(n_420),
.Y(n_4535)
);

INVx1_ASAP7_75t_L g4536 ( 
.A(n_4383),
.Y(n_4536)
);

BUFx6f_ASAP7_75t_L g4537 ( 
.A(n_4348),
.Y(n_4537)
);

NOR4xp25_ASAP7_75t_L g4538 ( 
.A(n_4421),
.B(n_4422),
.C(n_4444),
.D(n_4443),
.Y(n_4538)
);

OAI22xp33_ASAP7_75t_L g4539 ( 
.A1(n_4375),
.A2(n_424),
.B1(n_422),
.B2(n_423),
.Y(n_4539)
);

OAI22xp5_ASAP7_75t_L g4540 ( 
.A1(n_4344),
.A2(n_425),
.B1(n_422),
.B2(n_423),
.Y(n_4540)
);

INVx2_ASAP7_75t_L g4541 ( 
.A(n_4423),
.Y(n_4541)
);

AOI22xp33_ASAP7_75t_L g4542 ( 
.A1(n_4354),
.A2(n_427),
.B1(n_425),
.B2(n_426),
.Y(n_4542)
);

AOI211xp5_ASAP7_75t_L g4543 ( 
.A1(n_4363),
.A2(n_426),
.B(n_427),
.C(n_428),
.Y(n_4543)
);

AOI22xp33_ASAP7_75t_L g4544 ( 
.A1(n_4423),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_4544)
);

AND2x2_ASAP7_75t_L g4545 ( 
.A(n_4370),
.B(n_433),
.Y(n_4545)
);

AND2x2_ASAP7_75t_L g4546 ( 
.A(n_4389),
.B(n_433),
.Y(n_4546)
);

OA21x2_ASAP7_75t_L g4547 ( 
.A1(n_4380),
.A2(n_434),
.B(n_435),
.Y(n_4547)
);

INVx1_ASAP7_75t_L g4548 ( 
.A(n_4310),
.Y(n_4548)
);

OAI221xp5_ASAP7_75t_L g4549 ( 
.A1(n_4330),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.C(n_439),
.Y(n_4549)
);

AOI22xp33_ASAP7_75t_L g4550 ( 
.A1(n_4330),
.A2(n_436),
.B1(n_438),
.B2(n_439),
.Y(n_4550)
);

INVx6_ASAP7_75t_L g4551 ( 
.A(n_4388),
.Y(n_4551)
);

AND2x2_ASAP7_75t_L g4552 ( 
.A(n_4389),
.B(n_440),
.Y(n_4552)
);

OAI22xp5_ASAP7_75t_L g4553 ( 
.A1(n_4314),
.A2(n_440),
.B1(n_441),
.B2(n_442),
.Y(n_4553)
);

OAI22xp5_ASAP7_75t_L g4554 ( 
.A1(n_4440),
.A2(n_441),
.B1(n_443),
.B2(n_444),
.Y(n_4554)
);

OAI22xp5_ASAP7_75t_SL g4555 ( 
.A1(n_4424),
.A2(n_4357),
.B1(n_4391),
.B2(n_4388),
.Y(n_4555)
);

AOI21xp5_ASAP7_75t_L g4556 ( 
.A1(n_4329),
.A2(n_443),
.B(n_444),
.Y(n_4556)
);

NAND2xp5_ASAP7_75t_L g4557 ( 
.A(n_4446),
.B(n_445),
.Y(n_4557)
);

AND2x2_ASAP7_75t_L g4558 ( 
.A(n_4445),
.B(n_446),
.Y(n_4558)
);

NAND3xp33_ASAP7_75t_L g4559 ( 
.A(n_4329),
.B(n_447),
.C(n_448),
.Y(n_4559)
);

AOI21xp33_ASAP7_75t_SL g4560 ( 
.A1(n_4424),
.A2(n_449),
.B(n_450),
.Y(n_4560)
);

OAI22xp33_ASAP7_75t_L g4561 ( 
.A1(n_4415),
.A2(n_450),
.B1(n_451),
.B2(n_453),
.Y(n_4561)
);

OAI221xp5_ASAP7_75t_L g4562 ( 
.A1(n_4380),
.A2(n_451),
.B1(n_453),
.B2(n_454),
.C(n_455),
.Y(n_4562)
);

AOI22xp33_ASAP7_75t_L g4563 ( 
.A1(n_4307),
.A2(n_455),
.B1(n_456),
.B2(n_457),
.Y(n_4563)
);

OAI21xp33_ASAP7_75t_L g4564 ( 
.A1(n_4369),
.A2(n_456),
.B(n_457),
.Y(n_4564)
);

NAND2xp5_ASAP7_75t_L g4565 ( 
.A(n_4420),
.B(n_458),
.Y(n_4565)
);

NOR2xp33_ASAP7_75t_L g4566 ( 
.A(n_4309),
.B(n_458),
.Y(n_4566)
);

OAI21x1_ASAP7_75t_L g4567 ( 
.A1(n_4384),
.A2(n_459),
.B(n_460),
.Y(n_4567)
);

OA21x2_ASAP7_75t_L g4568 ( 
.A1(n_4384),
.A2(n_459),
.B(n_460),
.Y(n_4568)
);

AOI221xp5_ASAP7_75t_L g4569 ( 
.A1(n_4316),
.A2(n_461),
.B1(n_462),
.B2(n_464),
.C(n_465),
.Y(n_4569)
);

OAI22xp5_ASAP7_75t_L g4570 ( 
.A1(n_4431),
.A2(n_461),
.B1(n_464),
.B2(n_465),
.Y(n_4570)
);

INVx2_ASAP7_75t_SL g4571 ( 
.A(n_4309),
.Y(n_4571)
);

AOI221xp5_ASAP7_75t_L g4572 ( 
.A1(n_4316),
.A2(n_466),
.B1(n_467),
.B2(n_468),
.C(n_469),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4308),
.Y(n_4573)
);

AOI22xp33_ASAP7_75t_L g4574 ( 
.A1(n_4307),
.A2(n_467),
.B1(n_469),
.B2(n_471),
.Y(n_4574)
);

INVx1_ASAP7_75t_L g4575 ( 
.A(n_4318),
.Y(n_4575)
);

INVx1_ASAP7_75t_L g4576 ( 
.A(n_4319),
.Y(n_4576)
);

OAI22xp33_ASAP7_75t_L g4577 ( 
.A1(n_4415),
.A2(n_471),
.B1(n_472),
.B2(n_473),
.Y(n_4577)
);

INVx2_ASAP7_75t_L g4578 ( 
.A(n_4429),
.Y(n_4578)
);

AOI22xp33_ASAP7_75t_L g4579 ( 
.A1(n_4311),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.Y(n_4579)
);

AOI22xp33_ASAP7_75t_L g4580 ( 
.A1(n_4311),
.A2(n_475),
.B1(n_476),
.B2(n_477),
.Y(n_4580)
);

AND2x2_ASAP7_75t_L g4581 ( 
.A(n_4368),
.B(n_475),
.Y(n_4581)
);

AOI21xp5_ASAP7_75t_L g4582 ( 
.A1(n_4325),
.A2(n_477),
.B(n_478),
.Y(n_4582)
);

AOI22xp33_ASAP7_75t_L g4583 ( 
.A1(n_4429),
.A2(n_478),
.B1(n_479),
.B2(n_480),
.Y(n_4583)
);

HB1xp67_ASAP7_75t_L g4584 ( 
.A(n_4322),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_4326),
.Y(n_4585)
);

HB1xp67_ASAP7_75t_SL g4586 ( 
.A(n_4391),
.Y(n_4586)
);

INVx1_ASAP7_75t_L g4587 ( 
.A(n_4327),
.Y(n_4587)
);

OR2x6_ASAP7_75t_L g4588 ( 
.A(n_4435),
.B(n_479),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_4368),
.B(n_481),
.Y(n_4589)
);

AND2x4_ASAP7_75t_L g4590 ( 
.A(n_4470),
.B(n_4358),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4453),
.B(n_4376),
.Y(n_4591)
);

HB1xp67_ASAP7_75t_L g4592 ( 
.A(n_4479),
.Y(n_4592)
);

INVx2_ASAP7_75t_L g4593 ( 
.A(n_4468),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4474),
.Y(n_4594)
);

INVx1_ASAP7_75t_L g4595 ( 
.A(n_4584),
.Y(n_4595)
);

AND2x2_ASAP7_75t_L g4596 ( 
.A(n_4512),
.B(n_4358),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_4469),
.Y(n_4597)
);

INVx2_ASAP7_75t_L g4598 ( 
.A(n_4523),
.Y(n_4598)
);

INVx2_ASAP7_75t_L g4599 ( 
.A(n_4492),
.Y(n_4599)
);

INVx2_ASAP7_75t_L g4600 ( 
.A(n_4513),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4513),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_4513),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4512),
.B(n_4373),
.Y(n_4603)
);

OR2x2_ASAP7_75t_L g4604 ( 
.A(n_4461),
.B(n_4434),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4459),
.B(n_4373),
.Y(n_4605)
);

AND2x2_ASAP7_75t_L g4606 ( 
.A(n_4509),
.B(n_4449),
.Y(n_4606)
);

NAND2xp5_ASAP7_75t_L g4607 ( 
.A(n_4538),
.B(n_4454),
.Y(n_4607)
);

NAND2xp5_ASAP7_75t_L g4608 ( 
.A(n_4582),
.B(n_4400),
.Y(n_4608)
);

INVx1_ASAP7_75t_L g4609 ( 
.A(n_4521),
.Y(n_4609)
);

INVx3_ASAP7_75t_L g4610 ( 
.A(n_4478),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4463),
.B(n_4490),
.Y(n_4611)
);

OR2x2_ASAP7_75t_L g4612 ( 
.A(n_4516),
.B(n_4328),
.Y(n_4612)
);

AND2x4_ASAP7_75t_L g4613 ( 
.A(n_4531),
.B(n_4437),
.Y(n_4613)
);

BUFx2_ASAP7_75t_L g4614 ( 
.A(n_4483),
.Y(n_4614)
);

INVx2_ASAP7_75t_L g4615 ( 
.A(n_4513),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4477),
.B(n_4393),
.Y(n_4616)
);

AND2x4_ASAP7_75t_SL g4617 ( 
.A(n_4452),
.B(n_4432),
.Y(n_4617)
);

BUFx3_ASAP7_75t_L g4618 ( 
.A(n_4537),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4521),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4495),
.Y(n_4620)
);

INVx2_ASAP7_75t_L g4621 ( 
.A(n_4513),
.Y(n_4621)
);

AND2x2_ASAP7_75t_L g4622 ( 
.A(n_4458),
.B(n_4334),
.Y(n_4622)
);

AND2x2_ASAP7_75t_L g4623 ( 
.A(n_4520),
.B(n_4343),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4506),
.B(n_4351),
.Y(n_4624)
);

HB1xp67_ASAP7_75t_L g4625 ( 
.A(n_4507),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4510),
.Y(n_4626)
);

OR2x2_ASAP7_75t_L g4627 ( 
.A(n_4451),
.B(n_4353),
.Y(n_4627)
);

INVx2_ASAP7_75t_L g4628 ( 
.A(n_4547),
.Y(n_4628)
);

HB1xp67_ASAP7_75t_L g4629 ( 
.A(n_4536),
.Y(n_4629)
);

AND2x2_ASAP7_75t_L g4630 ( 
.A(n_4531),
.B(n_4359),
.Y(n_4630)
);

INVx3_ASAP7_75t_L g4631 ( 
.A(n_4452),
.Y(n_4631)
);

INVx5_ASAP7_75t_L g4632 ( 
.A(n_4537),
.Y(n_4632)
);

INVx1_ASAP7_75t_L g4633 ( 
.A(n_4517),
.Y(n_4633)
);

BUFx2_ASAP7_75t_L g4634 ( 
.A(n_4455),
.Y(n_4634)
);

INVx1_ASAP7_75t_L g4635 ( 
.A(n_4519),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4543),
.B(n_4362),
.Y(n_4636)
);

INVx2_ASAP7_75t_L g4637 ( 
.A(n_4547),
.Y(n_4637)
);

OR2x2_ASAP7_75t_L g4638 ( 
.A(n_4465),
.B(n_4565),
.Y(n_4638)
);

INVx1_ASAP7_75t_L g4639 ( 
.A(n_4575),
.Y(n_4639)
);

AND2x2_ASAP7_75t_L g4640 ( 
.A(n_4551),
.B(n_4466),
.Y(n_4640)
);

INVx1_ASAP7_75t_L g4641 ( 
.A(n_4576),
.Y(n_4641)
);

OR2x2_ASAP7_75t_L g4642 ( 
.A(n_4557),
.B(n_4364),
.Y(n_4642)
);

NAND2xp5_ASAP7_75t_L g4643 ( 
.A(n_4548),
.B(n_4367),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_4585),
.Y(n_4644)
);

HB1xp67_ASAP7_75t_L g4645 ( 
.A(n_4573),
.Y(n_4645)
);

HB1xp67_ASAP7_75t_L g4646 ( 
.A(n_4511),
.Y(n_4646)
);

HB1xp67_ASAP7_75t_L g4647 ( 
.A(n_4587),
.Y(n_4647)
);

INVxp67_ASAP7_75t_SL g4648 ( 
.A(n_4559),
.Y(n_4648)
);

NOR2xp33_ASAP7_75t_L g4649 ( 
.A(n_4537),
.B(n_4325),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_L g4650 ( 
.A(n_4541),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4568),
.Y(n_4651)
);

INVx1_ASAP7_75t_L g4652 ( 
.A(n_4578),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4558),
.Y(n_4653)
);

INVx2_ASAP7_75t_L g4654 ( 
.A(n_4568),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4527),
.Y(n_4655)
);

NAND2xp5_ASAP7_75t_SL g4656 ( 
.A(n_4462),
.B(n_4385),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4527),
.Y(n_4657)
);

OR2x2_ASAP7_75t_L g4658 ( 
.A(n_4467),
.B(n_4392),
.Y(n_4658)
);

INVx2_ASAP7_75t_SL g4659 ( 
.A(n_4551),
.Y(n_4659)
);

AND2x2_ASAP7_75t_L g4660 ( 
.A(n_4545),
.B(n_4395),
.Y(n_4660)
);

AND2x2_ASAP7_75t_L g4661 ( 
.A(n_4496),
.B(n_4396),
.Y(n_4661)
);

INVx1_ASAP7_75t_L g4662 ( 
.A(n_4501),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_4460),
.B(n_4399),
.Y(n_4663)
);

INVx2_ASAP7_75t_L g4664 ( 
.A(n_4489),
.Y(n_4664)
);

INVx1_ASAP7_75t_L g4665 ( 
.A(n_4540),
.Y(n_4665)
);

INVx1_ASAP7_75t_L g4666 ( 
.A(n_4581),
.Y(n_4666)
);

NAND2xp5_ASAP7_75t_L g4667 ( 
.A(n_4556),
.B(n_4410),
.Y(n_4667)
);

AND2x4_ASAP7_75t_L g4668 ( 
.A(n_4503),
.B(n_4385),
.Y(n_4668)
);

HB1xp67_ASAP7_75t_L g4669 ( 
.A(n_4456),
.Y(n_4669)
);

INVx1_ASAP7_75t_L g4670 ( 
.A(n_4589),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4533),
.B(n_4412),
.Y(n_4671)
);

INVxp67_ASAP7_75t_SL g4672 ( 
.A(n_4484),
.Y(n_4672)
);

AND2x2_ASAP7_75t_L g4673 ( 
.A(n_4571),
.B(n_4413),
.Y(n_4673)
);

INVx1_ASAP7_75t_L g4674 ( 
.A(n_4505),
.Y(n_4674)
);

BUFx3_ASAP7_75t_L g4675 ( 
.A(n_4588),
.Y(n_4675)
);

INVxp67_ASAP7_75t_L g4676 ( 
.A(n_4586),
.Y(n_4676)
);

INVx1_ASAP7_75t_L g4677 ( 
.A(n_4504),
.Y(n_4677)
);

INVx1_ASAP7_75t_L g4678 ( 
.A(n_4553),
.Y(n_4678)
);

INVx2_ASAP7_75t_L g4679 ( 
.A(n_4528),
.Y(n_4679)
);

HB1xp67_ASAP7_75t_L g4680 ( 
.A(n_4493),
.Y(n_4680)
);

OR2x2_ASAP7_75t_L g4681 ( 
.A(n_4471),
.B(n_4414),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_L g4682 ( 
.A(n_4457),
.B(n_4416),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_L g4683 ( 
.A(n_4486),
.B(n_4419),
.Y(n_4683)
);

NAND2xp5_ASAP7_75t_L g4684 ( 
.A(n_4482),
.B(n_4398),
.Y(n_4684)
);

INVx1_ASAP7_75t_L g4685 ( 
.A(n_4546),
.Y(n_4685)
);

CKINVDCx14_ASAP7_75t_R g4686 ( 
.A(n_4555),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4508),
.B(n_4398),
.Y(n_4687)
);

INVx2_ASAP7_75t_L g4688 ( 
.A(n_4530),
.Y(n_4688)
);

OR2x2_ASAP7_75t_L g4689 ( 
.A(n_4481),
.B(n_4335),
.Y(n_4689)
);

INVx2_ASAP7_75t_SL g4690 ( 
.A(n_4530),
.Y(n_4690)
);

INVx4_ASAP7_75t_L g4691 ( 
.A(n_4552),
.Y(n_4691)
);

AND2x2_ASAP7_75t_L g4692 ( 
.A(n_4476),
.B(n_4325),
.Y(n_4692)
);

INVx2_ASAP7_75t_L g4693 ( 
.A(n_4588),
.Y(n_4693)
);

INVx1_ASAP7_75t_L g4694 ( 
.A(n_4567),
.Y(n_4694)
);

AND2x4_ASAP7_75t_SL g4695 ( 
.A(n_4566),
.B(n_4401),
.Y(n_4695)
);

OR2x2_ASAP7_75t_L g4696 ( 
.A(n_4499),
.B(n_4335),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4485),
.Y(n_4697)
);

NAND2xp5_ASAP7_75t_L g4698 ( 
.A(n_4515),
.B(n_4338),
.Y(n_4698)
);

INVx1_ASAP7_75t_L g4699 ( 
.A(n_4502),
.Y(n_4699)
);

INVx2_ASAP7_75t_L g4700 ( 
.A(n_4628),
.Y(n_4700)
);

NOR2xp33_ASAP7_75t_L g4701 ( 
.A(n_4607),
.B(n_4464),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_4592),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4592),
.Y(n_4703)
);

INVx1_ASAP7_75t_L g4704 ( 
.A(n_4650),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4606),
.B(n_4480),
.Y(n_4705)
);

HB1xp67_ASAP7_75t_L g4706 ( 
.A(n_4607),
.Y(n_4706)
);

AND2x4_ASAP7_75t_L g4707 ( 
.A(n_4613),
.B(n_4401),
.Y(n_4707)
);

AND2x2_ASAP7_75t_L g4708 ( 
.A(n_4614),
.B(n_4494),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4672),
.B(n_4653),
.Y(n_4709)
);

INVx1_ASAP7_75t_L g4710 ( 
.A(n_4650),
.Y(n_4710)
);

BUFx2_ASAP7_75t_L g4711 ( 
.A(n_4613),
.Y(n_4711)
);

NAND2xp5_ASAP7_75t_SL g4712 ( 
.A(n_4669),
.B(n_4539),
.Y(n_4712)
);

NAND2xp5_ASAP7_75t_L g4713 ( 
.A(n_4672),
.B(n_4535),
.Y(n_4713)
);

HB1xp67_ASAP7_75t_L g4714 ( 
.A(n_4648),
.Y(n_4714)
);

INVx2_ASAP7_75t_L g4715 ( 
.A(n_4637),
.Y(n_4715)
);

OR2x2_ASAP7_75t_L g4716 ( 
.A(n_4591),
.B(n_4554),
.Y(n_4716)
);

OAI21xp33_ASAP7_75t_L g4717 ( 
.A1(n_4591),
.A2(n_4564),
.B(n_4472),
.Y(n_4717)
);

AND2x2_ASAP7_75t_L g4718 ( 
.A(n_4616),
.B(n_4402),
.Y(n_4718)
);

AOI21xp33_ASAP7_75t_L g4719 ( 
.A1(n_4669),
.A2(n_4408),
.B(n_4402),
.Y(n_4719)
);

INVx1_ASAP7_75t_L g4720 ( 
.A(n_4625),
.Y(n_4720)
);

AND2x2_ASAP7_75t_L g4721 ( 
.A(n_4617),
.B(n_4408),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4625),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4661),
.B(n_4491),
.Y(n_4723)
);

INVx1_ASAP7_75t_SL g4724 ( 
.A(n_4632),
.Y(n_4724)
);

INVx1_ASAP7_75t_L g4725 ( 
.A(n_4629),
.Y(n_4725)
);

HB1xp67_ASAP7_75t_L g4726 ( 
.A(n_4648),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4629),
.Y(n_4727)
);

INVx2_ASAP7_75t_SL g4728 ( 
.A(n_4632),
.Y(n_4728)
);

INVxp67_ASAP7_75t_SL g4729 ( 
.A(n_4676),
.Y(n_4729)
);

INVx2_ASAP7_75t_SL g4730 ( 
.A(n_4632),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4647),
.Y(n_4731)
);

AND2x2_ASAP7_75t_L g4732 ( 
.A(n_4640),
.B(n_4475),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4691),
.B(n_4560),
.Y(n_4733)
);

AND2x4_ASAP7_75t_SL g4734 ( 
.A(n_4590),
.B(n_4583),
.Y(n_4734)
);

HB1xp67_ASAP7_75t_L g4735 ( 
.A(n_4680),
.Y(n_4735)
);

AND2x2_ASAP7_75t_L g4736 ( 
.A(n_4691),
.B(n_4377),
.Y(n_4736)
);

AND2x2_ASAP7_75t_L g4737 ( 
.A(n_4660),
.B(n_4473),
.Y(n_4737)
);

NAND2xp5_ASAP7_75t_L g4738 ( 
.A(n_4680),
.B(n_4498),
.Y(n_4738)
);

NOR2xp67_ASAP7_75t_L g4739 ( 
.A(n_4676),
.B(n_4338),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4647),
.Y(n_4740)
);

INVx2_ASAP7_75t_L g4741 ( 
.A(n_4651),
.Y(n_4741)
);

OR2x2_ASAP7_75t_L g4742 ( 
.A(n_4593),
.B(n_4598),
.Y(n_4742)
);

INVx1_ASAP7_75t_L g4743 ( 
.A(n_4645),
.Y(n_4743)
);

AND2x4_ASAP7_75t_SL g4744 ( 
.A(n_4590),
.B(n_4487),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_4662),
.B(n_4518),
.Y(n_4745)
);

INVx2_ASAP7_75t_SL g4746 ( 
.A(n_4632),
.Y(n_4746)
);

OR2x6_ASAP7_75t_SL g4747 ( 
.A(n_4682),
.B(n_4570),
.Y(n_4747)
);

AND2x2_ASAP7_75t_L g4748 ( 
.A(n_4695),
.B(n_4339),
.Y(n_4748)
);

AOI22xp33_ASAP7_75t_L g4749 ( 
.A1(n_4677),
.A2(n_4544),
.B1(n_4526),
.B2(n_4549),
.Y(n_4749)
);

AND2x2_ASAP7_75t_L g4750 ( 
.A(n_4605),
.B(n_4618),
.Y(n_4750)
);

AND2x2_ASAP7_75t_L g4751 ( 
.A(n_4686),
.B(n_4409),
.Y(n_4751)
);

HB1xp67_ASAP7_75t_L g4752 ( 
.A(n_4645),
.Y(n_4752)
);

OR2x2_ASAP7_75t_L g4753 ( 
.A(n_4597),
.B(n_4339),
.Y(n_4753)
);

AND2x2_ASAP7_75t_L g4754 ( 
.A(n_4603),
.B(n_4342),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4594),
.Y(n_4755)
);

INVx1_ASAP7_75t_L g4756 ( 
.A(n_4646),
.Y(n_4756)
);

INVx1_ASAP7_75t_L g4757 ( 
.A(n_4646),
.Y(n_4757)
);

AND2x4_ASAP7_75t_L g4758 ( 
.A(n_4631),
.B(n_4342),
.Y(n_4758)
);

AND2x2_ASAP7_75t_L g4759 ( 
.A(n_4634),
.B(n_4622),
.Y(n_4759)
);

INVx1_ASAP7_75t_L g4760 ( 
.A(n_4643),
.Y(n_4760)
);

INVx2_ASAP7_75t_L g4761 ( 
.A(n_4654),
.Y(n_4761)
);

AND2x2_ASAP7_75t_L g4762 ( 
.A(n_4610),
.B(n_4433),
.Y(n_4762)
);

AND2x2_ASAP7_75t_L g4763 ( 
.A(n_4610),
.B(n_4403),
.Y(n_4763)
);

INVx1_ASAP7_75t_L g4764 ( 
.A(n_4643),
.Y(n_4764)
);

AND2x2_ASAP7_75t_L g4765 ( 
.A(n_4596),
.B(n_4659),
.Y(n_4765)
);

AOI22xp33_ASAP7_75t_L g4766 ( 
.A1(n_4633),
.A2(n_4417),
.B1(n_4572),
.B2(n_4569),
.Y(n_4766)
);

INVx1_ASAP7_75t_L g4767 ( 
.A(n_4611),
.Y(n_4767)
);

AND2x2_ASAP7_75t_L g4768 ( 
.A(n_4735),
.B(n_4630),
.Y(n_4768)
);

INVx1_ASAP7_75t_SL g4769 ( 
.A(n_4751),
.Y(n_4769)
);

AND2x2_ASAP7_75t_L g4770 ( 
.A(n_4711),
.B(n_4729),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4752),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_4752),
.Y(n_4772)
);

INVx1_ASAP7_75t_L g4773 ( 
.A(n_4729),
.Y(n_4773)
);

INVxp67_ASAP7_75t_L g4774 ( 
.A(n_4735),
.Y(n_4774)
);

INVx2_ASAP7_75t_L g4775 ( 
.A(n_4714),
.Y(n_4775)
);

AND2x2_ASAP7_75t_L g4776 ( 
.A(n_4750),
.B(n_4759),
.Y(n_4776)
);

AND2x2_ASAP7_75t_L g4777 ( 
.A(n_4765),
.B(n_4673),
.Y(n_4777)
);

INVxp67_ASAP7_75t_L g4778 ( 
.A(n_4714),
.Y(n_4778)
);

AND2x2_ASAP7_75t_L g4779 ( 
.A(n_4708),
.B(n_4690),
.Y(n_4779)
);

INVx2_ASAP7_75t_L g4780 ( 
.A(n_4726),
.Y(n_4780)
);

HB1xp67_ASAP7_75t_L g4781 ( 
.A(n_4726),
.Y(n_4781)
);

AND2x2_ASAP7_75t_L g4782 ( 
.A(n_4705),
.B(n_4623),
.Y(n_4782)
);

AOI221xp5_ASAP7_75t_L g4783 ( 
.A1(n_4706),
.A2(n_4663),
.B1(n_4682),
.B2(n_4649),
.C(n_4635),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4700),
.Y(n_4784)
);

INVxp67_ASAP7_75t_L g4785 ( 
.A(n_4706),
.Y(n_4785)
);

OR2x2_ASAP7_75t_L g4786 ( 
.A(n_4709),
.B(n_4738),
.Y(n_4786)
);

BUFx2_ASAP7_75t_L g4787 ( 
.A(n_4733),
.Y(n_4787)
);

OR2x2_ASAP7_75t_L g4788 ( 
.A(n_4742),
.B(n_4663),
.Y(n_4788)
);

HB1xp67_ASAP7_75t_L g4789 ( 
.A(n_4713),
.Y(n_4789)
);

NAND2xp5_ASAP7_75t_L g4790 ( 
.A(n_4739),
.B(n_4666),
.Y(n_4790)
);

INVx2_ASAP7_75t_SL g4791 ( 
.A(n_4728),
.Y(n_4791)
);

AND2x4_ASAP7_75t_L g4792 ( 
.A(n_4728),
.B(n_4631),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4747),
.Y(n_4793)
);

HB1xp67_ASAP7_75t_L g4794 ( 
.A(n_4720),
.Y(n_4794)
);

OR2x2_ASAP7_75t_L g4795 ( 
.A(n_4723),
.B(n_4642),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4700),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4747),
.B(n_4670),
.Y(n_4797)
);

INVx1_ASAP7_75t_L g4798 ( 
.A(n_4715),
.Y(n_4798)
);

OAI21xp33_ASAP7_75t_L g4799 ( 
.A1(n_4701),
.A2(n_4658),
.B(n_4692),
.Y(n_4799)
);

AND2x2_ASAP7_75t_L g4800 ( 
.A(n_4718),
.B(n_4685),
.Y(n_4800)
);

AND2x2_ASAP7_75t_L g4801 ( 
.A(n_4762),
.B(n_4638),
.Y(n_4801)
);

BUFx3_ASAP7_75t_L g4802 ( 
.A(n_4730),
.Y(n_4802)
);

INVxp67_ASAP7_75t_SL g4803 ( 
.A(n_4712),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4715),
.Y(n_4804)
);

INVx1_ASAP7_75t_L g4805 ( 
.A(n_4741),
.Y(n_4805)
);

OR2x2_ASAP7_75t_L g4806 ( 
.A(n_4702),
.B(n_4612),
.Y(n_4806)
);

BUFx3_ASAP7_75t_L g4807 ( 
.A(n_4730),
.Y(n_4807)
);

BUFx2_ASAP7_75t_L g4808 ( 
.A(n_4707),
.Y(n_4808)
);

AND2x2_ASAP7_75t_L g4809 ( 
.A(n_4763),
.B(n_4688),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_4741),
.Y(n_4810)
);

AND2x2_ASAP7_75t_L g4811 ( 
.A(n_4754),
.B(n_4599),
.Y(n_4811)
);

INVx1_ASAP7_75t_SL g4812 ( 
.A(n_4732),
.Y(n_4812)
);

OR2x2_ASAP7_75t_L g4813 ( 
.A(n_4703),
.B(n_4636),
.Y(n_4813)
);

INVx1_ASAP7_75t_L g4814 ( 
.A(n_4761),
.Y(n_4814)
);

NAND2xp5_ASAP7_75t_L g4815 ( 
.A(n_4754),
.B(n_4699),
.Y(n_4815)
);

OR2x2_ASAP7_75t_L g4816 ( 
.A(n_4756),
.B(n_4636),
.Y(n_4816)
);

AND2x4_ASAP7_75t_L g4817 ( 
.A(n_4746),
.B(n_4675),
.Y(n_4817)
);

AND2x2_ASAP7_75t_L g4818 ( 
.A(n_4721),
.B(n_4595),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_4761),
.Y(n_4819)
);

AND2x4_ASAP7_75t_L g4820 ( 
.A(n_4746),
.B(n_4674),
.Y(n_4820)
);

AND2x4_ASAP7_75t_L g4821 ( 
.A(n_4721),
.B(n_4724),
.Y(n_4821)
);

INVx1_ASAP7_75t_L g4822 ( 
.A(n_4757),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4704),
.Y(n_4823)
);

AND2x2_ASAP7_75t_L g4824 ( 
.A(n_4736),
.B(n_4627),
.Y(n_4824)
);

OAI221xp5_ASAP7_75t_L g4825 ( 
.A1(n_4803),
.A2(n_4712),
.B1(n_4717),
.B2(n_4701),
.C(n_4766),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_4803),
.B(n_4766),
.Y(n_4826)
);

AND2x4_ASAP7_75t_L g4827 ( 
.A(n_4821),
.B(n_4817),
.Y(n_4827)
);

INVx1_ASAP7_75t_L g4828 ( 
.A(n_4770),
.Y(n_4828)
);

OR2x2_ASAP7_75t_L g4829 ( 
.A(n_4793),
.B(n_4722),
.Y(n_4829)
);

INVx1_ASAP7_75t_L g4830 ( 
.A(n_4768),
.Y(n_4830)
);

AND2x4_ASAP7_75t_L g4831 ( 
.A(n_4821),
.B(n_4748),
.Y(n_4831)
);

AND2x4_ASAP7_75t_L g4832 ( 
.A(n_4821),
.B(n_4748),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4793),
.B(n_4725),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4781),
.B(n_4727),
.Y(n_4834)
);

AND2x2_ASAP7_75t_L g4835 ( 
.A(n_4776),
.B(n_4707),
.Y(n_4835)
);

AND2x2_ASAP7_75t_L g4836 ( 
.A(n_4782),
.B(n_4707),
.Y(n_4836)
);

OR2x2_ASAP7_75t_L g4837 ( 
.A(n_4795),
.B(n_4767),
.Y(n_4837)
);

AND2x2_ASAP7_75t_L g4838 ( 
.A(n_4779),
.B(n_4737),
.Y(n_4838)
);

OR2x2_ASAP7_75t_L g4839 ( 
.A(n_4797),
.B(n_4667),
.Y(n_4839)
);

INVx1_ASAP7_75t_L g4840 ( 
.A(n_4768),
.Y(n_4840)
);

INVx1_ASAP7_75t_L g4841 ( 
.A(n_4781),
.Y(n_4841)
);

AND2x2_ASAP7_75t_L g4842 ( 
.A(n_4777),
.B(n_4760),
.Y(n_4842)
);

OR2x2_ASAP7_75t_L g4843 ( 
.A(n_4786),
.B(n_4815),
.Y(n_4843)
);

AND2x2_ASAP7_75t_L g4844 ( 
.A(n_4800),
.B(n_4764),
.Y(n_4844)
);

INVx2_ASAP7_75t_SL g4845 ( 
.A(n_4817),
.Y(n_4845)
);

INVx3_ASAP7_75t_L g4846 ( 
.A(n_4802),
.Y(n_4846)
);

INVx1_ASAP7_75t_L g4847 ( 
.A(n_4808),
.Y(n_4847)
);

NAND2xp5_ASAP7_75t_L g4848 ( 
.A(n_4778),
.B(n_4731),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4804),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4787),
.B(n_4818),
.Y(n_4850)
);

INVx2_ASAP7_75t_L g4851 ( 
.A(n_4802),
.Y(n_4851)
);

OR2x2_ASAP7_75t_L g4852 ( 
.A(n_4806),
.B(n_4667),
.Y(n_4852)
);

OR2x2_ASAP7_75t_L g4853 ( 
.A(n_4816),
.B(n_4740),
.Y(n_4853)
);

INVx2_ASAP7_75t_L g4854 ( 
.A(n_4807),
.Y(n_4854)
);

NAND2xp5_ASAP7_75t_L g4855 ( 
.A(n_4778),
.B(n_4743),
.Y(n_4855)
);

AND2x2_ASAP7_75t_L g4856 ( 
.A(n_4801),
.B(n_4755),
.Y(n_4856)
);

OR2x2_ASAP7_75t_L g4857 ( 
.A(n_4813),
.B(n_4788),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4804),
.Y(n_4858)
);

HB1xp67_ASAP7_75t_L g4859 ( 
.A(n_4774),
.Y(n_4859)
);

AND2x2_ASAP7_75t_L g4860 ( 
.A(n_4817),
.B(n_4620),
.Y(n_4860)
);

AND2x2_ASAP7_75t_L g4861 ( 
.A(n_4811),
.B(n_4626),
.Y(n_4861)
);

BUFx3_ASAP7_75t_L g4862 ( 
.A(n_4792),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4819),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4819),
.Y(n_4864)
);

AND2x2_ASAP7_75t_L g4865 ( 
.A(n_4824),
.B(n_4744),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4773),
.Y(n_4866)
);

NAND2xp5_ASAP7_75t_L g4867 ( 
.A(n_4774),
.B(n_4710),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4794),
.Y(n_4868)
);

AND2x2_ASAP7_75t_L g4869 ( 
.A(n_4824),
.B(n_4744),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4794),
.Y(n_4870)
);

OR2x2_ASAP7_75t_L g4871 ( 
.A(n_4785),
.B(n_4753),
.Y(n_4871)
);

OR2x2_ASAP7_75t_L g4872 ( 
.A(n_4785),
.B(n_4683),
.Y(n_4872)
);

OAI21xp5_ASAP7_75t_L g4873 ( 
.A1(n_4789),
.A2(n_4783),
.B(n_4799),
.Y(n_4873)
);

NAND2xp5_ASAP7_75t_L g4874 ( 
.A(n_4789),
.B(n_4716),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4792),
.B(n_4734),
.Y(n_4875)
);

AND2x2_ASAP7_75t_L g4876 ( 
.A(n_4792),
.B(n_4734),
.Y(n_4876)
);

NAND2xp5_ASAP7_75t_L g4877 ( 
.A(n_4845),
.B(n_4769),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_4827),
.B(n_4807),
.Y(n_4878)
);

AND2x2_ASAP7_75t_L g4879 ( 
.A(n_4850),
.B(n_4809),
.Y(n_4879)
);

INVx2_ASAP7_75t_L g4880 ( 
.A(n_4862),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4862),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_L g4882 ( 
.A(n_4827),
.B(n_4820),
.Y(n_4882)
);

INVx2_ASAP7_75t_L g4883 ( 
.A(n_4831),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4859),
.Y(n_4884)
);

INVx2_ASAP7_75t_L g4885 ( 
.A(n_4831),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4846),
.B(n_4820),
.Y(n_4886)
);

OR2x2_ASAP7_75t_L g4887 ( 
.A(n_4857),
.B(n_4775),
.Y(n_4887)
);

NOR2xp33_ASAP7_75t_L g4888 ( 
.A(n_4846),
.B(n_4825),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4859),
.Y(n_4889)
);

AND2x4_ASAP7_75t_L g4890 ( 
.A(n_4832),
.B(n_4791),
.Y(n_4890)
);

AND2x2_ASAP7_75t_L g4891 ( 
.A(n_4875),
.B(n_4820),
.Y(n_4891)
);

BUFx3_ASAP7_75t_L g4892 ( 
.A(n_4851),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_SL g4893 ( 
.A(n_4826),
.B(n_4775),
.Y(n_4893)
);

NAND2xp5_ASAP7_75t_L g4894 ( 
.A(n_4832),
.B(n_4791),
.Y(n_4894)
);

INVx1_ASAP7_75t_L g4895 ( 
.A(n_4874),
.Y(n_4895)
);

INVx2_ASAP7_75t_L g4896 ( 
.A(n_4876),
.Y(n_4896)
);

AND2x4_ASAP7_75t_L g4897 ( 
.A(n_4835),
.B(n_4780),
.Y(n_4897)
);

AND2x4_ASAP7_75t_L g4898 ( 
.A(n_4836),
.B(n_4780),
.Y(n_4898)
);

INVx1_ASAP7_75t_L g4899 ( 
.A(n_4874),
.Y(n_4899)
);

NOR3xp33_ASAP7_75t_L g4900 ( 
.A(n_4825),
.B(n_4812),
.C(n_4719),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4842),
.B(n_4758),
.Y(n_4901)
);

OR2x2_ASAP7_75t_L g4902 ( 
.A(n_4843),
.B(n_4790),
.Y(n_4902)
);

AND2x2_ASAP7_75t_L g4903 ( 
.A(n_4865),
.B(n_4771),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4838),
.B(n_4772),
.Y(n_4904)
);

INVx1_ASAP7_75t_L g4905 ( 
.A(n_4830),
.Y(n_4905)
);

OR2x2_ASAP7_75t_L g4906 ( 
.A(n_4852),
.B(n_4840),
.Y(n_4906)
);

HB1xp67_ASAP7_75t_L g4907 ( 
.A(n_4869),
.Y(n_4907)
);

INVx2_ASAP7_75t_L g4908 ( 
.A(n_4826),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_4860),
.B(n_4822),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4844),
.B(n_4758),
.Y(n_4910)
);

AND2x2_ASAP7_75t_L g4911 ( 
.A(n_4856),
.B(n_4823),
.Y(n_4911)
);

AND2x2_ASAP7_75t_L g4912 ( 
.A(n_4861),
.B(n_4639),
.Y(n_4912)
);

HB1xp67_ASAP7_75t_L g4913 ( 
.A(n_4854),
.Y(n_4913)
);

NOR2xp33_ASAP7_75t_L g4914 ( 
.A(n_4828),
.B(n_4784),
.Y(n_4914)
);

AND2x2_ASAP7_75t_L g4915 ( 
.A(n_4847),
.B(n_4641),
.Y(n_4915)
);

AND2x2_ASAP7_75t_L g4916 ( 
.A(n_4891),
.B(n_4837),
.Y(n_4916)
);

INVxp67_ASAP7_75t_SL g4917 ( 
.A(n_4893),
.Y(n_4917)
);

INVx1_ASAP7_75t_SL g4918 ( 
.A(n_4879),
.Y(n_4918)
);

OR2x2_ASAP7_75t_L g4919 ( 
.A(n_4887),
.B(n_4839),
.Y(n_4919)
);

AND2x4_ASAP7_75t_SL g4920 ( 
.A(n_4878),
.B(n_4868),
.Y(n_4920)
);

INVx2_ASAP7_75t_L g4921 ( 
.A(n_4908),
.Y(n_4921)
);

BUFx6f_ASAP7_75t_L g4922 ( 
.A(n_4893),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4907),
.Y(n_4923)
);

INVx1_ASAP7_75t_L g4924 ( 
.A(n_4911),
.Y(n_4924)
);

NAND2xp5_ASAP7_75t_L g4925 ( 
.A(n_4900),
.B(n_4873),
.Y(n_4925)
);

OR2x2_ASAP7_75t_L g4926 ( 
.A(n_4883),
.B(n_4853),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4911),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4891),
.B(n_4870),
.Y(n_4928)
);

HB1xp67_ASAP7_75t_L g4929 ( 
.A(n_4888),
.Y(n_4929)
);

NAND4xp25_ASAP7_75t_L g4930 ( 
.A(n_4888),
.B(n_4873),
.C(n_4833),
.D(n_4872),
.Y(n_4930)
);

BUFx2_ASAP7_75t_L g4931 ( 
.A(n_4890),
.Y(n_4931)
);

BUFx2_ASAP7_75t_L g4932 ( 
.A(n_4890),
.Y(n_4932)
);

INVx2_ASAP7_75t_SL g4933 ( 
.A(n_4878),
.Y(n_4933)
);

INVx2_ASAP7_75t_L g4934 ( 
.A(n_4890),
.Y(n_4934)
);

OR2x2_ASAP7_75t_L g4935 ( 
.A(n_4883),
.B(n_4871),
.Y(n_4935)
);

INVx8_ASAP7_75t_L g4936 ( 
.A(n_4897),
.Y(n_4936)
);

AND2x2_ASAP7_75t_L g4937 ( 
.A(n_4903),
.B(n_4829),
.Y(n_4937)
);

HB1xp67_ASAP7_75t_L g4938 ( 
.A(n_4897),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4903),
.B(n_4841),
.Y(n_4939)
);

NAND2xp5_ASAP7_75t_L g4940 ( 
.A(n_4897),
.B(n_4796),
.Y(n_4940)
);

INVx2_ASAP7_75t_L g4941 ( 
.A(n_4898),
.Y(n_4941)
);

INVx1_ASAP7_75t_L g4942 ( 
.A(n_4909),
.Y(n_4942)
);

INVx2_ASAP7_75t_L g4943 ( 
.A(n_4908),
.Y(n_4943)
);

AND2x2_ASAP7_75t_L g4944 ( 
.A(n_4904),
.B(n_4866),
.Y(n_4944)
);

AND2x2_ASAP7_75t_L g4945 ( 
.A(n_4896),
.B(n_4833),
.Y(n_4945)
);

OR2x2_ASAP7_75t_L g4946 ( 
.A(n_4885),
.B(n_4867),
.Y(n_4946)
);

NOR2xp33_ASAP7_75t_L g4947 ( 
.A(n_4898),
.B(n_4798),
.Y(n_4947)
);

INVx2_ASAP7_75t_L g4948 ( 
.A(n_4898),
.Y(n_4948)
);

AND2x4_ASAP7_75t_L g4949 ( 
.A(n_4933),
.B(n_4892),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4938),
.Y(n_4950)
);

INVxp67_ASAP7_75t_SL g4951 ( 
.A(n_4922),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4936),
.B(n_4896),
.Y(n_4952)
);

AND2x2_ASAP7_75t_L g4953 ( 
.A(n_4937),
.B(n_4892),
.Y(n_4953)
);

OR2x2_ASAP7_75t_L g4954 ( 
.A(n_4919),
.B(n_4885),
.Y(n_4954)
);

AND2x4_ASAP7_75t_L g4955 ( 
.A(n_4941),
.B(n_4880),
.Y(n_4955)
);

HB1xp67_ASAP7_75t_L g4956 ( 
.A(n_4922),
.Y(n_4956)
);

INVx1_ASAP7_75t_L g4957 ( 
.A(n_4938),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4922),
.Y(n_4958)
);

NAND2xp5_ASAP7_75t_L g4959 ( 
.A(n_4936),
.B(n_4880),
.Y(n_4959)
);

O2A1O1Ixp5_ASAP7_75t_L g4960 ( 
.A1(n_4917),
.A2(n_4886),
.B(n_4882),
.C(n_4901),
.Y(n_4960)
);

NOR2x1p5_ASAP7_75t_L g4961 ( 
.A(n_4926),
.B(n_4910),
.Y(n_4961)
);

AND2x4_ASAP7_75t_L g4962 ( 
.A(n_4934),
.B(n_4948),
.Y(n_4962)
);

INVx2_ASAP7_75t_L g4963 ( 
.A(n_4922),
.Y(n_4963)
);

AOI22xp5_ASAP7_75t_L g4964 ( 
.A1(n_4917),
.A2(n_4805),
.B1(n_4814),
.B2(n_4810),
.Y(n_4964)
);

AOI211xp5_ASAP7_75t_L g4965 ( 
.A1(n_4930),
.A2(n_4914),
.B(n_4895),
.C(n_4899),
.Y(n_4965)
);

INVx1_ASAP7_75t_L g4966 ( 
.A(n_4931),
.Y(n_4966)
);

INVxp67_ASAP7_75t_SL g4967 ( 
.A(n_4929),
.Y(n_4967)
);

INVx1_ASAP7_75t_SL g4968 ( 
.A(n_4916),
.Y(n_4968)
);

INVx1_ASAP7_75t_L g4969 ( 
.A(n_4932),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4948),
.Y(n_4970)
);

NAND2xp5_ASAP7_75t_L g4971 ( 
.A(n_4936),
.B(n_4909),
.Y(n_4971)
);

OR2x2_ASAP7_75t_L g4972 ( 
.A(n_4918),
.B(n_4906),
.Y(n_4972)
);

INVx2_ASAP7_75t_L g4973 ( 
.A(n_4921),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4953),
.B(n_4939),
.Y(n_4974)
);

O2A1O1Ixp33_ASAP7_75t_L g4975 ( 
.A1(n_4967),
.A2(n_4925),
.B(n_4929),
.C(n_4884),
.Y(n_4975)
);

INVx1_ASAP7_75t_L g4976 ( 
.A(n_4956),
.Y(n_4976)
);

OR2x2_ASAP7_75t_L g4977 ( 
.A(n_4968),
.B(n_4935),
.Y(n_4977)
);

NOR2xp33_ASAP7_75t_R g4978 ( 
.A(n_4972),
.B(n_4923),
.Y(n_4978)
);

INVx2_ASAP7_75t_L g4979 ( 
.A(n_4949),
.Y(n_4979)
);

NOR2xp33_ASAP7_75t_L g4980 ( 
.A(n_4954),
.B(n_4902),
.Y(n_4980)
);

INVx1_ASAP7_75t_SL g4981 ( 
.A(n_4949),
.Y(n_4981)
);

OR2x2_ASAP7_75t_L g4982 ( 
.A(n_4971),
.B(n_4946),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4961),
.B(n_4928),
.Y(n_4983)
);

NOR3xp33_ASAP7_75t_L g4984 ( 
.A(n_4960),
.B(n_4925),
.C(n_4959),
.Y(n_4984)
);

INVx2_ASAP7_75t_SL g4985 ( 
.A(n_4955),
.Y(n_4985)
);

AOI22xp33_ASAP7_75t_L g4986 ( 
.A1(n_4973),
.A2(n_4921),
.B1(n_4943),
.B2(n_4696),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4955),
.B(n_4945),
.Y(n_4987)
);

INVx1_ASAP7_75t_SL g4988 ( 
.A(n_4962),
.Y(n_4988)
);

AND2x2_ASAP7_75t_L g4989 ( 
.A(n_4966),
.B(n_4944),
.Y(n_4989)
);

OR2x2_ASAP7_75t_L g4990 ( 
.A(n_4952),
.B(n_4942),
.Y(n_4990)
);

HB1xp67_ASAP7_75t_L g4991 ( 
.A(n_4962),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4969),
.B(n_4913),
.Y(n_4992)
);

NOR2xp33_ASAP7_75t_SL g4993 ( 
.A(n_4951),
.B(n_4881),
.Y(n_4993)
);

INVx2_ASAP7_75t_L g4994 ( 
.A(n_4963),
.Y(n_4994)
);

INVx1_ASAP7_75t_L g4995 ( 
.A(n_4991),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4987),
.Y(n_4996)
);

INVx2_ASAP7_75t_L g4997 ( 
.A(n_4977),
.Y(n_4997)
);

AND2x2_ASAP7_75t_L g4998 ( 
.A(n_4983),
.B(n_4924),
.Y(n_4998)
);

AND2x2_ASAP7_75t_L g4999 ( 
.A(n_4992),
.B(n_4927),
.Y(n_4999)
);

NAND2xp5_ASAP7_75t_L g5000 ( 
.A(n_4988),
.B(n_4947),
.Y(n_5000)
);

AND2x2_ASAP7_75t_L g5001 ( 
.A(n_4980),
.B(n_4920),
.Y(n_5001)
);

AND2x2_ASAP7_75t_L g5002 ( 
.A(n_4981),
.B(n_4920),
.Y(n_5002)
);

CKINVDCx16_ASAP7_75t_R g5003 ( 
.A(n_4978),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4988),
.B(n_4947),
.Y(n_5004)
);

CKINVDCx16_ASAP7_75t_R g5005 ( 
.A(n_4989),
.Y(n_5005)
);

INVx2_ASAP7_75t_L g5006 ( 
.A(n_4985),
.Y(n_5006)
);

AND2x2_ASAP7_75t_L g5007 ( 
.A(n_4979),
.B(n_4912),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4974),
.Y(n_5008)
);

INVx1_ASAP7_75t_SL g5009 ( 
.A(n_4982),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4975),
.Y(n_5010)
);

INVx4_ASAP7_75t_L g5011 ( 
.A(n_4994),
.Y(n_5011)
);

NOR2xp33_ASAP7_75t_L g5012 ( 
.A(n_5005),
.B(n_4993),
.Y(n_5012)
);

OAI21xp5_ASAP7_75t_L g5013 ( 
.A1(n_5000),
.A2(n_4984),
.B(n_4940),
.Y(n_5013)
);

INVx1_ASAP7_75t_L g5014 ( 
.A(n_5004),
.Y(n_5014)
);

INVx2_ASAP7_75t_L g5015 ( 
.A(n_5001),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_5007),
.Y(n_5016)
);

INVx1_ASAP7_75t_SL g5017 ( 
.A(n_5009),
.Y(n_5017)
);

OAI221xp5_ASAP7_75t_L g5018 ( 
.A1(n_4995),
.A2(n_4940),
.B1(n_4964),
.B2(n_4950),
.C(n_4957),
.Y(n_5018)
);

INVx2_ASAP7_75t_L g5019 ( 
.A(n_5011),
.Y(n_5019)
);

NOR2xp33_ASAP7_75t_L g5020 ( 
.A(n_5003),
.B(n_4993),
.Y(n_5020)
);

OAI21xp5_ASAP7_75t_L g5021 ( 
.A1(n_4995),
.A2(n_4914),
.B(n_4877),
.Y(n_5021)
);

CKINVDCx20_ASAP7_75t_R g5022 ( 
.A(n_5002),
.Y(n_5022)
);

AOI22xp5_ASAP7_75t_L g5023 ( 
.A1(n_5010),
.A2(n_4970),
.B1(n_4943),
.B2(n_4997),
.Y(n_5023)
);

INVx1_ASAP7_75t_SL g5024 ( 
.A(n_4999),
.Y(n_5024)
);

AND2x2_ASAP7_75t_L g5025 ( 
.A(n_4998),
.B(n_4912),
.Y(n_5025)
);

OAI22xp5_ASAP7_75t_L g5026 ( 
.A1(n_4996),
.A2(n_4965),
.B1(n_4990),
.B2(n_4958),
.Y(n_5026)
);

INVx2_ASAP7_75t_L g5027 ( 
.A(n_5011),
.Y(n_5027)
);

INVx1_ASAP7_75t_SL g5028 ( 
.A(n_5006),
.Y(n_5028)
);

OAI21xp5_ASAP7_75t_SL g5029 ( 
.A1(n_4996),
.A2(n_4976),
.B(n_4894),
.Y(n_5029)
);

INVx1_ASAP7_75t_L g5030 ( 
.A(n_5008),
.Y(n_5030)
);

OAI21xp5_ASAP7_75t_SL g5031 ( 
.A1(n_5009),
.A2(n_4889),
.B(n_4905),
.Y(n_5031)
);

AOI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_5012),
.A2(n_4834),
.B(n_4867),
.Y(n_5032)
);

AOI22xp5_ASAP7_75t_L g5033 ( 
.A1(n_5020),
.A2(n_4986),
.B1(n_4849),
.B2(n_4863),
.Y(n_5033)
);

AOI221xp5_ASAP7_75t_L g5034 ( 
.A1(n_5013),
.A2(n_4864),
.B1(n_4858),
.B2(n_4834),
.C(n_4855),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_5024),
.B(n_4848),
.Y(n_5035)
);

OAI22xp5_ASAP7_75t_L g5036 ( 
.A1(n_5017),
.A2(n_4855),
.B1(n_4848),
.B2(n_4915),
.Y(n_5036)
);

AOI22xp33_ASAP7_75t_L g5037 ( 
.A1(n_5014),
.A2(n_4758),
.B1(n_4655),
.B2(n_4657),
.Y(n_5037)
);

AOI32xp33_ASAP7_75t_L g5038 ( 
.A1(n_5025),
.A2(n_4915),
.A3(n_4609),
.B1(n_4619),
.B2(n_4602),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_L g5039 ( 
.A(n_5028),
.B(n_4693),
.Y(n_5039)
);

NAND2xp5_ASAP7_75t_L g5040 ( 
.A(n_5023),
.B(n_4664),
.Y(n_5040)
);

AOI22xp33_ASAP7_75t_SL g5041 ( 
.A1(n_5016),
.A2(n_4745),
.B1(n_4604),
.B2(n_4668),
.Y(n_5041)
);

AND2x2_ASAP7_75t_L g5042 ( 
.A(n_5015),
.B(n_5021),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_5023),
.B(n_4668),
.Y(n_5043)
);

OAI322xp33_ASAP7_75t_L g5044 ( 
.A1(n_5018),
.A2(n_4656),
.A3(n_4611),
.B1(n_4600),
.B2(n_4601),
.C1(n_4615),
.C2(n_4621),
.Y(n_5044)
);

INVxp67_ASAP7_75t_SL g5045 ( 
.A(n_5022),
.Y(n_5045)
);

INVx1_ASAP7_75t_SL g5046 ( 
.A(n_5019),
.Y(n_5046)
);

AND2x2_ASAP7_75t_L g5047 ( 
.A(n_5030),
.B(n_4644),
.Y(n_5047)
);

OAI221xp5_ASAP7_75t_L g5048 ( 
.A1(n_5031),
.A2(n_4681),
.B1(n_4608),
.B2(n_4671),
.C(n_4684),
.Y(n_5048)
);

AOI22xp5_ASAP7_75t_L g5049 ( 
.A1(n_5029),
.A2(n_4608),
.B1(n_4679),
.B2(n_4671),
.Y(n_5049)
);

INVx1_ASAP7_75t_L g5050 ( 
.A(n_5027),
.Y(n_5050)
);

NAND2xp5_ASAP7_75t_L g5051 ( 
.A(n_5026),
.B(n_4665),
.Y(n_5051)
);

NAND2xp5_ASAP7_75t_L g5052 ( 
.A(n_5025),
.B(n_4749),
.Y(n_5052)
);

OAI32xp33_ASAP7_75t_L g5053 ( 
.A1(n_5017),
.A2(n_4684),
.A3(n_4624),
.B1(n_4687),
.B2(n_4689),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_5025),
.B(n_4749),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_5025),
.Y(n_5055)
);

NAND2xp5_ASAP7_75t_L g5056 ( 
.A(n_5025),
.B(n_4678),
.Y(n_5056)
);

INVx2_ASAP7_75t_L g5057 ( 
.A(n_5022),
.Y(n_5057)
);

AND2x4_ASAP7_75t_L g5058 ( 
.A(n_5045),
.B(n_5057),
.Y(n_5058)
);

NOR2xp33_ASAP7_75t_L g5059 ( 
.A(n_5043),
.B(n_4652),
.Y(n_5059)
);

NAND2xp5_ASAP7_75t_L g5060 ( 
.A(n_5041),
.B(n_4697),
.Y(n_5060)
);

AOI22xp33_ASAP7_75t_L g5061 ( 
.A1(n_5040),
.A2(n_4694),
.B1(n_4698),
.B2(n_4687),
.Y(n_5061)
);

INVx1_ASAP7_75t_L g5062 ( 
.A(n_5042),
.Y(n_5062)
);

OR2x2_ASAP7_75t_L g5063 ( 
.A(n_5039),
.B(n_4624),
.Y(n_5063)
);

INVx1_ASAP7_75t_L g5064 ( 
.A(n_5052),
.Y(n_5064)
);

NOR2xp33_ASAP7_75t_L g5065 ( 
.A(n_5049),
.B(n_4698),
.Y(n_5065)
);

INVx1_ASAP7_75t_L g5066 ( 
.A(n_5054),
.Y(n_5066)
);

NAND2xp5_ASAP7_75t_L g5067 ( 
.A(n_5035),
.B(n_4683),
.Y(n_5067)
);

CKINVDCx20_ASAP7_75t_R g5068 ( 
.A(n_5036),
.Y(n_5068)
);

NAND2xp33_ASAP7_75t_R g5069 ( 
.A(n_5055),
.B(n_482),
.Y(n_5069)
);

INVx1_ASAP7_75t_L g5070 ( 
.A(n_5056),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_5032),
.B(n_5034),
.Y(n_5071)
);

BUFx2_ASAP7_75t_L g5072 ( 
.A(n_5047),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_5051),
.Y(n_5073)
);

NOR2xp33_ASAP7_75t_SL g5074 ( 
.A(n_5046),
.B(n_4562),
.Y(n_5074)
);

INVx2_ASAP7_75t_L g5075 ( 
.A(n_5050),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_5033),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_5037),
.B(n_5038),
.Y(n_5077)
);

NAND2x1p5_ASAP7_75t_L g5078 ( 
.A(n_5053),
.B(n_4347),
.Y(n_5078)
);

AND2x2_ASAP7_75t_L g5079 ( 
.A(n_5044),
.B(n_5048),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_5045),
.B(n_4561),
.Y(n_5080)
);

AND2x2_ASAP7_75t_L g5081 ( 
.A(n_5045),
.B(n_4347),
.Y(n_5081)
);

AND2x2_ASAP7_75t_L g5082 ( 
.A(n_5045),
.B(n_4349),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_5045),
.B(n_4577),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_5045),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_5045),
.B(n_4349),
.Y(n_5085)
);

NAND2xp5_ASAP7_75t_SL g5086 ( 
.A(n_5057),
.B(n_4514),
.Y(n_5086)
);

XOR2xp5_ASAP7_75t_L g5087 ( 
.A(n_5058),
.B(n_4488),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_5072),
.Y(n_5088)
);

NAND3xp33_ASAP7_75t_L g5089 ( 
.A(n_5062),
.B(n_4525),
.C(n_4500),
.Y(n_5089)
);

INVx1_ASAP7_75t_L g5090 ( 
.A(n_5058),
.Y(n_5090)
);

INVx4_ASAP7_75t_L g5091 ( 
.A(n_5075),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_5063),
.Y(n_5092)
);

INVxp67_ASAP7_75t_SL g5093 ( 
.A(n_5069),
.Y(n_5093)
);

NAND2xp5_ASAP7_75t_L g5094 ( 
.A(n_5064),
.B(n_4497),
.Y(n_5094)
);

INVx1_ASAP7_75t_SL g5095 ( 
.A(n_5081),
.Y(n_5095)
);

INVx1_ASAP7_75t_L g5096 ( 
.A(n_5082),
.Y(n_5096)
);

INVx1_ASAP7_75t_L g5097 ( 
.A(n_5085),
.Y(n_5097)
);

INVx1_ASAP7_75t_L g5098 ( 
.A(n_5084),
.Y(n_5098)
);

OR2x2_ASAP7_75t_L g5099 ( 
.A(n_5060),
.B(n_4365),
.Y(n_5099)
);

XOR2x2_ASAP7_75t_L g5100 ( 
.A(n_5066),
.B(n_5080),
.Y(n_5100)
);

NAND2xp5_ASAP7_75t_L g5101 ( 
.A(n_5061),
.B(n_4550),
.Y(n_5101)
);

INVx1_ASAP7_75t_L g5102 ( 
.A(n_5078),
.Y(n_5102)
);

INVx1_ASAP7_75t_L g5103 ( 
.A(n_5067),
.Y(n_5103)
);

INVx1_ASAP7_75t_SL g5104 ( 
.A(n_5068),
.Y(n_5104)
);

INVx1_ASAP7_75t_L g5105 ( 
.A(n_5083),
.Y(n_5105)
);

A2O1A1Ixp33_ASAP7_75t_L g5106 ( 
.A1(n_5065),
.A2(n_4580),
.B(n_4579),
.C(n_4574),
.Y(n_5106)
);

INVx1_ASAP7_75t_L g5107 ( 
.A(n_5071),
.Y(n_5107)
);

INVx1_ASAP7_75t_L g5108 ( 
.A(n_5074),
.Y(n_5108)
);

INVx2_ASAP7_75t_L g5109 ( 
.A(n_5070),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_5074),
.B(n_4522),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_5076),
.B(n_4524),
.Y(n_5111)
);

HB1xp67_ASAP7_75t_L g5112 ( 
.A(n_5090),
.Y(n_5112)
);

AOI21x1_ASAP7_75t_L g5113 ( 
.A1(n_5088),
.A2(n_5073),
.B(n_5077),
.Y(n_5113)
);

OA22x2_ASAP7_75t_L g5114 ( 
.A1(n_5104),
.A2(n_5086),
.B1(n_5079),
.B2(n_5059),
.Y(n_5114)
);

OAI21xp5_ASAP7_75t_L g5115 ( 
.A1(n_5093),
.A2(n_4532),
.B(n_4529),
.Y(n_5115)
);

AOI21xp5_ASAP7_75t_L g5116 ( 
.A1(n_5107),
.A2(n_4366),
.B(n_4365),
.Y(n_5116)
);

NAND3xp33_ASAP7_75t_L g5117 ( 
.A(n_5091),
.B(n_4542),
.C(n_4534),
.Y(n_5117)
);

AOI21xp5_ASAP7_75t_L g5118 ( 
.A1(n_5098),
.A2(n_4366),
.B(n_4563),
.Y(n_5118)
);

NOR2xp33_ASAP7_75t_L g5119 ( 
.A(n_5091),
.B(n_4441),
.Y(n_5119)
);

INVx1_ASAP7_75t_SL g5120 ( 
.A(n_5095),
.Y(n_5120)
);

AO21x1_ASAP7_75t_L g5121 ( 
.A1(n_5092),
.A2(n_482),
.B(n_483),
.Y(n_5121)
);

INVx2_ASAP7_75t_L g5122 ( 
.A(n_5100),
.Y(n_5122)
);

INVx1_ASAP7_75t_L g5123 ( 
.A(n_5087),
.Y(n_5123)
);

NOR2x1_ASAP7_75t_L g5124 ( 
.A(n_5109),
.B(n_483),
.Y(n_5124)
);

INVx1_ASAP7_75t_SL g5125 ( 
.A(n_5108),
.Y(n_5125)
);

OAI222xp33_ASAP7_75t_L g5126 ( 
.A1(n_5102),
.A2(n_4417),
.B1(n_4442),
.B2(n_4441),
.C1(n_488),
.C2(n_489),
.Y(n_5126)
);

NAND2xp5_ASAP7_75t_L g5127 ( 
.A(n_5096),
.B(n_4442),
.Y(n_5127)
);

AOI22xp5_ASAP7_75t_L g5128 ( 
.A1(n_5097),
.A2(n_484),
.B1(n_485),
.B2(n_486),
.Y(n_5128)
);

OAI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_5105),
.A2(n_484),
.B(n_485),
.Y(n_5129)
);

AOI22xp33_ASAP7_75t_L g5130 ( 
.A1(n_5122),
.A2(n_5103),
.B1(n_5110),
.B2(n_5099),
.Y(n_5130)
);

OAI211xp5_ASAP7_75t_L g5131 ( 
.A1(n_5120),
.A2(n_5094),
.B(n_5111),
.C(n_5101),
.Y(n_5131)
);

AOI22xp33_ASAP7_75t_L g5132 ( 
.A1(n_5112),
.A2(n_5089),
.B1(n_5106),
.B2(n_490),
.Y(n_5132)
);

AOI22xp5_ASAP7_75t_L g5133 ( 
.A1(n_5125),
.A2(n_486),
.B1(n_489),
.B2(n_492),
.Y(n_5133)
);

AOI22xp5_ASAP7_75t_L g5134 ( 
.A1(n_5114),
.A2(n_492),
.B1(n_494),
.B2(n_495),
.Y(n_5134)
);

NAND2xp33_ASAP7_75t_R g5135 ( 
.A(n_5123),
.B(n_494),
.Y(n_5135)
);

INVx1_ASAP7_75t_L g5136 ( 
.A(n_5121),
.Y(n_5136)
);

AOI22xp5_ASAP7_75t_L g5137 ( 
.A1(n_5119),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_5137)
);

OAI21xp33_ASAP7_75t_L g5138 ( 
.A1(n_5113),
.A2(n_496),
.B(n_497),
.Y(n_5138)
);

AOI221x1_ASAP7_75t_L g5139 ( 
.A1(n_5129),
.A2(n_5127),
.B1(n_5116),
.B2(n_5118),
.C(n_5115),
.Y(n_5139)
);

INVx2_ASAP7_75t_L g5140 ( 
.A(n_5124),
.Y(n_5140)
);

INVx1_ASAP7_75t_L g5141 ( 
.A(n_5128),
.Y(n_5141)
);

INVx2_ASAP7_75t_L g5142 ( 
.A(n_5117),
.Y(n_5142)
);

AOI221xp5_ASAP7_75t_L g5143 ( 
.A1(n_5126),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.C(n_501),
.Y(n_5143)
);

AOI22xp5_ASAP7_75t_L g5144 ( 
.A1(n_5120),
.A2(n_498),
.B1(n_499),
.B2(n_500),
.Y(n_5144)
);

O2A1O1Ixp33_ASAP7_75t_L g5145 ( 
.A1(n_5122),
.A2(n_501),
.B(n_502),
.C(n_503),
.Y(n_5145)
);

NAND4xp25_ASAP7_75t_L g5146 ( 
.A(n_5130),
.B(n_502),
.C(n_503),
.D(n_504),
.Y(n_5146)
);

AOI211xp5_ASAP7_75t_L g5147 ( 
.A1(n_5131),
.A2(n_5138),
.B(n_5145),
.C(n_5136),
.Y(n_5147)
);

AOI221xp5_ASAP7_75t_L g5148 ( 
.A1(n_5142),
.A2(n_504),
.B1(n_505),
.B2(n_506),
.C(n_507),
.Y(n_5148)
);

OAI211xp5_ASAP7_75t_L g5149 ( 
.A1(n_5134),
.A2(n_5132),
.B(n_5139),
.C(n_5143),
.Y(n_5149)
);

NAND3xp33_ASAP7_75t_L g5150 ( 
.A(n_5135),
.B(n_505),
.C(n_506),
.Y(n_5150)
);

INVx2_ASAP7_75t_SL g5151 ( 
.A(n_5140),
.Y(n_5151)
);

AOI221xp5_ASAP7_75t_L g5152 ( 
.A1(n_5141),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.C(n_510),
.Y(n_5152)
);

OAI22xp5_ASAP7_75t_L g5153 ( 
.A1(n_5144),
.A2(n_508),
.B1(n_509),
.B2(n_511),
.Y(n_5153)
);

OAI221xp5_ASAP7_75t_L g5154 ( 
.A1(n_5133),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.C(n_514),
.Y(n_5154)
);

AOI321xp33_ASAP7_75t_L g5155 ( 
.A1(n_5137),
.A2(n_512),
.A3(n_514),
.B1(n_515),
.B2(n_516),
.C(n_517),
.Y(n_5155)
);

AOI211xp5_ASAP7_75t_L g5156 ( 
.A1(n_5131),
.A2(n_515),
.B(n_516),
.C(n_517),
.Y(n_5156)
);

AOI31xp33_ASAP7_75t_L g5157 ( 
.A1(n_5130),
.A2(n_520),
.A3(n_521),
.B(n_522),
.Y(n_5157)
);

NAND4xp25_ASAP7_75t_L g5158 ( 
.A(n_5130),
.B(n_520),
.C(n_522),
.D(n_523),
.Y(n_5158)
);

AOI221xp5_ASAP7_75t_L g5159 ( 
.A1(n_5136),
.A2(n_523),
.B1(n_524),
.B2(n_526),
.C(n_527),
.Y(n_5159)
);

NOR3xp33_ASAP7_75t_L g5160 ( 
.A(n_5131),
.B(n_524),
.C(n_526),
.Y(n_5160)
);

NOR2xp33_ASAP7_75t_R g5161 ( 
.A(n_5135),
.B(n_529),
.Y(n_5161)
);

OAI21xp5_ASAP7_75t_L g5162 ( 
.A1(n_5136),
.A2(n_529),
.B(n_530),
.Y(n_5162)
);

OAI21xp33_ASAP7_75t_L g5163 ( 
.A1(n_5130),
.A2(n_531),
.B(n_532),
.Y(n_5163)
);

NAND4xp25_ASAP7_75t_L g5164 ( 
.A(n_5130),
.B(n_534),
.C(n_535),
.D(n_536),
.Y(n_5164)
);

NOR2x1_ASAP7_75t_L g5165 ( 
.A(n_5150),
.B(n_534),
.Y(n_5165)
);

NOR3xp33_ASAP7_75t_L g5166 ( 
.A(n_5151),
.B(n_536),
.C(n_538),
.Y(n_5166)
);

NOR3xp33_ASAP7_75t_L g5167 ( 
.A(n_5149),
.B(n_538),
.C(n_539),
.Y(n_5167)
);

NOR2x1_ASAP7_75t_L g5168 ( 
.A(n_5146),
.B(n_539),
.Y(n_5168)
);

OAI222xp33_ASAP7_75t_L g5169 ( 
.A1(n_5154),
.A2(n_540),
.B1(n_542),
.B2(n_543),
.C1(n_544),
.C2(n_545),
.Y(n_5169)
);

NAND4xp75_ASAP7_75t_L g5170 ( 
.A(n_5162),
.B(n_542),
.C(n_544),
.D(n_545),
.Y(n_5170)
);

OAI21xp5_ASAP7_75t_L g5171 ( 
.A1(n_5160),
.A2(n_546),
.B(n_547),
.Y(n_5171)
);

NOR3xp33_ASAP7_75t_L g5172 ( 
.A(n_5147),
.B(n_546),
.C(n_548),
.Y(n_5172)
);

NAND4xp75_ASAP7_75t_L g5173 ( 
.A(n_5148),
.B(n_550),
.C(n_551),
.D(n_552),
.Y(n_5173)
);

NAND3xp33_ASAP7_75t_SL g5174 ( 
.A(n_5161),
.B(n_551),
.C(n_552),
.Y(n_5174)
);

NOR3xp33_ASAP7_75t_L g5175 ( 
.A(n_5157),
.B(n_553),
.C(n_554),
.Y(n_5175)
);

NOR2x1_ASAP7_75t_L g5176 ( 
.A(n_5158),
.B(n_554),
.Y(n_5176)
);

AOI22xp5_ASAP7_75t_L g5177 ( 
.A1(n_5164),
.A2(n_555),
.B1(n_556),
.B2(n_557),
.Y(n_5177)
);

NOR3xp33_ASAP7_75t_L g5178 ( 
.A(n_5163),
.B(n_556),
.C(n_558),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_5155),
.Y(n_5179)
);

NOR2xp67_ASAP7_75t_L g5180 ( 
.A(n_5153),
.B(n_558),
.Y(n_5180)
);

HB1xp67_ASAP7_75t_L g5181 ( 
.A(n_5156),
.Y(n_5181)
);

NOR2x1_ASAP7_75t_L g5182 ( 
.A(n_5159),
.B(n_559),
.Y(n_5182)
);

NAND4xp25_ASAP7_75t_SL g5183 ( 
.A(n_5172),
.B(n_5152),
.C(n_561),
.D(n_562),
.Y(n_5183)
);

NAND3xp33_ASAP7_75t_L g5184 ( 
.A(n_5179),
.B(n_560),
.C(n_561),
.Y(n_5184)
);

OR2x2_ASAP7_75t_L g5185 ( 
.A(n_5174),
.B(n_560),
.Y(n_5185)
);

NAND3xp33_ASAP7_75t_SL g5186 ( 
.A(n_5167),
.B(n_563),
.C(n_564),
.Y(n_5186)
);

OAI221xp5_ASAP7_75t_L g5187 ( 
.A1(n_5166),
.A2(n_563),
.B1(n_564),
.B2(n_566),
.C(n_567),
.Y(n_5187)
);

AO22x1_ASAP7_75t_L g5188 ( 
.A1(n_5165),
.A2(n_566),
.B1(n_567),
.B2(n_568),
.Y(n_5188)
);

NAND4xp75_ASAP7_75t_L g5189 ( 
.A(n_5168),
.B(n_568),
.C(n_569),
.D(n_570),
.Y(n_5189)
);

AOI221xp5_ASAP7_75t_SL g5190 ( 
.A1(n_5171),
.A2(n_569),
.B1(n_570),
.B2(n_571),
.C(n_572),
.Y(n_5190)
);

NAND4xp25_ASAP7_75t_SL g5191 ( 
.A(n_5177),
.B(n_571),
.C(n_572),
.D(n_574),
.Y(n_5191)
);

NOR4xp25_ASAP7_75t_L g5192 ( 
.A(n_5169),
.B(n_574),
.C(n_575),
.D(n_576),
.Y(n_5192)
);

NOR3xp33_ASAP7_75t_L g5193 ( 
.A(n_5181),
.B(n_575),
.C(n_576),
.Y(n_5193)
);

XNOR2xp5_ASAP7_75t_L g5194 ( 
.A(n_5176),
.B(n_577),
.Y(n_5194)
);

INVx3_ASAP7_75t_L g5195 ( 
.A(n_5185),
.Y(n_5195)
);

NOR2x1_ASAP7_75t_L g5196 ( 
.A(n_5189),
.B(n_5170),
.Y(n_5196)
);

AND4x1_ASAP7_75t_L g5197 ( 
.A(n_5192),
.B(n_5175),
.C(n_5182),
.D(n_5178),
.Y(n_5197)
);

OR2x2_ASAP7_75t_L g5198 ( 
.A(n_5188),
.B(n_5180),
.Y(n_5198)
);

NOR2xp33_ASAP7_75t_L g5199 ( 
.A(n_5194),
.B(n_5173),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_SL g5200 ( 
.A(n_5193),
.B(n_577),
.Y(n_5200)
);

AOI211xp5_ASAP7_75t_L g5201 ( 
.A1(n_5199),
.A2(n_5184),
.B(n_5186),
.C(n_5183),
.Y(n_5201)
);

NOR3xp33_ASAP7_75t_SL g5202 ( 
.A(n_5200),
.B(n_5191),
.C(n_5187),
.Y(n_5202)
);

INVx1_ASAP7_75t_L g5203 ( 
.A(n_5198),
.Y(n_5203)
);

NAND2xp5_ASAP7_75t_L g5204 ( 
.A(n_5203),
.B(n_5195),
.Y(n_5204)
);

NOR3xp33_ASAP7_75t_L g5205 ( 
.A(n_5201),
.B(n_5196),
.C(n_5190),
.Y(n_5205)
);

OAI22xp5_ASAP7_75t_L g5206 ( 
.A1(n_5204),
.A2(n_5202),
.B1(n_5197),
.B2(n_582),
.Y(n_5206)
);

INVx1_ASAP7_75t_L g5207 ( 
.A(n_5206),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_5207),
.B(n_5205),
.Y(n_5208)
);

NAND3x1_ASAP7_75t_L g5209 ( 
.A(n_5208),
.B(n_579),
.C(n_581),
.Y(n_5209)
);

AOI21xp5_ASAP7_75t_L g5210 ( 
.A1(n_5209),
.A2(n_583),
.B(n_584),
.Y(n_5210)
);

XNOR2x2_ASAP7_75t_L g5211 ( 
.A(n_5210),
.B(n_583),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5211),
.Y(n_5212)
);

AO22x2_ASAP7_75t_L g5213 ( 
.A1(n_5212),
.A2(n_584),
.B1(n_606),
.B2(n_607),
.Y(n_5213)
);

AOI31xp33_ASAP7_75t_L g5214 ( 
.A1(n_5213),
.A2(n_683),
.A3(n_609),
.B(n_610),
.Y(n_5214)
);

OAI22xp5_ASAP7_75t_L g5215 ( 
.A1(n_5214),
.A2(n_608),
.B1(n_613),
.B2(n_617),
.Y(n_5215)
);

OR2x6_ASAP7_75t_L g5216 ( 
.A(n_5215),
.B(n_619),
.Y(n_5216)
);

OA21x2_ASAP7_75t_L g5217 ( 
.A1(n_5216),
.A2(n_620),
.B(n_621),
.Y(n_5217)
);

OAI221xp5_ASAP7_75t_R g5218 ( 
.A1(n_5217),
.A2(n_625),
.B1(n_626),
.B2(n_628),
.C(n_629),
.Y(n_5218)
);

AOI221xp5_ASAP7_75t_L g5219 ( 
.A1(n_5217),
.A2(n_631),
.B1(n_632),
.B2(n_633),
.C(n_634),
.Y(n_5219)
);

AOI22xp5_ASAP7_75t_L g5220 ( 
.A1(n_5219),
.A2(n_636),
.B1(n_642),
.B2(n_644),
.Y(n_5220)
);

AOI211xp5_ASAP7_75t_L g5221 ( 
.A1(n_5220),
.A2(n_5218),
.B(n_652),
.C(n_653),
.Y(n_5221)
);


endmodule