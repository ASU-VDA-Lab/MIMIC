module fake_jpeg_367_n_79 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx11_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_21),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_33),
.Y(n_37)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_23),
.B1(n_30),
.B2(n_28),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_32),
.B1(n_35),
.B2(n_27),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_36),
.C(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_25),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_42),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_26),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_41),
.A2(n_35),
.B(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_45),
.B(n_48),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_32),
.B1(n_27),
.B2(n_11),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_50),
.B1(n_12),
.B2(n_20),
.Y(n_53)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_0),
.Y(n_50)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_8),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_44),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_22),
.B1(n_13),
.B2(n_15),
.Y(n_67)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_47),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_58),
.B1(n_9),
.B2(n_10),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_57),
.B(n_7),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_8),
.Y(n_62)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_57),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_64),
.B(n_59),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_67),
.B1(n_59),
.B2(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_68),
.Y(n_74)
);

OAI21x1_ASAP7_75t_L g75 ( 
.A1(n_74),
.A2(n_62),
.B(n_71),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_63),
.B(n_72),
.Y(n_77)
);

OAI311xp33_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_69),
.A3(n_66),
.B1(n_72),
.C1(n_61),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_19),
.Y(n_79)
);


endmodule