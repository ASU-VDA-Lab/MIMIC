module fake_jpeg_11111_n_573 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_573);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_573;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_2),
.B(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_6),
.B(n_14),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_16),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_54),
.Y(n_110)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_57),
.Y(n_124)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_58),
.Y(n_148)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_59),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_61),
.Y(n_136)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_63),
.B(n_73),
.Y(n_127)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_64),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g167 ( 
.A(n_66),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_67),
.Y(n_119)
);

BUFx24_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g163 ( 
.A(n_69),
.B(n_32),
.Y(n_163)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_31),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_74),
.Y(n_126)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_75),
.Y(n_112)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx6_ASAP7_75t_SL g135 ( 
.A(n_77),
.Y(n_135)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_27),
.Y(n_81)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_81),
.Y(n_165)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_20),
.B(n_0),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_32),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_21),
.Y(n_86)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_86),
.Y(n_140)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_87),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g88 ( 
.A(n_26),
.Y(n_88)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_88),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_89),
.Y(n_113)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_0),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_91),
.B(n_95),
.Y(n_142)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_30),
.Y(n_92)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_26),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_24),
.B(n_52),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_28),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_99),
.Y(n_134)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_28),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_40),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_100),
.B(n_39),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

BUFx12_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_103),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_34),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_51),
.B(n_45),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_108),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_65),
.A2(n_38),
.B1(n_49),
.B2(n_48),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_65),
.B1(n_59),
.B2(n_42),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_118),
.B(n_161),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_57),
.B(n_20),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_128),
.B(n_137),
.Y(n_218)
);

AOI21xp33_ASAP7_75t_L g137 ( 
.A1(n_68),
.A2(n_23),
.B(n_37),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_70),
.B(n_27),
.C(n_51),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_143),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_57),
.B(n_22),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_164),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_104),
.B(n_22),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_29),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_64),
.B(n_23),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_86),
.Y(n_162)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_74),
.B(n_52),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_55),
.Y(n_166)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_58),
.Y(n_168)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_82),
.B(n_37),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_36),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_170),
.Y(n_209)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_107),
.B(n_68),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_172),
.B(n_213),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_174),
.Y(n_268)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_140),
.Y(n_175)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_175),
.Y(n_237)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_176),
.Y(n_238)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_177),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_179),
.B(n_203),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_45),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_182),
.B(n_193),
.Y(n_259)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_112),
.Y(n_183)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_183),
.Y(n_253)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_127),
.B(n_44),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_185),
.B(n_191),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_186),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_187),
.A2(n_222),
.B1(n_229),
.B2(n_172),
.Y(n_239)
);

CKINVDCx12_ASAP7_75t_R g189 ( 
.A(n_135),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_189),
.Y(n_267)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_190),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_44),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_147),
.A2(n_42),
.B1(n_87),
.B2(n_98),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_192),
.A2(n_138),
.B1(n_113),
.B2(n_122),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_33),
.Y(n_193)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_150),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_196),
.Y(n_277)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_136),
.Y(n_197)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_197),
.Y(n_285)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_198),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_134),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_129),
.Y(n_200)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_200),
.Y(n_245)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_202),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_153),
.B(n_33),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_153),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_150),
.Y(n_205)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_205),
.Y(n_283)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_111),
.A2(n_61),
.B1(n_66),
.B2(n_103),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_208),
.A2(n_132),
.B(n_160),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_210),
.B(n_215),
.Y(n_248)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_211),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_154),
.B(n_29),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_212),
.B(n_214),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_121),
.B(n_34),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_105),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_109),
.Y(n_215)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_117),
.Y(n_217)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_217),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_114),
.A2(n_62),
.B1(n_92),
.B2(n_88),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_220),
.A2(n_221),
.B1(n_231),
.B2(n_132),
.Y(n_235)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_115),
.A2(n_77),
.B1(n_54),
.B2(n_89),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_L g222 ( 
.A1(n_155),
.A2(n_56),
.B1(n_60),
.B2(n_79),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_111),
.B(n_39),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_226),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_159),
.Y(n_224)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_155),
.Y(n_225)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_136),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_234),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_119),
.A2(n_72),
.B1(n_67),
.B2(n_48),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_130),
.B1(n_149),
.B2(n_120),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_119),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_233),
.Y(n_252)
);

OA22x2_ASAP7_75t_L g231 ( 
.A1(n_159),
.A2(n_102),
.B1(n_47),
.B2(n_49),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_113),
.B(n_122),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_232),
.B(n_144),
.Y(n_271)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_124),
.B(n_145),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_136),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_235),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_219),
.B(n_148),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_265),
.C(n_278),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_239),
.B(n_241),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_244),
.B(n_263),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_216),
.A2(n_130),
.B1(n_149),
.B2(n_120),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_250),
.A2(n_288),
.B1(n_228),
.B2(n_208),
.Y(n_306)
);

MAJx2_ASAP7_75t_L g265 ( 
.A(n_173),
.B(n_139),
.C(n_102),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_178),
.B(n_167),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_269),
.B(n_270),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_218),
.B(n_167),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_273),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_182),
.B(n_144),
.Y(n_273)
);

NAND2xp33_ASAP7_75t_SL g274 ( 
.A(n_226),
.B(n_145),
.Y(n_274)
);

NAND2xp33_ASAP7_75t_SL g331 ( 
.A(n_274),
.B(n_205),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_193),
.B(n_1),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_282),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_209),
.B(n_201),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_276),
.B(n_286),
.Y(n_312)
);

AND2x2_ASAP7_75t_SL g278 ( 
.A(n_172),
.B(n_139),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_224),
.A2(n_124),
.B1(n_139),
.B2(n_167),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_279),
.A2(n_205),
.B1(n_181),
.B2(n_234),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g281 ( 
.A(n_213),
.B(n_93),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_233),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_232),
.B(n_1),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_176),
.B(n_48),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g287 ( 
.A1(n_213),
.A2(n_34),
.B(n_39),
.C(n_36),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_231),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_222),
.A2(n_49),
.B1(n_47),
.B2(n_36),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_291),
.Y(n_360)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_292),
.Y(n_364)
);

INVx4_ASAP7_75t_SL g294 ( 
.A(n_277),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_297),
.Y(n_351)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_259),
.B(n_236),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_296),
.B(n_299),
.Y(n_342)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_261),
.Y(n_298)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_298),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_254),
.B(n_177),
.Y(n_299)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_300),
.Y(n_345)
);

CKINVDCx12_ASAP7_75t_R g302 ( 
.A(n_267),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_302),
.Y(n_348)
);

INVx4_ASAP7_75t_SL g303 ( 
.A(n_267),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_243),
.Y(n_305)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_305),
.Y(n_380)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_243),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_308),
.B(n_310),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_309),
.A2(n_315),
.B1(n_318),
.B2(n_322),
.Y(n_341)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_313),
.B(n_260),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_254),
.B(n_195),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_316),
.B(n_324),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_259),
.B(n_183),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_333),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_258),
.A2(n_227),
.B1(n_197),
.B2(n_181),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_239),
.A2(n_221),
.B1(n_231),
.B2(n_225),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_319),
.A2(n_326),
.B1(n_244),
.B2(n_278),
.Y(n_340)
);

OR2x4_ASAP7_75t_L g320 ( 
.A(n_274),
.B(n_231),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g346 ( 
.A(n_320),
.B(n_325),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_265),
.B(n_180),
.C(n_230),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_245),
.C(n_251),
.Y(n_359)
);

INVx13_ASAP7_75t_L g322 ( 
.A(n_283),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_252),
.A2(n_221),
.B1(n_190),
.B2(n_211),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_323),
.A2(n_262),
.B1(n_256),
.B2(n_257),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_255),
.B(n_194),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_249),
.B(n_221),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_273),
.A2(n_184),
.B1(n_217),
.B2(n_207),
.Y(n_326)
);

INVx13_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_327),
.A2(n_330),
.B1(n_268),
.B2(n_285),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_247),
.B(n_202),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_328),
.B(n_332),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_263),
.A2(n_205),
.B(n_196),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_329),
.A2(n_331),
.B(n_281),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_284),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_255),
.B(n_188),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_282),
.B(n_175),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_238),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_334),
.B(n_336),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_186),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_337),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_245),
.B(n_174),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_237),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_339),
.A2(n_356),
.B(n_361),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_340),
.A2(n_367),
.B1(n_368),
.B2(n_370),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_240),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_343),
.B(n_359),
.C(n_379),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_313),
.B(n_278),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_344),
.B(n_352),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_292),
.A2(n_250),
.B1(n_240),
.B2(n_242),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_347),
.A2(n_369),
.B1(n_371),
.B2(n_376),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_289),
.B(n_317),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_289),
.B(n_248),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_355),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_293),
.B(n_240),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_329),
.A2(n_262),
.B(n_287),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_331),
.A2(n_262),
.B(n_258),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_306),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_328),
.B(n_238),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_363),
.B(n_294),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_319),
.A2(n_290),
.B1(n_325),
.B2(n_311),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_314),
.A2(n_256),
.B1(n_257),
.B2(n_268),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_290),
.A2(n_268),
.B1(n_251),
.B2(n_280),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g371 ( 
.A1(n_314),
.A2(n_280),
.B1(n_260),
.B2(n_253),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_293),
.B(n_237),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_310),
.Y(n_397)
);

NOR2x1_ASAP7_75t_L g387 ( 
.A(n_374),
.B(n_368),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_309),
.A2(n_266),
.B1(n_264),
.B2(n_272),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_375),
.A2(n_291),
.B(n_330),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_290),
.A2(n_301),
.B1(n_311),
.B2(n_335),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_301),
.A2(n_311),
.B1(n_320),
.B2(n_333),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_377),
.A2(n_330),
.B1(n_266),
.B2(n_264),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_321),
.B(n_253),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_307),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_381),
.B(n_393),
.C(n_396),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_384),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_312),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_385),
.B(n_386),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_348),
.B(n_312),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_387),
.B(n_405),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_339),
.B(n_303),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_388),
.A2(n_390),
.B(n_392),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_340),
.A2(n_304),
.B1(n_295),
.B2(n_305),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_374),
.B1(n_364),
.B2(n_354),
.Y(n_418)
);

AND2x6_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_302),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_303),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_308),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_358),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_395),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_353),
.B(n_326),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_409),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_377),
.B(n_298),
.C(n_272),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_415),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_346),
.A2(n_294),
.B(n_300),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_400),
.A2(n_412),
.B(n_356),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_345),
.Y(n_402)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_402),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_338),
.B(n_309),
.Y(n_403)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_403),
.Y(n_428)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_360),
.Y(n_404)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_373),
.Y(n_406)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_406),
.Y(n_440)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_407),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_408),
.A2(n_402),
.B1(n_357),
.B2(n_404),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_338),
.B(n_337),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_410),
.A2(n_357),
.B1(n_360),
.B2(n_6),
.Y(n_445)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_358),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_414),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g412 ( 
.A(n_344),
.B(n_327),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_349),
.B(n_322),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_18),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_1),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_352),
.B(n_1),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_378),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_417),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_3),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_418),
.A2(n_427),
.B1(n_435),
.B2(n_446),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_388),
.A2(n_346),
.B1(n_354),
.B2(n_374),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_420),
.A2(n_392),
.B1(n_387),
.B2(n_412),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_401),
.A2(n_364),
.B1(n_383),
.B2(n_410),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_422),
.A2(n_437),
.B1(n_411),
.B2(n_403),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_382),
.A2(n_354),
.B1(n_369),
.B2(n_350),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_393),
.B(n_355),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_429),
.B(n_9),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_430),
.A2(n_433),
.B(n_415),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_383),
.B(n_370),
.Y(n_431)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_431),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_394),
.A2(n_341),
.B(n_351),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_397),
.B(n_350),
.Y(n_434)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_434),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_389),
.A2(n_371),
.B1(n_351),
.B2(n_366),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_401),
.A2(n_380),
.B1(n_366),
.B2(n_365),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_391),
.B(n_380),
.Y(n_438)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

NOR4xp25_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_351),
.C(n_359),
.D(n_345),
.Y(n_443)
);

MAJx2_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_396),
.C(n_390),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_365),
.Y(n_444)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_444),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_445),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_407),
.A2(n_357),
.B1(n_5),
.B2(n_7),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_447),
.A2(n_408),
.B1(n_394),
.B2(n_400),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_448),
.B(n_417),
.Y(n_455)
);

INVxp33_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_452),
.B(n_455),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_441),
.B(n_381),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_453),
.B(n_469),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_449),
.B(n_398),
.C(n_399),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_462),
.C(n_473),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_459),
.A2(n_463),
.B1(n_428),
.B2(n_445),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_449),
.B(n_398),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_460),
.B(n_471),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_461),
.A2(n_470),
.B1(n_431),
.B2(n_446),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_426),
.B(n_388),
.C(n_392),
.Y(n_462)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_440),
.Y(n_464)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_465),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_466),
.A2(n_468),
.B(n_420),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_440),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_467),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_439),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_441),
.B(n_7),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_422),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_8),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_429),
.B(n_424),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_438),
.Y(n_474)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_474),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g475 ( 
.A(n_432),
.B(n_8),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_475),
.A2(n_478),
.B1(n_479),
.B2(n_448),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_429),
.C(n_450),
.Y(n_488)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_444),
.Y(n_477)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_477),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_432),
.B(n_9),
.Y(n_478)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_480),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_461),
.A2(n_431),
.B1(n_427),
.B2(n_418),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_483),
.A2(n_500),
.B1(n_451),
.B2(n_419),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_488),
.B(n_489),
.Y(n_513)
);

FAx1_ASAP7_75t_SL g490 ( 
.A(n_473),
.B(n_443),
.CI(n_434),
.CON(n_490),
.SN(n_490)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_490),
.B(n_501),
.Y(n_507)
);

AO221x1_ASAP7_75t_L g519 ( 
.A1(n_491),
.A2(n_471),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_457),
.B(n_450),
.C(n_425),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_492),
.B(n_498),
.C(n_499),
.Y(n_508)
);

NOR2x1_ASAP7_75t_L g494 ( 
.A(n_468),
.B(n_419),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_494),
.B(n_452),
.Y(n_511)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_464),
.Y(n_496)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_496),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_425),
.C(n_437),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_430),
.C(n_439),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_454),
.A2(n_428),
.B1(n_433),
.B2(n_447),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_470),
.A2(n_442),
.B1(n_435),
.B2(n_423),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_502),
.B(n_472),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_503),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g504 ( 
.A1(n_500),
.A2(n_459),
.B(n_451),
.Y(n_504)
);

XNOR2x1_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_512),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_497),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_506),
.A2(n_502),
.B1(n_486),
.B2(n_485),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_510),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_511),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_SL g512 ( 
.A(n_484),
.B(n_465),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_494),
.A2(n_466),
.B(n_456),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g530 ( 
.A(n_514),
.B(n_519),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_515),
.A2(n_518),
.B1(n_491),
.B2(n_486),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_482),
.B(n_436),
.Y(n_516)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_516),
.Y(n_534)
);

OA22x2_ASAP7_75t_L g517 ( 
.A1(n_485),
.A2(n_421),
.B1(n_436),
.B2(n_479),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_517),
.B(n_503),
.C(n_483),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g518 ( 
.A1(n_495),
.A2(n_421),
.B1(n_423),
.B2(n_476),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_520),
.A2(n_521),
.B1(n_480),
.B2(n_497),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_SL g521 ( 
.A1(n_495),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_492),
.B(n_13),
.C(n_14),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_482),
.C(n_496),
.Y(n_523)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_523),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_481),
.C(n_498),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_524),
.A2(n_527),
.B(n_529),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_536),
.Y(n_548)
);

AO21x1_ASAP7_75t_L g542 ( 
.A1(n_526),
.A2(n_516),
.B(n_509),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_481),
.C(n_513),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_499),
.C(n_493),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g540 ( 
.A1(n_531),
.A2(n_504),
.B1(n_506),
.B2(n_507),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_505),
.B(n_493),
.C(n_484),
.Y(n_532)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_532),
.A2(n_535),
.B(n_534),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_533),
.A2(n_507),
.B1(n_511),
.B2(n_510),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_515),
.B(n_488),
.C(n_490),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_522),
.B(n_487),
.Y(n_536)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_540),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_543),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g554 ( 
.A(n_542),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_504),
.C(n_514),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_525),
.A2(n_490),
.B1(n_512),
.B2(n_509),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_545),
.B(n_537),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_529),
.B(n_517),
.C(n_520),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_546),
.A2(n_547),
.B(n_550),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_517),
.C(n_519),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_549),
.B(n_538),
.C(n_530),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_535),
.B(n_517),
.C(n_15),
.Y(n_550)
);

AOI21x1_ASAP7_75t_SL g562 ( 
.A1(n_551),
.A2(n_555),
.B(n_556),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_548),
.Y(n_561)
);

O2A1O1Ixp33_ASAP7_75t_L g555 ( 
.A1(n_542),
.A2(n_528),
.B(n_530),
.C(n_538),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g556 ( 
.A1(n_539),
.A2(n_14),
.B(n_18),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_543),
.Y(n_559)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_559),
.A2(n_560),
.B(n_552),
.Y(n_564)
);

OAI21xp5_ASAP7_75t_SL g560 ( 
.A1(n_551),
.A2(n_544),
.B(n_550),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_561),
.B(n_548),
.C(n_558),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_554),
.A2(n_540),
.B1(n_546),
.B2(n_547),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_563),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_564),
.A2(n_562),
.B(n_555),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_566),
.B(n_561),
.C(n_562),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_567),
.B(n_568),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_569),
.B(n_565),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_570),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_571),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_545),
.B(n_18),
.Y(n_573)
);


endmodule