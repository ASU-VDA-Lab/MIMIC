module real_jpeg_17099_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_7),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_SL g64 ( 
.A(n_7),
.B(n_50),
.Y(n_64)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

A2O1A1Ixp33_ASAP7_75t_L g10 ( 
.A1(n_11),
.A2(n_34),
.B(n_99),
.C(n_103),
.Y(n_10)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_11),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_17),
.Y(n_11)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_45),
.B(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_13),
.A2(n_88),
.B1(n_89),
.B2(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_13),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_24),
.B1(n_25),
.B2(n_33),
.Y(n_17)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_18),
.A2(n_33),
.B1(n_104),
.B2(n_108),
.Y(n_103)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_24),
.A2(n_25),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_25),
.B(n_89),
.C(n_98),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_26),
.Y(n_92)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_SL g99 ( 
.A1(n_33),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_94),
.C(n_95),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_86),
.C(n_87),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_73),
.C(n_74),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_61),
.C(n_62),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_46),
.B(n_56),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_39),
.A2(n_40),
.B1(n_66),
.B2(n_71),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_39),
.B(n_64),
.C(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_66),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_78),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_55),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_50),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_65),
.B2(n_72),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_64),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_78),
.C(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_85),
.Y(n_74)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_75),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_89),
.C(n_92),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_104),
.Y(n_108)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);


endmodule