module fake_jpeg_10081_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_42),
.Y(n_51)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_32),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_29),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_16),
.B(n_0),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_20),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_60),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_27),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_55),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_20),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_40),
.A2(n_31),
.B1(n_26),
.B2(n_25),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_27),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_35),
.A2(n_26),
.B1(n_25),
.B2(n_24),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_35),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_28),
.B1(n_22),
.B2(n_37),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_21),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_23),
.B(n_18),
.C(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_21),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_22),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_72),
.Y(n_90)
);

AOI32xp33_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_19),
.A3(n_43),
.B1(n_41),
.B2(n_30),
.Y(n_66)
);

AOI21xp33_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_44),
.B(n_19),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_28),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_82),
.B1(n_84),
.B2(n_72),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_71),
.Y(n_105)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_83),
.Y(n_103)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_76),
.A2(n_56),
.B1(n_50),
.B2(n_39),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_19),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_54),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_62),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_30),
.B1(n_41),
.B2(n_43),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_46),
.A2(n_43),
.B1(n_41),
.B2(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_61),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_85),
.B(n_88),
.Y(n_118)
);

NOR2x1_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_51),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_89),
.B(n_94),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_87),
.A2(n_99),
.B1(n_73),
.B2(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_44),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_92),
.B(n_97),
.Y(n_120)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_101),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_54),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_71),
.B(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_106),
.B1(n_76),
.B2(n_51),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_46),
.B1(n_39),
.B2(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_79),
.Y(n_102)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_104),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_79),
.A2(n_56),
.B1(n_49),
.B2(n_25),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_115),
.B1(n_106),
.B2(n_97),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_108),
.A2(n_110),
.B(n_109),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_94),
.A2(n_71),
.B(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_94),
.Y(n_128)
);

AOI322xp5_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_15),
.A3(n_11),
.B1(n_10),
.B2(n_74),
.C1(n_71),
.C2(n_64),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_117),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_96),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_38),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_76),
.B(n_89),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_93),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_124),
.B(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_127),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_85),
.Y(n_129)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_130),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_134),
.B(n_140),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_135),
.A2(n_115),
.B1(n_112),
.B2(n_109),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_102),
.C(n_110),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_138),
.C(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_137),
.A2(n_139),
.B1(n_143),
.B2(n_113),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_103),
.C(n_86),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_119),
.B(n_103),
.C(n_101),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_89),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_146),
.B(n_151),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_135),
.A2(n_98),
.B1(n_111),
.B2(n_95),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_153),
.B(n_156),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_105),
.B(n_64),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_155),
.B1(n_158),
.B2(n_38),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_136),
.B1(n_130),
.B2(n_128),
.Y(n_155)
);

NAND3xp33_ASAP7_75t_L g156 ( 
.A(n_131),
.B(n_11),
.C(n_2),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_157),
.B(n_62),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_141),
.A2(n_105),
.B1(n_26),
.B2(n_25),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_143),
.A3(n_138),
.B1(n_129),
.B2(n_126),
.C1(n_19),
.C2(n_74),
.Y(n_159)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_159),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_62),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

AOI321xp33_ASAP7_75t_L g161 ( 
.A1(n_147),
.A2(n_19),
.A3(n_38),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_157),
.B(n_1),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_162),
.B(n_163),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_38),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_165),
.B(n_38),
.C(n_3),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_166),
.A2(n_168),
.B(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_148),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_19),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_1),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_171),
.A2(n_154),
.B1(n_144),
.B2(n_148),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_174),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_168),
.A2(n_145),
.B1(n_152),
.B2(n_62),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_177),
.A2(n_165),
.B1(n_161),
.B2(n_6),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_178),
.B(n_170),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_180),
.B(n_9),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_181),
.A2(n_187),
.B(n_188),
.Y(n_193)
);

NOR2xp67_ASAP7_75t_L g183 ( 
.A(n_179),
.B(n_171),
.Y(n_183)
);

OAI221xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_172),
.B1(n_180),
.B2(n_173),
.C(n_8),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_175),
.B(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_186),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_8),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_176),
.A2(n_2),
.B1(n_4),
.B2(n_7),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_2),
.B(n_7),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_187),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_192),
.Y(n_197)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_8),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_9),
.C(n_191),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_9),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_196),
.B(n_189),
.C(n_197),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_200),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_195),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_202),
.Y(n_204)
);


endmodule