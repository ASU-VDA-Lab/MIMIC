module fake_jpeg_24957_n_170 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_36),
.B(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_37),
.B(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_46),
.B(n_65),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_25),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_57),
.B(n_61),
.C(n_19),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_31),
.B1(n_17),
.B2(n_18),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_26),
.B1(n_17),
.B2(n_18),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_21),
.B1(n_30),
.B2(n_23),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_32),
.A2(n_21),
.B1(n_28),
.B2(n_24),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_53),
.A2(n_48),
.B(n_52),
.C(n_45),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_33),
.A2(n_23),
.B1(n_27),
.B2(n_16),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_27),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_43),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_38),
.A2(n_29),
.B(n_19),
.C(n_2),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_67),
.B(n_73),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_57),
.A2(n_33),
.B1(n_38),
.B2(n_42),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_85),
.B1(n_89),
.B2(n_61),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_34),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_53),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_62),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_74),
.A2(n_77),
.B(n_71),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_33),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_50),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_65),
.B(n_11),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_38),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_40),
.C(n_39),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_58),
.C(n_54),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_43),
.B1(n_42),
.B2(n_40),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_1),
.B1(n_8),
.B2(n_9),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_44),
.B(n_39),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_87),
.A2(n_10),
.B1(n_12),
.B2(n_13),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_72),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_88),
.B(n_64),
.C(n_59),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_100),
.C(n_101),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_103),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_49),
.C(n_50),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_102),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_1),
.C(n_6),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_107),
.A2(n_88),
.B1(n_74),
.B2(n_86),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_94),
.B1(n_93),
.B2(n_91),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_114),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_70),
.Y(n_112)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_112),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_81),
.C(n_66),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_120),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_82),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_73),
.B(n_71),
.Y(n_128)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_118),
.B(n_119),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_104),
.B(n_76),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_75),
.Y(n_124)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_124),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_100),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_104),
.C(n_103),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_129),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_102),
.B(n_81),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_116),
.A2(n_94),
.B1(n_93),
.B2(n_84),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_132),
.A2(n_137),
.B1(n_91),
.B2(n_79),
.Y(n_139)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_131),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_140),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_137),
.Y(n_140)
);

XOR2x1_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_115),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_134),
.A2(n_109),
.B1(n_113),
.B2(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_147),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_127),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_146),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_133),
.A2(n_122),
.B1(n_118),
.B2(n_120),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_126),
.C(n_117),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_152),
.C(n_153),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_129),
.C(n_135),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_143),
.B(n_136),
.C(n_112),
.Y(n_153)
);

BUFx12f_ASAP7_75t_SL g154 ( 
.A(n_141),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_154),
.A2(n_146),
.B(n_140),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_156),
.Y(n_164)
);

AOI322xp5_ASAP7_75t_L g157 ( 
.A1(n_149),
.A2(n_116),
.A3(n_142),
.B1(n_136),
.B2(n_125),
.C1(n_138),
.C2(n_114),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_157),
.Y(n_161)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_158),
.B(n_159),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g159 ( 
.A1(n_149),
.A2(n_95),
.A3(n_105),
.B1(n_110),
.B2(n_78),
.C1(n_14),
.C2(n_13),
.Y(n_159)
);

OR2x6_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_162),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_162),
.B(n_155),
.C(n_105),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_166),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_164),
.A2(n_110),
.B1(n_12),
.B2(n_9),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_163),
.B1(n_9),
.B2(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_169),
.Y(n_170)
);


endmodule