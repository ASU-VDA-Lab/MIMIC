module fake_aes_10608_n_671 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_671);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_671;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_455;
wire n_312;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx6f_ASAP7_75t_L g90 ( .A(n_30), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_1), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_11), .Y(n_92) );
NAND2xp5_ASAP7_75t_L g93 ( .A(n_52), .B(n_58), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_31), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_56), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_47), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_44), .Y(n_97) );
BUFx3_ASAP7_75t_L g98 ( .A(n_75), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_6), .Y(n_99) );
BUFx10_ASAP7_75t_L g100 ( .A(n_14), .Y(n_100) );
BUFx8_ASAP7_75t_SL g101 ( .A(n_11), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_12), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_64), .Y(n_103) );
HB1xp67_ASAP7_75t_L g104 ( .A(n_51), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_88), .Y(n_105) );
INVxp67_ASAP7_75t_SL g106 ( .A(n_60), .Y(n_106) );
BUFx10_ASAP7_75t_L g107 ( .A(n_87), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_85), .Y(n_108) );
INVxp67_ASAP7_75t_L g109 ( .A(n_74), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_4), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_29), .Y(n_111) );
INVx4_ASAP7_75t_R g112 ( .A(n_76), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_10), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_40), .Y(n_114) );
INVxp67_ASAP7_75t_SL g115 ( .A(n_27), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_14), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_34), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_49), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_38), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_43), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_7), .Y(n_122) );
CKINVDCx16_ASAP7_75t_R g123 ( .A(n_72), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_57), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_61), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_89), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_6), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_3), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_53), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_46), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_124), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_104), .B(n_0), .Y(n_133) );
AND2x6_ASAP7_75t_L g134 ( .A(n_98), .B(n_36), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_105), .B(n_0), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_90), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_90), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_90), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_90), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_110), .B(n_1), .Y(n_141) );
BUFx3_ASAP7_75t_L g142 ( .A(n_98), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_90), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_103), .Y(n_144) );
INVx4_ASAP7_75t_L g145 ( .A(n_107), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_103), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_126), .Y(n_147) );
OAI21x1_ASAP7_75t_L g148 ( .A1(n_126), .A2(n_39), .B(n_84), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_129), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_129), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_123), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_130), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_130), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_99), .B(n_2), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_100), .B(n_2), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_108), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_101), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_116), .Y(n_158) );
INVx2_ASAP7_75t_SL g159 ( .A(n_145), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_136), .Y(n_160) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_141), .B(n_111), .Y(n_161) );
INVxp67_ASAP7_75t_L g162 ( .A(n_155), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_145), .B(n_99), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g164 ( .A(n_145), .B(n_109), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_136), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_145), .B(n_102), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
INVx4_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_137), .B(n_102), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_151), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_141), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_155), .B(n_137), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_144), .B(n_107), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
INVx4_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
AND2x6_ASAP7_75t_SL g179 ( .A(n_141), .B(n_92), .Y(n_179) );
BUFx2_ASAP7_75t_L g180 ( .A(n_142), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_144), .B(n_114), .Y(n_182) );
NOR2xp33_ASAP7_75t_SL g183 ( .A(n_134), .B(n_94), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_132), .Y(n_184) );
NAND2xp33_ASAP7_75t_SL g185 ( .A(n_157), .B(n_127), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g186 ( .A1(n_133), .A2(n_127), .B1(n_91), .B2(n_122), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_134), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_149), .Y(n_188) );
OR2x6_ASAP7_75t_L g189 ( .A(n_135), .B(n_92), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_146), .B(n_119), .Y(n_190) );
AND2x4_ASAP7_75t_L g191 ( .A(n_146), .B(n_110), .Y(n_191) );
INVx5_ASAP7_75t_L g192 ( .A(n_134), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_147), .B(n_113), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_163), .B(n_147), .Y(n_194) );
BUFx2_ASAP7_75t_L g195 ( .A(n_189), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_173), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_161), .Y(n_197) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_175), .A2(n_150), .B1(n_156), .B2(n_153), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_177), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_175), .B(n_150), .Y(n_200) );
INVxp67_ASAP7_75t_L g201 ( .A(n_177), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_169), .B(n_94), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_181), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_159), .B(n_142), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_159), .B(n_142), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_181), .Y(n_206) );
AND2x6_ASAP7_75t_SL g207 ( .A(n_189), .B(n_158), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_169), .B(n_178), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_184), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_160), .Y(n_210) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_189), .A2(n_134), .B1(n_156), .B2(n_152), .Y(n_211) );
OAI22xp5_ASAP7_75t_L g212 ( .A1(n_161), .A2(n_131), .B1(n_152), .B2(n_149), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_167), .B(n_153), .Y(n_213) );
AND2x4_ASAP7_75t_SL g214 ( .A(n_169), .B(n_107), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_184), .Y(n_217) );
AOI221xp5_ASAP7_75t_SL g218 ( .A1(n_168), .A2(n_113), .B1(n_125), .B2(n_121), .C(n_120), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_189), .A2(n_134), .B1(n_100), .B2(n_97), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_178), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_164), .B(n_96), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_165), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_165), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g225 ( .A1(n_186), .A2(n_128), .B1(n_96), .B2(n_97), .Y(n_225) );
INVxp67_ASAP7_75t_L g226 ( .A(n_170), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_180), .B(n_118), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_188), .Y(n_228) );
INVx1_ASAP7_75t_SL g229 ( .A(n_173), .Y(n_229) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_161), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_178), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g232 ( .A1(n_183), .A2(n_100), .B1(n_118), .B2(n_117), .Y(n_232) );
INVxp67_ASAP7_75t_SL g233 ( .A(n_180), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_166), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_168), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_187), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_174), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_174), .B(n_148), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_226), .B(n_179), .Y(n_239) );
INVxp33_ASAP7_75t_SL g240 ( .A(n_229), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_238), .A2(n_187), .B(n_192), .Y(n_241) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_220), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_203), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_210), .Y(n_244) );
BUFx8_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_230), .B(n_187), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_199), .B(n_191), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_230), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_201), .A2(n_176), .B1(n_185), .B2(n_182), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_216), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_SL g252 ( .A1(n_194), .A2(n_190), .B(n_140), .C(n_138), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_216), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_238), .A2(n_192), .B(n_148), .Y(n_254) );
O2A1O1Ixp33_ASAP7_75t_SL g255 ( .A1(n_213), .A2(n_93), .B(n_106), .C(n_115), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_203), .Y(n_256) );
NAND2xp33_ASAP7_75t_L g257 ( .A(n_197), .B(n_192), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_223), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_206), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_230), .Y(n_260) );
INVx4_ASAP7_75t_L g261 ( .A(n_197), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_200), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_215), .B(n_193), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_238), .A2(n_192), .B(n_193), .Y(n_264) );
BUFx3_ASAP7_75t_L g265 ( .A(n_197), .Y(n_265) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_195), .A2(n_198), .B1(n_196), .B2(n_212), .Y(n_266) );
INVx4_ASAP7_75t_L g267 ( .A(n_214), .Y(n_267) );
NOR3xp33_ASAP7_75t_L g268 ( .A(n_225), .B(n_117), .C(n_191), .Y(n_268) );
INVx4_ASAP7_75t_L g269 ( .A(n_214), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_227), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_198), .B(n_193), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_233), .B(n_191), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_209), .Y(n_274) );
BUFx3_ASAP7_75t_L g275 ( .A(n_220), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_207), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_223), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_220), .Y(n_278) );
BUFx4f_ASAP7_75t_L g279 ( .A(n_214), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_238), .A2(n_192), .B(n_171), .Y(n_280) );
CKINVDCx11_ASAP7_75t_R g281 ( .A(n_207), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_225), .Y(n_282) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
BUFx8_ASAP7_75t_L g284 ( .A(n_260), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_254), .A2(n_237), .B(n_235), .Y(n_285) );
CKINVDCx6p67_ASAP7_75t_R g286 ( .A(n_260), .Y(n_286) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_279), .B(n_236), .Y(n_287) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_264), .A2(n_218), .B(n_237), .Y(n_288) );
BUFx8_ASAP7_75t_L g289 ( .A(n_248), .Y(n_289) );
AOI22xp33_ASAP7_75t_SL g290 ( .A1(n_240), .A2(n_222), .B1(n_217), .B2(n_209), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_280), .A2(n_235), .B(n_211), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_241), .A2(n_192), .B(n_205), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_262), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_244), .Y(n_294) );
AND2x4_ASAP7_75t_L g295 ( .A(n_248), .B(n_217), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_243), .A2(n_221), .B(n_228), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_247), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_252), .A2(n_228), .B(n_221), .Y(n_298) );
NOR2x1_ASAP7_75t_SL g299 ( .A(n_267), .B(n_269), .Y(n_299) );
AOI21xp33_ASAP7_75t_L g300 ( .A1(n_239), .A2(n_219), .B(n_232), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_243), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_242), .Y(n_302) );
AO31x2_ASAP7_75t_L g303 ( .A1(n_256), .A2(n_138), .A3(n_139), .B(n_140), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_244), .Y(n_304) );
OAI21x1_ASAP7_75t_L g305 ( .A1(n_256), .A2(n_204), .B(n_208), .Y(n_305) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_259), .A2(n_202), .B(n_234), .Y(n_306) );
OAI21x1_ASAP7_75t_L g307 ( .A1(n_259), .A2(n_234), .B(n_224), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_240), .B(n_231), .Y(n_308) );
BUFx8_ASAP7_75t_L g309 ( .A(n_271), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_272), .A2(n_224), .B(n_139), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_271), .B(n_218), .Y(n_311) );
OAI21x1_ASAP7_75t_L g312 ( .A1(n_272), .A2(n_139), .B(n_140), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_249), .A2(n_231), .B(n_236), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_282), .B(n_3), .Y(n_314) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_274), .A2(n_171), .B(n_166), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_245), .Y(n_316) );
OAI21x1_ASAP7_75t_L g317 ( .A1(n_274), .A2(n_112), .B(n_143), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_268), .A2(n_143), .B1(n_172), .B2(n_7), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_301), .A2(n_266), .B1(n_271), .B2(n_279), .Y(n_320) );
OAI22x1_ASAP7_75t_L g321 ( .A1(n_314), .A2(n_276), .B1(n_270), .B2(n_267), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_299), .B(n_301), .Y(n_322) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
OAI22xp33_ASAP7_75t_L g324 ( .A1(n_316), .A2(n_279), .B1(n_276), .B2(n_267), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_311), .A2(n_263), .B1(n_281), .B2(n_273), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_293), .B(n_245), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_289), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_292), .A2(n_251), .B(n_253), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_296), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_297), .B(n_319), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_307), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g332 ( .A1(n_290), .A2(n_245), .B1(n_269), .B2(n_261), .Y(n_332) );
AND2x2_ASAP7_75t_L g333 ( .A(n_311), .B(n_249), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_300), .A2(n_269), .B1(n_261), .B2(n_265), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_309), .A2(n_250), .B1(n_258), .B2(n_277), .Y(n_335) );
AOI22xp33_ASAP7_75t_L g336 ( .A1(n_309), .A2(n_261), .B1(n_265), .B2(n_278), .Y(n_336) );
BUFx2_ASAP7_75t_L g337 ( .A(n_309), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_284), .Y(n_338) );
INVx4_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_285), .A2(n_277), .B(n_251), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_308), .A2(n_278), .B1(n_275), .B2(n_283), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_296), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_295), .A2(n_275), .B1(n_242), .B2(n_283), .Y(n_344) );
AOI21xp5_ASAP7_75t_L g345 ( .A1(n_285), .A2(n_253), .B(n_258), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_316), .B(n_255), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_294), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_294), .B(n_283), .Y(n_348) );
AOI22xp33_ASAP7_75t_L g349 ( .A1(n_295), .A2(n_242), .B1(n_283), .B2(n_246), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_333), .B(n_304), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_331), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_339), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_333), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_320), .B(n_288), .Y(n_354) );
BUFx3_ASAP7_75t_L g355 ( .A(n_327), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_304), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_347), .B(n_286), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_329), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_347), .B(n_288), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_347), .Y(n_361) );
AO31x2_ASAP7_75t_L g362 ( .A1(n_329), .A2(n_299), .A3(n_315), .B(n_288), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_330), .B(n_322), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_322), .B(n_298), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_339), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_325), .B(n_286), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_331), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_330), .B(n_298), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_335), .A2(n_318), .B1(n_287), .B2(n_295), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_343), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_322), .B(n_298), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_343), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_348), .B(n_302), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_331), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_342), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_342), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_348), .B(n_302), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_371), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_367), .A2(n_337), .B1(n_325), .B2(n_327), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_364), .B(n_342), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_350), .B(n_340), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_355), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_376), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_350), .B(n_357), .Y(n_386) );
AOI22xp5_ASAP7_75t_L g387 ( .A1(n_363), .A2(n_337), .B1(n_335), .B2(n_327), .Y(n_387) );
INVx3_ASAP7_75t_L g388 ( .A(n_352), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_350), .B(n_340), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_376), .Y(n_390) );
INVx4_ASAP7_75t_L g391 ( .A(n_352), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_357), .B(n_339), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_353), .B(n_303), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_353), .B(n_334), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_363), .B(n_303), .Y(n_395) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_359), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_367), .A2(n_321), .B1(n_332), .B2(n_346), .Y(n_397) );
INVx1_ASAP7_75t_SL g398 ( .A(n_355), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_374), .B(n_378), .Y(n_399) );
OR2x6_ASAP7_75t_L g400 ( .A(n_356), .B(n_323), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_371), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_374), .B(n_303), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_374), .B(n_303), .Y(n_403) );
BUFx2_ASAP7_75t_SL g404 ( .A(n_355), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_373), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_378), .B(n_303), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_373), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_358), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_361), .B(n_345), .Y(n_409) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_370), .A2(n_321), .B(n_324), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_352), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_378), .B(n_323), .Y(n_412) );
NAND3xp33_ASAP7_75t_L g413 ( .A(n_369), .B(n_326), .C(n_341), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_359), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_385), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_399), .B(n_361), .Y(n_416) );
INVx1_ASAP7_75t_SL g417 ( .A(n_404), .Y(n_417) );
OAI31xp33_ASAP7_75t_L g418 ( .A1(n_410), .A2(n_338), .A3(n_370), .B(n_358), .Y(n_418) );
OR2x6_ASAP7_75t_L g419 ( .A(n_404), .B(n_352), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_399), .B(n_364), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_382), .B(n_364), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_380), .B(n_284), .Y(n_422) );
INVx1_ASAP7_75t_SL g423 ( .A(n_383), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_382), .B(n_372), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_408), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_396), .B(n_369), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_379), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_408), .B(n_365), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_379), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_401), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_401), .Y(n_431) );
BUFx2_ASAP7_75t_L g432 ( .A(n_391), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_385), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_391), .B(n_365), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_405), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_389), .B(n_372), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_385), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_405), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_386), .B(n_393), .Y(n_439) );
INVx4_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_386), .B(n_365), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_396), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_393), .B(n_365), .Y(n_443) );
OR2x2_ASAP7_75t_L g444 ( .A(n_414), .B(n_354), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_407), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_407), .B(n_366), .Y(n_446) );
NOR2x1_ASAP7_75t_L g447 ( .A(n_391), .B(n_366), .Y(n_447) );
NAND2xp33_ASAP7_75t_SL g448 ( .A(n_380), .B(n_366), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_414), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_389), .Y(n_450) );
INVxp67_ASAP7_75t_L g451 ( .A(n_383), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_402), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_395), .B(n_366), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_395), .B(n_360), .Y(n_454) );
OR2x6_ASAP7_75t_L g455 ( .A(n_388), .B(n_356), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_381), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_377), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_410), .A2(n_354), .B1(n_336), .B2(n_349), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_384), .B(n_377), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_402), .Y(n_460) );
AND2x6_ASAP7_75t_L g461 ( .A(n_392), .B(n_351), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_381), .Y(n_462) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_388), .B(n_351), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_397), .B(n_360), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_412), .B(n_368), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_430), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_430), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_452), .B(n_403), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_460), .B(n_403), .Y(n_469) );
NAND2x2_ASAP7_75t_L g470 ( .A(n_464), .B(n_397), .Y(n_470) );
OR2x2_ASAP7_75t_L g471 ( .A(n_439), .B(n_384), .Y(n_471) );
INVx2_ASAP7_75t_SL g472 ( .A(n_440), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_416), .B(n_390), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_449), .B(n_406), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_425), .B(n_406), .Y(n_475) );
NOR2xp67_ASAP7_75t_L g476 ( .A(n_440), .B(n_388), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_431), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_420), .B(n_381), .Y(n_479) );
AND3x2_ASAP7_75t_L g480 ( .A(n_432), .B(n_390), .C(n_392), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_450), .B(n_394), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_420), .B(n_381), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_445), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_450), .B(n_394), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_440), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_457), .B(n_398), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_457), .B(n_398), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_424), .B(n_388), .Y(n_488) );
INVxp67_ASAP7_75t_L g489 ( .A(n_432), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_427), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_442), .B(n_413), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_422), .B(n_387), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_429), .B(n_435), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_445), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_438), .B(n_413), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_446), .Y(n_496) );
NAND4xp25_ASAP7_75t_SL g497 ( .A(n_417), .B(n_387), .C(n_344), .D(n_284), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_459), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_415), .Y(n_499) );
NOR3xp33_ASAP7_75t_L g500 ( .A(n_448), .B(n_411), .C(n_409), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_454), .B(n_409), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_424), .B(n_411), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_421), .B(n_411), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_459), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_426), .Y(n_505) );
INVx2_ASAP7_75t_SL g506 ( .A(n_419), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_436), .B(n_411), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g508 ( .A1(n_448), .A2(n_143), .B1(n_360), .B2(n_368), .C(n_375), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_423), .B(n_4), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_421), .B(n_400), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_436), .B(n_362), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_453), .B(n_368), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_465), .B(n_400), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_415), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_465), .B(n_362), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_441), .B(n_400), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_451), .B(n_400), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_434), .A2(n_400), .B(n_375), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_426), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_443), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_456), .B(n_400), .Y(n_521) );
INVx1_ASAP7_75t_SL g522 ( .A(n_419), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_444), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_456), .B(n_375), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_428), .B(n_362), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_444), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_492), .A2(n_461), .B1(n_419), .B2(n_455), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_489), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_523), .B(n_418), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_485), .B(n_447), .Y(n_530) );
AOI21xp33_ASAP7_75t_L g531 ( .A1(n_509), .A2(n_434), .B(n_458), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_526), .B(n_505), .Y(n_532) );
O2A1O1Ixp33_ASAP7_75t_SL g533 ( .A1(n_472), .A2(n_419), .B(n_461), .C(n_462), .Y(n_533) );
OAI21xp33_ASAP7_75t_L g534 ( .A1(n_492), .A2(n_455), .B(n_462), .Y(n_534) );
INVx2_ASAP7_75t_SL g535 ( .A(n_472), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_479), .B(n_455), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_519), .Y(n_537) );
OAI32xp33_ASAP7_75t_L g538 ( .A1(n_470), .A2(n_461), .A3(n_437), .B1(n_433), .B2(n_287), .Y(n_538) );
INVx2_ASAP7_75t_SL g539 ( .A(n_485), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_489), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g541 ( .A1(n_509), .A2(n_461), .B(n_463), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_475), .B(n_455), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_520), .B(n_461), .Y(n_543) );
OAI21xp33_ASAP7_75t_L g544 ( .A1(n_491), .A2(n_437), .B(n_433), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_485), .B(n_461), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_496), .B(n_362), .Y(n_546) );
OAI222xp33_ASAP7_75t_L g547 ( .A1(n_506), .A2(n_328), .B1(n_362), .B2(n_9), .C1(n_10), .C2(n_12), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g548 ( .A1(n_470), .A2(n_317), .B1(n_289), .B2(n_302), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_479), .B(n_362), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_482), .B(n_362), .Y(n_550) );
OAI22xp33_ASAP7_75t_L g551 ( .A1(n_506), .A2(n_323), .B1(n_302), .B2(n_313), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_482), .B(n_323), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_471), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_497), .A2(n_317), .B1(n_289), .B2(n_143), .Y(n_554) );
INVx2_ASAP7_75t_SL g555 ( .A(n_486), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_501), .B(n_143), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_498), .B(n_5), .Y(n_557) );
AND2x2_ASAP7_75t_SL g558 ( .A(n_500), .B(n_323), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_504), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_490), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_473), .B(n_5), .Y(n_561) );
AOI21xp33_ASAP7_75t_L g562 ( .A1(n_495), .A2(n_8), .B(n_9), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_468), .B(n_8), .Y(n_563) );
AOI222xp33_ASAP7_75t_L g564 ( .A1(n_511), .A2(n_13), .B1(n_15), .B2(n_16), .C1(n_17), .C2(n_18), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_476), .A2(n_310), .B(n_291), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_499), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_469), .B(n_13), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_500), .A2(n_323), .B1(n_291), .B2(n_306), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_481), .B(n_15), .Y(n_569) );
NAND4xp25_ASAP7_75t_L g570 ( .A(n_508), .B(n_16), .C(n_17), .D(n_18), .Y(n_570) );
AOI322xp5_ASAP7_75t_L g571 ( .A1(n_522), .A2(n_257), .A3(n_283), .B1(n_242), .B2(n_310), .C1(n_23), .C2(n_24), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_493), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_484), .B(n_474), .Y(n_573) );
AOI211x1_ASAP7_75t_L g574 ( .A1(n_503), .A2(n_19), .B(n_20), .C(n_21), .Y(n_574) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_499), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_510), .A2(n_257), .B1(n_312), .B2(n_242), .Y(n_576) );
INVx1_ASAP7_75t_SL g577 ( .A(n_487), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_466), .B(n_305), .Y(n_578) );
OAI21xp33_ASAP7_75t_SL g579 ( .A1(n_510), .A2(n_312), .B(n_305), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_556), .Y(n_580) );
XNOR2xp5_ASAP7_75t_L g581 ( .A(n_577), .B(n_507), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_536), .B(n_502), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_529), .B(n_488), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_560), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_564), .B(n_525), .C(n_518), .D(n_517), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_549), .B(n_513), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g587 ( .A1(n_527), .A2(n_515), .B1(n_512), .B2(n_513), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_555), .A2(n_516), .B1(n_521), .B2(n_467), .Y(n_588) );
INVxp33_ASAP7_75t_L g589 ( .A(n_530), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_566), .Y(n_590) );
INVx1_ASAP7_75t_L g591 ( .A(n_572), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_532), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_528), .Y(n_593) );
XNOR2x1_ASAP7_75t_L g594 ( .A(n_561), .B(n_480), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_575), .Y(n_595) );
OAI22xp33_ASAP7_75t_L g596 ( .A1(n_541), .A2(n_480), .B1(n_478), .B2(n_477), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_553), .B(n_494), .Y(n_597) );
O2A1O1Ixp33_ASAP7_75t_L g598 ( .A1(n_570), .A2(n_494), .B(n_483), .C(n_514), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_559), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_537), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_550), .B(n_483), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_570), .A2(n_514), .B1(n_524), .B2(n_26), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_573), .B(n_524), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g604 ( .A1(n_545), .A2(n_172), .B1(n_25), .B2(n_28), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_535), .Y(n_605) );
AOI222xp33_ASAP7_75t_L g606 ( .A1(n_557), .A2(n_306), .B1(n_172), .B2(n_33), .C1(n_35), .C2(n_37), .Y(n_606) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_567), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_540), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_531), .B(n_22), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_542), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_546), .B(n_32), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_552), .B(n_539), .Y(n_612) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_534), .A2(n_172), .B1(n_42), .B2(n_45), .Y(n_613) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_547), .A2(n_41), .B(n_48), .C(n_54), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_545), .B(n_55), .Y(n_615) );
OAI22xp5_ASAP7_75t_SL g616 ( .A1(n_607), .A2(n_574), .B1(n_558), .B2(n_576), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_608), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_607), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_597), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_593), .Y(n_620) );
NAND4xp25_ASAP7_75t_L g621 ( .A(n_598), .B(n_548), .C(n_562), .D(n_534), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g622 ( .A1(n_585), .A2(n_538), .B1(n_563), .B2(n_569), .C(n_544), .Y(n_622) );
OAI32xp33_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_543), .A3(n_579), .B1(n_544), .B2(n_533), .Y(n_623) );
INVx2_ASAP7_75t_L g624 ( .A(n_595), .Y(n_624) );
OAI21xp5_ASAP7_75t_L g625 ( .A1(n_598), .A2(n_571), .B(n_551), .Y(n_625) );
OAI321xp33_ASAP7_75t_L g626 ( .A1(n_596), .A2(n_554), .A3(n_568), .B1(n_565), .B2(n_578), .C(n_571), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_583), .B(n_59), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g628 ( .A(n_594), .B(n_62), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_605), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_602), .A2(n_63), .B(n_65), .C(n_66), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_591), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_580), .B(n_67), .Y(n_632) );
AOI22xp5_ASAP7_75t_L g633 ( .A1(n_587), .A2(n_172), .B1(n_69), .B2(n_70), .Y(n_633) );
INVx3_ASAP7_75t_SL g634 ( .A(n_615), .Y(n_634) );
OAI322xp33_ASAP7_75t_L g635 ( .A1(n_596), .A2(n_68), .A3(n_71), .B1(n_73), .B2(n_77), .C1(n_78), .C2(n_79), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g636 ( .A1(n_589), .A2(n_80), .B(n_81), .C(n_82), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_584), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_618), .B(n_592), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_629), .B(n_586), .Y(n_639) );
OAI21xp33_ASAP7_75t_L g640 ( .A1(n_623), .A2(n_588), .B(n_610), .Y(n_640) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_634), .Y(n_641) );
NOR4xp25_ASAP7_75t_L g642 ( .A(n_626), .B(n_602), .C(n_614), .D(n_599), .Y(n_642) );
BUFx2_ASAP7_75t_L g643 ( .A(n_629), .Y(n_643) );
A2O1A1Ixp33_ASAP7_75t_L g644 ( .A1(n_630), .A2(n_614), .B(n_609), .C(n_613), .Y(n_644) );
NAND4xp25_ASAP7_75t_L g645 ( .A(n_625), .B(n_606), .C(n_609), .D(n_604), .Y(n_645) );
NAND4xp25_ASAP7_75t_L g646 ( .A(n_621), .B(n_611), .C(n_601), .D(n_600), .Y(n_646) );
AOI221x1_ASAP7_75t_L g647 ( .A1(n_621), .A2(n_603), .B1(n_590), .B2(n_612), .C(n_582), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_619), .Y(n_648) );
AOI211xp5_ASAP7_75t_SL g649 ( .A1(n_616), .A2(n_581), .B(n_83), .C(n_86), .Y(n_649) );
AOI211xp5_ASAP7_75t_L g650 ( .A1(n_622), .A2(n_635), .B(n_627), .C(n_620), .Y(n_650) );
OAI21xp5_ASAP7_75t_L g651 ( .A1(n_642), .A2(n_628), .B(n_636), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_643), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_639), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_641), .B(n_637), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_648), .B(n_617), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_650), .B(n_631), .Y(n_656) );
NOR4xp75_ASAP7_75t_SL g657 ( .A(n_638), .B(n_632), .C(n_624), .D(n_633), .Y(n_657) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_651), .B(n_645), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_652), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_654), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_653), .B(n_646), .Y(n_661) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_659), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_660), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_661), .Y(n_664) );
AO22x1_ASAP7_75t_L g665 ( .A1(n_663), .A2(n_658), .B1(n_651), .B2(n_656), .Y(n_665) );
AOI22x1_ASAP7_75t_L g666 ( .A1(n_663), .A2(n_649), .B1(n_657), .B2(n_655), .Y(n_666) );
INVx2_ASAP7_75t_L g667 ( .A(n_666), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_665), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_668), .A2(n_664), .B1(n_662), .B2(n_640), .C1(n_644), .C2(n_647), .Y(n_669) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_669), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_670), .A2(n_667), .B(n_644), .Y(n_671) );
endmodule