module fake_jpeg_15223_n_319 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_0),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g40 ( 
.A(n_33),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_40),
.Y(n_46)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_56),
.Y(n_77)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_31),
.B1(n_29),
.B2(n_32),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_54),
.A2(n_59),
.B1(n_39),
.B2(n_26),
.Y(n_94)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_36),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_63),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_31),
.B1(n_32),
.B2(n_18),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_31),
.B1(n_20),
.B2(n_32),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_60),
.B(n_28),
.Y(n_91)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_66),
.Y(n_86)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_22),
.Y(n_95)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_17),
.B1(n_21),
.B2(n_33),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_40),
.B1(n_43),
.B2(n_44),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_74),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_40),
.C(n_37),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_37),
.B1(n_42),
.B2(n_41),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_71),
.A2(n_81),
.B1(n_92),
.B2(n_88),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_37),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_83),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_42),
.B1(n_41),
.B2(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_39),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_47),
.Y(n_108)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_39),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_16),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_93),
.B(n_16),
.Y(n_97)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_68),
.B(n_66),
.C(n_65),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_22),
.B1(n_20),
.B2(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_22),
.Y(n_104)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_101),
.B(n_95),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_74),
.A2(n_47),
.B1(n_61),
.B2(n_38),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_58),
.B1(n_72),
.B2(n_73),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_R g101 ( 
.A1(n_91),
.A2(n_68),
.B1(n_23),
.B2(n_21),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_109),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_45),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_91),
.B(n_82),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_70),
.A2(n_38),
.B1(n_43),
.B2(n_44),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_114),
.A2(n_121),
.B1(n_123),
.B2(n_96),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_40),
.C(n_35),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_81),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_90),
.B(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_120),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_69),
.B(n_24),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_24),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_79),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_92),
.A2(n_44),
.B1(n_43),
.B2(n_52),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_92),
.A2(n_43),
.B1(n_48),
.B2(n_56),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_124),
.A2(n_80),
.B1(n_89),
.B2(n_78),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_127),
.B(n_128),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_126),
.B(n_114),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_80),
.B(n_86),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_131),
.A2(n_133),
.B1(n_135),
.B2(n_115),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_89),
.B1(n_78),
.B2(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_134),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_138),
.B1(n_141),
.B2(n_145),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_106),
.A2(n_73),
.B1(n_87),
.B2(n_58),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_106),
.A2(n_103),
.B(n_117),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_148),
.B(n_150),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_40),
.B1(n_76),
.B2(n_28),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_142),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_102),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_144),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_106),
.A2(n_30),
.B1(n_28),
.B2(n_19),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_30),
.B1(n_27),
.B2(n_19),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_146),
.A2(n_147),
.B1(n_110),
.B2(n_120),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_101),
.A2(n_30),
.B1(n_27),
.B2(n_76),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_113),
.A2(n_26),
.B(n_40),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_103),
.A2(n_35),
.B(n_21),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_100),
.C(n_112),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_164),
.C(n_25),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_143),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_154),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_155),
.A2(n_148),
.B1(n_127),
.B2(n_146),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_167),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_100),
.Y(n_158)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_113),
.B1(n_123),
.B2(n_121),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_159),
.A2(n_162),
.B1(n_128),
.B2(n_136),
.Y(n_183)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_35),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_119),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_104),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_166),
.B(n_168),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_139),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_115),
.Y(n_168)
);

NOR3xp33_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_99),
.C(n_118),
.Y(n_172)
);

OAI21xp33_ASAP7_75t_L g199 ( 
.A1(n_172),
.A2(n_23),
.B(n_21),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_142),
.A2(n_99),
.B1(n_105),
.B2(n_107),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_168),
.B(n_175),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_144),
.B(n_122),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_174),
.Y(n_184)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_176),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_176),
.A2(n_133),
.B1(n_135),
.B2(n_137),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_179),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_170),
.A2(n_137),
.B1(n_125),
.B2(n_141),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_162),
.A2(n_128),
.B1(n_138),
.B2(n_148),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_145),
.Y(n_189)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_189),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_173),
.A2(n_99),
.B1(n_150),
.B2(n_147),
.Y(n_190)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_159),
.A2(n_99),
.B1(n_105),
.B2(n_107),
.Y(n_191)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_153),
.B(n_25),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_164),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_165),
.A2(n_153),
.B(n_175),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_194),
.A2(n_197),
.B(n_199),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_196),
.C(n_200),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_161),
.B(n_35),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_170),
.A2(n_105),
.B1(n_111),
.B2(n_102),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_111),
.B1(n_118),
.B2(n_85),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_201),
.A2(n_166),
.B(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_23),
.Y(n_202)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_205),
.B(n_209),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_186),
.A2(n_160),
.B1(n_154),
.B2(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_206),
.A2(n_180),
.B1(n_188),
.B2(n_202),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_185),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_215),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_221),
.B(n_225),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_151),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_155),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_211),
.C(n_212),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_152),
.C(n_156),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_192),
.B(n_156),
.C(n_169),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_194),
.B(n_163),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_218),
.C(n_222),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_178),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_216),
.A2(n_197),
.B1(n_188),
.B2(n_178),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_171),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_169),
.B(n_15),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_183),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_184),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_186),
.A2(n_14),
.B(n_13),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_218),
.B(n_214),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_227),
.B(n_229),
.Y(n_262)
);

AO22x1_ASAP7_75t_L g228 ( 
.A1(n_208),
.A2(n_191),
.B1(n_190),
.B2(n_193),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_209),
.B(n_198),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_217),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_231),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_219),
.A2(n_177),
.B1(n_193),
.B2(n_179),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_242),
.B1(n_223),
.B2(n_204),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_234),
.B(n_235),
.Y(n_258)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_210),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_237),
.B(n_245),
.C(n_247),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_239),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_221),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_243),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_213),
.A2(n_184),
.B(n_189),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_177),
.C(n_180),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_85),
.C(n_23),
.Y(n_247)
);

NAND2xp67_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_213),
.Y(n_248)
);

AOI21x1_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_227),
.B(n_237),
.Y(n_265)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_252),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_245),
.A2(n_222),
.B1(n_220),
.B2(n_212),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_259),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_228),
.A2(n_220),
.B1(n_205),
.B2(n_225),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_255),
.A2(n_3),
.B(n_5),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_240),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_244),
.A2(n_232),
.B(n_239),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_238),
.A2(n_240),
.B1(n_229),
.B2(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_260),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_264),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_265),
.A2(n_262),
.B1(n_12),
.B2(n_7),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_249),
.A2(n_246),
.B1(n_13),
.B2(n_12),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_268),
.A2(n_273),
.B1(n_277),
.B2(n_266),
.Y(n_288)
);

NOR2xp67_ASAP7_75t_SL g269 ( 
.A(n_248),
.B(n_246),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_6),
.B(n_7),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_13),
.Y(n_270)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_270),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_12),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_275),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_253),
.B(n_25),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_278),
.C(n_262),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_11),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_3),
.C(n_5),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_249),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_279),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_274),
.A2(n_261),
.B1(n_257),
.B2(n_258),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_280),
.B(n_283),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_257),
.Y(n_283)
);

OAI221xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_256),
.B1(n_254),
.B2(n_261),
.C(n_263),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_284),
.B(n_286),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_287),
.B(n_288),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_5),
.C(n_6),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_277),
.C(n_7),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_8),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_276),
.B(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_294),
.B(n_298),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_6),
.C(n_8),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_296),
.A2(n_299),
.B(n_282),
.Y(n_303)
);

NOR2xp67_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_281),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_8),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_9),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_301),
.B(n_305),
.Y(n_312)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_280),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_289),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_295),
.B(n_296),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_310),
.B(n_311),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_301),
.C(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_312),
.B(n_294),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_313),
.Y(n_316)
);

O2A1O1Ixp33_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_314),
.B(n_309),
.C(n_10),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_317),
.B(n_9),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_9),
.Y(n_319)
);


endmodule