module fake_jpeg_18212_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx3_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_7),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_13),
.B(n_1),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_6),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_12),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_22),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_28),
.B(n_15),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_31),
.Y(n_37)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_21),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

BUFx24_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_24),
.B1(n_12),
.B2(n_8),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_39),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_43),
.Y(n_47)
);

AO22x1_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_40),
.B1(n_37),
.B2(n_35),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_38),
.A2(n_19),
.B(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_45),
.B(n_9),
.Y(n_46)
);

A2O1A1Ixp33_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_35),
.B(n_9),
.C(n_5),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_48),
.B(n_24),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_49),
.B(n_47),
.C(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_14),
.B(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_4),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_52),
.Y(n_55)
);


endmodule