module fake_jpeg_11127_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_19),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_52),
.Y(n_149)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_22),
.B(n_9),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_54),
.B(n_63),
.Y(n_114)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_24),
.A2(n_29),
.B1(n_36),
.B2(n_47),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_56),
.A2(n_29),
.B1(n_31),
.B2(n_47),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_19),
.Y(n_59)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_9),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_61),
.B(n_64),
.Y(n_111)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_62),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_9),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_65),
.Y(n_158)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_66),
.Y(n_141)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_23),
.B(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_69),
.B(n_95),
.Y(n_131)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_76),
.Y(n_132)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_28),
.Y(n_78)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_79),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_23),
.B(n_8),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_80),
.B(n_89),
.Y(n_151)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_81),
.Y(n_152)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_87),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_26),
.B(n_8),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

CKINVDCx6p67_ASAP7_75t_R g155 ( 
.A(n_92),
.Y(n_155)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g94 ( 
.A(n_31),
.B(n_0),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_SL g139 ( 
.A1(n_94),
.A2(n_44),
.B(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_26),
.B(n_10),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_38),
.B(n_10),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_98),
.B(n_25),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_101),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_29),
.Y(n_103)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_105),
.A2(n_76),
.B1(n_92),
.B2(n_86),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_85),
.A2(n_47),
.B1(n_31),
.B2(n_50),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_107),
.A2(n_117),
.B1(n_120),
.B2(n_145),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_35),
.B1(n_27),
.B2(n_31),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_113),
.A2(n_44),
.B(n_25),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_52),
.A2(n_59),
.B1(n_72),
.B2(n_84),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_38),
.B1(n_35),
.B2(n_31),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_61),
.A2(n_51),
.B1(n_32),
.B2(n_49),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_122),
.A2(n_136),
.B1(n_32),
.B2(n_49),
.Y(n_204)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_138),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_55),
.A2(n_25),
.B1(n_39),
.B2(n_20),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_0),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_50),
.B1(n_21),
.B2(n_33),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_82),
.B(n_39),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_157),
.B(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_160),
.B(n_131),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_73),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_101),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_75),
.B(n_39),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_105),
.A2(n_102),
.B1(n_103),
.B2(n_100),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_164),
.A2(n_167),
.B1(n_181),
.B2(n_209),
.Y(n_264)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_94),
.C(n_60),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_166),
.B(n_169),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_122),
.A2(n_53),
.B1(n_67),
.B2(n_97),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_161),
.Y(n_168)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_168),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_134),
.B(n_94),
.C(n_74),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_171),
.B(n_173),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g172 ( 
.A(n_114),
.B(n_81),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_172),
.B(n_183),
.Y(n_224)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_110),
.Y(n_174)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_174),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_104),
.B(n_96),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_175),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_44),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_178),
.B(n_185),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_180),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_107),
.A2(n_78),
.B1(n_68),
.B2(n_57),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_65),
.B1(n_62),
.B2(n_66),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_32),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_189),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_99),
.B1(n_33),
.B2(n_42),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_190),
.A2(n_198),
.B1(n_200),
.B2(n_203),
.Y(n_225)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_118),
.Y(n_191)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_191),
.Y(n_258)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_126),
.Y(n_192)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_192),
.Y(n_268)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_106),
.Y(n_193)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_193),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_108),
.B(n_93),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_166),
.Y(n_241)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_151),
.A2(n_20),
.B1(n_50),
.B2(n_45),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_149),
.A2(n_21),
.B1(n_33),
.B2(n_42),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

INVx13_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_202),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_129),
.A2(n_21),
.B1(n_42),
.B2(n_45),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_204),
.A2(n_221),
.B1(n_153),
.B2(n_150),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_129),
.A2(n_20),
.B1(n_45),
.B2(n_90),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_205),
.A2(n_210),
.B1(n_130),
.B2(n_133),
.Y(n_250)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_206),
.Y(n_251)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_207),
.Y(n_260)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_146),
.Y(n_208)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_208),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_145),
.A2(n_83),
.B1(n_88),
.B2(n_87),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_140),
.A2(n_91),
.B1(n_49),
.B2(n_79),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_147),
.Y(n_211)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_152),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_217),
.Y(n_236)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_116),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_213),
.Y(n_242)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_116),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_214),
.B(n_188),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_112),
.B(n_0),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_215),
.B(n_218),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_216),
.A2(n_123),
.B1(n_132),
.B2(n_130),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_117),
.B(n_11),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_48),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_222),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_121),
.B(n_0),
.Y(n_220)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_153),
.A3(n_150),
.B1(n_143),
.B2(n_137),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_121),
.A2(n_40),
.B1(n_3),
.B2(n_4),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_144),
.B(n_159),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_229),
.A2(n_238),
.B1(n_248),
.B2(n_255),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_231),
.B(n_252),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_241),
.B(n_165),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_143),
.B1(n_137),
.B2(n_133),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_256),
.B1(n_195),
.B2(n_187),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_201),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_217),
.A2(n_119),
.B1(n_40),
.B2(n_5),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_172),
.A2(n_40),
.B1(n_4),
.B2(n_5),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_164),
.A2(n_40),
.B1(n_4),
.B2(n_6),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_177),
.A2(n_40),
.B1(n_6),
.B2(n_7),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_257),
.A2(n_265),
.B1(n_267),
.B2(n_269),
.Y(n_297)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_173),
.B(n_2),
.C(n_7),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_263),
.B(n_173),
.C(n_175),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_216),
.A2(n_2),
.B1(n_7),
.B2(n_10),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_169),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_199),
.A2(n_185),
.B1(n_215),
.B2(n_220),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_270),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_264),
.A2(n_181),
.B1(n_196),
.B2(n_183),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_274),
.A2(n_276),
.B1(n_288),
.B2(n_300),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_259),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_275),
.B(n_303),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_264),
.A2(n_178),
.B1(n_171),
.B2(n_218),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_294),
.Y(n_326)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_278),
.Y(n_332)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

BUFx5_ASAP7_75t_L g280 ( 
.A(n_251),
.Y(n_280)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_282),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_175),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_283),
.A2(n_287),
.B(n_290),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_284),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_234),
.B(n_247),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_285),
.B(n_289),
.C(n_291),
.Y(n_359)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_232),
.Y(n_286)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_286),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_170),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_269),
.A2(n_247),
.B1(n_253),
.B2(n_225),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_234),
.B(n_180),
.C(n_197),
.Y(n_289)
);

AO22x1_ASAP7_75t_L g290 ( 
.A1(n_231),
.A2(n_211),
.B1(n_208),
.B2(n_207),
.Y(n_290)
);

MAJx2_ASAP7_75t_L g291 ( 
.A(n_237),
.B(n_224),
.C(n_253),
.Y(n_291)
);

AOI22x1_ASAP7_75t_L g292 ( 
.A1(n_238),
.A2(n_272),
.B1(n_265),
.B2(n_237),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_292),
.A2(n_296),
.B(n_305),
.Y(n_330)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_273),
.Y(n_293)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_293),
.Y(n_357)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_295),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_237),
.A2(n_189),
.B(n_191),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_168),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_298),
.B(n_301),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_248),
.A2(n_227),
.B1(n_272),
.B2(n_267),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_299),
.A2(n_273),
.B1(n_233),
.B2(n_223),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_227),
.A2(n_174),
.B1(n_184),
.B2(n_193),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_230),
.B(n_192),
.C(n_212),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_266),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_235),
.B(n_213),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_246),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_230),
.A2(n_214),
.B(n_202),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_239),
.B(n_206),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_307),
.B(n_308),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_240),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_235),
.Y(n_309)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_226),
.B(n_186),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_318),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_271),
.B(n_176),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g347 ( 
.A1(n_311),
.A2(n_315),
.B(n_268),
.Y(n_347)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_244),
.Y(n_312)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_271),
.A2(n_201),
.B1(n_14),
.B2(n_15),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_313),
.A2(n_268),
.B1(n_258),
.B2(n_249),
.Y(n_336)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_262),
.Y(n_314)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_314),
.Y(n_360)
);

A2O1A1O1Ixp25_ASAP7_75t_L g315 ( 
.A1(n_257),
.A2(n_262),
.B(n_251),
.C(n_240),
.D(n_245),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_242),
.B(n_252),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_316),
.B(n_317),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_242),
.B(n_12),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_226),
.B(n_201),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_240),
.B(n_12),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_18),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_306),
.A2(n_244),
.B1(n_232),
.B2(n_245),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_323),
.B1(n_337),
.B2(n_341),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_288),
.B(n_223),
.Y(n_325)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_311),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_327),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_311),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_329),
.B(n_343),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_297),
.A2(n_233),
.B1(n_246),
.B2(n_243),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_297),
.A2(n_299),
.B1(n_281),
.B2(n_274),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_243),
.Y(n_342)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_342),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_300),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_345),
.B(n_298),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_292),
.A2(n_228),
.B(n_258),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_346),
.A2(n_358),
.B(n_296),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g380 ( 
.A(n_347),
.B(n_315),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_304),
.B(n_249),
.Y(n_348)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_301),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_350),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_302),
.A2(n_228),
.B1(n_15),
.B2(n_16),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_351),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_281),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_352),
.A2(n_355),
.B1(n_313),
.B2(n_287),
.Y(n_376)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_353),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_292),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_302),
.A2(n_18),
.B(n_284),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_361),
.B(n_321),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_363),
.A2(n_365),
.B(n_336),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_330),
.A2(n_283),
.B(n_290),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_326),
.B(n_294),
.C(n_289),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_366),
.B(n_370),
.C(n_379),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_356),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g411 ( 
.A(n_367),
.B(n_382),
.Y(n_411)
);

OAI21xp33_ASAP7_75t_SL g368 ( 
.A1(n_330),
.A2(n_290),
.B(n_276),
.Y(n_368)
);

AOI21xp33_ASAP7_75t_L g427 ( 
.A1(n_368),
.A2(n_389),
.B(n_357),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_283),
.C(n_291),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_376),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_375),
.B(n_360),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_277),
.C(n_287),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_380),
.A2(n_347),
.B(n_346),
.Y(n_399)
);

A2O1A1Ixp33_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_320),
.B(n_309),
.C(n_280),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_381),
.B(n_388),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_362),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_321),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_384),
.B(n_392),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_359),
.B(n_312),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_385),
.B(n_386),
.C(n_387),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_335),
.B(n_293),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_286),
.C(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_332),
.Y(n_388)
);

NAND2xp33_ASAP7_75t_SL g389 ( 
.A(n_332),
.B(n_360),
.Y(n_389)
);

INVxp33_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_341),
.A2(n_322),
.B1(n_325),
.B2(n_355),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_391),
.A2(n_395),
.B1(n_396),
.B2(n_358),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_331),
.B(n_342),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_343),
.A2(n_354),
.B1(n_352),
.B2(n_337),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_354),
.A2(n_323),
.B1(n_333),
.B2(n_329),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_334),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_397),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_372),
.A2(n_394),
.B1(n_380),
.B2(n_374),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_398),
.A2(n_401),
.B1(n_412),
.B2(n_421),
.Y(n_435)
);

XNOR2x2_ASAP7_75t_SL g430 ( 
.A(n_399),
.B(n_365),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_333),
.B1(n_327),
.B2(n_348),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_383),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_402),
.B(n_417),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_366),
.B(n_345),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_405),
.B(n_414),
.Y(n_443)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_383),
.B(n_340),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_408),
.B(n_369),
.Y(n_449)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_397),
.Y(n_409)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_373),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_410),
.B(n_364),
.Y(n_452)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_388),
.Y(n_413)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_413),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_386),
.B(n_334),
.Y(n_414)
);

INVx13_ASAP7_75t_L g416 ( 
.A(n_393),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_416),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_391),
.A2(n_338),
.B1(n_339),
.B2(n_340),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_338),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_418),
.B(n_428),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_385),
.B(n_339),
.C(n_344),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_419),
.B(n_393),
.C(n_377),
.Y(n_432)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_374),
.Y(n_420)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_394),
.A2(n_344),
.B1(n_328),
.B2(n_349),
.Y(n_421)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_424),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_380),
.A2(n_328),
.B1(n_349),
.B2(n_357),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_426),
.A2(n_424),
.B1(n_421),
.B2(n_398),
.Y(n_453)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_427),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_387),
.B(n_375),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_405),
.B(n_379),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_430),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_432),
.B(n_440),
.C(n_450),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_418),
.B(n_377),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_433),
.B(n_441),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_378),
.C(n_371),
.Y(n_440)
);

MAJx2_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_378),
.C(n_381),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_402),
.B(n_396),
.Y(n_442)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_442),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_407),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_445),
.B(n_423),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_449),
.B(n_408),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_369),
.C(n_363),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_403),
.B(n_376),
.C(n_364),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_403),
.C(n_419),
.Y(n_463)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_453),
.A2(n_400),
.B1(n_409),
.B2(n_416),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_407),
.B(n_417),
.Y(n_454)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_454),
.Y(n_472)
);

A2O1A1Ixp33_ASAP7_75t_SL g455 ( 
.A1(n_430),
.A2(n_412),
.B(n_399),
.C(n_423),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_455),
.B(n_435),
.C(n_449),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_439),
.A2(n_422),
.B1(n_425),
.B2(n_411),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_457),
.A2(n_461),
.B1(n_466),
.B2(n_435),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_458),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_439),
.A2(n_422),
.B1(n_401),
.B2(n_420),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_462),
.B(n_444),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_469),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_437),
.Y(n_465)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_465),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_447),
.A2(n_426),
.B1(n_406),
.B2(n_413),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_438),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_468),
.B(n_470),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_429),
.B(n_414),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_448),
.B(n_404),
.C(n_400),
.Y(n_470)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_471),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_434),
.Y(n_473)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_473),
.Y(n_489)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_431),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_474),
.B(n_475),
.Y(n_484)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_446),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_478),
.A2(n_461),
.B1(n_491),
.B2(n_466),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_443),
.Y(n_481)
);

XNOR2x1_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_486),
.Y(n_498)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_482),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_463),
.B(n_448),
.C(n_440),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_485),
.B(n_488),
.Y(n_503)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_464),
.B(n_443),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_464),
.B(n_450),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_487),
.B(n_491),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_451),
.C(n_432),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_441),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_456),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_470),
.B(n_433),
.C(n_436),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_492),
.B(n_462),
.Y(n_504)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_477),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_494),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_480),
.A2(n_444),
.B(n_436),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_476),
.A2(n_467),
.B1(n_472),
.B2(n_471),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_500),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_499),
.B(n_504),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_489),
.A2(n_442),
.B1(n_459),
.B2(n_483),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_473),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_501),
.B(n_502),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_478),
.B(n_454),
.Y(n_502)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_487),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_506),
.B(n_479),
.Y(n_511)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_507),
.Y(n_520)
);

BUFx24_ASAP7_75t_SL g509 ( 
.A(n_503),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_509),
.B(n_497),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_511),
.B(n_481),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_495),
.B(n_488),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_512),
.B(n_515),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_SL g513 ( 
.A(n_502),
.B(n_485),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_513),
.A2(n_499),
.B(n_494),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_493),
.B(n_465),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_514),
.B(n_501),
.Y(n_518)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_518),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_519),
.B(n_521),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_522),
.A2(n_523),
.B(n_514),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_508),
.B(n_498),
.C(n_486),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_517),
.B(n_520),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g527 ( 
.A1(n_518),
.A2(n_516),
.B1(n_510),
.B2(n_455),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g529 ( 
.A1(n_527),
.A2(n_455),
.B(n_456),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_529),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_525),
.B(n_524),
.Y(n_531)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_531),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_498),
.C(n_455),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_492),
.Y(n_534)
);


endmodule