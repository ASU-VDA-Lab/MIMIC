module real_jpeg_1683_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_1),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_105),
.Y(n_104)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_2),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_3),
.A2(n_29),
.B1(n_31),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_3),
.A2(n_34),
.B1(n_42),
.B2(n_45),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_34),
.B1(n_58),
.B2(n_59),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_3),
.B(n_42),
.C(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_34),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_53),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_3),
.B(n_29),
.C(n_39),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_3),
.B(n_73),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_21),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_3),
.B(n_22),
.C(n_24),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_37),
.Y(n_149)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_5),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_5),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_44),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_5),
.A2(n_29),
.B1(n_31),
.B2(n_44),
.Y(n_101)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g12 ( 
.A1(n_13),
.A2(n_109),
.B1(n_167),
.B2(n_168),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_13),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_108),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_86),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_15),
.B(n_86),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_67),
.C(n_77),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_16),
.B(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_51),
.B2(n_66),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_35),
.B1(n_36),
.B2(n_50),
.Y(n_18)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_19),
.B(n_36),
.C(n_66),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_32),
.B(n_33),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_20),
.A2(n_32),
.B1(n_33),
.B2(n_101),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_20),
.A2(n_32),
.B1(n_33),
.B2(n_101),
.Y(n_119)
);

OR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

AO22x1_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_21)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g28 ( 
.A1(n_22),
.A2(n_27),
.B1(n_29),
.B2(n_31),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_23),
.B(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_24),
.B(n_135),
.Y(n_134)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

AOI22x1_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_29),
.B(n_142),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_35),
.A2(n_36),
.B1(n_99),
.B2(n_100),
.Y(n_157)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_36),
.B(n_99),
.C(n_158),
.Y(n_164)
);

AO21x1_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B(n_46),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_37),
.A2(n_41),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_39),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_45),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_42),
.Y(n_45)
);

AO22x1_ASAP7_75t_SL g53 ( 
.A1(n_42),
.A2(n_45),
.B1(n_54),
.B2(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_42),
.B(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

OA21x2_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_57),
.B(n_62),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

O2A1O1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_54),
.B(n_58),
.C(n_65),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_63),
.B1(n_64),
.B2(n_93),
.Y(n_92)
);

INVx4_ASAP7_75t_SL g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_58),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_69),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_77),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_76),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_76),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_70),
.A2(n_71),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_71),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_71),
.B(n_137),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_71),
.B(n_119),
.C(n_149),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_75),
.B(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.C(n_82),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_78),
.A2(n_91),
.B1(n_92),
.B2(n_94),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_78),
.A2(n_94),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_81),
.A2(n_82),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_82),
.B(n_134),
.Y(n_133)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B(n_85),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_85),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_83),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_95),
.B2(n_96),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_SL g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_106),
.B2(n_107),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_99),
.A2(n_100),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_143),
.Y(n_152)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

OAI21x1_ASAP7_75t_SL g109 ( 
.A1(n_110),
.A2(n_128),
.B(n_166),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_113),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_111),
.B(n_113),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_119),
.C(n_120),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_114),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

NOR2xp67_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_140),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_119),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_148)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_119),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_119),
.A2(n_120),
.B1(n_150),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_120),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_124),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_121),
.A2(n_122),
.B1(n_124),
.B2(n_125),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_160),
.B(n_165),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_154),
.B(n_159),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_145),
.B(n_153),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_139),
.B(n_144),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_136),
.B(n_138),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_141),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_152),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_146),
.B(n_152),
.Y(n_153)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_156),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_164),
.Y(n_165)
);


endmodule