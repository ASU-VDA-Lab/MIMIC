module fake_jpeg_20963_n_67 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_67);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_67;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_48;
wire n_35;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_24;
wire n_38;
wire n_26;
wire n_28;
wire n_36;
wire n_62;
wire n_25;
wire n_56;
wire n_31;
wire n_43;
wire n_37;
wire n_29;
wire n_50;
wire n_32;
wire n_66;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_20),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_0),
.B(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_3),
.Y(n_30)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_1),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_52)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_35),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_23),
.B(n_41),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_42),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_49),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_53),
.B1(n_41),
.B2(n_33),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_57),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_24),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_36),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_26),
.B(n_34),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_30),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_61),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_64),
.A2(n_29),
.B1(n_50),
.B2(n_31),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_65),
.A2(n_28),
.B1(n_50),
.B2(n_40),
.Y(n_66)
);

BUFx24_ASAP7_75t_SL g67 ( 
.A(n_66),
.Y(n_67)
);


endmodule