module real_jpeg_26252_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_1),
.A2(n_40),
.B1(n_42),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_47),
.B1(n_54),
.B2(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_1),
.A2(n_22),
.B1(n_25),
.B2(n_47),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_47),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_2),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_2),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_40),
.B1(n_42),
.B2(n_141),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_2),
.A2(n_22),
.B1(n_25),
.B2(n_141),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_2),
.A2(n_27),
.B1(n_28),
.B2(n_141),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_4),
.A2(n_22),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_32),
.B1(n_40),
.B2(n_42),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_4),
.A2(n_32),
.B1(n_54),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_32),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_4),
.A2(n_57),
.B(n_142),
.C(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_4),
.B(n_55),
.Y(n_220)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_4),
.A2(n_36),
.B(n_42),
.C(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_4),
.B(n_24),
.C(n_27),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_4),
.B(n_85),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_4),
.B(n_11),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_4),
.B(n_26),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_7),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_52),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_7),
.A2(n_22),
.B1(n_25),
.B2(n_52),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_52),
.Y(n_167)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_11),
.Y(n_105)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_11),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_78),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_76),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_71),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_15),
.B(n_71),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_65),
.C(n_66),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_16),
.A2(n_17),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_33),
.C(n_48),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_18),
.A2(n_95),
.B1(n_96),
.B2(n_99),
.Y(n_94)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_18),
.A2(n_33),
.B1(n_99),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_18),
.A2(n_99),
.B1(n_189),
.B2(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_29),
.B(n_30),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_19),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_20),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_20),
.B(n_31),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_20),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_26),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_25),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_22),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_23),
.A2(n_24),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_25),
.A2(n_32),
.B(n_37),
.Y(n_231)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_26),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_26),
.B(n_235),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_27),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_27),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_27),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_29),
.B(n_30),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_29),
.A2(n_89),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g205 ( 
.A1(n_32),
.A2(n_42),
.B(n_56),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_33),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_43),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_34),
.B(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_45),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_35),
.A2(n_38),
.B(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_35),
.B(n_46),
.Y(n_98)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_36),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_40),
.B2(n_42),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_39),
.B(n_97),
.Y(n_135)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_43),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_43),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_44),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_48),
.B(n_149),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_55),
.B(n_58),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_49),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_50),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_61)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_51),
.Y(n_140)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_55),
.B(n_139),
.Y(n_175)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_72),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_59),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_62),
.Y(n_59)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_60),
.B(n_74),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_139),
.Y(n_138)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_65),
.B(n_164),
.C(n_174),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_65),
.A2(n_174),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_65),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_306),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_68),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_70),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_70),
.B(n_138),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_319),
.B(n_324),
.Y(n_78)
);

OAI211xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_143),
.B(n_153),
.C(n_318),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_118),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_81),
.B(n_118),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_81),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_91),
.CI(n_102),
.CON(n_81),
.SN(n_81)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_82),
.A2(n_83),
.B(n_86),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_91),
.C(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_85),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_87),
.B(n_233),
.Y(n_232)
);

INVxp33_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_89),
.B(n_245),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_94),
.B1(n_100),
.B2(n_101),
.Y(n_91)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_92),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_92),
.A2(n_100),
.B1(n_148),
.B2(n_151),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_96),
.C(n_99),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_92),
.B(n_148),
.C(n_152),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_93),
.B(n_175),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_98),
.B(n_198),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_99),
.B(n_187),
.C(n_189),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_110),
.B(n_114),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_114),
.B1(n_115),
.B2(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_103),
.A2(n_111),
.B1(n_122),
.B2(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_103),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_103),
.A2(n_122),
.B1(n_230),
.B2(n_289),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_106),
.B(n_109),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_104),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_104),
.B(n_109),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_104),
.B(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_108),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_111),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_113),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_113),
.B(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_123),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_124),
.B(n_177),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.C(n_136),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_126),
.B(n_132),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_127),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_130),
.A2(n_167),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_130),
.B(n_265),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_131),
.B(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_133),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_135),
.B(n_191),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_140),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

NAND3xp33_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_154),
.C(n_155),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_145),
.B(n_146),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.Y(n_146)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_148),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_179),
.B(n_317),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_176),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_157),
.B(n_176),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_163),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_158),
.B(n_161),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_163),
.B(n_315),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_164),
.A2(n_165),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_172),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_172),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_169),
.B(n_258),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_173),
.B(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_174),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_312),
.B(n_316),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_223),
.B(n_298),
.C(n_311),
.Y(n_180)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_211),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_182),
.B(n_211),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_184),
.B1(n_195),
.B2(n_210),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_193),
.B2(n_194),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_185),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_185),
.B(n_194),
.C(n_210),
.Y(n_299)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_186),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_188),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_192),
.Y(n_199)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_203),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_196)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_197),
.B(n_202),
.C(n_203),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_206),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_206),
.Y(n_217)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.C(n_218),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_212),
.A2(n_213),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.C(n_221),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_220),
.B(n_221),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_222),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_297),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_239),
.B(n_296),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_236),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_226),
.B(n_236),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.C(n_232),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_227),
.B(n_294),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_229),
.B(n_232),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_230),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_291),
.B(n_295),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_282),
.B(n_290),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_262),
.B(n_281),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_249),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_243),
.B(n_249),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_244),
.A2(n_246),
.B1(n_247),
.B2(n_269),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_256),
.B2(n_261),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_255),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_252),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_252),
.B(n_255),
.C(n_261),
.Y(n_283)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_253),
.Y(n_255)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_256),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_260),
.B(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_270),
.B(n_280),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_268),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_276),
.B(n_279),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_283),
.B(n_284),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_288),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_287),
.C(n_288),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_299),
.B(n_300),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_310),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_308),
.B2(n_309),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_309),
.C(n_310),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_313),
.B(n_314),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_323),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_320),
.B(n_323),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_321),
.Y(n_322)
);


endmodule