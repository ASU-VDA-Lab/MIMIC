module real_jpeg_16520_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_1),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_1),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_1),
.B(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_1),
.B(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_1),
.B(n_152),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_1),
.B(n_314),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_1),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_3),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_4),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_4),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_4),
.B(n_137),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_4),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_4),
.B(n_107),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_4),
.B(n_217),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_5),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_5),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_5),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_6),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_6),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_6),
.B(n_28),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_7),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

NAND2x1_ASAP7_75t_SL g49 ( 
.A(n_8),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_8),
.B(n_95),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_8),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_8),
.B(n_251),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_8),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_8),
.B(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_9),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_9),
.Y(n_157)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_10),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_10),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_10),
.Y(n_219)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_11),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_11),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_12),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_12),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g186 ( 
.A(n_12),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_12),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_12),
.B(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_14),
.Y(n_131)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_14),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_14),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_14),
.B(n_71),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_14),
.B(n_234),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_15),
.Y(n_127)
);

BUFx4f_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_15),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_27),
.Y(n_26)
);

NAND2x2_ASAP7_75t_SL g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_16),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_16),
.B(n_107),
.Y(n_106)
);

AND2x4_ASAP7_75t_SL g197 ( 
.A(n_16),
.B(n_198),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_16),
.B(n_137),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_16),
.B(n_340),
.Y(n_339)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_17),
.Y(n_170)
);

BUFx12f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_116),
.B(n_339),
.C(n_407),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_39),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_24),
.A2(n_25),
.B1(n_62),
.B2(n_74),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_26),
.A2(n_30),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_26),
.B(n_54),
.C(n_58),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_26),
.A2(n_46),
.B1(n_58),
.B2(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_26),
.A2(n_46),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_26),
.B(n_155),
.C(n_160),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_29),
.Y(n_133)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_30),
.A2(n_70),
.B(n_73),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_30),
.B(n_70),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_30),
.A2(n_47),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g296 ( 
.A(n_30),
.B(n_247),
.C(n_250),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_33),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_33),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_33),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

INVxp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_34),
.B(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_75),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_40),
.B(n_75),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_61),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_48),
.C(n_53),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_43),
.B(n_155),
.C(n_361),
.Y(n_372)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_49),
.B1(n_53),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_54),
.B(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_57),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_106),
.C(n_110),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_58),
.Y(n_115)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_58),
.B(n_168),
.C(n_171),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_58),
.A2(n_106),
.B1(n_115),
.B2(n_272),
.Y(n_370)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_60),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_59),
.Y(n_283)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_63),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_63),
.A2(n_64),
.B1(n_378),
.B2(n_379),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_81),
.C(n_88),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_64),
.B(n_73),
.Y(n_407)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g211 ( 
.A(n_66),
.Y(n_211)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_66),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_70),
.B(n_305),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_70),
.B(n_197),
.C(n_307),
.Y(n_342)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_72),
.Y(n_129)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_72),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.C(n_101),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_76),
.B(n_79),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_93),
.C(n_97),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_103),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_82),
.B(n_88),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_84),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_83),
.B(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_86),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_88),
.A2(n_89),
.B1(n_241),
.B2(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_88),
.B(n_239),
.C(n_241),
.Y(n_301)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_91),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_92),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_94),
.B1(n_97),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_96),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_97),
.A2(n_104),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_97),
.A2(n_104),
.B1(n_339),
.B2(n_341),
.Y(n_338)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_100),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_100),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_101),
.B(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.C(n_113),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_102),
.B(n_367),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_104),
.B(n_300),
.C(n_301),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_104),
.B(n_339),
.C(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_105),
.B(n_113),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_147),
.C(n_149),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_106),
.A2(n_147),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_106),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_106),
.A2(n_272),
.B1(n_306),
.B2(n_307),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_SL g371 ( 
.A(n_106),
.B(n_307),
.C(n_346),
.Y(n_371)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_110),
.B(n_370),
.Y(n_369)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_115),
.B(n_184),
.Y(n_183)
);

O2A1O1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_363),
.B(n_401),
.C(n_406),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_286),
.B(n_324),
.C(n_325),
.D(n_362),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_257),
.B(n_285),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_224),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_120),
.B(n_224),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_181),
.C(n_208),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_121),
.B(n_259),
.Y(n_258)
);

XOR2x2_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_153),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_122),
.B(n_154),
.C(n_166),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_134),
.C(n_146),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_123),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

MAJx3_ASAP7_75t_L g223 ( 
.A(n_125),
.B(n_128),
.C(n_130),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_134),
.A2(n_135),
.B1(n_146),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_136),
.B(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_136),
.A2(n_197),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_136),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_136),
.A2(n_139),
.B1(n_140),
.B2(n_236),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g310 ( 
.A1(n_136),
.A2(n_197),
.B(n_231),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_146),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_147),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_149),
.B(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_151),
.Y(n_317)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_166),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_158),
.B1(n_159),
.B2(n_165),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_155),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_155),
.A2(n_165),
.B1(n_357),
.B2(n_361),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_172),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_167),
.B(n_173),
.C(n_178),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_168),
.B(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_171),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_171),
.B(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_178),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_181),
.B(n_208),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_194),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_182),
.B(n_185),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_184),
.B(n_316),
.C(n_318),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_193),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_190),
.Y(n_193)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_193),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_194),
.B(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.C(n_203),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_196),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_197),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_197),
.A2(n_237),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_220),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_209),
.B(n_221),
.C(n_223),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_210),
.B(n_213),
.C(n_216),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_225),
.B(n_227),
.C(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_243),
.Y(n_226)
);

XOR2x2_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_229),
.B(n_230),
.C(n_238),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_241),
.Y(n_242)
);

INVxp33_ASAP7_75t_L g323 ( 
.A(n_243),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

INVxp33_ASAP7_75t_SL g290 ( 
.A(n_244),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_245)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_246),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_254),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_255),
.C(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.C(n_268),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.C(n_274),
.Y(n_268)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.C(n_284),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_279),
.Y(n_278)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_322),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_322),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_291),
.Y(n_288)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_289),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_303),
.B1(n_320),
.B2(n_321),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_295),
.C(n_302),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_302),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_297),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_301),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_303),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_303),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_309),
.C(n_311),
.Y(n_334)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_306),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_316),
.B1(n_318),
.B2(n_319),
.Y(n_312)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_313),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_316),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_328),
.C(n_329),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_330),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_330),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_331),
.B(n_333),
.C(n_343),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_343),
.Y(n_332)
);

XOR2x1_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_334),
.B(n_336),
.C(n_337),
.Y(n_395)
);

XNOR2x1_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

XNOR2x1_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_342),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_339),
.Y(n_341)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

XNOR2x2_ASAP7_75t_SL g343 ( 
.A(n_344),
.B(n_353),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_344),
.B(n_354),
.C(n_355),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_352),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_357),
.Y(n_361)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_SL g363 ( 
.A(n_364),
.B(n_384),
.C(n_396),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_364),
.A2(n_402),
.B(n_405),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_382),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_365),
.B(n_382),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_368),
.C(n_373),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_366),
.B(n_368),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.C(n_372),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_369),
.B(n_390),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_372),
.Y(n_390)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_399),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.C(n_380),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_375),
.B(n_393),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_376),
.A2(n_377),
.B1(n_380),
.B2(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_385),
.B(n_386),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_395),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_391),
.B2(n_392),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_389),
.B(n_391),
.C(n_395),
.Y(n_400)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_397),
.A2(n_403),
.B(n_404),
.Y(n_402)
);

NOR2x1_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_400),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_400),
.Y(n_404)
);


endmodule