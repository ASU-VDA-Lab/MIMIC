module fake_jpeg_11638_n_526 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_526);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_526;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx8_ASAP7_75t_SL g39 ( 
.A(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_27),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_52),
.B(n_62),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_58),
.B(n_74),
.Y(n_106)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_18),
.B(n_15),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_63),
.Y(n_122)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_68),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_14),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_69),
.B(n_96),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_0),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_86),
.Y(n_120)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_80),
.Y(n_130)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_81),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_82),
.Y(n_157)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_44),
.Y(n_83)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_30),
.B(n_0),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_87),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_31),
.Y(n_110)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_92),
.Y(n_152)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_21),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_93),
.B(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_39),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_97),
.Y(n_142)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_28),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g153 ( 
.A(n_99),
.Y(n_153)
);

INVx4_ASAP7_75t_SL g100 ( 
.A(n_47),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_100),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_58),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_103),
.B(n_104),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_74),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_89),
.A2(n_50),
.B1(n_30),
.B2(n_31),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_105),
.A2(n_135),
.B1(n_61),
.B2(n_42),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_53),
.A2(n_50),
.B1(n_48),
.B2(n_46),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_109),
.A2(n_20),
.B1(n_40),
.B2(n_36),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_110),
.B(n_22),
.Y(n_204)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_40),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_114),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_100),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_67),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_126),
.B(n_145),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_78),
.A2(n_37),
.B1(n_50),
.B2(n_22),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_133),
.A2(n_42),
.B1(n_22),
.B2(n_19),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_54),
.A2(n_43),
.B1(n_41),
.B2(n_37),
.Y(n_135)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx3_ASAP7_75t_SL g163 ( 
.A(n_140),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_67),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_88),
.B(n_41),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_149),
.B(n_151),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_88),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_42),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_91),
.B(n_43),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_56),
.B(n_48),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_160),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_56),
.B(n_46),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_161),
.A2(n_182),
.B1(n_185),
.B2(n_159),
.Y(n_241)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_158),
.B(n_112),
.C(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_174),
.Y(n_211)
);

AO22x2_ASAP7_75t_L g164 ( 
.A1(n_152),
.A2(n_98),
.B1(n_92),
.B2(n_87),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_SL g215 ( 
.A(n_164),
.B(n_165),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_154),
.Y(n_165)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_108),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_166),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_142),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_167),
.B(n_203),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_170),
.Y(n_247)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_171),
.Y(n_224)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_120),
.Y(n_174)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_125),
.Y(n_180)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_133),
.A2(n_85),
.B1(n_82),
.B2(n_73),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_143),
.A2(n_35),
.B(n_33),
.Y(n_183)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_183),
.B(n_140),
.C(n_137),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_102),
.B(n_35),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_184),
.B(n_187),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_109),
.A2(n_72),
.B1(n_63),
.B2(n_55),
.Y(n_185)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_124),
.B(n_36),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_130),
.B(n_42),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_188),
.B(n_202),
.Y(n_226)
);

BUFx16f_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_190),
.Y(n_243)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_192),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_141),
.B(n_1),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_193),
.B(n_197),
.Y(n_227)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_146),
.Y(n_196)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_196),
.Y(n_238)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_198),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_101),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_199),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_200),
.A2(n_209),
.B1(n_210),
.B2(n_117),
.Y(n_249)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_128),
.B(n_22),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_128),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_206),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_19),
.B1(n_16),
.B2(n_3),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_159),
.B1(n_116),
.B2(n_117),
.Y(n_245)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_138),
.Y(n_207)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_208),
.B(n_116),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_107),
.A2(n_19),
.B1(n_16),
.B2(n_3),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_101),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_185),
.A2(n_148),
.B1(n_157),
.B2(n_121),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_214),
.A2(n_218),
.B1(n_241),
.B2(n_197),
.Y(n_263)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_166),
.Y(n_217)
);

INVx3_ASAP7_75t_SL g257 ( 
.A(n_217),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_164),
.A2(n_148),
.B1(n_157),
.B2(n_121),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_231),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_227),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_173),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_245),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_169),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_132),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_190),
.B(n_191),
.Y(n_277)
);

INVx8_ASAP7_75t_L g251 ( 
.A(n_234),
.Y(n_251)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_253),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_177),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_254),
.A2(n_260),
.B(n_255),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_212),
.B(n_168),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_255),
.B(n_268),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_216),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_256),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_204),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_258),
.B(n_260),
.C(n_261),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_259),
.B(n_269),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_162),
.C(n_119),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_115),
.C(n_129),
.Y(n_261)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_118),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_221),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_264),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_265),
.B(n_245),
.Y(n_288)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_230),
.Y(n_266)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_222),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_180),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_213),
.B(n_175),
.Y(n_271)
);

INVxp33_ASAP7_75t_L g317 ( 
.A(n_271),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_241),
.A2(n_200),
.B1(n_164),
.B2(n_209),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_215),
.B(n_164),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_274),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_236),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_236),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_276),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_277),
.A2(n_280),
.B(n_283),
.Y(n_310)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_237),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_215),
.A2(n_210),
.B(n_113),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_281),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g283 ( 
.A(n_243),
.B(n_153),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_213),
.B(n_179),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_254),
.A2(n_233),
.B1(n_217),
.B2(n_201),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_287),
.A2(n_292),
.B1(n_293),
.B2(n_297),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_288),
.B(n_228),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_254),
.A2(n_195),
.B1(n_181),
.B2(n_196),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_219),
.B1(n_216),
.B2(n_223),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_295),
.B(n_266),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_282),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_298),
.A2(n_301),
.B(n_277),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_242),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_258),
.C(n_261),
.Y(n_322)
);

AO22x1_ASAP7_75t_L g301 ( 
.A1(n_252),
.A2(n_242),
.B1(n_229),
.B2(n_238),
.Y(n_301)
);

OAI32xp33_ASAP7_75t_L g303 ( 
.A1(n_250),
.A2(n_283),
.A3(n_252),
.B1(n_272),
.B2(n_267),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_303),
.B(n_243),
.Y(n_345)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_270),
.Y(n_308)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_264),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_318),
.Y(n_323)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_316),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_274),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_321),
.B(n_310),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_332),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_291),
.B(n_259),
.Y(n_324)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_324),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_320),
.A2(n_257),
.B1(n_251),
.B2(n_276),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_326),
.A2(n_343),
.B(n_353),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_311),
.B(n_247),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_329),
.B(n_340),
.Y(n_370)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_L g331 ( 
.A1(n_290),
.A2(n_263),
.B1(n_256),
.B2(n_278),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_331),
.A2(n_335),
.B1(n_299),
.B2(n_294),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_285),
.C(n_281),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_291),
.B(n_275),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_333),
.B(n_309),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_290),
.A2(n_303),
.B1(n_288),
.B2(n_297),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_228),
.C(n_224),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_336),
.B(n_346),
.Y(n_364)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_286),
.Y(n_337)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_337),
.Y(n_361)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_286),
.Y(n_338)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_339),
.B(n_347),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_307),
.B(n_317),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_302),
.Y(n_341)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_296),
.B(n_247),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_342),
.B(n_344),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_298),
.A2(n_262),
.B(n_253),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_295),
.B(n_229),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_305),
.B(n_234),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_297),
.A2(n_257),
.B1(n_256),
.B2(n_223),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_348),
.A2(n_349),
.B1(n_355),
.B2(n_163),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_298),
.A2(n_257),
.B1(n_219),
.B2(n_224),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_302),
.Y(n_350)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_350),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_309),
.B(n_192),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_319),
.Y(n_369)
);

INVx13_ASAP7_75t_L g352 ( 
.A(n_320),
.Y(n_352)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_352),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_310),
.A2(n_238),
.B(n_165),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_304),
.Y(n_354)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_354),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_300),
.A2(n_122),
.B1(n_131),
.B2(n_134),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_323),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_387),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_357),
.A2(n_377),
.B1(n_379),
.B2(n_331),
.Y(n_397)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_360),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_365),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_324),
.B(n_304),
.Y(n_366)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_306),
.Y(n_367)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_367),
.Y(n_400)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

AO21x2_ASAP7_75t_L g373 ( 
.A1(n_345),
.A2(n_301),
.B(n_316),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_373),
.A2(n_380),
.B1(n_163),
.B2(n_134),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_315),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_374),
.B(n_378),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_328),
.A2(n_306),
.B1(n_308),
.B2(n_301),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_344),
.B(n_332),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_328),
.A2(n_319),
.B1(n_299),
.B2(n_294),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_336),
.B(n_289),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_382),
.B(n_107),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_325),
.B(n_289),
.Y(n_383)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_383),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_325),
.B(n_312),
.Y(n_385)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_343),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_334),
.B(n_207),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_388),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_322),
.C(n_346),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_394),
.C(n_398),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_335),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_391),
.B(n_412),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_389),
.B(n_353),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_393),
.B(n_401),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_365),
.C(n_376),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_365),
.A2(n_321),
.B(n_349),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_396),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_373),
.B1(n_372),
.B2(n_371),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_366),
.B(n_355),
.C(n_354),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_360),
.B(n_338),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_330),
.Y(n_402)
);

CKINVDCx14_ASAP7_75t_R g422 ( 
.A(n_402),
.Y(n_422)
);

XNOR2x1_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_348),
.Y(n_403)
);

XNOR2x1_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_414),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_368),
.B(n_350),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_383),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_379),
.B(n_341),
.C(n_337),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_361),
.C(n_384),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_334),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_410),
.B(n_411),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_352),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_381),
.A2(n_352),
.B(n_327),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_413),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_377),
.B(n_199),
.Y(n_414)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_415),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_359),
.Y(n_416)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_416),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_367),
.B(n_189),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_417),
.B(n_388),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_404),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_421),
.B(n_441),
.Y(n_451)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_400),
.Y(n_426)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_426),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_357),
.B1(n_362),
.B2(n_384),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_432),
.Y(n_456)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_401),
.Y(n_429)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_436),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_390),
.B(n_373),
.Y(n_432)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_433),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_434),
.B(n_438),
.C(n_440),
.Y(n_447)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_437),
.A2(n_414),
.B1(n_417),
.B2(n_403),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_393),
.B(n_394),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_361),
.C(n_372),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_358),
.Y(n_441)
);

FAx1_ASAP7_75t_SL g442 ( 
.A(n_408),
.B(n_373),
.CI(n_385),
.CON(n_442),
.SN(n_442)
);

NOR2xp33_ASAP7_75t_SL g460 ( 
.A(n_442),
.B(n_414),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_439),
.A2(n_408),
.B(n_414),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_444),
.A2(n_450),
.B(n_172),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_439),
.A2(n_373),
.B1(n_399),
.B2(n_431),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_448),
.A2(n_453),
.B1(n_435),
.B2(n_420),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_443),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_455),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_432),
.A2(n_411),
.B(n_402),
.Y(n_450)
);

BUFx12f_ASAP7_75t_SL g452 ( 
.A(n_435),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g480 ( 
.A(n_452),
.B(n_153),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_440),
.A2(n_398),
.B1(n_406),
.B2(n_418),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_430),
.B(n_419),
.Y(n_454)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_454),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_434),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_409),
.Y(n_457)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_457),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_458),
.A2(n_420),
.B1(n_427),
.B2(n_358),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_460),
.A2(n_363),
.B1(n_113),
.B2(n_170),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_425),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_445),
.B1(n_454),
.B2(n_459),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_371),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_463),
.B(n_423),
.Y(n_469)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_464),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_447),
.B(n_424),
.C(n_427),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_466),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_424),
.C(n_455),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_474),
.Y(n_488)
);

CKINVDCx14_ASAP7_75t_R g490 ( 
.A(n_469),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_359),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_470),
.B(n_471),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_363),
.C(n_362),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_462),
.Y(n_493)
);

INVx11_ASAP7_75t_L g473 ( 
.A(n_449),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_473),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_444),
.A2(n_171),
.B(n_208),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_475),
.A2(n_480),
.B(n_450),
.Y(n_487)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_476),
.B(n_446),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_463),
.A2(n_131),
.B1(n_122),
.B2(n_136),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_478),
.B(n_448),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_479),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_466),
.B(n_453),
.C(n_456),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_486),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_476),
.A2(n_461),
.B1(n_458),
.B2(n_445),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_485),
.A2(n_495),
.B1(n_136),
.B2(n_153),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_487),
.B(n_492),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_481),
.A2(n_460),
.B(n_459),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_491),
.A2(n_478),
.B(n_189),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_493),
.B(n_488),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_468),
.A2(n_446),
.B1(n_462),
.B2(n_452),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_483),
.B(n_465),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_499),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_484),
.A2(n_481),
.B1(n_468),
.B2(n_473),
.Y(n_498)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_482),
.B(n_471),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_490),
.B(n_477),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_500),
.A2(n_501),
.B1(n_505),
.B2(n_508),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_494),
.A2(n_467),
.B1(n_464),
.B2(n_474),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_504),
.A2(n_507),
.B1(n_1),
.B2(n_2),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_491),
.A2(n_472),
.B(n_475),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_495),
.C(n_493),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_489),
.C(n_496),
.Y(n_509)
);

AOI21x1_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_501),
.B(n_4),
.Y(n_517)
);

AOI322xp5_ASAP7_75t_L g512 ( 
.A1(n_502),
.A2(n_487),
.A3(n_19),
.B1(n_16),
.B2(n_6),
.C1(n_7),
.C2(n_10),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_512),
.A2(n_514),
.B1(n_16),
.B2(n_11),
.Y(n_519)
);

OAI31xp33_ASAP7_75t_L g515 ( 
.A1(n_503),
.A2(n_1),
.A3(n_2),
.B(n_4),
.Y(n_515)
);

NAND3xp33_ASAP7_75t_SL g518 ( 
.A(n_515),
.B(n_2),
.C(n_6),
.Y(n_518)
);

AOI21xp33_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_507),
.B(n_506),
.Y(n_516)
);

AOI322xp5_ASAP7_75t_L g520 ( 
.A1(n_516),
.A2(n_518),
.A3(n_519),
.B1(n_513),
.B2(n_511),
.C1(n_514),
.C2(n_12),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_509),
.C(n_12),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_520),
.A2(n_521),
.B(n_6),
.Y(n_522)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_522),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g524 ( 
.A(n_523),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_12),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_525),
.A2(n_12),
.B(n_14),
.Y(n_526)
);


endmodule