module fake_jpeg_13206_n_386 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_386);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_386;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_42),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_43),
.B(n_51),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_14),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_46),
.Y(n_80)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_14),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_R g50 ( 
.A(n_25),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_50),
.B(n_41),
.CON(n_105),
.SN(n_105)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_29),
.B(n_11),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_29),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_11),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_63),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_25),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_29),
.B(n_0),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_58),
.Y(n_123)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_59),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_62),
.B(n_20),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_10),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_70),
.Y(n_118)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_71),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_20),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_33),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_74),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_65),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_82),
.B(n_92),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_48),
.A2(n_23),
.B1(n_35),
.B2(n_27),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_86),
.A2(n_87),
.B1(n_101),
.B2(n_103),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_23),
.B1(n_35),
.B2(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_43),
.B(n_23),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_52),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_93),
.B(n_109),
.Y(n_143)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_96),
.B(n_107),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_56),
.A2(n_38),
.B1(n_15),
.B2(n_39),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_125),
.B1(n_31),
.B2(n_41),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_51),
.A2(n_38),
.B1(n_27),
.B2(n_26),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_64),
.A2(n_49),
.B1(n_26),
.B2(n_35),
.Y(n_103)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_105),
.B(n_1),
.C(n_2),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_68),
.A2(n_15),
.B1(n_38),
.B2(n_34),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_108),
.A2(n_22),
.B1(n_41),
.B2(n_34),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_17),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_67),
.A2(n_15),
.B1(n_18),
.B2(n_16),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_110),
.A2(n_117),
.B1(n_74),
.B2(n_70),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_57),
.B(n_18),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_111),
.B(n_126),
.Y(n_136)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_113),
.Y(n_176)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_42),
.A2(n_26),
.B1(n_18),
.B2(n_16),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_45),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_119),
.B(n_128),
.Y(n_145)
);

CKINVDCx12_ASAP7_75t_R g122 ( 
.A(n_62),
.Y(n_122)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_75),
.A2(n_40),
.B1(n_37),
.B2(n_24),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_50),
.B(n_16),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_50),
.A2(n_55),
.B(n_37),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_40),
.B(n_37),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_42),
.B(n_17),
.Y(n_128)
);

CKINVDCx12_ASAP7_75t_R g129 ( 
.A(n_42),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g172 ( 
.A(n_129),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_31),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_131),
.B(n_162),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_132),
.A2(n_164),
.B(n_97),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_112),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_133),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_134),
.B(n_137),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_139),
.A2(n_179),
.B1(n_182),
.B2(n_171),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_141),
.B(n_147),
.Y(n_212)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_81),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_160),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_72),
.B1(n_40),
.B2(n_24),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_149),
.A2(n_85),
.B1(n_76),
.B2(n_78),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_93),
.B(n_74),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_150),
.B(n_154),
.C(n_163),
.Y(n_208)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_90),
.B(n_74),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_152),
.B(n_156),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_95),
.B(n_70),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_155),
.A2(n_76),
.B1(n_78),
.B2(n_85),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_80),
.B(n_70),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_105),
.A2(n_60),
.B(n_34),
.C(n_31),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_168),
.B(n_179),
.C(n_8),
.Y(n_211)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_81),
.Y(n_160)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_106),
.Y(n_161)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_22),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_89),
.B(n_94),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_88),
.B(n_99),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_91),
.B(n_22),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_166),
.B(n_6),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_100),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_167),
.B(n_183),
.Y(n_221)
);

OA22x2_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_60),
.B1(n_58),
.B2(n_4),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_169),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_60),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_170),
.B(n_180),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_121),
.A2(n_1),
.B(n_2),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_171),
.A2(n_182),
.B(n_6),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_79),
.B(n_1),
.C(n_2),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_173),
.B(n_83),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_79),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_115),
.A2(n_124),
.B1(n_116),
.B2(n_118),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_177),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

AO22x2_ASAP7_75t_SL g179 ( 
.A1(n_114),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_5),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_100),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_181),
.B(n_160),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_113),
.A2(n_6),
.B(n_7),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_97),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_130),
.Y(n_186)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_130),
.Y(n_191)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_191),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_192),
.A2(n_137),
.B1(n_141),
.B2(n_168),
.Y(n_244)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_193),
.Y(n_240)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g245 ( 
.A(n_194),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_147),
.A2(n_84),
.B1(n_118),
.B2(n_124),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_196),
.A2(n_200),
.B(n_144),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_198),
.B(n_227),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_199),
.A2(n_192),
.B1(n_196),
.B2(n_228),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_131),
.B(n_116),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_203),
.B(n_205),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_143),
.B(n_8),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_139),
.A2(n_8),
.B1(n_83),
.B2(n_179),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_209),
.A2(n_151),
.B1(n_161),
.B2(n_165),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_226),
.B1(n_155),
.B2(n_207),
.Y(n_247)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_153),
.Y(n_213)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_164),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_218),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_132),
.A2(n_166),
.B(n_162),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_216),
.A2(n_168),
.B(n_172),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_217),
.B(n_223),
.C(n_176),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_164),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_138),
.Y(n_219)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_219),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_224),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_150),
.B(n_136),
.C(n_154),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_163),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_148),
.B(n_135),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_163),
.Y(n_228)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_145),
.B(n_169),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_159),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_157),
.B(n_173),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_208),
.Y(n_249)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_231),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

BUFx12_ASAP7_75t_L g237 ( 
.A(n_190),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_237),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_195),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_239),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_244),
.A2(n_268),
.B1(n_258),
.B2(n_261),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_168),
.B(n_158),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_246),
.A2(n_254),
.B(n_240),
.Y(n_294)
);

OAI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_247),
.A2(n_251),
.B1(n_260),
.B2(n_256),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_248),
.A2(n_264),
.B(n_265),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_249),
.B(n_239),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_250),
.B(n_252),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_176),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_140),
.B(n_165),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_184),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_261),
.Y(n_271)
);

INVx13_ASAP7_75t_L g257 ( 
.A(n_184),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_257),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_258),
.A2(n_267),
.B1(n_234),
.B2(n_238),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_266),
.C(n_225),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_185),
.A2(n_140),
.B1(n_172),
.B2(n_207),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_184),
.Y(n_261)
);

CKINVDCx12_ASAP7_75t_R g262 ( 
.A(n_221),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_214),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_188),
.B(n_205),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_263),
.B(n_253),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_R g264 ( 
.A(n_208),
.B(n_216),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_185),
.A2(n_211),
.B1(n_203),
.B2(n_187),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_217),
.C(n_188),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_200),
.A2(n_189),
.B1(n_198),
.B2(n_206),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_197),
.A2(n_187),
.B(n_204),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_269),
.A2(n_202),
.B(n_214),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_275),
.C(n_282),
.Y(n_302)
);

A2O1A1O1Ixp25_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_201),
.B(n_193),
.C(n_213),
.D(n_191),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_273),
.A2(n_274),
.B(n_278),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_204),
.C(n_219),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_234),
.A2(n_195),
.B(n_202),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_276),
.A2(n_290),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_277),
.B(n_288),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_210),
.C(n_194),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_210),
.B(n_235),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_283),
.A2(n_284),
.B(n_289),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_265),
.B(n_246),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_286),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_292),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_243),
.B(n_269),
.Y(n_288)
);

A2O1A1O1Ixp25_ASAP7_75t_L g289 ( 
.A1(n_264),
.A2(n_241),
.B(n_236),
.C(n_268),
.D(n_267),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_251),
.A2(n_257),
.B(n_241),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_232),
.C(n_233),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_245),
.C(n_237),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_232),
.A2(n_240),
.B1(n_233),
.B2(n_242),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_242),
.B(n_253),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_231),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_298),
.B(n_273),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_299),
.B(n_270),
.Y(n_312)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_312),
.C(n_282),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_292),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_306),
.B(n_310),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_272),
.B(n_231),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_307),
.B(n_313),
.Y(n_339)
);

OAI32xp33_ASAP7_75t_L g310 ( 
.A1(n_280),
.A2(n_231),
.A3(n_237),
.B1(n_245),
.B2(n_289),
.Y(n_310)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_296),
.Y(n_314)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_314),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_315),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_281),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_316),
.B(n_317),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_285),
.B(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_271),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_319),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_294),
.A2(n_283),
.B(n_284),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_320),
.A2(n_301),
.B(n_326),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_291),
.B(n_297),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_324),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_285),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_276),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_300),
.B(n_290),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_326),
.A2(n_319),
.B1(n_324),
.B2(n_301),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_293),
.B1(n_280),
.B2(n_286),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_327),
.A2(n_332),
.B1(n_308),
.B2(n_323),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_329),
.B(n_334),
.C(n_335),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_293),
.B1(n_295),
.B2(n_279),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_302),
.B(n_295),
.C(n_279),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_302),
.B(n_312),
.C(n_304),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_340),
.B(n_341),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_322),
.B(n_315),
.C(n_314),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_343),
.A2(n_320),
.B(n_309),
.Y(n_349)
);

BUFx12_ASAP7_75t_L g345 ( 
.A(n_310),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_316),
.Y(n_357)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_336),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_346),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_347),
.A2(n_328),
.B1(n_330),
.B2(n_338),
.Y(n_370)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_349),
.A2(n_358),
.B(n_359),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_343),
.A2(n_309),
.B(n_305),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_357),
.B(n_342),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_306),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_351),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_311),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_355),
.Y(n_362)
);

NOR3xp33_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_313),
.C(n_325),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_354),
.B(n_356),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_335),
.B(n_305),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_344),
.B(n_325),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_334),
.B(n_307),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_341),
.B(n_329),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_318),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_360),
.A2(n_336),
.B(n_337),
.Y(n_365)
);

FAx1_ASAP7_75t_SL g361 ( 
.A(n_348),
.B(n_331),
.CI(n_338),
.CON(n_361),
.SN(n_361)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_361),
.B(n_368),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_364),
.A2(n_349),
.B(n_350),
.Y(n_373)
);

OAI221xp5_ASAP7_75t_L g375 ( 
.A1(n_365),
.A2(n_328),
.B1(n_351),
.B2(n_330),
.C(n_303),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_348),
.B(n_327),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_370),
.B(n_352),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_368),
.B(n_353),
.C(n_355),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_372),
.B(n_375),
.Y(n_378)
);

AO21x1_ASAP7_75t_L g379 ( 
.A1(n_373),
.A2(n_374),
.B(n_369),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_367),
.B(n_332),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_376),
.B(n_369),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_371),
.A2(n_363),
.B(n_364),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_377),
.B(n_380),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

AOI322xp5_ASAP7_75t_L g383 ( 
.A1(n_382),
.A2(n_378),
.A3(n_345),
.B1(n_361),
.B2(n_303),
.C1(n_366),
.C2(n_362),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_383),
.B(n_384),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_381),
.B(n_372),
.C(n_362),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_385),
.B(n_345),
.Y(n_386)
);


endmodule