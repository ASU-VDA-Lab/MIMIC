module fake_netlist_5_875_n_122 (n_29, n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_30, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_122);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_122;

wire n_91;
wire n_82;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_114;
wire n_57;
wire n_96;
wire n_37;
wire n_111;
wire n_108;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_43;
wire n_107;
wire n_58;
wire n_69;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_105;
wire n_80;
wire n_35;
wire n_73;
wire n_92;
wire n_120;
wire n_33;
wire n_84;
wire n_79;
wire n_47;
wire n_53;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_71;
wire n_109;
wire n_112;
wire n_85;
wire n_95;
wire n_119;
wire n_59;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_64;
wire n_77;
wire n_102;
wire n_106;
wire n_81;
wire n_118;
wire n_89;
wire n_70;
wire n_115;
wire n_68;
wire n_93;
wire n_72;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_56;
wire n_51;
wire n_63;
wire n_97;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_6),
.B(n_19),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

NAND3xp33_ASAP7_75t_L g36 ( 
.A(n_15),
.B(n_27),
.C(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_4),
.B(n_23),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_18),
.B(n_14),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_10),
.B(n_11),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_22),
.B(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_1),
.B(n_16),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_7),
.B(n_1),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_2),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_40),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_51),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_31),
.B1(n_47),
.B2(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_31),
.B(n_47),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_49),
.C(n_36),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_47),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_59),
.A2(n_49),
.B(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_63),
.A2(n_36),
.B1(n_41),
.B2(n_45),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_42),
.B(n_33),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_65),
.A2(n_33),
.B(n_41),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_32),
.B(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g75 ( 
.A(n_56),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_67),
.B(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_58),
.A2(n_32),
.B(n_53),
.C(n_35),
.Y(n_80)
);

OR2x6_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_58),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_L g83 ( 
.A1(n_69),
.A2(n_32),
.B1(n_53),
.B2(n_63),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_60),
.B1(n_38),
.B2(n_39),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_81),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_95),
.B(n_84),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_93),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_101),
.Y(n_103)
);

OAI221xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_94),
.B1(n_81),
.B2(n_89),
.C(n_84),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_105),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_SL g109 ( 
.A(n_104),
.B(n_99),
.C(n_96),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_109),
.A2(n_110),
.B1(n_60),
.B2(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_107),
.Y(n_112)
);

NOR2xp67_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_108),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_112),
.B(n_105),
.Y(n_114)
);

NAND4xp75_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_83),
.C(n_74),
.D(n_92),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_98),
.Y(n_116)
);

AOI22x1_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_117)
);

OAI22x1_ASAP7_75t_L g118 ( 
.A1(n_116),
.A2(n_115),
.B1(n_90),
.B2(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

AOI21x1_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_118),
.B(n_38),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_118),
.B(n_37),
.Y(n_121)
);

OR2x6_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_120),
.Y(n_122)
);


endmodule