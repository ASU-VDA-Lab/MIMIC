module real_aes_18037_n_98 (n_17, n_28, n_76, n_56, n_34, n_866, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_866;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_148;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_0), .Y(n_575) );
AND2x4_ASAP7_75t_L g104 ( .A(n_1), .B(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_2), .A2(n_117), .B1(n_118), .B2(n_477), .Y(n_116) );
INVx1_ASAP7_75t_SL g117 ( .A(n_2), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g232 ( .A1(n_3), .A2(n_4), .B1(n_233), .B2(n_234), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_5), .A2(n_22), .B1(n_134), .B2(n_146), .Y(n_305) );
AOI22xp33_ASAP7_75t_L g165 ( .A1(n_6), .A2(n_51), .B1(n_166), .B2(n_167), .Y(n_165) );
BUFx3_ASAP7_75t_L g532 ( .A(n_7), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g198 ( .A1(n_8), .A2(n_14), .B1(n_143), .B2(n_183), .Y(n_198) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_10), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_11), .B(n_190), .Y(n_517) );
OR2x2_ASAP7_75t_L g112 ( .A(n_12), .B(n_31), .Y(n_112) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_13), .Y(n_135) );
OAI22xp33_ASAP7_75t_SL g485 ( .A1(n_15), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_15), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_15), .A2(n_486), .B1(n_500), .B2(n_837), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_16), .B(n_173), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_17), .B(n_211), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_18), .A2(n_83), .B1(n_146), .B2(n_173), .Y(n_581) );
CKINVDCx20_ASAP7_75t_R g480 ( .A(n_19), .Y(n_480) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_20), .A2(n_47), .B(n_129), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_21), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_23), .B(n_134), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_24), .B(n_141), .Y(n_257) );
INVx4_ASAP7_75t_R g219 ( .A(n_25), .Y(n_219) );
AO32x2_ASAP7_75t_L g578 ( .A1(n_26), .A2(n_152), .A3(n_153), .B1(n_579), .B2(n_582), .Y(n_578) );
AO32x1_ASAP7_75t_L g615 ( .A1(n_26), .A2(n_152), .A3(n_153), .B1(n_579), .B2(n_582), .Y(n_615) );
INVx1_ASAP7_75t_L g238 ( .A(n_27), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_28), .B(n_134), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_SL g142 ( .A1(n_29), .A2(n_143), .B(n_144), .C(n_147), .Y(n_142) );
AOI22xp33_ASAP7_75t_L g306 ( .A1(n_30), .A2(n_44), .B1(n_143), .B2(n_201), .Y(n_306) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_32), .Y(n_138) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_33), .A2(n_50), .B1(n_134), .B2(n_220), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g580 ( .A1(n_34), .A2(n_88), .B1(n_146), .B2(n_201), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_35), .B(n_519), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_36), .B(n_554), .Y(n_604) );
INVx1_ASAP7_75t_L g260 ( .A(n_37), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_38), .B(n_143), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_39), .A2(n_65), .B1(n_201), .B2(n_587), .Y(n_586) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_40), .Y(n_184) );
INVx2_ASAP7_75t_L g483 ( .A(n_41), .Y(n_483) );
INVx1_ASAP7_75t_L g110 ( .A(n_42), .Y(n_110) );
BUFx3_ASAP7_75t_L g498 ( .A(n_42), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_43), .B(n_606), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_45), .Y(n_221) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_46), .A2(n_82), .B1(n_143), .B2(n_201), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g571 ( .A(n_48), .Y(n_571) );
CKINVDCx5p33_ASAP7_75t_R g558 ( .A(n_49), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_52), .A2(n_76), .B1(n_175), .B2(n_554), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_53), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_54), .A2(n_80), .B1(n_146), .B2(n_173), .Y(n_528) );
INVx1_ASAP7_75t_L g129 ( .A(n_55), .Y(n_129) );
AND2x4_ASAP7_75t_L g149 ( .A(n_56), .B(n_150), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g230 ( .A1(n_57), .A2(n_87), .B1(n_201), .B2(n_231), .Y(n_230) );
AO22x1_ASAP7_75t_L g171 ( .A1(n_58), .A2(n_70), .B1(n_172), .B2(n_174), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_59), .B(n_146), .Y(n_516) );
INVx1_ASAP7_75t_L g150 ( .A(n_60), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_61), .B(n_152), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_62), .B(n_152), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g573 ( .A1(n_63), .A2(n_163), .B(n_166), .C(n_574), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g522 ( .A(n_64), .B(n_146), .C(n_521), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_66), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_67), .B(n_166), .Y(n_191) );
AND2x2_ASAP7_75t_L g576 ( .A(n_68), .B(n_224), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_69), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_71), .B(n_134), .Y(n_185) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_72), .A2(n_93), .B1(n_173), .B2(n_175), .Y(n_556) );
INVx2_ASAP7_75t_L g141 ( .A(n_73), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_74), .B(n_186), .Y(n_540) );
CKINVDCx5p33_ASAP7_75t_R g843 ( .A(n_75), .Y(n_843) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_77), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_78), .B(n_152), .Y(n_254) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_79), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_81), .B(n_127), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_84), .B(n_521), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_85), .A2(n_97), .B1(n_201), .B2(n_220), .Y(n_529) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_86), .B(n_554), .Y(n_601) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_89), .B(n_152), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g108 ( .A(n_90), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g493 ( .A(n_90), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_91), .B(n_211), .Y(n_607) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_92), .A2(n_166), .B(n_203), .C(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g223 ( .A(n_94), .B(n_224), .Y(n_223) );
NAND2xp33_ASAP7_75t_L g189 ( .A(n_95), .B(n_190), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_96), .Y(n_537) );
AOI21xp33_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_113), .B(n_850), .Y(n_98) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_100), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_102), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx2_ASAP7_75t_SL g860 ( .A(n_104), .Y(n_860) );
INVx5_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_107), .Y(n_115) );
INVx3_ASAP7_75t_L g479 ( .A(n_107), .Y(n_479) );
AND2x6_ASAP7_75t_SL g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_111), .B(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
NOR2x1_ASAP7_75t_L g849 ( .A(n_112), .B(n_498), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_481), .B(n_484), .Y(n_113) );
OAI22xp33_ASAP7_75t_SL g850 ( .A1(n_114), .A2(n_117), .B1(n_851), .B2(n_861), .Y(n_850) );
AOI21x1_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_116), .B(n_478), .Y(n_114) );
INVx1_ASAP7_75t_L g477 ( .A(n_118), .Y(n_477) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g488 ( .A(n_119), .Y(n_488) );
OR2x2_ASAP7_75t_L g119 ( .A(n_120), .B(n_377), .Y(n_119) );
NAND3xp33_ASAP7_75t_SL g120 ( .A(n_121), .B(n_279), .C(n_339), .Y(n_120) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_154), .B1(n_266), .B2(n_272), .Y(n_121) );
HB1xp67_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g336 ( .A(n_123), .B(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_123), .B(n_253), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_123), .B(n_299), .Y(n_447) );
AND2x2_ASAP7_75t_L g453 ( .A(n_123), .B(n_278), .Y(n_453) );
INVxp67_ASAP7_75t_L g458 ( .A(n_123), .Y(n_458) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
INVx2_ASAP7_75t_L g270 ( .A(n_124), .Y(n_270) );
AOI21x1_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_130), .B(n_151), .Y(n_124) );
AO31x2_ASAP7_75t_L g228 ( .A1(n_125), .A2(n_229), .A3(n_235), .B(n_237), .Y(n_228) );
BUFx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_126), .B(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g224 ( .A(n_126), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_126), .B(n_238), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_126), .B(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_126), .B(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
OAI21xp33_ASAP7_75t_L g177 ( .A1(n_127), .A2(n_148), .B(n_169), .Y(n_177) );
INVx2_ASAP7_75t_L g204 ( .A(n_127), .Y(n_204) );
INVx2_ASAP7_75t_L g212 ( .A(n_127), .Y(n_212) );
INVx2_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_128), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_142), .B(n_148), .Y(n_130) );
OAI21xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_136), .B(n_139), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
OAI22xp5_ASAP7_75t_L g569 ( .A1(n_134), .A2(n_220), .B1(n_570), .B2(n_571), .Y(n_569) );
INVx2_ASAP7_75t_L g587 ( .A(n_134), .Y(n_587) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g137 ( .A(n_135), .Y(n_137) );
INVx3_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx2_ASAP7_75t_L g146 ( .A(n_135), .Y(n_146) );
INVx1_ASAP7_75t_L g166 ( .A(n_135), .Y(n_166) );
INVx1_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_135), .Y(n_173) );
INVx1_ASAP7_75t_L g175 ( .A(n_135), .Y(n_175) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_135), .Y(n_201) );
INVx1_ASAP7_75t_L g220 ( .A(n_135), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
INVx2_ASAP7_75t_L g234 ( .A(n_137), .Y(n_234) );
O2A1O1Ixp5_ASAP7_75t_L g536 ( .A1(n_139), .A2(n_234), .B(n_537), .C(n_538), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_139), .A2(n_147), .B1(n_580), .B2(n_581), .Y(n_579) );
BUFx4f_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_140), .B(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g521 ( .A(n_140), .Y(n_521) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx8_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx2_ASAP7_75t_L g164 ( .A(n_141), .Y(n_164) );
INVx1_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
INVx4_ASAP7_75t_L g183 ( .A(n_143), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
INVx2_ASAP7_75t_SL g554 ( .A(n_146), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_147), .B(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_147), .A2(n_189), .B(n_191), .Y(n_188) );
INVx6_ASAP7_75t_L g199 ( .A(n_147), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_147), .A2(n_161), .B(n_171), .C(n_177), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_147), .A2(n_516), .B(n_517), .Y(n_515) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_147), .A2(n_199), .B1(n_528), .B2(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_148), .A2(n_568), .B(n_573), .Y(n_567) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx10_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
BUFx10_ASAP7_75t_L g205 ( .A(n_149), .Y(n_205) );
INVx1_ASAP7_75t_L g236 ( .A(n_149), .Y(n_236) );
AO31x2_ASAP7_75t_L g584 ( .A1(n_149), .A2(n_551), .A3(n_585), .B(n_589), .Y(n_584) );
NOR2x1_ASAP7_75t_L g192 ( .A(n_152), .B(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g307 ( .A(n_152), .Y(n_307) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g264 ( .A(n_153), .B(n_194), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_153), .B(n_531), .Y(n_530) );
INVx2_ASAP7_75t_L g534 ( .A(n_153), .Y(n_534) );
BUFx3_ASAP7_75t_L g551 ( .A(n_153), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_153), .B(n_590), .Y(n_589) );
INVx2_ASAP7_75t_SL g598 ( .A(n_153), .Y(n_598) );
OAI21xp5_ASAP7_75t_SL g154 ( .A1(n_155), .A2(n_225), .B(n_239), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_195), .Y(n_156) );
INVx1_ASAP7_75t_L g374 ( .A(n_157), .Y(n_374) );
AND2x2_ASAP7_75t_L g403 ( .A(n_157), .B(n_365), .Y(n_403) );
AND2x2_ASAP7_75t_L g157 ( .A(n_158), .B(n_178), .Y(n_157) );
AND2x2_ASAP7_75t_L g296 ( .A(n_158), .B(n_209), .Y(n_296) );
INVx1_ASAP7_75t_L g352 ( .A(n_158), .Y(n_352) );
AND2x2_ASAP7_75t_L g402 ( .A(n_158), .B(n_208), .Y(n_402) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
AND2x2_ASAP7_75t_L g276 ( .A(n_159), .B(n_208), .Y(n_276) );
AND2x4_ASAP7_75t_L g421 ( .A(n_159), .B(n_209), .Y(n_421) );
AOI21x1_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_170), .B(n_176), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
OAI21x1_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_169), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_162), .A2(n_262), .B(n_263), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_162), .A2(n_199), .B1(n_305), .B2(n_306), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_162), .A2(n_199), .B1(n_586), .B2(n_588), .Y(n_585) );
AOI21x1_ASAP7_75t_L g600 ( .A1(n_162), .A2(n_601), .B(n_602), .Y(n_600) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g187 ( .A(n_164), .Y(n_187) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_168), .B(n_216), .Y(n_215) );
INVxp67_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
INVx3_ASAP7_75t_L g606 ( .A(n_173), .Y(n_606) );
OAI21xp33_ASAP7_75t_SL g256 ( .A1(n_174), .A2(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_175), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
BUFx2_ASAP7_75t_L g346 ( .A(n_178), .Y(n_346) );
AND2x2_ASAP7_75t_L g415 ( .A(n_178), .B(n_209), .Y(n_415) );
AND2x2_ASAP7_75t_L g422 ( .A(n_178), .B(n_247), .Y(n_422) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g243 ( .A(n_179), .Y(n_243) );
BUFx3_ASAP7_75t_L g278 ( .A(n_179), .Y(n_278) );
AND2x2_ASAP7_75t_L g289 ( .A(n_179), .B(n_275), .Y(n_289) );
AND2x2_ASAP7_75t_L g353 ( .A(n_179), .B(n_196), .Y(n_353) );
AND2x2_ASAP7_75t_L g358 ( .A(n_179), .B(n_209), .Y(n_358) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
OAI21x1_ASAP7_75t_L g181 ( .A1(n_182), .A2(n_188), .B(n_192), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_185), .C(n_186), .Y(n_182) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_187), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_539) );
OAI22xp33_ASAP7_75t_L g218 ( .A1(n_190), .A2(n_219), .B1(n_220), .B2(n_221), .Y(n_218) );
INVx2_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AO31x2_ASAP7_75t_L g303 ( .A1(n_194), .A2(n_304), .A3(n_307), .B(n_308), .Y(n_303) );
OAI21x1_ASAP7_75t_L g514 ( .A1(n_194), .A2(n_515), .B(n_518), .Y(n_514) );
AOI31xp67_ASAP7_75t_L g526 ( .A1(n_194), .A2(n_307), .A3(n_527), .B(n_530), .Y(n_526) );
OAI21x1_ASAP7_75t_L g535 ( .A1(n_194), .A2(n_536), .B(n_539), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_195), .B(n_364), .Y(n_466) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_208), .Y(n_195) );
INVx2_ASAP7_75t_L g247 ( .A(n_196), .Y(n_247) );
OR2x2_ASAP7_75t_L g250 ( .A(n_196), .B(n_209), .Y(n_250) );
INVx2_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_196), .B(n_245), .Y(n_291) );
AND2x2_ASAP7_75t_L g365 ( .A(n_196), .B(n_209), .Y(n_365) );
AO31x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_204), .A3(n_205), .B(n_206), .Y(n_196) );
OAI22x1_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B1(n_200), .B2(n_202), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_199), .A2(n_202), .B1(n_230), .B2(n_232), .Y(n_229) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_199), .A2(n_553), .B1(n_555), .B2(n_556), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_199), .A2(n_604), .B(n_605), .Y(n_603) );
INVx2_ASAP7_75t_L g233 ( .A(n_201), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_201), .B(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g519 ( .A(n_201), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_202), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_SL g555 ( .A(n_203), .Y(n_555) );
INVx1_ASAP7_75t_L g572 ( .A(n_203), .Y(n_572) );
INVx2_ASAP7_75t_L g513 ( .A(n_204), .Y(n_513) );
INVx2_ASAP7_75t_L g222 ( .A(n_205), .Y(n_222) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g292 ( .A(n_209), .Y(n_292) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_213), .B(n_223), .Y(n_209) );
AOI21x1_ASAP7_75t_L g566 ( .A1(n_210), .A2(n_567), .B(n_576), .Y(n_566) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_217), .B(n_222), .Y(n_213) );
INVx1_ASAP7_75t_L g541 ( .A(n_220), .Y(n_541) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_226), .B(n_328), .Y(n_474) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g285 ( .A(n_227), .Y(n_285) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g265 ( .A(n_228), .Y(n_265) );
AND2x2_ASAP7_75t_L g271 ( .A(n_228), .B(n_253), .Y(n_271) );
INVx1_ASAP7_75t_L g320 ( .A(n_228), .Y(n_320) );
OR2x2_ASAP7_75t_L g325 ( .A(n_228), .B(n_303), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_228), .B(n_303), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_228), .B(n_302), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_228), .B(n_270), .Y(n_410) );
AO31x2_ASAP7_75t_L g550 ( .A1(n_235), .A2(n_551), .A3(n_552), .B(n_557), .Y(n_550) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
INVx2_ASAP7_75t_SL g582 ( .A(n_236), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_240), .A2(n_248), .B(n_251), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_244), .Y(n_241) );
OR2x2_ASAP7_75t_L g249 ( .A(n_242), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g401 ( .A(n_242), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g431 ( .A(n_242), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_243), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g399 ( .A(n_243), .Y(n_399) );
OR2x2_ASAP7_75t_L g312 ( .A(n_244), .B(n_313), .Y(n_312) );
INVxp33_ASAP7_75t_L g430 ( .A(n_244), .Y(n_430) );
OR2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
INVx2_ASAP7_75t_L g334 ( .A(n_245), .Y(n_334) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g287 ( .A(n_247), .Y(n_287) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OAI221xp5_ASAP7_75t_SL g396 ( .A1(n_249), .A2(n_321), .B1(n_326), .B2(n_397), .C(n_400), .Y(n_396) );
OR2x2_ASAP7_75t_L g383 ( .A(n_250), .B(n_334), .Y(n_383) );
INVx2_ASAP7_75t_L g432 ( .A(n_250), .Y(n_432) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g332 ( .A(n_252), .Y(n_332) );
OR2x2_ASAP7_75t_L g335 ( .A(n_252), .B(n_336), .Y(n_335) );
INVxp67_ASAP7_75t_SL g376 ( .A(n_252), .Y(n_376) );
OR2x2_ASAP7_75t_L g389 ( .A(n_252), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_265), .Y(n_252) );
NAND2x1p5_ASAP7_75t_SL g284 ( .A(n_253), .B(n_269), .Y(n_284) );
INVx3_ASAP7_75t_L g299 ( .A(n_253), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_253), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g323 ( .A(n_253), .Y(n_323) );
AND2x2_ASAP7_75t_L g404 ( .A(n_253), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g411 ( .A(n_253), .B(n_318), .Y(n_411) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_261), .B(n_264), .Y(n_255) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_271), .Y(n_266) );
AND2x2_ASAP7_75t_L g463 ( .A(n_267), .B(n_322), .Y(n_463) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g367 ( .A(n_269), .B(n_337), .Y(n_367) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g301 ( .A(n_270), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g328 ( .A(n_270), .B(n_303), .Y(n_328) );
AND2x4_ASAP7_75t_L g425 ( .A(n_271), .B(n_395), .Y(n_425) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_277), .Y(n_272) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_277), .B(n_365), .Y(n_449) );
AND2x2_ASAP7_75t_L g456 ( .A(n_277), .B(n_416), .Y(n_456) );
INVx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
BUFx2_ASAP7_75t_L g381 ( .A(n_278), .Y(n_381) );
AOI321xp33_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_293), .A3(n_310), .B1(n_311), .B2(n_314), .C(n_329), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_281), .B(n_290), .Y(n_280) );
AOI21xp33_ASAP7_75t_SL g281 ( .A1(n_282), .A2(n_286), .B(n_288), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OAI21xp33_ASAP7_75t_L g293 ( .A1(n_283), .A2(n_294), .B(n_297), .Y(n_293) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
OR2x2_ASAP7_75t_L g393 ( .A(n_284), .B(n_325), .Y(n_393) );
INVx1_ASAP7_75t_L g385 ( .A(n_285), .Y(n_385) );
INVx2_ASAP7_75t_L g370 ( .A(n_286), .Y(n_370) );
OAI32xp33_ASAP7_75t_L g473 ( .A1(n_286), .A2(n_435), .A3(n_446), .B1(n_474), .B2(n_475), .Y(n_473) );
INVx1_ASAP7_75t_L g388 ( .A(n_287), .Y(n_388) );
INVx1_ASAP7_75t_L g338 ( .A(n_288), .Y(n_338) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_SL g426 ( .A(n_289), .B(n_333), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_290), .B(n_294), .Y(n_310) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_290), .A2(n_367), .B1(n_428), .B2(n_449), .Y(n_448) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g416 ( .A(n_291), .Y(n_416) );
INVx1_ASAP7_75t_L g313 ( .A(n_292), .Y(n_313) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx2_ASAP7_75t_L g398 ( .A(n_296), .Y(n_398) );
NAND4xp25_ASAP7_75t_L g314 ( .A(n_297), .B(n_315), .C(n_321), .D(n_326), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
INVxp67_ASAP7_75t_L g340 ( .A(n_298), .Y(n_340) );
AND2x2_ASAP7_75t_L g419 ( .A(n_298), .B(n_328), .Y(n_419) );
OR2x2_ASAP7_75t_L g428 ( .A(n_298), .B(n_301), .Y(n_428) );
AND2x2_ASAP7_75t_L g452 ( .A(n_298), .B(n_324), .Y(n_452) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g366 ( .A(n_299), .B(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g373 ( .A(n_299), .B(n_320), .Y(n_373) );
INVx1_ASAP7_75t_L g437 ( .A(n_300), .Y(n_437) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g345 ( .A(n_301), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g395 ( .A(n_301), .Y(n_395) );
INVx1_ASAP7_75t_L g337 ( .A(n_302), .Y(n_337) );
INVx2_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g318 ( .A(n_303), .Y(n_318) );
INVx3_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NOR2xp33_ASAP7_75t_L g316 ( .A(n_317), .B(n_319), .Y(n_316) );
AND2x4_ASAP7_75t_L g331 ( .A(n_317), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g372 ( .A(n_317), .Y(n_372) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_319), .Y(n_436) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g327 ( .A(n_323), .B(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g413 ( .A(n_325), .Y(n_413) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g390 ( .A(n_328), .Y(n_390) );
AND2x2_ASAP7_75t_L g433 ( .A(n_328), .B(n_373), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_SL g329 ( .A1(n_330), .A2(n_333), .B(n_335), .C(n_338), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g444 ( .A(n_333), .B(n_422), .Y(n_444) );
INVx2_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g348 ( .A(n_336), .Y(n_348) );
AOI211xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B(n_354), .C(n_368), .Y(n_339) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_345), .B(n_347), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_343), .A2(n_451), .B(n_454), .Y(n_450) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g364 ( .A(n_346), .Y(n_364) );
AND2x2_ASAP7_75t_L g424 ( .A(n_346), .B(n_421), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g443 ( .A(n_351), .Y(n_443) );
AND2x2_ASAP7_75t_L g469 ( .A(n_351), .B(n_432), .Y(n_469) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g357 ( .A(n_352), .Y(n_357) );
INVx2_ASAP7_75t_L g408 ( .A(n_353), .Y(n_408) );
NAND2x1_ASAP7_75t_L g442 ( .A(n_353), .B(n_443), .Y(n_442) );
AOI33xp33_ASAP7_75t_L g460 ( .A1(n_353), .A2(n_373), .A3(n_411), .B1(n_421), .B2(n_453), .B3(n_866), .Y(n_460) );
OAI22xp33_ASAP7_75t_SL g354 ( .A1(n_355), .A2(n_359), .B1(n_362), .B2(n_366), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g387 ( .A(n_358), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_359), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
OR2x2_ASAP7_75t_L g472 ( .A(n_361), .B(n_406), .Y(n_472) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OAI22xp33_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_371), .B1(n_374), .B2(n_375), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_372), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_372), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g394 ( .A(n_373), .B(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g459 ( .A(n_373), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_438), .Y(n_377) );
NOR4xp25_ASAP7_75t_L g378 ( .A(n_379), .B(n_396), .C(n_417), .D(n_434), .Y(n_378) );
OAI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_384), .B1(n_386), .B2(n_389), .C(n_391), .Y(n_379) );
O2A1O1Ixp33_ASAP7_75t_SL g434 ( .A1(n_380), .A2(n_435), .B(n_436), .C(n_437), .Y(n_434) );
NAND2x1_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g467 ( .A(n_383), .Y(n_467) );
INVx2_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_387), .A2(n_392), .B(n_394), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
O2A1O1Ixp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_404), .C(n_407), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g446 ( .A(n_406), .B(n_447), .Y(n_446) );
INVxp67_ASAP7_75t_SL g470 ( .A(n_406), .Y(n_470) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_409), .B1(n_412), .B2(n_414), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_411), .Y(n_409) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
OAI211xp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_420), .B(n_423), .C(n_429), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AOI221xp5_ASAP7_75t_L g468 ( .A1(n_421), .A2(n_469), .B1(n_470), .B2(n_471), .C(n_473), .Y(n_468) );
INVx3_ASAP7_75t_L g476 ( .A(n_421), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_425), .B1(n_426), .B2(n_427), .Y(n_423) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_433), .Y(n_429) );
INVx1_ASAP7_75t_L g435 ( .A(n_432), .Y(n_435) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_461), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_450), .Y(n_439) );
O2A1O1Ixp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_444), .B(n_445), .C(n_448), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_444), .B(n_465), .C(n_467), .Y(n_464) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
OAI21xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_457), .B(n_460), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_459), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_462), .A2(n_464), .B(n_468), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_SL g478 ( .A(n_479), .B(n_480), .Y(n_478) );
OR2x6_ASAP7_75t_L g855 ( .A(n_479), .B(n_856), .Y(n_855) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_479), .B(n_483), .Y(n_864) );
BUFx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x6_ASAP7_75t_SL g495 ( .A(n_482), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g846 ( .A(n_483), .B(n_847), .Y(n_846) );
INVx3_ASAP7_75t_L g858 ( .A(n_483), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_489), .B1(n_499), .B2(n_839), .C(n_842), .Y(n_484) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
NOR2xp67_ASAP7_75t_SL g489 ( .A(n_490), .B(n_494), .Y(n_489) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g848 ( .A(n_492), .B(n_849), .Y(n_848) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g841 ( .A(n_493), .Y(n_841) );
NOR2x1_ASAP7_75t_R g839 ( .A(n_494), .B(n_840), .Y(n_839) );
INVx5_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
HB1xp67_ASAP7_75t_L g838 ( .A(n_502), .Y(n_838) );
OR2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_747), .Y(n_502) );
NAND4xp25_ASAP7_75t_L g503 ( .A(n_504), .B(n_652), .C(n_679), .D(n_715), .Y(n_503) );
AOI221x1_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_563), .B1(n_591), .B2(n_627), .C(n_631), .Y(n_504) );
NAND3xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_544), .C(n_561), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_524), .Y(n_508) );
INVx2_ASAP7_75t_L g592 ( .A(n_509), .Y(n_592) );
AND2x2_ASAP7_75t_L g765 ( .A(n_509), .B(n_709), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_509), .B(n_562), .Y(n_774) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g780 ( .A(n_510), .Y(n_780) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g625 ( .A(n_511), .Y(n_625) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OR2x2_ASAP7_75t_L g708 ( .A(n_512), .B(n_560), .Y(n_708) );
OAI21x1_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_523), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g637 ( .A1(n_513), .A2(n_514), .B(n_523), .Y(n_637) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_522), .Y(n_518) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_524), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_524), .B(n_736), .Y(n_735) );
INVxp67_ASAP7_75t_L g778 ( .A(n_524), .Y(n_778) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_533), .Y(n_524) );
AND2x2_ASAP7_75t_L g562 ( .A(n_525), .B(n_550), .Y(n_562) );
INVx2_ASAP7_75t_L g634 ( .A(n_525), .Y(n_634) );
AND2x2_ASAP7_75t_L g699 ( .A(n_525), .B(n_637), .Y(n_699) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g560 ( .A(n_526), .Y(n_560) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g626 ( .A(n_533), .Y(n_626) );
AND2x2_ASAP7_75t_L g636 ( .A(n_533), .B(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g698 ( .A(n_533), .B(n_550), .Y(n_698) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_535), .B(n_543), .Y(n_533) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_534), .A2(n_535), .B(n_543), .Y(n_547) );
INVx1_ASAP7_75t_L g663 ( .A(n_544), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_546), .B(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_546), .B(n_678), .Y(n_677) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_546), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_546), .B(n_733), .Y(n_740) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g709 ( .A(n_547), .B(n_684), .Y(n_709) );
OR2x2_ASAP7_75t_L g711 ( .A(n_547), .B(n_637), .Y(n_711) );
INVx1_ASAP7_75t_L g770 ( .A(n_547), .Y(n_770) );
BUFx2_ASAP7_75t_L g784 ( .A(n_547), .Y(n_784) );
OR2x2_ASAP7_75t_L g812 ( .A(n_547), .B(n_550), .Y(n_812) );
INVx1_ASAP7_75t_L g831 ( .A(n_548), .Y(n_831) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g678 ( .A(n_549), .Y(n_678) );
OR2x2_ASAP7_75t_L g691 ( .A(n_549), .B(n_692), .Y(n_691) );
OR2x2_ASAP7_75t_L g710 ( .A(n_549), .B(n_711), .Y(n_710) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_559), .Y(n_549) );
INVx2_ASAP7_75t_L g630 ( .A(n_550), .Y(n_630) );
AND2x2_ASAP7_75t_L g646 ( .A(n_550), .B(n_559), .Y(n_646) );
INVx1_ASAP7_75t_L g684 ( .A(n_550), .Y(n_684) );
INVx1_ASAP7_75t_L g727 ( .A(n_550), .Y(n_727) );
AND2x2_ASAP7_75t_L g769 ( .A(n_550), .B(n_770), .Y(n_769) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g825 ( .A(n_561), .Y(n_825) );
AND2x4_ASAP7_75t_L g763 ( .A(n_562), .B(n_623), .Y(n_763) );
INVx2_ASAP7_75t_L g792 ( .A(n_562), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_562), .B(n_784), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_563), .B(n_782), .Y(n_781) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_577), .Y(n_563) );
AND2x2_ASAP7_75t_L g703 ( .A(n_564), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g724 ( .A(n_564), .B(n_725), .Y(n_724) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x2_ASAP7_75t_L g595 ( .A(n_565), .B(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g619 ( .A(n_565), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g650 ( .A(n_565), .Y(n_650) );
AND2x2_ASAP7_75t_L g690 ( .A(n_565), .B(n_583), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_565), .B(n_674), .Y(n_731) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_L g643 ( .A(n_566), .Y(n_643) );
NAND2xp5_ASAP7_75t_SL g568 ( .A(n_569), .B(n_572), .Y(n_568) );
INVx3_ASAP7_75t_L g609 ( .A(n_577), .Y(n_609) );
AND2x2_ASAP7_75t_L g654 ( .A(n_577), .B(n_649), .Y(n_654) );
AND2x2_ASAP7_75t_L g809 ( .A(n_577), .B(n_613), .Y(n_809) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_583), .Y(n_577) );
INVx1_ASAP7_75t_L g660 ( .A(n_578), .Y(n_660) );
AND2x2_ASAP7_75t_L g688 ( .A(n_578), .B(n_596), .Y(n_688) );
OAI21x1_ASAP7_75t_L g599 ( .A1(n_582), .A2(n_600), .B(n_603), .Y(n_599) );
AND2x4_ASAP7_75t_L g641 ( .A(n_583), .B(n_642), .Y(n_641) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g614 ( .A(n_584), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g651 ( .A(n_584), .B(n_615), .Y(n_651) );
AND2x2_ASAP7_75t_L g661 ( .A(n_584), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_584), .B(n_596), .Y(n_713) );
AND2x2_ASAP7_75t_L g719 ( .A(n_584), .B(n_643), .Y(n_719) );
OAI21xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_610), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g752 ( .A1(n_592), .A2(n_753), .B(n_757), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g830 ( .A(n_592), .B(n_783), .Y(n_830) );
NAND2x1_ASAP7_75t_SL g593 ( .A(n_594), .B(n_608), .Y(n_593) );
INVx1_ASAP7_75t_L g836 ( .A(n_594), .Y(n_836) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx2_ASAP7_75t_L g613 ( .A(n_596), .Y(n_613) );
INVx2_ASAP7_75t_L g618 ( .A(n_596), .Y(n_618) );
INVxp67_ASAP7_75t_L g639 ( .A(n_596), .Y(n_639) );
AND2x2_ASAP7_75t_L g659 ( .A(n_596), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g670 ( .A(n_596), .B(n_671), .Y(n_670) );
INVx3_ASAP7_75t_L g674 ( .A(n_596), .Y(n_674) );
INVx1_ASAP7_75t_L g692 ( .A(n_596), .Y(n_692) );
OR2x2_ASAP7_75t_L g725 ( .A(n_596), .B(n_660), .Y(n_725) );
INVx1_ASAP7_75t_L g796 ( .A(n_596), .Y(n_796) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
OAI21x1_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_607), .Y(n_597) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_616), .B(n_621), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g734 ( .A1(n_612), .A2(n_735), .B1(n_737), .B2(n_740), .Y(n_734) );
OR2x2_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_613), .B(n_661), .Y(n_695) );
BUFx2_ASAP7_75t_L g754 ( .A(n_613), .Y(n_754) );
INVx2_ASAP7_75t_L g704 ( .A(n_614), .Y(n_704) );
OR2x2_ASAP7_75t_L g788 ( .A(n_614), .B(n_618), .Y(n_788) );
INVx1_ASAP7_75t_L g620 ( .A(n_615), .Y(n_620) );
INVx1_ASAP7_75t_L g669 ( .A(n_615), .Y(n_669) );
NOR2x1p5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVxp67_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
HB1xp67_ASAP7_75t_L g739 ( .A(n_618), .Y(n_739) );
OR2x2_ASAP7_75t_L g823 ( .A(n_618), .B(n_824), .Y(n_823) );
AND2x2_ASAP7_75t_L g826 ( .A(n_618), .B(n_661), .Y(n_826) );
INVxp67_ASAP7_75t_SL g789 ( .A(n_619), .Y(n_789) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_623), .B(n_683), .Y(n_745) );
AND2x2_ASAP7_75t_L g835 ( .A(n_623), .B(n_633), .Y(n_835) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
OR2x2_ASAP7_75t_L g744 ( .A(n_624), .B(n_633), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g701 ( .A(n_625), .B(n_634), .Y(n_701) );
AND2x2_ASAP7_75t_L g736 ( .A(n_625), .B(n_630), .Y(n_736) );
INVxp67_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
AND2x2_ASAP7_75t_L g655 ( .A(n_628), .B(n_636), .Y(n_655) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g795 ( .A(n_630), .B(n_796), .Y(n_795) );
OAI22xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_638), .B1(n_644), .B2(n_647), .Y(n_631) );
O2A1O1Ixp33_ASAP7_75t_L g832 ( .A1(n_632), .A2(n_833), .B(n_834), .C(n_836), .Y(n_832) );
OR2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g683 ( .A(n_634), .B(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g751 ( .A(n_634), .Y(n_751) );
OR2x2_ASAP7_75t_L g798 ( .A(n_635), .B(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
AND2x2_ASAP7_75t_L g653 ( .A(n_639), .B(n_654), .Y(n_653) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g756 ( .A(n_642), .Y(n_756) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g662 ( .A(n_643), .Y(n_662) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_643), .Y(n_671) );
INVx1_ASAP7_75t_L g743 ( .A(n_643), .Y(n_743) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g799 ( .A(n_646), .Y(n_799) );
AND2x2_ASAP7_75t_L g821 ( .A(n_646), .B(n_784), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_647), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g673 ( .A(n_651), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g729 ( .A(n_651), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_SL g824 ( .A(n_651), .Y(n_824) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_656), .B2(n_663), .C(n_664), .Y(n_652) );
INVxp67_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVx2_ASAP7_75t_L g746 ( .A(n_659), .Y(n_746) );
BUFx2_ASAP7_75t_L g766 ( .A(n_661), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_672), .B(n_675), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_667), .B(n_670), .Y(n_666) );
AND2x2_ASAP7_75t_L g808 ( .A(n_667), .B(n_730), .Y(n_808) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g714 ( .A(n_669), .Y(n_714) );
AND2x2_ASAP7_75t_L g804 ( .A(n_669), .B(n_674), .Y(n_804) );
INVx1_ASAP7_75t_L g687 ( .A(n_671), .Y(n_687) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_680), .A2(n_681), .B(n_693), .C(n_705), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B1(n_689), .B2(n_691), .Y(n_681) );
INVx2_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_688), .Y(n_686) );
BUFx2_ASAP7_75t_L g721 ( .A(n_688), .Y(n_721) );
AND2x2_ASAP7_75t_L g814 ( .A(n_688), .B(n_756), .Y(n_814) );
OAI21xp33_ASAP7_75t_L g817 ( .A1(n_689), .A2(n_818), .B(n_820), .Y(n_817) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_696), .B1(n_700), .B2(n_702), .Y(n_693) );
HB1xp67_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_696), .B(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVxp67_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g768 ( .A(n_701), .B(n_769), .Y(n_768) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
AND2x4_ASAP7_75t_L g755 ( .A(n_704), .B(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g771 ( .A(n_704), .Y(n_771) );
AOI21xp33_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_710), .B(n_712), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
AND2x2_ASAP7_75t_L g782 ( .A(n_707), .B(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g819 ( .A(n_707), .B(n_784), .Y(n_819) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g733 ( .A(n_708), .Y(n_733) );
OR2x2_ASAP7_75t_L g811 ( .A(n_708), .B(n_812), .Y(n_811) );
OR2x2_ASAP7_75t_L g726 ( .A(n_711), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g758 ( .A(n_711), .Y(n_758) );
OR2x2_ASAP7_75t_L g791 ( .A(n_711), .B(n_792), .Y(n_791) );
INVx2_ASAP7_75t_L g762 ( .A(n_712), .Y(n_762) );
OR2x2_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NOR3xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_734), .C(n_741), .Y(n_715) );
OAI322xp33_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_720), .A3(n_722), .B1(n_724), .B2(n_726), .C1(n_728), .C2(n_732), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g793 ( .A1(n_718), .A2(n_758), .B(n_794), .C(n_797), .Y(n_793) );
BUFx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g738 ( .A(n_719), .B(n_739), .Y(n_738) );
INVx2_ASAP7_75t_L g775 ( .A(n_719), .Y(n_775) );
AND2x4_ASAP7_75t_L g803 ( .A(n_719), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AOI32xp33_ASAP7_75t_L g772 ( .A1(n_721), .A2(n_759), .A3(n_773), .B1(n_775), .B2(n_776), .Y(n_772) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g759 ( .A(n_725), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_727), .B(n_780), .Y(n_779) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
O2A1O1Ixp33_ASAP7_75t_L g741 ( .A1(n_742), .A2(n_744), .B(n_745), .C(n_746), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_SL g747 ( .A(n_748), .B(n_805), .Y(n_747) );
AOI211xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_752), .B(n_760), .C(n_785), .Y(n_748) );
INVxp67_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_SL g827 ( .A1(n_753), .A2(n_828), .B(n_829), .C(n_831), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
OAI31xp33_ASAP7_75t_L g807 ( .A1(n_755), .A2(n_808), .A3(n_809), .B(n_810), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
INVx2_ASAP7_75t_L g767 ( .A(n_759), .Y(n_767) );
NAND4xp25_ASAP7_75t_SL g760 ( .A(n_761), .B(n_764), .C(n_772), .D(n_781), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
AOI32xp33_ASAP7_75t_L g764 ( .A1(n_765), .A2(n_766), .A3(n_767), .B1(n_768), .B2(n_771), .Y(n_764) );
INVx1_ASAP7_75t_L g816 ( .A(n_768), .Y(n_816) );
INVx1_ASAP7_75t_L g828 ( .A(n_771), .Y(n_828) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_786), .B(n_793), .C(n_800), .Y(n_785) );
OAI21xp5_ASAP7_75t_SL g786 ( .A1(n_787), .A2(n_789), .B(n_790), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx3_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_794), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_803), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NOR4xp25_ASAP7_75t_L g805 ( .A(n_806), .B(n_817), .C(n_827), .D(n_832), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_807), .B(n_813), .Y(n_806) );
OAI21xp33_ASAP7_75t_L g813 ( .A1(n_808), .A2(n_814), .B(n_815), .Y(n_813) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_821), .A2(n_822), .B1(n_825), .B2(n_826), .Y(n_820) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
HB1xp67_ASAP7_75t_L g833 ( .A(n_824), .Y(n_833) );
INVxp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
BUFx6f_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
NOR2xp33_ASAP7_75t_L g842 ( .A(n_843), .B(n_844), .Y(n_842) );
INVx6_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
BUFx10_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
CKINVDCx20_ASAP7_75t_R g851 ( .A(n_852), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g852 ( .A(n_853), .Y(n_852) );
CKINVDCx20_ASAP7_75t_R g853 ( .A(n_854), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .Y(n_857) );
OR2x4_ASAP7_75t_L g863 ( .A(n_859), .B(n_864), .Y(n_863) );
BUFx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx4_ASAP7_75t_L g861 ( .A(n_862), .Y(n_861) );
BUFx3_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
endmodule