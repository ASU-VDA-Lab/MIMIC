module fake_netlist_5_1180_n_488 (n_137, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_488);

input n_137;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_488;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_451;
wire n_408;
wire n_376;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_483;
wire n_467;
wire n_423;
wire n_284;
wire n_245;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_275;
wire n_252;
wire n_295;
wire n_330;
wire n_373;
wire n_307;
wire n_439;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_191;
wire n_171;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_470;
wire n_325;
wire n_449;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_457;
wire n_297;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_192;
wire n_223;
wire n_392;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_344;
wire n_287;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_485;
wire n_355;
wire n_486;
wire n_336;
wire n_337;
wire n_430;
wire n_313;
wire n_479;
wire n_216;
wire n_168;
wire n_395;
wire n_432;
wire n_311;
wire n_208;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_468;
wire n_213;
wire n_342;
wire n_482;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_309;
wire n_462;
wire n_322;
wire n_258;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_463;
wire n_239;
wire n_466;
wire n_420;
wire n_310;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_345;
wire n_210;
wire n_365;
wire n_176;
wire n_182;
wire n_354;
wire n_480;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_410;
wire n_269;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_426;
wire n_409;
wire n_300;
wire n_435;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

INVx1_ASAP7_75t_L g168 ( 
.A(n_21),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_88),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_130),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_121),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_53),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_10),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_92),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_8),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_0),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_27),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_102),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_43),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_58),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_134),
.Y(n_193)
);

INVxp67_ASAP7_75t_SL g194 ( 
.A(n_70),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_75),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_94),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_86),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_76),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_6),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_69),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_41),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_99),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_50),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_23),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g207 ( 
.A(n_26),
.Y(n_207)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_9),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_89),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_135),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_155),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_49),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_95),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_30),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_19),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_74),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_12),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_100),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_47),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_13),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_128),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_103),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_105),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_66),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_17),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_148),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_127),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_0),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_153),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_39),
.Y(n_232)
);

INVxp33_ASAP7_75t_SL g233 ( 
.A(n_40),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_120),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_126),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_108),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_98),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_137),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_111),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_71),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_110),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_77),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_73),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_31),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_4),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_48),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_20),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_64),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_37),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_25),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_2),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_96),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_18),
.Y(n_255)
);

INVxp33_ASAP7_75t_SL g256 ( 
.A(n_42),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_104),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g258 ( 
.A(n_124),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_106),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_163),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_55),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_32),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_81),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_44),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_118),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_157),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_56),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_146),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_63),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_149),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_136),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_147),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_35),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_33),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_68),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_28),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_62),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_132),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_140),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_7),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_46),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_79),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_61),
.Y(n_283)
);

INVxp67_ASAP7_75t_SL g284 ( 
.A(n_85),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_143),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_51),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_52),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_129),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_144),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_109),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_1),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_230),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_207),
.B(n_221),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_205),
.B(n_5),
.Y(n_295)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_184),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_232),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_168),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_214),
.B(n_14),
.C(n_15),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_169),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_179),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_172),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_173),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_176),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_177),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_178),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_187),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_180),
.A2(n_16),
.B(n_22),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_181),
.Y(n_313)
);

AND2x6_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_290),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_198),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_203),
.B(n_211),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_182),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_183),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_233),
.A2(n_24),
.B1(n_29),
.B2(n_34),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_185),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_186),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_189),
.Y(n_322)
);

BUFx2_ASAP7_75t_L g323 ( 
.A(n_190),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_196),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_200),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_202),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_285),
.B(n_36),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_204),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_240),
.A2(n_38),
.B1(n_45),
.B2(n_54),
.Y(n_329)
);

INVxp33_ASAP7_75t_L g330 ( 
.A(n_206),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_212),
.B(n_224),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_210),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_213),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_216),
.B(n_57),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_265),
.B(n_59),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_256),
.A2(n_60),
.B1(n_65),
.B2(n_67),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_217),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_199),
.A2(n_72),
.B1(n_78),
.B2(n_80),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_250),
.B(n_82),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_170),
.B(n_83),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_171),
.B(n_84),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_219),
.B(n_87),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_222),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_225),
.B(n_91),
.Y(n_344)
);

NAND2xp33_ASAP7_75t_L g345 ( 
.A(n_174),
.B(n_93),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_226),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_227),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_228),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_231),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_234),
.Y(n_350)
);

AOI21x1_ASAP7_75t_L g351 ( 
.A1(n_235),
.A2(n_97),
.B(n_101),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_238),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_239),
.B(n_241),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_188),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_301),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_294),
.B(n_192),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_355),
.B(n_244),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_330),
.B(n_245),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_246),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_303),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_297),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_352),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_293),
.B(n_292),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_323),
.Y(n_365)
);

NOR3xp33_ASAP7_75t_SL g366 ( 
.A(n_354),
.B(n_272),
.C(n_269),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_309),
.Y(n_367)
);

INVx2_ASAP7_75t_SL g368 ( 
.A(n_307),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_310),
.Y(n_369)
);

OAI21xp33_ASAP7_75t_L g370 ( 
.A1(n_299),
.A2(n_289),
.B(n_247),
.Y(n_370)
);

NAND2x1p5_ASAP7_75t_L g371 ( 
.A(n_295),
.B(n_248),
.Y(n_371)
);

AND2x4_ASAP7_75t_L g372 ( 
.A(n_298),
.B(n_191),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_313),
.Y(n_373)
);

NOR3xp33_ASAP7_75t_SL g374 ( 
.A(n_316),
.B(n_193),
.C(n_255),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_296),
.B(n_262),
.Y(n_375)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_323),
.A2(n_243),
.B1(n_281),
.B2(n_276),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_318),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_327),
.B(n_331),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_335),
.B(n_252),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_320),
.Y(n_381)
);

BUFx12f_ASAP7_75t_SL g382 ( 
.A(n_349),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g383 ( 
.A(n_349),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_321),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_305),
.A2(n_236),
.B1(n_223),
.B2(n_218),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_311),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

NOR3xp33_ASAP7_75t_SL g388 ( 
.A(n_342),
.B(n_242),
.C(n_263),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_334),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_314),
.B(n_273),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_337),
.Y(n_391)
);

AND3x2_ASAP7_75t_SL g392 ( 
.A(n_343),
.B(n_251),
.C(n_220),
.Y(n_392)
);

AND2x6_ASAP7_75t_SL g393 ( 
.A(n_344),
.B(n_288),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_315),
.B(n_338),
.Y(n_394)
);

AO31x2_ASAP7_75t_L g395 ( 
.A1(n_378),
.A2(n_346),
.A3(n_308),
.B(n_348),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_314),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_380),
.A2(n_312),
.B(n_351),
.Y(n_397)
);

OAI21x1_ASAP7_75t_L g398 ( 
.A1(n_371),
.A2(n_339),
.B(n_341),
.Y(n_398)
);

INVx3_ASAP7_75t_SL g399 ( 
.A(n_386),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_368),
.B(n_365),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_314),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_357),
.B(n_306),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_389),
.B(n_253),
.Y(n_403)
);

O2A1O1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_317),
.B(n_322),
.C(n_347),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_372),
.B(n_270),
.Y(n_405)
);

AOI31xp33_ASAP7_75t_L g406 ( 
.A1(n_376),
.A2(n_319),
.A3(n_336),
.B(n_329),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_364),
.A2(n_345),
.B(n_340),
.Y(n_407)
);

A2O1A1Ixp33_ASAP7_75t_L g408 ( 
.A1(n_359),
.A2(n_328),
.B(n_326),
.C(n_302),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_361),
.B(n_353),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_383),
.Y(n_410)
);

OAI21x1_ASAP7_75t_L g411 ( 
.A1(n_390),
.A2(n_350),
.B(n_333),
.Y(n_411)
);

AOI221xp5_ASAP7_75t_SL g412 ( 
.A1(n_370),
.A2(n_268),
.B1(n_254),
.B2(n_257),
.C(n_287),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_381),
.Y(n_413)
);

AOI21x1_ASAP7_75t_L g414 ( 
.A1(n_360),
.A2(n_249),
.B(n_259),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_362),
.B(n_332),
.Y(n_416)
);

AOI211x1_ASAP7_75t_L g417 ( 
.A1(n_367),
.A2(n_275),
.B(n_260),
.C(n_286),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_324),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_375),
.A2(n_271),
.B(n_284),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_385),
.B(n_304),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g421 ( 
.A1(n_356),
.A2(n_194),
.B(n_267),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_369),
.B(n_283),
.Y(n_422)
);

AND3x1_ASAP7_75t_L g423 ( 
.A(n_366),
.B(n_282),
.C(n_279),
.Y(n_423)
);

INVxp67_ASAP7_75t_SL g424 ( 
.A(n_413),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_407),
.A2(n_208),
.B(n_215),
.Y(n_425)
);

AOI21x1_ASAP7_75t_SL g426 ( 
.A1(n_396),
.A2(n_388),
.B(n_392),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_402),
.B(n_374),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_406),
.A2(n_258),
.B1(n_266),
.B2(n_264),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_395),
.B(n_391),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_409),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_401),
.A2(n_384),
.B(n_377),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_395),
.B(n_420),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_416),
.Y(n_434)
);

AOI21x1_ASAP7_75t_SL g435 ( 
.A1(n_422),
.A2(n_393),
.B(n_277),
.Y(n_435)
);

O2A1O1Ixp5_ASAP7_75t_L g436 ( 
.A1(n_419),
.A2(n_278),
.B(n_373),
.C(n_363),
.Y(n_436)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_261),
.B(n_229),
.Y(n_437)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_405),
.A2(n_209),
.B1(n_201),
.B2(n_197),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_404),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_195),
.B1(n_382),
.B2(n_114),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_421),
.A2(n_112),
.B(n_113),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_427),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_434),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_395),
.Y(n_445)
);

INVxp67_ASAP7_75t_SL g446 ( 
.A(n_424),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_410),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_430),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_418),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_399),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_433),
.B(n_400),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_432),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_437),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_439),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_443),
.Y(n_457)
);

NAND3xp33_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_423),
.C(n_441),
.Y(n_458)
);

INVx4_ASAP7_75t_L g459 ( 
.A(n_447),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_447),
.Y(n_460)
);

INVx4_ASAP7_75t_SL g461 ( 
.A(n_450),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_445),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_448),
.Y(n_465)
);

AND2x4_ASAP7_75t_L g466 ( 
.A(n_453),
.B(n_398),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_459),
.B(n_451),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_465),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_464),
.B(n_456),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_463),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_457),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_462),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_469),
.A2(n_458),
.B1(n_461),
.B2(n_460),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_467),
.A2(n_466),
.B1(n_452),
.B2(n_425),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_468),
.Y(n_475)
);

OAI21xp33_ASAP7_75t_L g476 ( 
.A1(n_473),
.A2(n_472),
.B(n_471),
.Y(n_476)
);

AOI32xp33_ASAP7_75t_L g477 ( 
.A1(n_475),
.A2(n_470),
.A3(n_435),
.B1(n_426),
.B2(n_454),
.Y(n_477)
);

AOI221xp5_ASAP7_75t_L g478 ( 
.A1(n_474),
.A2(n_442),
.B1(n_417),
.B2(n_412),
.C(n_455),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_477),
.Y(n_479)
);

NAND3xp33_ASAP7_75t_L g480 ( 
.A(n_476),
.B(n_437),
.C(n_414),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_479),
.B(n_116),
.Y(n_481)
);

AND2x2_ASAP7_75t_SL g482 ( 
.A(n_480),
.B(n_478),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_482),
.Y(n_483)
);

OAI322xp33_ASAP7_75t_L g484 ( 
.A1(n_481),
.A2(n_119),
.A3(n_123),
.B1(n_125),
.B2(n_131),
.C1(n_138),
.C2(n_150),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_483),
.B(n_151),
.Y(n_485)
);

OAI21x1_ASAP7_75t_SL g486 ( 
.A1(n_485),
.A2(n_484),
.B(n_154),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_486),
.A2(n_411),
.B(n_156),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_487),
.A2(n_152),
.B1(n_164),
.B2(n_165),
.Y(n_488)
);


endmodule