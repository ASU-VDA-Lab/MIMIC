module real_jpeg_23072_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_1),
.A2(n_34),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_1),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_70),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_54),
.B1(n_55),
.B2(n_70),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_1),
.A2(n_39),
.B1(n_43),
.B2(n_70),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_2),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_3),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_44),
.B1(n_54),
.B2(n_55),
.Y(n_98)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_62),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_5),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_5),
.A2(n_62),
.B1(n_78),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_62),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_5),
.A2(n_39),
.B1(n_43),
.B2(n_62),
.Y(n_200)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_8),
.A2(n_39),
.B1(n_43),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_8),
.Y(n_85)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_10),
.A2(n_65),
.B1(n_77),
.B2(n_78),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_10),
.A2(n_54),
.B1(n_55),
.B2(n_65),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_39),
.B1(n_43),
.B2(n_65),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_11),
.A2(n_54),
.B1(n_55),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_11),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_97),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_11),
.A2(n_39),
.B1(n_43),
.B2(n_97),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_12),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_12),
.B(n_73),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_55),
.C(n_57),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_109),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_12),
.B(n_66),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_12),
.A2(n_54),
.B1(n_55),
.B2(n_109),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_12),
.B(n_39),
.C(n_93),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_12),
.A2(n_38),
.B(n_201),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_14),
.A2(n_39),
.B1(n_43),
.B2(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_14),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_15),
.A2(n_39),
.B1(n_43),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_15),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_124)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_16),
.Y(n_88)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_16),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_141),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_140),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_112),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_21),
.B(n_112),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_99),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_22),
.B(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_50),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_23),
.B(n_51),
.C(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_24),
.B(n_36),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.A3(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_25),
.A2(n_26),
.B1(n_57),
.B2(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_73)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_26),
.B(n_32),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_26),
.B(n_167),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_29),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_78),
.Y(n_80)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp33_ASAP7_75t_L g110 ( 
.A(n_33),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_45),
.B2(n_48),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_37),
.A2(n_121),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_38),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_38),
.A2(n_84),
.B1(n_118),
.B2(n_120),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_38),
.A2(n_42),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_38),
.B(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_38),
.A2(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_39),
.A2(n_43),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_40),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_43),
.B(n_225),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_45),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_67),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_60),
.B(n_63),
.Y(n_51)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_52),
.A2(n_63),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_53),
.A2(n_137),
.B(n_138),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_53),
.A2(n_138),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_54),
.A2(n_55),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_55),
.B(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_66),
.B1(n_105),
.B2(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_64),
.B(n_106),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_72),
.B(n_74),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_69),
.A2(n_73),
.B1(n_79),
.B2(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_72),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_76),
.Y(n_111)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_79),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_79),
.A2(n_108),
.B(n_111),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_81),
.B(n_99),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_89),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_82),
.B(n_89),
.Y(n_139)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_88),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_88),
.B(n_109),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_95),
.B1(n_96),
.B2(n_98),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_90),
.A2(n_188),
.B(n_189),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_90),
.A2(n_189),
.B(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_91),
.B(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_91),
.A2(n_125),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_96),
.B(n_102),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_95),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_95),
.A2(n_102),
.B(n_174),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_95),
.B(n_109),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.C(n_107),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_103),
.B(n_125),
.Y(n_189)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_105),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_116),
.B1(n_128),
.B2(n_129),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_117),
.A2(n_122),
.B1(n_126),
.B2(n_127),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_139),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_243),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_161),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_159),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_145),
.B(n_159),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_146),
.A2(n_147),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_150),
.B(n_151),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_156),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_152),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_183),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_156),
.Y(n_183)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_158),
.A2(n_214),
.B(n_222),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_237),
.B(n_242),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_190),
.B(n_236),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_179),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_164),
.B(n_179),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_172),
.C(n_176),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_168),
.Y(n_186)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_172),
.A2(n_176),
.B1(n_177),
.B2(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_172),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_186),
.C(n_187),
.Y(n_241)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_230),
.B(n_235),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_210),
.B(n_229),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_204),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_204),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_199),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_234)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_208),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_218),
.B(n_228),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_216),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_216),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_223),
.B(n_227),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_221),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_231),
.B(n_234),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_231),
.B(n_234),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_241),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_241),
.Y(n_242)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);


endmodule