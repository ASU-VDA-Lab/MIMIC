module fake_ibex_994_n_1702 (n_151, n_85, n_84, n_64, n_171, n_103, n_204, n_274, n_130, n_177, n_76, n_273, n_309, n_9, n_293, n_124, n_37, n_256, n_193, n_108, n_165, n_86, n_70, n_255, n_175, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_312, n_239, n_94, n_134, n_88, n_142, n_226, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_15, n_24, n_189, n_280, n_317, n_105, n_187, n_1, n_154, n_182, n_196, n_89, n_50, n_144, n_170, n_270, n_113, n_117, n_265, n_158, n_259, n_276, n_210, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_244, n_73, n_310, n_143, n_106, n_8, n_224, n_183, n_67, n_110, n_306, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_60, n_7, n_109, n_127, n_121, n_48, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_0, n_289, n_12, n_150, n_286, n_133, n_51, n_215, n_279, n_49, n_235, n_22, n_136, n_261, n_30, n_221, n_102, n_52, n_99, n_269, n_156, n_126, n_25, n_104, n_45, n_141, n_222, n_186, n_295, n_230, n_96, n_185, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_82, n_263, n_27, n_299, n_87, n_262, n_75, n_137, n_173, n_180, n_201, n_14, n_257, n_77, n_44, n_66, n_305, n_307, n_192, n_140, n_4, n_6, n_100, n_179, n_206, n_26, n_188, n_200, n_199, n_308, n_135, n_283, n_111, n_36, n_18, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_214, n_238, n_211, n_218, n_314, n_132, n_277, n_225, n_272, n_23, n_223, n_95, n_285, n_288, n_247, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_233, n_118, n_164, n_38, n_198, n_264, n_217, n_78, n_20, n_69, n_39, n_178, n_303, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_119, n_72, n_195, n_212, n_311, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_297, n_41, n_252, n_83, n_32, n_107, n_149, n_254, n_213, n_271, n_241, n_68, n_292, n_79, n_81, n_35, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_281, n_1702);

input n_151;
input n_85;
input n_84;
input n_64;
input n_171;
input n_103;
input n_204;
input n_274;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_9;
input n_293;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_312;
input n_239;
input n_94;
input n_134;
input n_88;
input n_142;
input n_226;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_210;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_244;
input n_73;
input n_310;
input n_143;
input n_106;
input n_8;
input n_224;
input n_183;
input n_67;
input n_110;
input n_306;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_221;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_295;
input n_230;
input n_96;
input n_185;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_82;
input n_263;
input n_27;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_173;
input n_180;
input n_201;
input n_14;
input n_257;
input n_77;
input n_44;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_4;
input n_6;
input n_100;
input n_179;
input n_206;
input n_26;
input n_188;
input n_200;
input n_199;
input n_308;
input n_135;
input n_283;
input n_111;
input n_36;
input n_18;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_214;
input n_238;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_225;
input n_272;
input n_23;
input n_223;
input n_95;
input n_285;
input n_288;
input n_247;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_233;
input n_118;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_78;
input n_20;
input n_69;
input n_39;
input n_178;
input n_303;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_119;
input n_72;
input n_195;
input n_212;
input n_311;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_297;
input n_41;
input n_252;
input n_83;
input n_32;
input n_107;
input n_149;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_79;
input n_81;
input n_35;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_281;

output n_1702;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_452;
wire n_1234;
wire n_1594;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_678;
wire n_969;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_872;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1614;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_500;
wire n_963;
wire n_376;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_375;
wire n_1391;
wire n_667;
wire n_884;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_346;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_504;
wire n_948;
wire n_1338;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_671;
wire n_989;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_550;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_441;
wire n_694;
wire n_523;
wire n_787;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_321;
wire n_1081;
wire n_374;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_904;
wire n_355;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1618;
wire n_1648;
wire n_857;
wire n_765;
wire n_1070;
wire n_777;
wire n_331;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_352;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_359;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_338;
wire n_1401;
wire n_369;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1252;
wire n_1170;
wire n_605;
wire n_539;
wire n_630;
wire n_567;
wire n_745;
wire n_447;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_397;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_1326;
wire n_971;
wire n_451;
wire n_1350;
wire n_906;
wire n_1093;
wire n_978;
wire n_579;
wire n_899;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_382;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_379;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1609;
wire n_324;
wire n_391;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_390;
wire n_1467;
wire n_544;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_870;
wire n_1610;
wire n_1298;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_345;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_406;
wire n_606;
wire n_737;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1003;
wire n_889;
wire n_435;
wire n_396;
wire n_816;
wire n_1058;
wire n_399;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1441;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_743;
wire n_754;
wire n_395;
wire n_1319;
wire n_389;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_330;
wire n_1182;
wire n_1271;
wire n_1031;
wire n_372;
wire n_981;
wire n_350;
wire n_398;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_371;
wire n_974;
wire n_1036;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1634;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1189;
wire n_761;
wire n_748;
wire n_901;
wire n_1577;
wire n_340;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_471;
wire n_846;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_384;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1032;
wire n_936;
wire n_469;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1510;
wire n_1201;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_590;
wire n_1568;
wire n_325;
wire n_1184;
wire n_1477;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1075;
wire n_1249;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_669;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_388;
wire n_1522;
wire n_1279;
wire n_931;
wire n_607;
wire n_827;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1146;
wire n_358;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_472;
wire n_347;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_363;
wire n_1628;
wire n_725;
wire n_596;
wire n_1545;
wire n_351;
wire n_456;
wire n_1471;
wire n_998;
wire n_1115;
wire n_1395;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_365;
wire n_814;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1470;
wire n_444;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1599;
wire n_650;
wire n_409;
wire n_1575;
wire n_332;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_337;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_633;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_486;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_344;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_380;
wire n_947;
wire n_1004;
wire n_831;
wire n_778;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_328;
wire n_418;
wire n_510;
wire n_972;
wire n_601;
wire n_610;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_545;
wire n_887;
wire n_1162;
wire n_334;
wire n_634;
wire n_961;
wire n_991;
wire n_1223;
wire n_1331;
wire n_1349;
wire n_1323;
wire n_578;
wire n_432;
wire n_403;
wire n_1353;
wire n_423;
wire n_357;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1286;
wire n_1657;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_377;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_326;
wire n_1629;
wire n_1662;
wire n_1340;
wire n_339;
wire n_348;
wire n_1626;
wire n_674;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_400;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_404;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_719;
wire n_370;
wire n_1491;
wire n_716;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1037;
wire n_464;
wire n_1289;
wire n_838;
wire n_1348;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1587;
wire n_636;
wire n_1259;
wire n_407;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_356;
wire n_1538;
wire n_487;
wire n_349;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_851;
wire n_993;
wire n_1135;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_353;
wire n_1604;
wire n_1639;
wire n_826;
wire n_1337;
wire n_1647;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_402;
wire n_1415;
wire n_1238;
wire n_976;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_804;
wire n_1455;
wire n_484;
wire n_1642;
wire n_480;
wire n_354;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_329;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_624;
wire n_463;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_360;
wire n_1107;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_320;
wire n_1411;
wire n_1139;
wire n_858;
wire n_1018;
wire n_385;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_833;
wire n_1343;
wire n_1371;
wire n_1513;
wire n_728;
wire n_786;
wire n_362;
wire n_505;
wire n_1621;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_393;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1060;
wire n_1372;
wire n_756;
wire n_1565;
wire n_1257;
wire n_387;
wire n_1632;
wire n_688;
wire n_1547;
wire n_946;
wire n_1542;
wire n_707;
wire n_1362;
wire n_1586;
wire n_1097;
wire n_341;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_593;
wire n_1212;
wire n_1199;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1564;
wire n_1631;
wire n_336;
wire n_1623;
wire n_861;
wire n_1389;
wire n_1131;
wire n_547;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_828;
wire n_1438;
wire n_753;
wire n_645;
wire n_747;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_327;
wire n_1302;
wire n_383;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1572;
wire n_1635;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_373;
wire n_854;
wire n_343;
wire n_714;
wire n_1297;
wire n_1369;
wire n_323;
wire n_740;
wire n_386;
wire n_549;
wire n_533;
wire n_928;
wire n_898;
wire n_333;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1597;
wire n_1103;
wire n_1161;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_367;
wire n_880;
wire n_654;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_689;
wire n_960;
wire n_1022;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1020;
wire n_783;
wire n_1142;
wire n_1385;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_335;
wire n_1499;
wire n_1500;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_699;
wire n_368;
wire n_918;
wire n_672;
wire n_1039;
wire n_401;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_581;
wire n_416;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_392;
wire n_1536;
wire n_1049;
wire n_548;
wire n_1158;
wire n_763;
wire n_940;
wire n_1404;
wire n_546;
wire n_788;
wire n_410;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1026;
wire n_366;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_322;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_653;
wire n_1205;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_511;
wire n_381;
wire n_1414;
wire n_1002;
wire n_1111;
wire n_1341;
wire n_405;
wire n_1310;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_342;
wire n_414;
wire n_378;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_519;
wire n_408;
wire n_361;
wire n_1665;
wire n_319;
wire n_1091;
wire n_1678;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_661;
wire n_848;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_1674;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_394;
wire n_364;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_492;
wire n_649;
wire n_866;
wire n_559;
wire n_425;

HB1xp67_ASAP7_75t_L g319 ( 
.A(n_210),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_238),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_65),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_291),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_241),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_113),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_75),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_158),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_287),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_35),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_242),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_264),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_299),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_37),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_195),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_307),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_30),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_266),
.Y(n_337)
);

INVx1_ASAP7_75t_SL g338 ( 
.A(n_95),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_34),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_268),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_278),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_61),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_165),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_0),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_106),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_59),
.Y(n_346)
);

BUFx10_ASAP7_75t_L g347 ( 
.A(n_239),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_286),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_114),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_181),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_137),
.Y(n_351)
);

CKINVDCx11_ASAP7_75t_R g352 ( 
.A(n_230),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g354 ( 
.A(n_54),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_38),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_96),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_309),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_1),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_196),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_259),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_171),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_223),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_273),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_80),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_127),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_209),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_315),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_216),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_219),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_290),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_77),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_274),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_141),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_314),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_213),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_142),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_159),
.Y(n_378)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_31),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_189),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_221),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_302),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_117),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_151),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_318),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_275),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_211),
.Y(n_387)
);

BUFx10_ASAP7_75t_L g388 ( 
.A(n_214),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_218),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_316),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_99),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_85),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_166),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_222),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_243),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_306),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_310),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_253),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_202),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_160),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_280),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_188),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_10),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_89),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_312),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_108),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_261),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_89),
.Y(n_408)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_187),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_226),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_78),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_207),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_301),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_67),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_277),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_244),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_60),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_185),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_305),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_162),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_38),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_276),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_265),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_28),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_251),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_245),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_4),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_249),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_283),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_267),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_49),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_145),
.Y(n_432)
);

CKINVDCx16_ASAP7_75t_R g433 ( 
.A(n_93),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_97),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_5),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_228),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_47),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_161),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_254),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_13),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_10),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_101),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_132),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_212),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_17),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_169),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g447 ( 
.A(n_146),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_231),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_197),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_46),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_82),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_12),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_300),
.Y(n_453)
);

CKINVDCx14_ASAP7_75t_R g454 ( 
.A(n_317),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_257),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_206),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_263),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_49),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_118),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_6),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_260),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_148),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_37),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_282),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_236),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_272),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_23),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_182),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_80),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_269),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_76),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_220),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_34),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_57),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_144),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_289),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_156),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_15),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_247),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_296),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_48),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_48),
.Y(n_482)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_186),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_126),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_191),
.Y(n_485)
);

BUFx2_ASAP7_75t_R g486 ( 
.A(n_58),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_1),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_234),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_82),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_139),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_17),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_198),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_298),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_233),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_224),
.Y(n_495)
);

INVx1_ASAP7_75t_SL g496 ( 
.A(n_217),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_313),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_88),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_26),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_285),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_225),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_281),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_240),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_271),
.Y(n_504)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_297),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_86),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_65),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_13),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_94),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_75),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_53),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_295),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_57),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_119),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_255),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_270),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_246),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_120),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_130),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_258),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_96),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_174),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_227),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_279),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_27),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_92),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_288),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_55),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_256),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_248),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_293),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_215),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_54),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_9),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_304),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_14),
.Y(n_536)
);

INVx4_ASAP7_75t_R g537 ( 
.A(n_131),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_262),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_111),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_31),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_237),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_7),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_308),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_205),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_232),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_235),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_67),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_292),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_204),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_252),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_250),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_294),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_229),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_110),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_91),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_319),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_352),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_349),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_383),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_351),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_502),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_433),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_359),
.Y(n_563)
);

INVxp67_ASAP7_75t_SL g564 ( 
.A(n_391),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_447),
.Y(n_565)
);

CKINVDCx20_ASAP7_75t_R g566 ( 
.A(n_421),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_391),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_408),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_329),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_374),
.B(n_0),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_329),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_417),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_472),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_480),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_417),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_520),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_554),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_389),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_354),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_354),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_427),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_445),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_354),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_478),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_322),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_405),
.B(n_2),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_354),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_354),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_354),
.Y(n_590)
);

NOR2xp67_ASAP7_75t_L g591 ( 
.A(n_326),
.B(n_2),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_379),
.Y(n_592)
);

INVxp33_ASAP7_75t_SL g593 ( 
.A(n_333),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_379),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_508),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_339),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_379),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_379),
.Y(n_598)
);

BUFx2_ASAP7_75t_SL g599 ( 
.A(n_347),
.Y(n_599)
);

INVxp67_ASAP7_75t_SL g600 ( 
.A(n_442),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_379),
.Y(n_601)
);

INVxp67_ASAP7_75t_SL g602 ( 
.A(n_509),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_379),
.Y(n_603)
);

NOR2xp67_ASAP7_75t_L g604 ( 
.A(n_336),
.B(n_3),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_404),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_342),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_414),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_454),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_437),
.Y(n_609)
);

CKINVDCx20_ASAP7_75t_R g610 ( 
.A(n_344),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_346),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_355),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_440),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_441),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_469),
.Y(n_615)
);

CKINVDCx14_ASAP7_75t_R g616 ( 
.A(n_347),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_358),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_473),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_555),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_488),
.B(n_3),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_482),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_364),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_392),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_403),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_411),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

NOR2xp67_ASAP7_75t_L g627 ( 
.A(n_499),
.B(n_4),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_424),
.Y(n_628)
);

INVxp67_ASAP7_75t_SL g629 ( 
.A(n_513),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_431),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_533),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_353),
.B(n_5),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_434),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_540),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_435),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_451),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_590),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_556),
.B(n_547),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_590),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_566),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_600),
.B(n_353),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_566),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_568),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_557),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_569),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_580),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_558),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_R g648 ( 
.A(n_616),
.B(n_324),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_570),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_581),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_563),
.B(n_320),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_565),
.B(n_320),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_636),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_582),
.Y(n_654)
);

CKINVDCx20_ASAP7_75t_R g655 ( 
.A(n_582),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_560),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_584),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_588),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_R g659 ( 
.A(n_608),
.B(n_325),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_589),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_625),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_574),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_602),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_559),
.B(n_388),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_575),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

NOR2xp67_ASAP7_75t_L g667 ( 
.A(n_609),
.B(n_321),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_592),
.Y(n_668)
);

XOR2xp5_ASAP7_75t_L g669 ( 
.A(n_562),
.B(n_486),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_573),
.Y(n_670)
);

CKINVDCx20_ASAP7_75t_R g671 ( 
.A(n_583),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_594),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_598),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_R g675 ( 
.A(n_608),
.B(n_327),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_577),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_564),
.B(n_363),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_601),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g679 ( 
.A(n_610),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_603),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_576),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_578),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_561),
.B(n_372),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_567),
.B(n_363),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_605),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_607),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_614),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_599),
.B(n_388),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_615),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_593),
.B(n_330),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_618),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_586),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_610),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_631),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_611),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_634),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_613),
.Y(n_698)
);

NAND2xp33_ASAP7_75t_L g699 ( 
.A(n_579),
.B(n_332),
.Y(n_699)
);

INVx3_ASAP7_75t_L g700 ( 
.A(n_632),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_621),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_629),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_611),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_604),
.Y(n_704)
);

BUFx6f_ASAP7_75t_L g705 ( 
.A(n_571),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_627),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_593),
.B(n_553),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_617),
.Y(n_708)
);

INVx5_ASAP7_75t_L g709 ( 
.A(n_587),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_620),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_635),
.B(n_373),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_635),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_596),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_SL g714 ( 
.A(n_636),
.B(n_452),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_R g715 ( 
.A(n_606),
.B(n_458),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_591),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_612),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_619),
.Y(n_718)
);

CKINVDCx20_ASAP7_75t_R g719 ( 
.A(n_583),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_617),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_622),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_623),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_628),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_624),
.B(n_323),
.Y(n_724)
);

INVx3_ASAP7_75t_L g725 ( 
.A(n_630),
.Y(n_725)
);

XOR2xp5_ASAP7_75t_L g726 ( 
.A(n_562),
.B(n_460),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_633),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_628),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_585),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_585),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_595),
.B(n_553),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_595),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_556),
.B(n_337),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_636),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_636),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_590),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_590),
.Y(n_737)
);

BUFx2_ASAP7_75t_L g738 ( 
.A(n_636),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_568),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_557),
.Y(n_740)
);

INVx6_ASAP7_75t_L g741 ( 
.A(n_632),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_564),
.B(n_373),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_568),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_R g744 ( 
.A(n_557),
.B(n_340),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_568),
.Y(n_745)
);

HB1xp67_ASAP7_75t_L g746 ( 
.A(n_625),
.Y(n_746)
);

CKINVDCx20_ASAP7_75t_R g747 ( 
.A(n_566),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_568),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_564),
.B(n_386),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_590),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_557),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_557),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_568),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_568),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_557),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_557),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_590),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_590),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_568),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_557),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_557),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_566),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_556),
.B(n_372),
.Y(n_763)
);

CKINVDCx20_ASAP7_75t_R g764 ( 
.A(n_566),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_557),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_564),
.B(n_386),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_568),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_557),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_568),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_590),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_590),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_568),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_564),
.B(n_401),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_566),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_563),
.B(n_401),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_556),
.B(n_343),
.Y(n_776)
);

INVx3_ASAP7_75t_L g777 ( 
.A(n_590),
.Y(n_777)
);

AND2x4_ASAP7_75t_L g778 ( 
.A(n_556),
.B(n_372),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_557),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_557),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_590),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_568),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_564),
.B(n_407),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_636),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_590),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_590),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_R g787 ( 
.A(n_644),
.B(n_463),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_649),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_638),
.B(n_338),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_746),
.Y(n_790)
);

INVxp67_ASAP7_75t_SL g791 ( 
.A(n_746),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_741),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_R g793 ( 
.A(n_740),
.B(n_467),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_683),
.Y(n_794)
);

NAND2x1p5_ASAP7_75t_L g795 ( 
.A(n_713),
.B(n_356),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_741),
.Y(n_796)
);

AND2x6_ASAP7_75t_L g797 ( 
.A(n_713),
.B(n_335),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_683),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_653),
.B(n_372),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_661),
.B(n_471),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_763),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_638),
.B(n_507),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_663),
.B(n_378),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_663),
.B(n_409),
.Y(n_804)
);

INVx4_ASAP7_75t_SL g805 ( 
.A(n_722),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_661),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_649),
.Y(n_807)
);

NAND2xp33_ASAP7_75t_SL g808 ( 
.A(n_648),
.B(n_474),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_705),
.B(n_345),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_700),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_698),
.A2(n_528),
.B1(n_450),
.B2(n_331),
.Y(n_811)
);

INVx1_ASAP7_75t_SL g812 ( 
.A(n_712),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_763),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_649),
.Y(n_814)
);

AO22x2_ASAP7_75t_L g815 ( 
.A1(n_669),
.A2(n_726),
.B1(n_732),
.B2(n_728),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_734),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_710),
.B(n_348),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_687),
.B(n_350),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_701),
.A2(n_481),
.B1(n_489),
.B2(n_487),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_778),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_778),
.Y(n_821)
);

AOI22xp33_ASAP7_75t_L g822 ( 
.A1(n_702),
.A2(n_686),
.B1(n_692),
.B2(n_685),
.Y(n_822)
);

INVx3_ASAP7_75t_L g823 ( 
.A(n_666),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_666),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_666),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_735),
.B(n_491),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_670),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_670),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_705),
.B(n_690),
.Y(n_829)
);

INVx3_ASAP7_75t_L g830 ( 
.A(n_670),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_645),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_645),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_643),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_679),
.B(n_506),
.Y(n_834)
);

OR2x6_ASAP7_75t_L g835 ( 
.A(n_738),
.B(n_450),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_784),
.B(n_641),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_739),
.Y(n_837)
);

INVx5_ASAP7_75t_L g838 ( 
.A(n_736),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_743),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_681),
.Y(n_840)
);

AND2x6_ASAP7_75t_L g841 ( 
.A(n_725),
.B(n_335),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_640),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_700),
.B(n_510),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_736),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_724),
.B(n_511),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_725),
.B(n_521),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_736),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_715),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_750),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_733),
.B(n_426),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_695),
.Y(n_851)
);

NAND2x1p5_ASAP7_75t_L g852 ( 
.A(n_722),
.B(n_727),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_689),
.B(n_357),
.Y(n_853)
);

BUFx3_ASAP7_75t_L g854 ( 
.A(n_722),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_750),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_750),
.Y(n_856)
);

BUFx6f_ASAP7_75t_L g857 ( 
.A(n_771),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_771),
.Y(n_858)
);

AND2x6_ASAP7_75t_L g859 ( 
.A(n_664),
.B(n_455),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_688),
.B(n_525),
.Y(n_860)
);

AND2x4_ASAP7_75t_L g861 ( 
.A(n_717),
.B(n_526),
.Y(n_861)
);

AND2x6_ASAP7_75t_L g862 ( 
.A(n_727),
.B(n_455),
.Y(n_862)
);

INVx4_ASAP7_75t_L g863 ( 
.A(n_727),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_771),
.Y(n_864)
);

BUFx10_ASAP7_75t_L g865 ( 
.A(n_751),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_757),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_691),
.B(n_360),
.Y(n_867)
);

AND2x6_ASAP7_75t_L g868 ( 
.A(n_718),
.B(n_476),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_745),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_697),
.B(n_361),
.Y(n_870)
);

INVx5_ASAP7_75t_L g871 ( 
.A(n_757),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_721),
.B(n_534),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_777),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_711),
.B(n_677),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_752),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_705),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_748),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_711),
.B(n_362),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_755),
.Y(n_879)
);

BUFx3_ASAP7_75t_L g880 ( 
.A(n_756),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_753),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_776),
.B(n_438),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_777),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_707),
.B(n_483),
.Y(n_884)
);

AOI22xp33_ASAP7_75t_L g885 ( 
.A1(n_651),
.A2(n_528),
.B1(n_450),
.B2(n_341),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_754),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_759),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_677),
.B(n_684),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_690),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_741),
.B(n_536),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_716),
.B(n_476),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_767),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_667),
.B(n_542),
.Y(n_893)
);

BUFx6f_ASAP7_75t_L g894 ( 
.A(n_769),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_772),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_709),
.B(n_365),
.Y(n_896)
);

INVxp67_ASAP7_75t_SL g897 ( 
.A(n_684),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_709),
.B(n_366),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_744),
.B(n_450),
.Y(n_899)
);

AND2x4_ASAP7_75t_L g900 ( 
.A(n_704),
.B(n_505),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_742),
.B(n_369),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_782),
.Y(n_902)
);

INVx4_ASAP7_75t_L g903 ( 
.A(n_657),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_742),
.B(n_370),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_749),
.B(n_371),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_709),
.B(n_496),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_693),
.B(n_528),
.Y(n_907)
);

INVxp33_ASAP7_75t_L g908 ( 
.A(n_659),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_749),
.Y(n_909)
);

INVx1_ASAP7_75t_SL g910 ( 
.A(n_694),
.Y(n_910)
);

INVx2_ASAP7_75t_SL g911 ( 
.A(n_766),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_637),
.Y(n_912)
);

NOR3xp33_ASAP7_75t_SL g913 ( 
.A(n_647),
.B(n_381),
.C(n_377),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_639),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_714),
.A2(n_367),
.B1(n_368),
.B2(n_328),
.Y(n_915)
);

AND2x2_ASAP7_75t_SL g916 ( 
.A(n_728),
.B(n_528),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_737),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_696),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_758),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_766),
.Y(n_920)
);

INVx8_ASAP7_75t_L g921 ( 
.A(n_760),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_703),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_770),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_708),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_773),
.B(n_382),
.Y(n_925)
);

INVx4_ASAP7_75t_L g926 ( 
.A(n_660),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_709),
.B(n_384),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_706),
.B(n_505),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_675),
.B(n_385),
.Y(n_929)
);

BUFx4f_ASAP7_75t_L g930 ( 
.A(n_761),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_773),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_783),
.B(n_651),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_786),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_783),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_781),
.Y(n_935)
);

BUFx4f_ASAP7_75t_L g936 ( 
.A(n_765),
.Y(n_936)
);

AND2x6_ASAP7_75t_L g937 ( 
.A(n_652),
.B(n_375),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_785),
.Y(n_938)
);

CKINVDCx20_ASAP7_75t_R g939 ( 
.A(n_642),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_652),
.B(n_387),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_775),
.B(n_376),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_775),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_768),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_699),
.A2(n_380),
.B1(n_393),
.B2(n_390),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_731),
.B(n_394),
.Y(n_945)
);

INVx3_ASAP7_75t_L g946 ( 
.A(n_668),
.Y(n_946)
);

OAI22xp33_ASAP7_75t_L g947 ( 
.A1(n_656),
.A2(n_399),
.B1(n_402),
.B2(n_398),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_646),
.B(n_395),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_672),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_720),
.B(n_6),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_662),
.B(n_552),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_779),
.B(n_396),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_723),
.Y(n_953)
);

NOR2x1p5_ASAP7_75t_L g954 ( 
.A(n_780),
.B(n_397),
.Y(n_954)
);

NOR2xp33_ASAP7_75t_L g955 ( 
.A(n_650),
.B(n_400),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_673),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_658),
.B(n_410),
.Y(n_957)
);

BUFx10_ASAP7_75t_L g958 ( 
.A(n_665),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_676),
.B(n_416),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_674),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_682),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_654),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_678),
.Y(n_963)
);

OR2x6_ASAP7_75t_L g964 ( 
.A(n_655),
.B(n_413),
.Y(n_964)
);

BUFx10_ASAP7_75t_L g965 ( 
.A(n_729),
.Y(n_965)
);

AND2x4_ASAP7_75t_L g966 ( 
.A(n_680),
.B(n_415),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_671),
.B(n_420),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_719),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_730),
.Y(n_969)
);

NAND2xp33_ASAP7_75t_L g970 ( 
.A(n_747),
.B(n_422),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_762),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_764),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_774),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_683),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_746),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_649),
.Y(n_976)
);

AND2x2_ASAP7_75t_SL g977 ( 
.A(n_653),
.B(n_418),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_638),
.B(n_419),
.Y(n_978)
);

NOR2x1p5_ASAP7_75t_L g979 ( 
.A(n_644),
.B(n_423),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_649),
.Y(n_980)
);

INVx4_ASAP7_75t_L g981 ( 
.A(n_683),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_645),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_683),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_663),
.B(n_428),
.Y(n_984)
);

INVx2_ASAP7_75t_SL g985 ( 
.A(n_746),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_683),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_663),
.B(n_429),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_746),
.B(n_430),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_663),
.B(n_439),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_649),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_649),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_649),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_705),
.B(n_443),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_683),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_663),
.B(n_444),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_746),
.B(n_453),
.Y(n_996)
);

NAND3x1_ASAP7_75t_L g997 ( 
.A(n_728),
.B(n_432),
.C(n_425),
.Y(n_997)
);

INVx2_ASAP7_75t_SL g998 ( 
.A(n_746),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_683),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_683),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_663),
.B(n_461),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_649),
.Y(n_1002)
);

BUFx10_ASAP7_75t_L g1003 ( 
.A(n_644),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_683),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_649),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_649),
.Y(n_1006)
);

AND2x6_ASAP7_75t_L g1007 ( 
.A(n_713),
.B(n_446),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_644),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_746),
.B(n_462),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_649),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_746),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_638),
.B(n_456),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_894),
.Y(n_1013)
);

INVx2_ASAP7_75t_SL g1014 ( 
.A(n_816),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_911),
.B(n_459),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_897),
.B(n_464),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_975),
.B(n_806),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_874),
.A2(n_493),
.B(n_500),
.C(n_484),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_909),
.B(n_465),
.Y(n_1019)
);

INVxp67_ASAP7_75t_L g1020 ( 
.A(n_1011),
.Y(n_1020)
);

AND2x6_ASAP7_75t_SL g1021 ( 
.A(n_964),
.B(n_518),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_894),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_985),
.B(n_468),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_920),
.B(n_931),
.Y(n_1024)
);

NAND2x1_ASAP7_75t_L g1025 ( 
.A(n_866),
.B(n_537),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_998),
.B(n_470),
.Y(n_1026)
);

NOR2xp33_ASAP7_75t_L g1027 ( 
.A(n_790),
.B(n_475),
.Y(n_1027)
);

NAND3xp33_ASAP7_75t_SL g1028 ( 
.A(n_812),
.B(n_479),
.C(n_477),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_894),
.Y(n_1029)
);

OR2x6_ASAP7_75t_L g1030 ( 
.A(n_921),
.B(n_522),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_902),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_810),
.Y(n_1032)
);

AOI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_934),
.A2(n_524),
.B1(n_532),
.B2(n_523),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_842),
.A2(n_490),
.B1(n_492),
.B2(n_485),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_960),
.A2(n_538),
.B(n_539),
.C(n_535),
.Y(n_1035)
);

INVx2_ASAP7_75t_SL g1036 ( 
.A(n_835),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_866),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_963),
.Y(n_1038)
);

AND2x6_ASAP7_75t_SL g1039 ( 
.A(n_964),
.B(n_541),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_888),
.B(n_932),
.Y(n_1040)
);

INVx8_ASAP7_75t_L g1041 ( 
.A(n_835),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_794),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_860),
.B(n_494),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_966),
.B(n_495),
.Y(n_1044)
);

INVx3_ASAP7_75t_L g1045 ( 
.A(n_903),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_966),
.B(n_497),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_942),
.B(n_503),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_833),
.A2(n_546),
.B(n_551),
.C(n_543),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_860),
.B(n_504),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_L g1050 ( 
.A1(n_937),
.A2(n_412),
.B1(n_436),
.B2(n_407),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_902),
.Y(n_1051)
);

AOI22xp33_ASAP7_75t_L g1052 ( 
.A1(n_937),
.A2(n_1012),
.B1(n_978),
.B2(n_941),
.Y(n_1052)
);

OAI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_791),
.A2(n_514),
.B1(n_515),
.B2(n_512),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_798),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_795),
.Y(n_1055)
);

AND2x2_ASAP7_75t_L g1056 ( 
.A(n_836),
.B(n_7),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_968),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_787),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_937),
.A2(n_436),
.B1(n_449),
.B2(n_412),
.Y(n_1059)
);

AOI22xp33_ASAP7_75t_L g1060 ( 
.A1(n_937),
.A2(n_457),
.B1(n_449),
.B2(n_516),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_800),
.A2(n_517),
.B1(n_527),
.B2(n_519),
.Y(n_1061)
);

AND2x6_ASAP7_75t_L g1062 ( 
.A(n_982),
.B(n_457),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_903),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_789),
.B(n_8),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_859),
.B(n_529),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_801),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_813),
.Y(n_1067)
);

NAND2xp33_ASAP7_75t_L g1068 ( 
.A(n_797),
.B(n_530),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_859),
.B(n_531),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_977),
.A2(n_545),
.B1(n_548),
.B2(n_544),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_967),
.B(n_549),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_974),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_859),
.B(n_550),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_859),
.B(n_8),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_889),
.B(n_334),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_822),
.B(n_978),
.Y(n_1076)
);

OR2x4_ASAP7_75t_L g1077 ( 
.A(n_834),
.B(n_334),
.Y(n_1077)
);

INVx2_ASAP7_75t_SL g1078 ( 
.A(n_789),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1012),
.B(n_9),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_941),
.A2(n_406),
.B1(n_448),
.B2(n_334),
.Y(n_1080)
);

NOR2x1_ASAP7_75t_R g1081 ( 
.A(n_879),
.B(n_334),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_803),
.B(n_804),
.Y(n_1082)
);

NOR2xp67_ASAP7_75t_SL g1083 ( 
.A(n_929),
.B(n_406),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_982),
.A2(n_448),
.B(n_406),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_983),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_799),
.A2(n_448),
.B1(n_466),
.B2(n_406),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_837),
.B(n_11),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_843),
.A2(n_466),
.B1(n_501),
.B2(n_448),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_921),
.B(n_466),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_802),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_839),
.B(n_11),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_869),
.B(n_12),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_802),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_902),
.Y(n_1094)
);

NOR2xp67_ASAP7_75t_L g1095 ( 
.A(n_876),
.B(n_107),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_986),
.Y(n_1096)
);

OAI221xp5_ASAP7_75t_L g1097 ( 
.A1(n_915),
.A2(n_501),
.B1(n_466),
.B2(n_16),
.C(n_18),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_994),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_SL g1099 ( 
.A1(n_916),
.A2(n_501),
.B1(n_16),
.B2(n_14),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_877),
.B(n_15),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_881),
.B(n_18),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_887),
.B(n_19),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_999),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_892),
.B(n_19),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_901),
.B(n_20),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1007),
.A2(n_820),
.B1(n_981),
.B2(n_821),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1007),
.A2(n_501),
.B1(n_22),
.B2(n_20),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_861),
.B(n_21),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_904),
.B(n_21),
.Y(n_1109)
);

NAND2xp33_ASAP7_75t_L g1110 ( 
.A(n_797),
.B(n_109),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_846),
.B(n_926),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1000),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_886),
.Y(n_1113)
);

INVx1_ASAP7_75t_SL g1114 ( 
.A(n_910),
.Y(n_1114)
);

HB1xp67_ASAP7_75t_L g1115 ( 
.A(n_918),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_905),
.B(n_22),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_925),
.B(n_23),
.Y(n_1117)
);

NOR3x1_ASAP7_75t_L g1118 ( 
.A(n_953),
.B(n_24),
.C(n_25),
.Y(n_1118)
);

NAND2x1p5_ASAP7_75t_L g1119 ( 
.A(n_875),
.B(n_24),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_926),
.B(n_25),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_949),
.B(n_26),
.Y(n_1121)
);

AOI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_861),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_949),
.B(n_29),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_846),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_895),
.Y(n_1125)
);

AO22x1_ASAP7_75t_L g1126 ( 
.A1(n_943),
.A2(n_33),
.B1(n_30),
.B2(n_32),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_984),
.B(n_32),
.Y(n_1127)
);

BUFx6f_ASAP7_75t_L g1128 ( 
.A(n_788),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_851),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_987),
.B(n_995),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_988),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_872),
.B(n_33),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_851),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_996),
.B(n_35),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1009),
.B(n_36),
.Y(n_1135)
);

AOI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1007),
.A2(n_40),
.B1(n_36),
.B2(n_39),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_917),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_878),
.B(n_39),
.Y(n_1138)
);

BUFx3_ASAP7_75t_L g1139 ( 
.A(n_854),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_788),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_1007),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_788),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_817),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_958),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_SL g1145 ( 
.A(n_845),
.B(n_43),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_989),
.B(n_1001),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_893),
.B(n_44),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_820),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_893),
.B(n_45),
.Y(n_1149)
);

INVx2_ASAP7_75t_SL g1150 ( 
.A(n_958),
.Y(n_1150)
);

INVxp67_ASAP7_75t_L g1151 ( 
.A(n_826),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_840),
.B(n_47),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_940),
.B(n_50),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_876),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_1008),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_831),
.Y(n_1156)
);

OR2x6_ASAP7_75t_L g1157 ( 
.A(n_880),
.B(n_961),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_845),
.B(n_50),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_872),
.B(n_51),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_907),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_832),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_821),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_797),
.B(n_52),
.Y(n_1163)
);

INVx3_ASAP7_75t_L g1164 ( 
.A(n_946),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_956),
.A2(n_115),
.B(n_112),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_976),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_981),
.A2(n_58),
.B1(n_55),
.B2(n_56),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_793),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_884),
.B(n_56),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_797),
.B(n_59),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_841),
.B(n_60),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_L g1172 ( 
.A(n_871),
.B(n_116),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_792),
.B(n_796),
.Y(n_1173)
);

INVxp67_ASAP7_75t_L g1174 ( 
.A(n_924),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1004),
.A2(n_63),
.B1(n_61),
.B2(n_62),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1004),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_841),
.B(n_62),
.Y(n_1177)
);

NOR2x1p5_ASAP7_75t_L g1178 ( 
.A(n_962),
.B(n_63),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_841),
.A2(n_68),
.B1(n_64),
.B2(n_66),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_805),
.B(n_64),
.Y(n_1180)
);

AND2x2_ASAP7_75t_L g1181 ( 
.A(n_951),
.B(n_66),
.Y(n_1181)
);

INVx5_ASAP7_75t_L g1182 ( 
.A(n_862),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_946),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_939),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_917),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_917),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_841),
.B(n_68),
.Y(n_1187)
);

AOI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_819),
.A2(n_71),
.B1(n_69),
.B2(n_70),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_933),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_890),
.B(n_69),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_959),
.B(n_70),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_900),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_818),
.B(n_71),
.Y(n_1193)
);

AND2x4_ASAP7_75t_L g1194 ( 
.A(n_805),
.B(n_72),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_853),
.B(n_72),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_867),
.B(n_73),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_870),
.B(n_73),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_944),
.B(n_74),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_865),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1024),
.Y(n_1200)
);

NOR3xp33_ASAP7_75t_SL g1201 ( 
.A(n_1155),
.B(n_808),
.C(n_947),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1040),
.B(n_848),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1128),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1128),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1017),
.A2(n_922),
.B1(n_970),
.B2(n_936),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1184),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1038),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1020),
.A2(n_930),
.B1(n_972),
.B2(n_865),
.Y(n_1208)
);

NOR2xp33_ASAP7_75t_R g1209 ( 
.A(n_1168),
.B(n_1003),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1128),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1078),
.A2(n_950),
.B1(n_815),
.B2(n_891),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1115),
.Y(n_1212)
);

INVx1_ASAP7_75t_SL g1213 ( 
.A(n_1114),
.Y(n_1213)
);

INVx3_ASAP7_75t_SL g1214 ( 
.A(n_1157),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1055),
.B(n_954),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1113),
.Y(n_1216)
);

BUFx2_ASAP7_75t_L g1217 ( 
.A(n_1089),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1144),
.B(n_979),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1015),
.B(n_900),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1125),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_1014),
.Y(n_1221)
);

AND2x6_ASAP7_75t_L g1222 ( 
.A(n_1180),
.B(n_1194),
.Y(n_1222)
);

BUFx3_ASAP7_75t_L g1223 ( 
.A(n_1057),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1042),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1054),
.Y(n_1225)
);

CKINVDCx16_ASAP7_75t_R g1226 ( 
.A(n_1030),
.Y(n_1226)
);

OR2x6_ASAP7_75t_L g1227 ( 
.A(n_1041),
.B(n_815),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_SL g1228 ( 
.A(n_1081),
.B(n_1003),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1015),
.B(n_928),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1087),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1066),
.Y(n_1231)
);

INVx5_ASAP7_75t_L g1232 ( 
.A(n_1041),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1052),
.B(n_928),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_1053),
.B(n_952),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1091),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1092),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1157),
.Y(n_1237)
);

BUFx6f_ASAP7_75t_L g1238 ( 
.A(n_1140),
.Y(n_1238)
);

BUFx12f_ASAP7_75t_L g1239 ( 
.A(n_1057),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1100),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1151),
.A2(n_997),
.B1(n_973),
.B2(n_969),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1058),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1146),
.A2(n_829),
.B(n_948),
.Y(n_1243)
);

INVx3_ASAP7_75t_L g1244 ( 
.A(n_1045),
.Y(n_1244)
);

OR2x2_ASAP7_75t_L g1245 ( 
.A(n_1174),
.B(n_971),
.Y(n_1245)
);

BUFx4f_ASAP7_75t_L g1246 ( 
.A(n_1030),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1067),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1150),
.B(n_863),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1072),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1056),
.B(n_850),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1101),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1102),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1085),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1104),
.Y(n_1254)
);

BUFx4f_ASAP7_75t_L g1255 ( 
.A(n_1041),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_1021),
.Y(n_1256)
);

INVx3_ASAP7_75t_L g1257 ( 
.A(n_1045),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1096),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1098),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1103),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_1039),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_1036),
.B(n_908),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1131),
.B(n_863),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1112),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1090),
.B(n_971),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1082),
.B(n_882),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1156),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1076),
.B(n_945),
.Y(n_1268)
);

NOR2xp33_ASAP7_75t_L g1269 ( 
.A(n_1124),
.B(n_965),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1161),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1199),
.B(n_871),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1032),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_L g1273 ( 
.A(n_1140),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1181),
.B(n_1191),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_1089),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1093),
.A2(n_1064),
.B1(n_1132),
.B2(n_1108),
.Y(n_1276)
);

NOR3xp33_ASAP7_75t_SL g1277 ( 
.A(n_1028),
.B(n_993),
.C(n_809),
.Y(n_1277)
);

INVx3_ASAP7_75t_L g1278 ( 
.A(n_1063),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1063),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1018),
.B(n_868),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1180),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1192),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1033),
.B(n_1134),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1129),
.Y(n_1284)
);

AND3x1_ASAP7_75t_SL g1285 ( 
.A(n_1178),
.B(n_965),
.C(n_913),
.Y(n_1285)
);

NAND2x1p5_ASAP7_75t_L g1286 ( 
.A(n_1139),
.B(n_871),
.Y(n_1286)
);

NOR3xp33_ASAP7_75t_SL g1287 ( 
.A(n_1034),
.B(n_898),
.C(n_896),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1160),
.B(n_899),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1120),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1121),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1123),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1133),
.Y(n_1292)
);

INVx5_ASAP7_75t_L g1293 ( 
.A(n_1182),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1077),
.Y(n_1294)
);

NOR2xp33_ASAP7_75t_L g1295 ( 
.A(n_1111),
.B(n_852),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1183),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_1164),
.Y(n_1297)
);

NOR2xp33_ASAP7_75t_R g1298 ( 
.A(n_1068),
.B(n_862),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_SL g1299 ( 
.A(n_1119),
.B(n_1136),
.C(n_1122),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1079),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1152),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1081),
.Y(n_1302)
);

XNOR2xp5_ASAP7_75t_L g1303 ( 
.A(n_1070),
.B(n_885),
.Y(n_1303)
);

OR2x6_ASAP7_75t_L g1304 ( 
.A(n_1194),
.B(n_927),
.Y(n_1304)
);

CKINVDCx14_ASAP7_75t_R g1305 ( 
.A(n_1136),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1164),
.Y(n_1306)
);

NAND2x1p5_ASAP7_75t_L g1307 ( 
.A(n_1182),
.B(n_838),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1037),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1135),
.B(n_868),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1130),
.A2(n_914),
.B(n_912),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1198),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1037),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_SL g1313 ( 
.A(n_1182),
.B(n_862),
.Y(n_1313)
);

CKINVDCx8_ASAP7_75t_R g1314 ( 
.A(n_1062),
.Y(n_1314)
);

AND2x4_ASAP7_75t_L g1315 ( 
.A(n_1176),
.B(n_873),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1190),
.B(n_1147),
.Y(n_1316)
);

INVx5_ASAP7_75t_L g1317 ( 
.A(n_1140),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1149),
.B(n_1158),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1159),
.B(n_868),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1016),
.B(n_868),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1143),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1169),
.B(n_891),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1105),
.A2(n_906),
.B(n_883),
.C(n_811),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1035),
.B(n_891),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1062),
.Y(n_1325)
);

BUFx12f_ASAP7_75t_L g1326 ( 
.A(n_1062),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1023),
.B(n_838),
.Y(n_1327)
);

NOR3xp33_ASAP7_75t_SL g1328 ( 
.A(n_1145),
.B(n_957),
.C(n_955),
.Y(n_1328)
);

NOR3xp33_ASAP7_75t_SL g1329 ( 
.A(n_1043),
.B(n_862),
.C(n_891),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1048),
.B(n_919),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1109),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1026),
.B(n_1106),
.Y(n_1332)
);

NAND3xp33_ASAP7_75t_SL g1333 ( 
.A(n_1188),
.B(n_935),
.C(n_923),
.Y(n_1333)
);

AO22x1_ASAP7_75t_L g1334 ( 
.A1(n_1118),
.A2(n_838),
.B1(n_991),
.B2(n_976),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_SL g1335 ( 
.A(n_1126),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1116),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1117),
.Y(n_1337)
);

NAND2xp33_ASAP7_75t_L g1338 ( 
.A(n_1142),
.B(n_1166),
.Y(n_1338)
);

NOR2xp33_ASAP7_75t_L g1339 ( 
.A(n_1049),
.B(n_938),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1266),
.A2(n_1250),
.B(n_1283),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1316),
.A2(n_1059),
.B(n_1050),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1334),
.A2(n_1095),
.B(n_1075),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1213),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1239),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1200),
.B(n_1044),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_1232),
.B(n_1154),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1280),
.A2(n_1110),
.B(n_1165),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1243),
.A2(n_1138),
.B(n_1127),
.C(n_1153),
.Y(n_1348)
);

AOI21xp5_ASAP7_75t_L g1349 ( 
.A1(n_1320),
.A2(n_1166),
.B(n_1142),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1275),
.A2(n_1074),
.B(n_1163),
.Y(n_1350)
);

NAND2x1_ASAP7_75t_L g1351 ( 
.A(n_1222),
.B(n_1142),
.Y(n_1351)
);

INVx4_ASAP7_75t_L g1352 ( 
.A(n_1232),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1202),
.B(n_1046),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1305),
.B(n_1212),
.Y(n_1354)
);

AND2x2_ASAP7_75t_L g1355 ( 
.A(n_1226),
.B(n_1027),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1310),
.A2(n_1084),
.B(n_1095),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1203),
.Y(n_1357)
);

BUFx3_ASAP7_75t_L g1358 ( 
.A(n_1223),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1309),
.A2(n_1022),
.B(n_1013),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1307),
.A2(n_1031),
.B(n_1029),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1207),
.B(n_1071),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1302),
.B(n_1025),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1203),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1216),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1299),
.A2(n_1099),
.B1(n_1060),
.B2(n_1062),
.Y(n_1365)
);

OAI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1268),
.A2(n_1019),
.B(n_1047),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_L g1367 ( 
.A(n_1311),
.B(n_1061),
.Y(n_1367)
);

NAND2xp5_ASAP7_75t_L g1368 ( 
.A(n_1259),
.B(n_1193),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1246),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1245),
.B(n_1241),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1323),
.A2(n_1196),
.B(n_1195),
.Y(n_1371)
);

INVxp67_ASAP7_75t_SL g1372 ( 
.A(n_1281),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1330),
.A2(n_1094),
.B(n_1051),
.Y(n_1373)
);

NOR4xp25_ASAP7_75t_L g1374 ( 
.A(n_1211),
.B(n_1097),
.C(n_1162),
.D(n_1148),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1214),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1318),
.A2(n_1197),
.B(n_1088),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1289),
.A2(n_1185),
.B(n_1137),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1260),
.B(n_1173),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1314),
.A2(n_1274),
.B1(n_1229),
.B2(n_1219),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1290),
.A2(n_1189),
.B(n_1186),
.Y(n_1380)
);

AOI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1322),
.A2(n_1166),
.B(n_1170),
.Y(n_1381)
);

AOI22x1_ASAP7_75t_SL g1382 ( 
.A1(n_1256),
.A2(n_1118),
.B1(n_1141),
.B2(n_1179),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1264),
.B(n_1086),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1325),
.A2(n_1107),
.B1(n_1175),
.B2(n_1167),
.Y(n_1384)
);

BUFx2_ASAP7_75t_L g1385 ( 
.A(n_1222),
.Y(n_1385)
);

BUFx12f_ASAP7_75t_L g1386 ( 
.A(n_1206),
.Y(n_1386)
);

AOI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1334),
.A2(n_1083),
.B(n_1172),
.Y(n_1387)
);

AO21x2_ASAP7_75t_L g1388 ( 
.A1(n_1333),
.A2(n_1177),
.B(n_1171),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1331),
.A2(n_1187),
.B(n_1069),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1321),
.A2(n_1080),
.B(n_1172),
.C(n_1154),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1272),
.B(n_1073),
.Y(n_1391)
);

INVxp67_ASAP7_75t_L g1392 ( 
.A(n_1228),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1291),
.A2(n_824),
.A3(n_825),
.B(n_814),
.Y(n_1393)
);

BUFx6f_ASAP7_75t_L g1394 ( 
.A(n_1203),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1244),
.A2(n_1002),
.B(n_980),
.Y(n_1395)
);

AOI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1336),
.A2(n_1065),
.B(n_858),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1222),
.B(n_933),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1222),
.B(n_933),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1244),
.A2(n_1006),
.B(n_823),
.Y(n_1399)
);

NAND3xp33_ASAP7_75t_L g1400 ( 
.A(n_1328),
.B(n_991),
.C(n_976),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1257),
.A2(n_823),
.B(n_807),
.Y(n_1401)
);

AO31x2_ASAP7_75t_L g1402 ( 
.A1(n_1337),
.A2(n_864),
.A3(n_844),
.B(n_991),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1232),
.B(n_807),
.Y(n_1403)
);

AOI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1301),
.A2(n_849),
.B(n_847),
.Y(n_1404)
);

BUFx6f_ASAP7_75t_L g1405 ( 
.A(n_1204),
.Y(n_1405)
);

AND3x1_ASAP7_75t_L g1406 ( 
.A(n_1201),
.B(n_74),
.C(n_76),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1230),
.A2(n_828),
.B(n_830),
.C(n_827),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1233),
.B(n_1010),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1235),
.A2(n_849),
.B(n_847),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1234),
.A2(n_828),
.B(n_830),
.C(n_827),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1267),
.B(n_1270),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1224),
.B(n_990),
.Y(n_1412)
);

BUFx12f_ASAP7_75t_L g1413 ( 
.A(n_1261),
.Y(n_1413)
);

OAI22x1_ASAP7_75t_L g1414 ( 
.A1(n_1205),
.A2(n_79),
.B1(n_77),
.B2(n_78),
.Y(n_1414)
);

AO31x2_ASAP7_75t_L g1415 ( 
.A1(n_1236),
.A2(n_992),
.A3(n_849),
.B(n_855),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1326),
.A2(n_992),
.B1(n_855),
.B2(n_856),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1255),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1255),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1220),
.B(n_79),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1225),
.B(n_990),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1231),
.B(n_1010),
.Y(n_1421)
);

NAND2x1_ASAP7_75t_L g1422 ( 
.A(n_1204),
.B(n_992),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1257),
.A2(n_1005),
.B(n_855),
.Y(n_1423)
);

BUFx10_ASAP7_75t_L g1424 ( 
.A(n_1271),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1227),
.B(n_81),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1240),
.A2(n_856),
.B(n_847),
.Y(n_1426)
);

AO32x2_ASAP7_75t_L g1427 ( 
.A1(n_1335),
.A2(n_81),
.A3(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_1427)
);

NAND2xp5_ASAP7_75t_L g1428 ( 
.A(n_1247),
.B(n_1005),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1227),
.B(n_1221),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1294),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1364),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1411),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1340),
.A2(n_1353),
.B1(n_1370),
.B2(n_1276),
.C(n_1366),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1343),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1354),
.B(n_1248),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1345),
.B(n_1367),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_SL g1437 ( 
.A1(n_1350),
.A2(n_1387),
.B(n_1379),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_SL g1438 ( 
.A1(n_1352),
.A2(n_1324),
.B(n_1319),
.Y(n_1438)
);

AOI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1342),
.A2(n_1252),
.B(n_1251),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1344),
.Y(n_1440)
);

NAND2xp5_ASAP7_75t_L g1441 ( 
.A(n_1361),
.B(n_1249),
.Y(n_1441)
);

BUFx8_ASAP7_75t_L g1442 ( 
.A(n_1417),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1373),
.A2(n_1278),
.B(n_1254),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1348),
.A2(n_1338),
.B(n_1210),
.Y(n_1444)
);

AOI332xp33_ASAP7_75t_L g1445 ( 
.A1(n_1425),
.A2(n_1282),
.A3(n_1215),
.B1(n_1218),
.B2(n_1253),
.B3(n_1258),
.C1(n_1300),
.C2(n_1208),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1356),
.A2(n_1278),
.B(n_1297),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1377),
.Y(n_1447)
);

OR3x4_ASAP7_75t_SL g1448 ( 
.A(n_1372),
.B(n_1285),
.C(n_1209),
.Y(n_1448)
);

AO31x2_ASAP7_75t_L g1449 ( 
.A1(n_1347),
.A2(n_1390),
.A3(n_1389),
.B(n_1381),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1419),
.B(n_1248),
.Y(n_1450)
);

NOR2x1_ASAP7_75t_R g1451 ( 
.A(n_1386),
.B(n_1242),
.Y(n_1451)
);

INVx2_ASAP7_75t_SL g1452 ( 
.A(n_1424),
.Y(n_1452)
);

INVx8_ASAP7_75t_L g1453 ( 
.A(n_1346),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1359),
.A2(n_1306),
.B(n_1308),
.Y(n_1454)
);

OAI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1385),
.A2(n_1217),
.B1(n_1304),
.B2(n_1237),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1380),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1349),
.A2(n_1312),
.B(n_1279),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1404),
.A2(n_1292),
.B(n_1284),
.Y(n_1458)
);

OA21x2_ASAP7_75t_L g1459 ( 
.A1(n_1376),
.A2(n_1329),
.B(n_1296),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1355),
.B(n_1303),
.Y(n_1460)
);

AOI21xp33_ASAP7_75t_L g1461 ( 
.A1(n_1365),
.A2(n_1332),
.B(n_1304),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1357),
.B(n_1317),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1378),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1409),
.A2(n_1263),
.B(n_1286),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1415),
.Y(n_1465)
);

OAI21x1_ASAP7_75t_L g1466 ( 
.A1(n_1426),
.A2(n_1295),
.B(n_1210),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1271),
.Y(n_1467)
);

NAND2x1p5_ASAP7_75t_L g1468 ( 
.A(n_1352),
.B(n_1293),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1351),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1382),
.B(n_1265),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1341),
.A2(n_1384),
.B(n_1368),
.C(n_1383),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1358),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1415),
.Y(n_1473)
);

NOR2xp33_ASAP7_75t_L g1474 ( 
.A(n_1382),
.B(n_1332),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1470),
.B(n_1369),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1474),
.A2(n_1406),
.B1(n_1392),
.B2(n_1430),
.Y(n_1476)
);

OAI221xp5_ASAP7_75t_L g1477 ( 
.A1(n_1433),
.A2(n_1339),
.B1(n_1374),
.B2(n_1269),
.C(n_1277),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1465),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1465),
.Y(n_1479)
);

OR2x6_ASAP7_75t_L g1480 ( 
.A(n_1437),
.B(n_1414),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1432),
.B(n_1463),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1474),
.A2(n_1429),
.B1(n_1288),
.B2(n_1391),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1440),
.Y(n_1483)
);

INVx2_ASAP7_75t_SL g1484 ( 
.A(n_1453),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1470),
.B(n_1375),
.Y(n_1485)
);

BUFx3_ASAP7_75t_L g1486 ( 
.A(n_1453),
.Y(n_1486)
);

OR2x6_ASAP7_75t_L g1487 ( 
.A(n_1453),
.B(n_1362),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1473),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1436),
.B(n_1215),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1473),
.A2(n_1388),
.B(n_1396),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1447),
.Y(n_1491)
);

BUFx3_ASAP7_75t_L g1492 ( 
.A(n_1453),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1431),
.B(n_1418),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1462),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1440),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1461),
.A2(n_1288),
.B1(n_1362),
.B2(n_1327),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1460),
.A2(n_1327),
.B1(n_1371),
.B2(n_1346),
.Y(n_1497)
);

INVx3_ASAP7_75t_L g1498 ( 
.A(n_1469),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1441),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1471),
.B(n_1218),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1447),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1468),
.A2(n_1313),
.B1(n_1398),
.B2(n_1397),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_SL g1503 ( 
.A1(n_1442),
.A2(n_1298),
.B1(n_1293),
.B2(n_1371),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_SL g1504 ( 
.A1(n_1442),
.A2(n_1293),
.B1(n_1427),
.B2(n_1363),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1487),
.A2(n_1486),
.B1(n_1492),
.B2(n_1484),
.Y(n_1505)
);

AO21x2_ASAP7_75t_L g1506 ( 
.A1(n_1500),
.A2(n_1439),
.B(n_1490),
.Y(n_1506)
);

AOI221xp5_ASAP7_75t_L g1507 ( 
.A1(n_1477),
.A2(n_1455),
.B1(n_1434),
.B2(n_1471),
.C(n_1262),
.Y(n_1507)
);

OAI221xp5_ASAP7_75t_L g1508 ( 
.A1(n_1476),
.A2(n_1452),
.B1(n_1287),
.B2(n_1472),
.C(n_1445),
.Y(n_1508)
);

OR2x2_ASAP7_75t_L g1509 ( 
.A(n_1499),
.B(n_1449),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1481),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1494),
.Y(n_1511)
);

AOI222xp33_ASAP7_75t_L g1512 ( 
.A1(n_1489),
.A2(n_1442),
.B1(n_1451),
.B2(n_1450),
.C1(n_1435),
.C2(n_1467),
.Y(n_1512)
);

AOI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1482),
.A2(n_1315),
.B1(n_1438),
.B2(n_1408),
.C(n_1469),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1493),
.B(n_1469),
.Y(n_1514)
);

AOI21xp5_ASAP7_75t_L g1515 ( 
.A1(n_1502),
.A2(n_1444),
.B(n_1459),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1504),
.A2(n_1459),
.B1(n_1400),
.B2(n_1468),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1485),
.A2(n_1459),
.B1(n_1464),
.B2(n_1462),
.Y(n_1517)
);

INVx1_ASAP7_75t_SL g1518 ( 
.A(n_1486),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1475),
.A2(n_1464),
.B1(n_1462),
.B2(n_1458),
.Y(n_1519)
);

BUFx4f_ASAP7_75t_SL g1520 ( 
.A(n_1492),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_SL g1521 ( 
.A1(n_1484),
.A2(n_1448),
.B1(n_1427),
.B2(n_1357),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1497),
.A2(n_1458),
.B1(n_1456),
.B2(n_1466),
.Y(n_1522)
);

AOI21xp33_ASAP7_75t_SL g1523 ( 
.A1(n_1483),
.A2(n_1448),
.B(n_83),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1478),
.Y(n_1524)
);

AO21x1_ASAP7_75t_L g1525 ( 
.A1(n_1479),
.A2(n_1427),
.B(n_1443),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1494),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1490),
.A2(n_1456),
.B(n_1443),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1496),
.A2(n_1466),
.B1(n_1457),
.B2(n_1315),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1483),
.Y(n_1529)
);

OAI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1480),
.A2(n_1407),
.B1(n_1428),
.B2(n_1421),
.C(n_1420),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1524),
.Y(n_1531)
);

HB1xp67_ASAP7_75t_L g1532 ( 
.A(n_1511),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1509),
.B(n_1478),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1524),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1509),
.B(n_1488),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1510),
.B(n_1498),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1525),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1525),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1526),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1506),
.B(n_1488),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1506),
.B(n_1501),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1526),
.B(n_1501),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_L g1543 ( 
.A1(n_1521),
.A2(n_1508),
.B1(n_1507),
.B2(n_1513),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1512),
.A2(n_1480),
.B1(n_1487),
.B2(n_1503),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1527),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1514),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1518),
.Y(n_1547)
);

NAND4xp25_ASAP7_75t_L g1548 ( 
.A(n_1523),
.B(n_1498),
.C(n_1410),
.D(n_1412),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1505),
.B(n_1498),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_1506),
.B(n_1490),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1527),
.Y(n_1551)
);

AOI322xp5_ASAP7_75t_L g1552 ( 
.A1(n_1543),
.A2(n_1517),
.A3(n_1516),
.B1(n_1529),
.B2(n_1519),
.C1(n_1495),
.C2(n_1522),
.Y(n_1552)
);

BUFx2_ASAP7_75t_L g1553 ( 
.A(n_1547),
.Y(n_1553)
);

AOI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1537),
.A2(n_1529),
.B1(n_1530),
.B2(n_1515),
.C(n_1495),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1547),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1546),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1532),
.B(n_1480),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1544),
.A2(n_1546),
.B1(n_1520),
.B2(n_1549),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1536),
.Y(n_1559)
);

OAI211xp5_ASAP7_75t_L g1560 ( 
.A1(n_1537),
.A2(n_1528),
.B(n_1487),
.C(n_1317),
.Y(n_1560)
);

NOR2xp67_ASAP7_75t_L g1561 ( 
.A(n_1539),
.B(n_84),
.Y(n_1561)
);

NOR2x1_ASAP7_75t_L g1562 ( 
.A(n_1548),
.B(n_1487),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1533),
.B(n_1480),
.Y(n_1563)
);

OAI33xp33_ASAP7_75t_L g1564 ( 
.A1(n_1538),
.A2(n_1416),
.A3(n_87),
.B1(n_88),
.B2(n_90),
.B3(n_91),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1556),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1553),
.B(n_1555),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1557),
.B(n_1559),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1563),
.Y(n_1568)
);

BUFx2_ASAP7_75t_L g1569 ( 
.A(n_1563),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1558),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1562),
.B(n_1413),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1561),
.Y(n_1572)
);

BUFx2_ASAP7_75t_L g1573 ( 
.A(n_1554),
.Y(n_1573)
);

INVx3_ASAP7_75t_L g1574 ( 
.A(n_1560),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1552),
.B(n_1541),
.Y(n_1575)
);

NOR2x1_ASAP7_75t_L g1576 ( 
.A(n_1560),
.B(n_1538),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1554),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1564),
.B(n_1541),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1556),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1565),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1565),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1570),
.B(n_1542),
.Y(n_1582)
);

NAND2xp67_ASAP7_75t_L g1583 ( 
.A(n_1575),
.B(n_1540),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1575),
.B(n_1533),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1579),
.Y(n_1585)
);

NOR3xp33_ASAP7_75t_L g1586 ( 
.A(n_1584),
.B(n_1573),
.C(n_1577),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1582),
.B(n_1569),
.Y(n_1587)
);

BUFx2_ASAP7_75t_L g1588 ( 
.A(n_1580),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1587),
.Y(n_1589)
);

NOR2x1_ASAP7_75t_SL g1590 ( 
.A(n_1588),
.B(n_1578),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1589),
.B(n_1586),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1590),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1589),
.Y(n_1594)
);

OAI22xp5_ASAP7_75t_L g1595 ( 
.A1(n_1591),
.A2(n_1577),
.B1(n_1574),
.B2(n_1582),
.Y(n_1595)
);

XNOR2x2_ASAP7_75t_L g1596 ( 
.A(n_1594),
.B(n_1571),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1593),
.B(n_1574),
.Y(n_1597)
);

BUFx4f_ASAP7_75t_SL g1598 ( 
.A(n_1592),
.Y(n_1598)
);

AOI31xp33_ASAP7_75t_SL g1599 ( 
.A1(n_1591),
.A2(n_1568),
.A3(n_1583),
.B(n_1574),
.Y(n_1599)
);

NOR4xp25_ASAP7_75t_SL g1600 ( 
.A(n_1594),
.B(n_1572),
.C(n_1569),
.D(n_1581),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1594),
.Y(n_1601)
);

OAI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1597),
.A2(n_1600),
.B(n_1601),
.C(n_1595),
.Y(n_1602)
);

AOI221xp5_ASAP7_75t_L g1603 ( 
.A1(n_1596),
.A2(n_1578),
.B1(n_1566),
.B2(n_1585),
.C(n_1579),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1598),
.B(n_1566),
.Y(n_1604)
);

AOI211x1_ASAP7_75t_L g1605 ( 
.A1(n_1599),
.A2(n_1567),
.B(n_1576),
.C(n_1540),
.Y(n_1605)
);

XOR2xp5_ASAP7_75t_L g1606 ( 
.A(n_1596),
.B(n_86),
.Y(n_1606)
);

AOI311xp33_ASAP7_75t_L g1607 ( 
.A1(n_1597),
.A2(n_1534),
.A3(n_90),
.B(n_92),
.C(n_93),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1597),
.B(n_1567),
.Y(n_1608)
);

XNOR2x2_ASAP7_75t_L g1609 ( 
.A(n_1596),
.B(n_1568),
.Y(n_1609)
);

NOR4xp25_ASAP7_75t_L g1610 ( 
.A(n_1601),
.B(n_1551),
.C(n_1545),
.D(n_95),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1598),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1595),
.A2(n_1551),
.B(n_1545),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1610),
.A2(n_1550),
.B1(n_1534),
.B2(n_1403),
.C(n_1531),
.Y(n_1613)
);

AOI211xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1611),
.A2(n_1403),
.B(n_97),
.C(n_87),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1608),
.B(n_1542),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1604),
.Y(n_1616)
);

OAI21xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1606),
.A2(n_1535),
.B(n_1531),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1602),
.A2(n_1550),
.B(n_1457),
.Y(n_1618)
);

AOI21xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1609),
.A2(n_94),
.B(n_98),
.Y(n_1619)
);

O2A1O1Ixp5_ASAP7_75t_L g1620 ( 
.A1(n_1612),
.A2(n_1550),
.B(n_1422),
.C(n_100),
.Y(n_1620)
);

NOR2x1_ASAP7_75t_SL g1621 ( 
.A(n_1607),
.B(n_1317),
.Y(n_1621)
);

NAND2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1605),
.B(n_1550),
.Y(n_1622)
);

AOI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1603),
.A2(n_100),
.B(n_98),
.C(n_99),
.Y(n_1623)
);

NOR2xp67_ASAP7_75t_L g1624 ( 
.A(n_1611),
.B(n_101),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_SL g1625 ( 
.A1(n_1611),
.A2(n_1535),
.B1(n_103),
.B2(n_104),
.C(n_105),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1606),
.A2(n_1446),
.B(n_102),
.Y(n_1626)
);

OA21x2_ASAP7_75t_L g1627 ( 
.A1(n_1611),
.A2(n_1360),
.B(n_1401),
.Y(n_1627)
);

CKINVDCx16_ASAP7_75t_R g1628 ( 
.A(n_1616),
.Y(n_1628)
);

OAI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1617),
.A2(n_102),
.B(n_103),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1624),
.Y(n_1630)
);

INVx1_ASAP7_75t_SL g1631 ( 
.A(n_1626),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1621),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1620),
.Y(n_1633)
);

NAND4xp25_ASAP7_75t_SL g1634 ( 
.A(n_1625),
.B(n_104),
.C(n_105),
.D(n_1491),
.Y(n_1634)
);

AOI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1619),
.A2(n_1446),
.B(n_1363),
.Y(n_1635)
);

CKINVDCx20_ASAP7_75t_R g1636 ( 
.A(n_1614),
.Y(n_1636)
);

AOI22xp33_ASAP7_75t_L g1637 ( 
.A1(n_1622),
.A2(n_1527),
.B1(n_1394),
.B2(n_1357),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1615),
.Y(n_1638)
);

OAI211xp5_ASAP7_75t_SL g1639 ( 
.A1(n_1623),
.A2(n_121),
.B(n_122),
.C(n_123),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1613),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_R g1641 ( 
.A(n_1618),
.B(n_124),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1627),
.A2(n_1394),
.B(n_1363),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1632),
.B(n_1627),
.Y(n_1643)
);

NAND4xp25_ASAP7_75t_L g1644 ( 
.A(n_1633),
.B(n_1631),
.C(n_1629),
.D(n_1640),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1636),
.A2(n_1628),
.B1(n_1630),
.B2(n_1638),
.Y(n_1645)
);

NOR2xp67_ASAP7_75t_L g1646 ( 
.A(n_1634),
.B(n_125),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1641),
.B(n_1449),
.Y(n_1647)
);

AND2x2_ASAP7_75t_SL g1648 ( 
.A(n_1637),
.B(n_1394),
.Y(n_1648)
);

NAND3xp33_ASAP7_75t_L g1649 ( 
.A(n_1639),
.B(n_1405),
.C(n_1210),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1635),
.B(n_1449),
.Y(n_1650)
);

BUFx6f_ASAP7_75t_L g1651 ( 
.A(n_1642),
.Y(n_1651)
);

NOR4xp75_ASAP7_75t_L g1652 ( 
.A(n_1629),
.B(n_128),
.C(n_129),
.D(n_133),
.Y(n_1652)
);

OAI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1632),
.A2(n_1405),
.B(n_1273),
.C(n_1238),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1632),
.B(n_1491),
.Y(n_1654)
);

NOR2x1_ASAP7_75t_L g1655 ( 
.A(n_1632),
.B(n_1405),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1628),
.B(n_1449),
.Y(n_1656)
);

NOR4xp75_ASAP7_75t_SL g1657 ( 
.A(n_1636),
.B(n_134),
.C(n_135),
.D(n_136),
.Y(n_1657)
);

NOR2x1_ASAP7_75t_L g1658 ( 
.A(n_1632),
.B(n_1204),
.Y(n_1658)
);

NOR2x1_ASAP7_75t_L g1659 ( 
.A(n_1632),
.B(n_1238),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1644),
.B(n_1646),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1655),
.A2(n_138),
.B(n_140),
.C(n_143),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_SL g1662 ( 
.A(n_1657),
.B(n_1238),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1645),
.Y(n_1663)
);

OA22x2_ASAP7_75t_L g1664 ( 
.A1(n_1643),
.A2(n_1454),
.B1(n_1399),
.B2(n_1395),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1651),
.B(n_147),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_SL g1666 ( 
.A(n_1656),
.B(n_149),
.C(n_150),
.D(n_152),
.Y(n_1666)
);

OAI321xp33_ASAP7_75t_L g1667 ( 
.A1(n_1651),
.A2(n_1273),
.A3(n_1393),
.B1(n_155),
.B2(n_157),
.C(n_163),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1658),
.B(n_1393),
.Y(n_1668)
);

NOR3xp33_ASAP7_75t_L g1669 ( 
.A(n_1659),
.B(n_1423),
.C(n_153),
.Y(n_1669)
);

NOR3xp33_ASAP7_75t_SL g1670 ( 
.A(n_1653),
.B(n_154),
.C(n_164),
.Y(n_1670)
);

NOR4xp25_ASAP7_75t_L g1671 ( 
.A(n_1647),
.B(n_167),
.C(n_168),
.D(n_170),
.Y(n_1671)
);

OA22x2_ASAP7_75t_L g1672 ( 
.A1(n_1654),
.A2(n_1454),
.B1(n_1393),
.B2(n_175),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1663),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1665),
.Y(n_1674)
);

NOR3xp33_ASAP7_75t_L g1675 ( 
.A(n_1660),
.B(n_1649),
.C(n_1652),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1662),
.B(n_1648),
.Y(n_1676)
);

NOR2x1_ASAP7_75t_L g1677 ( 
.A(n_1666),
.B(n_1650),
.Y(n_1677)
);

XNOR2xp5_ASAP7_75t_L g1678 ( 
.A(n_1670),
.B(n_172),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1671),
.B(n_173),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1661),
.B(n_176),
.Y(n_1680)
);

INVx1_ASAP7_75t_SL g1681 ( 
.A(n_1668),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1673),
.B(n_1667),
.Y(n_1682)
);

OR5x1_ASAP7_75t_L g1683 ( 
.A(n_1675),
.B(n_1672),
.C(n_1664),
.D(n_1669),
.E(n_180),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1676),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1681),
.B(n_177),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1679),
.Y(n_1686)
);

XNOR2x1_ASAP7_75t_L g1687 ( 
.A(n_1678),
.B(n_178),
.Y(n_1687)
);

XNOR2x1_ASAP7_75t_L g1688 ( 
.A(n_1687),
.B(n_1677),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1684),
.A2(n_1674),
.B1(n_1680),
.B2(n_1273),
.Y(n_1689)
);

XNOR2x1_ASAP7_75t_L g1690 ( 
.A(n_1686),
.B(n_179),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1685),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1691),
.Y(n_1692)
);

NAND2xp33_ASAP7_75t_SL g1693 ( 
.A(n_1688),
.B(n_1683),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1690),
.A2(n_1682),
.B1(n_857),
.B2(n_856),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1692),
.Y(n_1695)
);

AO22x2_ASAP7_75t_SL g1696 ( 
.A1(n_1693),
.A2(n_1689),
.B1(n_184),
.B2(n_190),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1695),
.Y(n_1697)
);

OAI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1696),
.A2(n_1694),
.B(n_183),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_SL g1699 ( 
.A1(n_1697),
.A2(n_192),
.B1(n_193),
.B2(n_194),
.Y(n_1699)
);

AOI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1698),
.A2(n_1402),
.B1(n_857),
.B2(n_1415),
.Y(n_1700)
);

OAI221xp5_ASAP7_75t_R g1701 ( 
.A1(n_1700),
.A2(n_1402),
.B1(n_199),
.B2(n_200),
.C(n_201),
.Y(n_1701)
);

AOI211xp5_ASAP7_75t_L g1702 ( 
.A1(n_1701),
.A2(n_1699),
.B(n_203),
.C(n_208),
.Y(n_1702)
);


endmodule