module real_jpeg_33594_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g99 ( 
.A(n_0),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_0),
.Y(n_299)
);

BUFx12f_ASAP7_75t_L g344 ( 
.A(n_0),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_1),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_1),
.B(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_1),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_1),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_1),
.B(n_224),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_2),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_4),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_4),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_4),
.B(n_349),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_5),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_6),
.Y(n_306)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_7),
.Y(n_165)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_7),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_8),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_8),
.B(n_43),
.Y(n_42)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_8),
.B(n_51),
.Y(n_50)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_8),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_8),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_8),
.B(n_108),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_8),
.B(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_8),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_9),
.B(n_45),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_9),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_9),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_9),
.B(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_10),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_10),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_11),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_12),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_12),
.B(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g275 ( 
.A(n_12),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g308 ( 
.A(n_12),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_12),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_13),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_13),
.B(n_127),
.Y(n_126)
);

AND2x6_ASAP7_75t_SL g136 ( 
.A(n_13),
.B(n_137),
.Y(n_136)
);

NAND2x1_ASAP7_75t_L g171 ( 
.A(n_13),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g281 ( 
.A(n_13),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_13),
.B(n_297),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_13),
.B(n_371),
.Y(n_370)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_14),
.Y(n_85)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_14),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_15),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_16),
.B(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_16),
.B(n_93),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_16),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_16),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_16),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_16),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_16),
.B(n_133),
.Y(n_132)
);

NAND2x1_ASAP7_75t_L g223 ( 
.A(n_16),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_17),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_17),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_17),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_17),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_17),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_17),
.B(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1O1Ixp25_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_103),
.B(n_267),
.C(n_430),
.D(n_439),
.Y(n_23)
);

NOR3xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_231),
.C(n_258),
.Y(n_24)
);

NAND2x1_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_188),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_27),
.A2(n_433),
.B(n_434),
.Y(n_432)
);

AOI21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_146),
.B(n_149),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_109),
.Y(n_28)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_29),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_29),
.B(n_110),
.C(n_141),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_29),
.A2(n_109),
.B1(n_147),
.B2(n_148),
.Y(n_435)
);

MAJx2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_47),
.C(n_95),
.Y(n_29)
);

XNOR2x1_ASAP7_75t_SL g187 ( 
.A(n_30),
.B(n_95),
.Y(n_187)
);

XOR2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_42),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_31)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_R g112 ( 
.A(n_32),
.B(n_35),
.C(n_42),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_32),
.B(n_171),
.C(n_174),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_32),
.A2(n_41),
.B1(n_174),
.B2(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_34),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_34),
.Y(n_321)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_39),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_42),
.B(n_262),
.CI(n_263),
.CON(n_261),
.SN(n_261)
);

NOR3xp33_ASAP7_75t_L g439 ( 
.A(n_42),
.B(n_222),
.C(n_264),
.Y(n_439)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_44),
.Y(n_252)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_46),
.Y(n_161)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_48),
.B(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_65),
.C(n_78),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_49),
.B(n_65),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_54),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_50),
.B(n_55),
.C(n_64),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_50),
.A2(n_222),
.B1(n_223),
.B2(n_244),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_50),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_50),
.B(n_135),
.C(n_222),
.Y(n_262)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_53),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_53),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_63),
.B2(n_64),
.Y(n_54)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_55),
.A2(n_63),
.B1(n_376),
.B2(n_378),
.Y(n_375)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_63),
.B(n_135),
.C(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_69),
.C(n_73),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_66),
.A2(n_73),
.B1(n_74),
.B2(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_66),
.Y(n_156)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_69),
.A2(n_70),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_69),
.A2(n_70),
.B1(n_348),
.B2(n_351),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_69),
.B(n_122),
.C(n_348),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g195 ( 
.A(n_78),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_91),
.B2(n_92),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_R g143 ( 
.A1(n_81),
.A2(n_82),
.B1(n_122),
.B2(n_123),
.Y(n_143)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_122),
.C(n_126),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_86),
.C(n_91),
.Y(n_145)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_82),
.B(n_302),
.C(n_308),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_82),
.B(n_302),
.Y(n_314)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_85),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_89),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_90),
.Y(n_369)
);

MAJx2_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_97),
.C(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_92),
.B(n_100),
.Y(n_168)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_94),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_103),
.C(n_106),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_96),
.B(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_97),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_97),
.B(n_163),
.Y(n_166)
);

XOR2x2_ASAP7_75t_SL g167 ( 
.A(n_97),
.B(n_168),
.Y(n_167)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_97),
.B(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_99),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_100),
.A2(n_222),
.B1(n_223),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_100),
.Y(n_264)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_103),
.A2(n_106),
.B1(n_107),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_103),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_105),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_105),
.Y(n_177)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_105),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_107),
.B1(n_114),
.B2(n_117),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_170),
.C(n_176),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_106),
.A2(n_107),
.B1(n_176),
.B2(n_228),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_106),
.B(n_114),
.C(n_118),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_108),
.Y(n_325)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_140),
.Y(n_109)
);

XNOR2x1_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_120),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_111),
.B(n_130),
.C(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_113),
.B1(n_118),
.B2(n_119),
.Y(n_111)
);

INVxp67_ASAP7_75t_SL g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_114),
.Y(n_117)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2x1_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_130),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_121),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_123),
.B1(n_132),
.B2(n_135),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_122),
.B(n_246),
.C(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_122),
.B(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_124),
.Y(n_318)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_143),
.Y(n_142)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_136),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_132),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_132),
.A2(n_242),
.B1(n_243),
.B2(n_245),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_132),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_132),
.A2(n_135),
.B1(n_204),
.B2(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_136),
.Y(n_255)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.C(n_145),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_145),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_149),
.B(n_435),
.Y(n_434)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_182),
.C(n_185),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_151),
.B(n_230),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_169),
.C(n_178),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_192),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.C(n_167),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_154),
.B(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_158),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B(n_166),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_160),
.B1(n_163),
.B2(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_163),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_163),
.B(n_295),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_163),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_166),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_167),
.B(n_416),
.Y(n_415)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_171),
.B(n_201),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_173),
.Y(n_310)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_175),
.Y(n_339)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_183),
.B(n_186),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_229),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_189),
.B(n_229),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.C(n_197),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_191),
.B(n_194),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_197),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_211),
.C(n_225),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_198),
.A2(n_199),
.B1(n_411),
.B2(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_203),
.C(n_208),
.Y(n_199)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_200),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_203),
.B(n_208),
.Y(n_395)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_204),
.Y(n_377)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_211),
.A2(n_225),
.B1(n_226),
.B2(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_211),
.Y(n_413)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_218),
.C(n_222),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_212),
.B(n_390),
.Y(n_389)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_216),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_213),
.B(n_215),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_216),
.B(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_219),
.B(n_223),
.Y(n_390)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_232),
.Y(n_231)
);

A2O1A1O1Ixp25_ASAP7_75t_L g431 ( 
.A1(n_232),
.A2(n_259),
.B(n_432),
.C(n_436),
.D(n_437),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_257),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_233),
.B(n_257),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_234),
.B(n_238),
.C(n_239),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_247),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_254),
.C(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_247)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_248),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_266),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_260),
.B(n_266),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

BUFx24_ASAP7_75t_SL g440 ( 
.A(n_261),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_262),
.B(n_438),
.Y(n_437)
);

INVxp33_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_399),
.B1(n_424),
.B2(n_429),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_379),
.B(n_396),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_352),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_312),
.C(n_329),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_292),
.B2(n_311),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_273),
.B(n_293),
.C(n_301),
.Y(n_361)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

MAJx2_ASAP7_75t_L g359 ( 
.A(n_275),
.B(n_281),
.C(n_286),
.Y(n_359)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_286),
.B2(n_287),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_292),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_300),
.B2(n_301),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_295),
.A2(n_296),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_308),
.B(n_314),
.Y(n_313)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_315),
.C(n_326),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.C(n_322),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_340),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_341),
.C(n_346),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.C(n_336),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_346),
.Y(n_340)
);

OA21x2_ASAP7_75t_L g341 ( 
.A1(n_342),
.A2(n_343),
.B(n_345),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_342),
.B(n_343),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_345),
.B(n_359),
.Y(n_358)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_345),
.B(n_356),
.C(n_359),
.Y(n_387)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_348),
.Y(n_351)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_360),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJx2_ASAP7_75t_L g380 ( 
.A(n_354),
.B(n_355),
.C(n_360),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_358),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_362),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_363),
.C(n_375),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_375),
.Y(n_362)
);

XNOR2x2_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_373),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_370),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_370),
.C(n_392),
.Y(n_391)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_376),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_381),
.Y(n_379)
);

AOI21x1_ASAP7_75t_L g396 ( 
.A1(n_380),
.A2(n_397),
.B(n_398),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_382),
.A2(n_383),
.B1(n_384),
.B2(n_385),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_382),
.B(n_384),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_402),
.C(n_403),
.Y(n_401)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_383),
.B(n_385),
.Y(n_397)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_393),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_388),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_387),
.B(n_389),
.C(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_391),
.Y(n_408)
);

HB1xp67_ASAP7_75t_L g402 ( 
.A(n_393),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_395),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_419),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_405),
.Y(n_400)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_401),
.Y(n_427)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_405),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_409),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_410),
.C(n_414),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_410),
.A2(n_414),
.B1(n_415),
.B2(n_418),
.Y(n_409)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_410),
.Y(n_418)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_419),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_420),
.Y(n_426)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_421),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_427),
.B2(n_428),
.Y(n_424)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);


endmodule