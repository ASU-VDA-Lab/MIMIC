module fake_aes_8352_n_15 (n_1, n_2, n_0, n_15);
input n_1;
input n_2;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
NAND2xp33_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .Y(n_4) );
AND2x4_ASAP7_75t_L g5 ( .A(n_2), .B(n_1), .Y(n_5) );
AO21x2_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_6) );
OAI22xp5_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_5), .Y(n_8) );
AOI33xp33_ASAP7_75t_L g9 ( .A1(n_7), .A2(n_5), .A3(n_4), .B1(n_3), .B2(n_1), .B3(n_0), .Y(n_9) );
A2O1A1Ixp33_ASAP7_75t_L g10 ( .A1(n_8), .A2(n_6), .B(n_2), .C(n_1), .Y(n_10) );
INVx1_ASAP7_75t_SL g11 ( .A(n_8), .Y(n_11) );
OAI31xp33_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_8), .A3(n_9), .B(n_0), .Y(n_12) );
AO221x1_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_2), .B1(n_9), .B2(n_7), .C(n_10), .Y(n_13) );
INVx4_ASAP7_75t_L g14 ( .A(n_13), .Y(n_14) );
AOI22xp33_ASAP7_75t_SL g15 ( .A1(n_14), .A2(n_13), .B1(n_11), .B2(n_12), .Y(n_15) );
endmodule