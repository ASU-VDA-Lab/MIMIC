module fake_ariane_1112_n_1421 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_16, n_273, n_305, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1421);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_16;
input n_273;
input n_305;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1421;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1026;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_967;
wire n_437;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_321;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1370;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1368;
wire n_1211;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_206),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_189),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_143),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_175),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_252),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_14),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_26),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_229),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_89),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_292),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_222),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_283),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_19),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_38),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_258),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_56),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_44),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_97),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_133),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_215),
.Y(n_331)
);

BUFx2_ASAP7_75t_SL g332 ( 
.A(n_242),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_87),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_51),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_137),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_254),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_91),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_102),
.Y(n_338)
);

BUFx10_ASAP7_75t_L g339 ( 
.A(n_232),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_272),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_161),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_81),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_63),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_135),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_36),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_76),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_166),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_149),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_15),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_288),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_224),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_85),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_253),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_219),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_243),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_289),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_297),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_301),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_273),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_120),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_154),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_129),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_95),
.Y(n_363)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_174),
.Y(n_364)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_205),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_73),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_162),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_41),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_230),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_5),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_4),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_279),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_310),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_302),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_168),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_216),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_286),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_66),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_159),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_103),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_52),
.Y(n_381)
);

BUFx10_ASAP7_75t_L g382 ( 
.A(n_96),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_194),
.Y(n_383)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_247),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_241),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_282),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_259),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_126),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_179),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_132),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_300),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_153),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_57),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_92),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_244),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_65),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_48),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_52),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_233),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_107),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_151),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_67),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_240),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_304),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_116),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_148),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_207),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_17),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_280),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_271),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_285),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_181),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_142),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_192),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_198),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_197),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_141),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_227),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_163),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_269),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_193),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_19),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_77),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_18),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_270),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_226),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_200),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_94),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_59),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_121),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_191),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_139),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_209),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_249),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_46),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_71),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_248),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_293),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_245),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_93),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_261),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_235),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_61),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_290),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_239),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_262),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_204),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_28),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_83),
.Y(n_449)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_184),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_18),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_64),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_145),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_86),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_62),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_255),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_44),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_217),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_196),
.Y(n_459)
);

BUFx10_ASAP7_75t_L g460 ( 
.A(n_183),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_13),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_12),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_32),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_40),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_131),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_30),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_214),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_124),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_53),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_178),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_47),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_2),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_260),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_54),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_28),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_264),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_7),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_144),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_90),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_51),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_257),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_23),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_136),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_115),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_265),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_238),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_140),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_256),
.Y(n_488)
);

BUFx5_ASAP7_75t_L g489 ( 
.A(n_246),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_70),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_138),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_84),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_50),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_318),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_341),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_349),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_370),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_451),
.Y(n_499)
);

NOR2xp67_ASAP7_75t_L g500 ( 
.A(n_371),
.B(n_0),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_330),
.Y(n_501)
);

CKINVDCx16_ASAP7_75t_R g502 ( 
.A(n_319),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_457),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_463),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_350),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_317),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_457),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_466),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_336),
.B(n_0),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_324),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g511 ( 
.A(n_475),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_441),
.B(n_1),
.Y(n_512)
);

INVxp33_ASAP7_75t_SL g513 ( 
.A(n_396),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_354),
.Y(n_514)
);

INVxp67_ASAP7_75t_SL g515 ( 
.A(n_368),
.Y(n_515)
);

INVxp67_ASAP7_75t_SL g516 ( 
.A(n_368),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_328),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_371),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_368),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_368),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_442),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_473),
.Y(n_523)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_325),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_339),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_339),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_394),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_464),
.Y(n_528)
);

BUFx6f_ASAP7_75t_SL g529 ( 
.A(n_339),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_382),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_403),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_330),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_407),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_351),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_334),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_438),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_345),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_382),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_382),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_397),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_367),
.B(n_1),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_460),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_460),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_398),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_313),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_408),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_422),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_315),
.Y(n_549)
);

NOR2xp67_ASAP7_75t_L g550 ( 
.A(n_367),
.B(n_2),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_316),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_424),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_461),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_438),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_462),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_323),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_469),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_337),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_338),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_456),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_367),
.B(n_3),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_340),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_471),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_346),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_472),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_347),
.Y(n_567)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_456),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_477),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_480),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_358),
.B(n_4),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_361),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_366),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_375),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_378),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_386),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_400),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_352),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_385),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_493),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_402),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_312),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_351),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_384),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_314),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_365),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_406),
.Y(n_587)
);

NOR2xp67_ASAP7_75t_L g588 ( 
.A(n_348),
.B(n_5),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_320),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_415),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g591 ( 
.A(n_381),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_417),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_321),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_384),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_418),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_322),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_423),
.B(n_6),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_430),
.Y(n_598)
);

HB1xp67_ASAP7_75t_L g599 ( 
.A(n_405),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_432),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_433),
.Y(n_601)
);

NOR2xp67_ASAP7_75t_L g602 ( 
.A(n_348),
.B(n_6),
.Y(n_602)
);

INVxp33_ASAP7_75t_SL g603 ( 
.A(n_332),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_436),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_520),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_515),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_516),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_494),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_542),
.B(n_365),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_496),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_497),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_498),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_571),
.A2(n_458),
.B(n_444),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_499),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_521),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_504),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_542),
.B(n_405),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_542),
.B(n_419),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_584),
.B(n_459),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_517),
.Y(n_620)
);

INVx5_ASAP7_75t_L g621 ( 
.A(n_532),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_532),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_525),
.B(n_484),
.Y(n_623)
);

BUFx2_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_594),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_594),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_501),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_599),
.B(n_419),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_604),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_546),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_501),
.B(n_474),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_549),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_551),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_557),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_534),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_519),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_559),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_603),
.B(n_474),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_560),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_563),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_534),
.B(n_364),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_565),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_583),
.B(n_567),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_572),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_591),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_583),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_573),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_526),
.B(n_530),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_574),
.B(n_450),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_575),
.B(n_490),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_576),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_577),
.B(n_440),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_581),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_587),
.B(n_387),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_538),
.B(n_486),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_590),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_592),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_595),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_512),
.B(n_488),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_539),
.B(n_326),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_598),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_543),
.B(n_327),
.Y(n_662)
);

AND2x6_ASAP7_75t_L g663 ( 
.A(n_541),
.B(n_387),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_329),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_600),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_603),
.B(n_331),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_601),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_582),
.B(n_333),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_513),
.A2(n_342),
.B1(n_343),
.B2(n_335),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_562),
.Y(n_670)
);

INVx5_ASAP7_75t_L g671 ( 
.A(n_506),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_522),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_597),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_509),
.Y(n_674)
);

BUFx8_ASAP7_75t_L g675 ( 
.A(n_529),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_508),
.B(n_387),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_570),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_511),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_550),
.Y(n_679)
);

INVx3_ASAP7_75t_L g680 ( 
.A(n_523),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_585),
.Y(n_681)
);

AND2x4_ASAP7_75t_L g682 ( 
.A(n_588),
.B(n_387),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_589),
.Y(n_683)
);

HB1xp67_ASAP7_75t_L g684 ( 
.A(n_535),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_500),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_602),
.A2(n_489),
.B(n_353),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_553),
.B(n_344),
.Y(n_687)
);

OA21x2_ASAP7_75t_L g688 ( 
.A1(n_510),
.A2(n_356),
.B(n_355),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_537),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_569),
.B(n_357),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_529),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_540),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_593),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_596),
.B(n_359),
.Y(n_694)
);

AND2x6_ASAP7_75t_L g695 ( 
.A(n_586),
.B(n_489),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_645),
.B(n_502),
.Y(n_696)
);

NAND2xp33_ASAP7_75t_SL g697 ( 
.A(n_683),
.B(n_578),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_622),
.Y(n_698)
);

AOI22xp33_ASAP7_75t_L g699 ( 
.A1(n_673),
.A2(n_513),
.B1(n_524),
.B2(n_586),
.Y(n_699)
);

OR2x6_ASAP7_75t_L g700 ( 
.A(n_624),
.B(n_495),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_670),
.B(n_489),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_622),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_608),
.Y(n_703)
);

NOR3xp33_ASAP7_75t_L g704 ( 
.A(n_638),
.B(n_648),
.C(n_672),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_673),
.A2(n_524),
.B1(n_547),
.B2(n_545),
.Y(n_705)
);

INVxp67_ASAP7_75t_SL g706 ( 
.A(n_672),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_610),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_611),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_670),
.B(n_548),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_617),
.B(n_489),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_612),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_672),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_609),
.B(n_660),
.Y(n_713)
);

INVx2_ASAP7_75t_SL g714 ( 
.A(n_641),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_690),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_663),
.Y(n_716)
);

BUFx4f_ASAP7_75t_L g717 ( 
.A(n_683),
.Y(n_717)
);

INVxp67_ASAP7_75t_SL g718 ( 
.A(n_680),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_662),
.B(n_552),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_677),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_625),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_625),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_626),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_678),
.B(n_579),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_626),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_661),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_636),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_635),
.Y(n_728)
);

INVxp33_ASAP7_75t_L g729 ( 
.A(n_628),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_617),
.B(n_489),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_636),
.Y(n_731)
);

INVx5_ASAP7_75t_L g732 ( 
.A(n_663),
.Y(n_732)
);

NAND2x1p5_ASAP7_75t_L g733 ( 
.A(n_683),
.B(n_554),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_614),
.Y(n_734)
);

AND2x2_ASAP7_75t_SL g735 ( 
.A(n_659),
.B(n_505),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_615),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_683),
.B(n_578),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_635),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_690),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_616),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_620),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_661),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_678),
.B(n_514),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_615),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_661),
.Y(n_745)
);

BUFx8_ASAP7_75t_SL g746 ( 
.A(n_677),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_L g747 ( 
.A(n_663),
.B(n_556),
.Y(n_747)
);

BUFx10_ASAP7_75t_L g748 ( 
.A(n_694),
.Y(n_748)
);

INVx8_ASAP7_75t_L g749 ( 
.A(n_695),
.Y(n_749)
);

NOR2x1p5_ASAP7_75t_L g750 ( 
.A(n_693),
.B(n_558),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_615),
.Y(n_751)
);

AND2x6_ASAP7_75t_L g752 ( 
.A(n_691),
.B(n_618),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_635),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_615),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_635),
.Y(n_755)
);

BUFx3_ASAP7_75t_L g756 ( 
.A(n_627),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_680),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_693),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_661),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_639),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_674),
.B(n_564),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_646),
.Y(n_762)
);

INVx4_ASAP7_75t_SL g763 ( 
.A(n_663),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_646),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_639),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_655),
.A2(n_674),
.B1(n_669),
.B2(n_680),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_691),
.B(n_489),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_675),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_664),
.B(n_666),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_647),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_675),
.Y(n_772)
);

INVx3_ASAP7_75t_L g773 ( 
.A(n_646),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_606),
.B(n_566),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_646),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_649),
.B(n_580),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_663),
.A2(n_489),
.B1(n_362),
.B2(n_363),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_653),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_SL g779 ( 
.A(n_675),
.B(n_527),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_605),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_649),
.B(n_531),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_627),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_674),
.B(n_360),
.Y(n_783)
);

INVx3_ASAP7_75t_L g784 ( 
.A(n_621),
.Y(n_784)
);

A2O1A1Ixp33_ASAP7_75t_L g785 ( 
.A1(n_709),
.A2(n_613),
.B(n_659),
.C(n_681),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_776),
.B(n_684),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_770),
.B(n_681),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_709),
.B(n_650),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_726),
.Y(n_789)
);

INVx3_ASAP7_75t_L g790 ( 
.A(n_728),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_758),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_706),
.B(n_650),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_713),
.B(n_618),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_706),
.B(n_712),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_703),
.Y(n_795)
);

XOR2xp5_ASAP7_75t_L g796 ( 
.A(n_769),
.B(n_533),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_707),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_781),
.B(n_689),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_708),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_770),
.B(n_692),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_698),
.Y(n_801)
);

NOR2x1p5_ASAP7_75t_L g802 ( 
.A(n_772),
.B(n_691),
.Y(n_802)
);

OAI22xp33_ASAP7_75t_L g803 ( 
.A1(n_766),
.A2(n_674),
.B1(n_655),
.B2(n_671),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_711),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_726),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_746),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_702),
.Y(n_807)
);

NOR2x1p5_ASAP7_75t_L g808 ( 
.A(n_696),
.B(n_694),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_717),
.B(n_694),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_724),
.B(n_628),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_712),
.B(n_687),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_721),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_720),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_734),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_728),
.Y(n_815)
);

AOI22xp5_ASAP7_75t_L g816 ( 
.A1(n_766),
.A2(n_663),
.B1(n_695),
.B2(n_659),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_717),
.B(n_687),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_718),
.B(n_687),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_740),
.Y(n_819)
);

AOI22xp5_ASAP7_75t_L g820 ( 
.A1(n_713),
.A2(n_695),
.B1(n_655),
.B2(n_676),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_748),
.B(n_671),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_722),
.Y(n_822)
);

INVx4_ASAP7_75t_L g823 ( 
.A(n_749),
.Y(n_823)
);

AOI22xp33_ASAP7_75t_L g824 ( 
.A1(n_714),
.A2(n_695),
.B1(n_688),
.B2(n_682),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_723),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_718),
.B(n_668),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_725),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_748),
.B(n_671),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_756),
.B(n_655),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_757),
.B(n_695),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_761),
.B(n_671),
.Y(n_831)
);

NAND3xp33_ASAP7_75t_L g832 ( 
.A(n_704),
.B(n_623),
.C(n_629),
.Y(n_832)
);

INVx8_ASAP7_75t_L g833 ( 
.A(n_752),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_743),
.B(n_643),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_733),
.B(n_671),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_741),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_733),
.B(n_679),
.Y(n_837)
);

AOI22xp33_ASAP7_75t_L g838 ( 
.A1(n_729),
.A2(n_688),
.B1(n_682),
.B2(n_631),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_757),
.B(n_676),
.Y(n_839)
);

BUFx12f_ASAP7_75t_SL g840 ( 
.A(n_700),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_726),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_760),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_719),
.B(n_619),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_699),
.B(n_685),
.Y(n_844)
);

NOR2xp67_ASAP7_75t_L g845 ( 
.A(n_716),
.B(n_621),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_765),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_727),
.Y(n_847)
);

INVx2_ASAP7_75t_SL g848 ( 
.A(n_715),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_719),
.B(n_652),
.Y(n_849)
);

OAI221xp5_ASAP7_75t_L g850 ( 
.A1(n_699),
.A2(n_644),
.B1(n_667),
.B2(n_630),
.C(n_632),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_729),
.B(n_739),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_767),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_704),
.A2(n_752),
.B1(n_735),
.B2(n_777),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_705),
.B(n_774),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_774),
.B(n_607),
.Y(n_855)
);

INVxp67_ASAP7_75t_L g856 ( 
.A(n_746),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_705),
.B(n_633),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_752),
.A2(n_654),
.B1(n_688),
.B2(n_658),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_735),
.B(n_634),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_731),
.Y(n_860)
);

AO22x2_ASAP7_75t_L g861 ( 
.A1(n_783),
.A2(n_555),
.B1(n_561),
.B2(n_536),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_752),
.A2(n_777),
.B1(n_747),
.B2(n_783),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_782),
.B(n_536),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_752),
.B(n_654),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_782),
.B(n_697),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_771),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_780),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_778),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_710),
.B(n_631),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_738),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_710),
.B(n_631),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_730),
.B(n_637),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_726),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_738),
.B(n_640),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_750),
.B(n_763),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_700),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_730),
.A2(n_658),
.B1(n_665),
.B2(n_653),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_800),
.B(n_555),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_847),
.Y(n_879)
);

INVx4_ASAP7_75t_L g880 ( 
.A(n_833),
.Y(n_880)
);

OAI21xp5_ASAP7_75t_L g881 ( 
.A1(n_785),
.A2(n_613),
.B(n_701),
.Y(n_881)
);

NAND2x1_ASAP7_75t_L g882 ( 
.A(n_823),
.B(n_753),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_813),
.Y(n_883)
);

AND2x4_ASAP7_75t_SL g884 ( 
.A(n_875),
.B(n_700),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_787),
.B(n_737),
.Y(n_885)
);

OAI21xp5_ASAP7_75t_L g886 ( 
.A1(n_830),
.A2(n_701),
.B(n_686),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_843),
.B(n_768),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_793),
.A2(n_749),
.B1(n_568),
.B2(n_561),
.Y(n_888)
);

AND2x4_ASAP7_75t_L g889 ( 
.A(n_875),
.B(n_763),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_833),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_826),
.A2(n_749),
.B(n_732),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_794),
.A2(n_732),
.B(n_716),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_833),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_793),
.A2(n_732),
.B(n_716),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_854),
.B(n_568),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_788),
.B(n_768),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_872),
.A2(n_732),
.B(n_716),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_795),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_811),
.A2(n_818),
.B(n_839),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_791),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_806),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_860),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_797),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_832),
.A2(n_686),
.B(n_742),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_849),
.B(n_768),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_853),
.A2(n_759),
.B(n_745),
.C(n_642),
.Y(n_906)
);

O2A1O1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_792),
.A2(n_651),
.B(n_657),
.C(n_656),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_817),
.A2(n_773),
.B(n_762),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_867),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_809),
.A2(n_773),
.B(n_764),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_803),
.B(n_779),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_786),
.B(n_518),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_863),
.B(n_518),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_799),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_804),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_810),
.B(n_528),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_801),
.Y(n_917)
);

AO21x1_ASAP7_75t_L g918 ( 
.A1(n_862),
.A2(n_682),
.B(n_755),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_855),
.B(n_768),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_807),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_814),
.B(n_768),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_832),
.A2(n_862),
.B(n_857),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_798),
.B(n_528),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_853),
.A2(n_665),
.B(n_775),
.C(n_744),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_819),
.B(n_736),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_836),
.B(n_751),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_820),
.A2(n_754),
.B1(n_507),
.B2(n_503),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_851),
.B(n_763),
.Y(n_928)
);

OAI22x1_ASAP7_75t_L g929 ( 
.A1(n_808),
.A2(n_507),
.B1(n_503),
.B2(n_605),
.Y(n_929)
);

O2A1O1Ixp5_ASAP7_75t_L g930 ( 
.A1(n_865),
.A2(n_784),
.B(n_621),
.C(n_9),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_859),
.B(n_784),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_869),
.A2(n_372),
.B(n_369),
.Y(n_932)
);

NOR2xp33_ASAP7_75t_L g933 ( 
.A(n_844),
.B(n_621),
.Y(n_933)
);

INVx4_ASAP7_75t_L g934 ( 
.A(n_829),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_871),
.B(n_621),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_842),
.Y(n_936)
);

AOI21x1_ASAP7_75t_L g937 ( 
.A1(n_864),
.A2(n_374),
.B(n_373),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_874),
.A2(n_377),
.B(n_376),
.Y(n_938)
);

AOI22xp5_ASAP7_75t_L g939 ( 
.A1(n_820),
.A2(n_816),
.B1(n_829),
.B2(n_831),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_840),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_796),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_816),
.B(n_379),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_848),
.B(n_380),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_834),
.B(n_383),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_846),
.B(n_388),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_790),
.A2(n_390),
.B(n_389),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_852),
.B(n_391),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_866),
.B(n_392),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_850),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_877),
.A2(n_492),
.B(n_395),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_877),
.B(n_393),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_L g952 ( 
.A(n_856),
.B(n_401),
.C(n_399),
.Y(n_952)
);

NAND2x1p5_ASAP7_75t_L g953 ( 
.A(n_823),
.B(n_55),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_949),
.B(n_838),
.Y(n_954)
);

AO21x1_ASAP7_75t_L g955 ( 
.A1(n_922),
.A2(n_858),
.B(n_837),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_898),
.Y(n_956)
);

NAND2xp33_ASAP7_75t_SL g957 ( 
.A(n_885),
.B(n_802),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_878),
.A2(n_858),
.B(n_868),
.C(n_824),
.Y(n_958)
);

INVx4_ASAP7_75t_L g959 ( 
.A(n_934),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_895),
.B(n_861),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_912),
.B(n_861),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_903),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_914),
.B(n_815),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_915),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_907),
.A2(n_835),
.B(n_828),
.C(n_821),
.Y(n_965)
);

OAI21xp33_ASAP7_75t_SL g966 ( 
.A1(n_939),
.A2(n_870),
.B(n_815),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_889),
.Y(n_967)
);

OAI21xp33_ASAP7_75t_SL g968 ( 
.A1(n_887),
.A2(n_870),
.B(n_873),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_879),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_913),
.A2(n_876),
.B(n_822),
.C(n_825),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_883),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_899),
.A2(n_805),
.B(n_789),
.Y(n_972)
);

INVx4_ASAP7_75t_L g973 ( 
.A(n_934),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_916),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_889),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_902),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_923),
.B(n_812),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_909),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_880),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_881),
.A2(n_827),
.B(n_845),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_919),
.A2(n_805),
.B(n_789),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_936),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_905),
.A2(n_896),
.B(n_881),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_888),
.B(n_789),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_896),
.A2(n_841),
.B(n_805),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_911),
.B(n_841),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_880),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_927),
.B(n_841),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_888),
.B(n_404),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_893),
.B(n_940),
.Y(n_990)
);

AO32x1_ASAP7_75t_L g991 ( 
.A1(n_918),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_991)
);

OR2x6_ASAP7_75t_L g992 ( 
.A(n_901),
.B(n_845),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_893),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_884),
.B(n_8),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_917),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_944),
.B(n_10),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_SL g997 ( 
.A1(n_921),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_900),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_922),
.A2(n_410),
.B(n_411),
.C(n_409),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_886),
.A2(n_413),
.B(n_412),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_941),
.B(n_11),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_890),
.Y(n_1002)
);

AOI22xp33_ASAP7_75t_L g1003 ( 
.A1(n_929),
.A2(n_491),
.B1(n_487),
.B2(n_485),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_945),
.A2(n_947),
.B1(n_948),
.B2(n_951),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_931),
.A2(n_483),
.B(n_481),
.C(n_479),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_886),
.A2(n_416),
.B(n_414),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_920),
.Y(n_1007)
);

NAND3xp33_ASAP7_75t_L g1008 ( 
.A(n_906),
.B(n_421),
.C(n_420),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_925),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_952),
.B(n_14),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_890),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_928),
.B(n_478),
.Y(n_1012)
);

NOR2xp67_ASAP7_75t_SL g1013 ( 
.A(n_943),
.B(n_425),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_950),
.B(n_476),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_942),
.A2(n_470),
.B(n_468),
.C(n_467),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_891),
.A2(n_894),
.B(n_935),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_977),
.B(n_971),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_1016),
.A2(n_904),
.B(n_924),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_972),
.A2(n_904),
.B(n_892),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_974),
.B(n_926),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_983),
.A2(n_933),
.B(n_908),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_998),
.Y(n_1022)
);

OAI21x1_ASAP7_75t_L g1023 ( 
.A1(n_980),
.A2(n_910),
.B(n_953),
.Y(n_1023)
);

CKINVDCx20_ASAP7_75t_R g1024 ( 
.A(n_992),
.Y(n_1024)
);

AOI31xp67_ASAP7_75t_L g1025 ( 
.A1(n_984),
.A2(n_937),
.A3(n_930),
.B(n_953),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_1004),
.A2(n_897),
.B(n_932),
.Y(n_1026)
);

AOI221x1_ASAP7_75t_L g1027 ( 
.A1(n_989),
.A2(n_946),
.B1(n_938),
.B2(n_20),
.C(n_21),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_966),
.A2(n_882),
.B(n_427),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_960),
.B(n_15),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_956),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_994),
.Y(n_1031)
);

AOI221xp5_ASAP7_75t_L g1032 ( 
.A1(n_961),
.A2(n_465),
.B1(n_455),
.B2(n_454),
.C(n_453),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_985),
.A2(n_60),
.B(n_58),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_986),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_996),
.A2(n_452),
.B(n_449),
.C(n_447),
.Y(n_1035)
);

AOI31xp67_ASAP7_75t_L g1036 ( 
.A1(n_1014),
.A2(n_446),
.A3(n_445),
.B(n_443),
.Y(n_1036)
);

AO31x2_ASAP7_75t_L g1037 ( 
.A1(n_955),
.A2(n_155),
.A3(n_311),
.B(n_309),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1009),
.B(n_16),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_969),
.Y(n_1039)
);

O2A1O1Ixp5_ASAP7_75t_L g1040 ( 
.A1(n_957),
.A2(n_16),
.B(n_20),
.C(n_21),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_976),
.Y(n_1041)
);

AO21x2_ASAP7_75t_L g1042 ( 
.A1(n_958),
.A2(n_428),
.B(n_426),
.Y(n_1042)
);

OA21x2_ASAP7_75t_L g1043 ( 
.A1(n_981),
.A2(n_431),
.B(n_429),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_978),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_954),
.B(n_22),
.Y(n_1045)
);

INVx3_ASAP7_75t_SL g1046 ( 
.A(n_1001),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_967),
.Y(n_1047)
);

AO32x2_ASAP7_75t_L g1048 ( 
.A1(n_991),
.A2(n_22),
.A3(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_SL g1049 ( 
.A1(n_999),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_962),
.B(n_27),
.Y(n_1050)
);

NOR2x1_ASAP7_75t_L g1051 ( 
.A(n_992),
.B(n_434),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_968),
.A2(n_439),
.B(n_437),
.Y(n_1052)
);

AO32x2_ASAP7_75t_L g1053 ( 
.A1(n_991),
.A2(n_27),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1000),
.A2(n_29),
.B(n_31),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_964),
.B(n_32),
.Y(n_1055)
);

NOR2xp67_ASAP7_75t_SL g1056 ( 
.A(n_959),
.B(n_33),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_982),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_970),
.A2(n_33),
.B(n_34),
.C(n_35),
.Y(n_1058)
);

AO32x2_ASAP7_75t_L g1059 ( 
.A1(n_959),
.A2(n_34),
.A3(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_995),
.Y(n_1060)
);

AND2x6_ASAP7_75t_L g1061 ( 
.A(n_967),
.B(n_68),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_967),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1007),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_975),
.B(n_994),
.Y(n_1064)
);

OR2x2_ASAP7_75t_L g1065 ( 
.A(n_988),
.B(n_37),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_1006),
.A2(n_167),
.A3(n_307),
.B(n_306),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_975),
.B(n_973),
.Y(n_1067)
);

AO31x2_ASAP7_75t_L g1068 ( 
.A1(n_1005),
.A2(n_164),
.A3(n_305),
.B(n_303),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_975),
.B(n_38),
.Y(n_1069)
);

BUFx12f_ASAP7_75t_L g1070 ( 
.A(n_979),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_963),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1012),
.A2(n_160),
.B(n_299),
.Y(n_1072)
);

AOI21x1_ASAP7_75t_SL g1073 ( 
.A1(n_1010),
.A2(n_39),
.B(n_40),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_1015),
.A2(n_165),
.A3(n_298),
.B(n_296),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_965),
.A2(n_157),
.B(n_295),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_1002),
.A2(n_156),
.B(n_294),
.Y(n_1076)
);

CKINVDCx11_ASAP7_75t_R g1077 ( 
.A(n_979),
.Y(n_1077)
);

AO32x2_ASAP7_75t_L g1078 ( 
.A1(n_973),
.A2(n_997),
.A3(n_993),
.B1(n_1003),
.B2(n_1008),
.Y(n_1078)
);

NOR2x1_ASAP7_75t_R g1079 ( 
.A(n_993),
.B(n_39),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1011),
.Y(n_1080)
);

INVx5_ASAP7_75t_L g1081 ( 
.A(n_979),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1030),
.Y(n_1082)
);

OAI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1017),
.A2(n_987),
.B1(n_990),
.B2(n_1011),
.Y(n_1083)
);

INVx6_ASAP7_75t_L g1084 ( 
.A(n_1070),
.Y(n_1084)
);

OR2x2_ASAP7_75t_SL g1085 ( 
.A(n_1065),
.B(n_987),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1045),
.A2(n_1002),
.B1(n_1011),
.B2(n_987),
.Y(n_1086)
);

OAI21xp33_ASAP7_75t_L g1087 ( 
.A1(n_1054),
.A2(n_1013),
.B(n_42),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_1022),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1039),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1057),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_1060),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1046),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_1092)
);

INVxp67_ASAP7_75t_L g1093 ( 
.A(n_1020),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1041),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_1094)
);

INVx6_ASAP7_75t_L g1095 ( 
.A(n_1081),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_1077),
.Y(n_1096)
);

INVx2_ASAP7_75t_L g1097 ( 
.A(n_1044),
.Y(n_1097)
);

CKINVDCx11_ASAP7_75t_R g1098 ( 
.A(n_1024),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1063),
.Y(n_1099)
);

AND2x2_ASAP7_75t_L g1100 ( 
.A(n_1064),
.B(n_45),
.Y(n_1100)
);

INVx6_ASAP7_75t_L g1101 ( 
.A(n_1081),
.Y(n_1101)
);

AO22x1_ASAP7_75t_L g1102 ( 
.A1(n_1061),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_1102)
);

CKINVDCx20_ASAP7_75t_R g1103 ( 
.A(n_1047),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1031),
.A2(n_49),
.B1(n_53),
.B2(n_69),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1071),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1034),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1032),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1050),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_1062),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_SL g1110 ( 
.A1(n_1027),
.A2(n_78),
.B(n_79),
.Y(n_1110)
);

CKINVDCx6p67_ASAP7_75t_R g1111 ( 
.A(n_1081),
.Y(n_1111)
);

OAI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1029),
.A2(n_80),
.B1(n_82),
.B2(n_88),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_1064),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_1080),
.Y(n_1114)
);

OAI22xp5_ASAP7_75t_L g1115 ( 
.A1(n_1035),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_1061),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_1116)
);

BUFx10_ASAP7_75t_L g1117 ( 
.A(n_1069),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1058),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1055),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1061),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_SL g1121 ( 
.A1(n_1079),
.A2(n_110),
.B1(n_111),
.B2(n_112),
.Y(n_1121)
);

INVx6_ASAP7_75t_L g1122 ( 
.A(n_1051),
.Y(n_1122)
);

AOI22xp33_ASAP7_75t_L g1123 ( 
.A1(n_1042),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_1038),
.Y(n_1124)
);

INVx2_ASAP7_75t_SL g1125 ( 
.A(n_1067),
.Y(n_1125)
);

OAI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_1026),
.A2(n_118),
.B1(n_119),
.B2(n_122),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1049),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1056),
.A2(n_128),
.B1(n_130),
.B2(n_134),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_SL g1129 ( 
.A1(n_1059),
.A2(n_146),
.B1(n_147),
.B2(n_150),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1078),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1059),
.Y(n_1131)
);

CKINVDCx14_ASAP7_75t_R g1132 ( 
.A(n_1073),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1043),
.A2(n_152),
.B1(n_158),
.B2(n_169),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_1078),
.Y(n_1134)
);

CKINVDCx11_ASAP7_75t_R g1135 ( 
.A(n_1036),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1040),
.Y(n_1136)
);

INVx1_ASAP7_75t_SL g1137 ( 
.A(n_1072),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1066),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1052),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1048),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1037),
.Y(n_1141)
);

AOI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1075),
.A2(n_173),
.B1(n_176),
.B2(n_177),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1018),
.A2(n_180),
.B1(n_182),
.B2(n_185),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1037),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_1105),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1082),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1090),
.B(n_1053),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1134),
.B(n_1053),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1130),
.B(n_1048),
.Y(n_1149)
);

OAI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1110),
.A2(n_1028),
.B1(n_1021),
.B2(n_1019),
.Y(n_1150)
);

INVx2_ASAP7_75t_SL g1151 ( 
.A(n_1106),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1140),
.B(n_1068),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1140),
.B(n_1068),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1091),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1099),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1138),
.A2(n_1023),
.B(n_1033),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_1131),
.B(n_1074),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_1088),
.B(n_1098),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1141),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1144),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1089),
.Y(n_1161)
);

AO21x2_ASAP7_75t_L g1162 ( 
.A1(n_1087),
.A2(n_1127),
.B(n_1136),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1120),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1097),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1108),
.Y(n_1165)
);

BUFx2_ASAP7_75t_L g1166 ( 
.A(n_1120),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1119),
.Y(n_1167)
);

AOI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1126),
.A2(n_1076),
.B(n_1025),
.Y(n_1168)
);

INVx3_ASAP7_75t_L g1169 ( 
.A(n_1137),
.Y(n_1169)
);

HB1xp67_ASAP7_75t_L g1170 ( 
.A(n_1093),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1142),
.A2(n_1074),
.B(n_187),
.Y(n_1171)
);

OAI21x1_ASAP7_75t_L g1172 ( 
.A1(n_1142),
.A2(n_186),
.B(n_188),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1124),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1127),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1125),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_1109),
.Y(n_1176)
);

AO21x2_ASAP7_75t_L g1177 ( 
.A1(n_1087),
.A2(n_190),
.B(n_195),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1083),
.B(n_308),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1084),
.B(n_199),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1086),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1132),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1085),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1143),
.A2(n_201),
.B(n_202),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1135),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_1129),
.B(n_203),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1095),
.Y(n_1186)
);

HB1xp67_ASAP7_75t_L g1187 ( 
.A(n_1114),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1118),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1133),
.A2(n_212),
.B(n_213),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1102),
.Y(n_1190)
);

AND2x2_ASAP7_75t_SL g1191 ( 
.A(n_1128),
.B(n_218),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1096),
.B(n_220),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1095),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1117),
.B(n_291),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1101),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1101),
.Y(n_1196)
);

AND2x2_ASAP7_75t_L g1197 ( 
.A(n_1100),
.B(n_221),
.Y(n_1197)
);

INVx4_ASAP7_75t_L g1198 ( 
.A(n_1111),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1117),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1123),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1103),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1122),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_1115),
.A2(n_223),
.A3(n_225),
.B(n_228),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1112),
.Y(n_1204)
);

OR2x6_ASAP7_75t_L g1205 ( 
.A(n_1182),
.B(n_1096),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1145),
.Y(n_1206)
);

NOR2x1_ASAP7_75t_SL g1207 ( 
.A(n_1199),
.B(n_1182),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1199),
.B(n_1096),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1191),
.A2(n_1121),
.B1(n_1092),
.B2(n_1094),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1199),
.B(n_1084),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1182),
.B(n_1113),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1187),
.B(n_1176),
.Y(n_1212)
);

OR2x2_ASAP7_75t_L g1213 ( 
.A(n_1170),
.B(n_1104),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1184),
.B(n_1122),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1151),
.B(n_1139),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1194),
.B(n_1116),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1165),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1201),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1184),
.B(n_1107),
.Y(n_1219)
);

OR2x6_ASAP7_75t_L g1220 ( 
.A(n_1163),
.B(n_231),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1165),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1169),
.Y(n_1222)
);

NOR2x1_ASAP7_75t_SL g1223 ( 
.A(n_1196),
.B(n_234),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1184),
.B(n_236),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1149),
.B(n_287),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1151),
.B(n_237),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1194),
.B(n_1181),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1165),
.Y(n_1228)
);

AND2x2_ASAP7_75t_L g1229 ( 
.A(n_1149),
.B(n_284),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1164),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1181),
.B(n_250),
.Y(n_1231)
);

O2A1O1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1174),
.A2(n_251),
.B(n_263),
.C(n_266),
.Y(n_1232)
);

OR2x2_ASAP7_75t_L g1233 ( 
.A(n_1146),
.B(n_267),
.Y(n_1233)
);

NOR2x1_ASAP7_75t_SL g1234 ( 
.A(n_1196),
.B(n_268),
.Y(n_1234)
);

AO32x2_ASAP7_75t_L g1235 ( 
.A1(n_1202),
.A2(n_274),
.A3(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1157),
.Y(n_1236)
);

INVxp67_ASAP7_75t_L g1237 ( 
.A(n_1169),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1146),
.B(n_278),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1163),
.B(n_281),
.Y(n_1239)
);

OAI211xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1174),
.A2(n_1150),
.B(n_1204),
.C(n_1190),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1166),
.B(n_1175),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1147),
.B(n_1167),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1147),
.B(n_1167),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1166),
.B(n_1152),
.Y(n_1244)
);

NOR2x1_ASAP7_75t_SL g1245 ( 
.A(n_1196),
.B(n_1177),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1191),
.A2(n_1204),
.B1(n_1190),
.B2(n_1200),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_1158),
.Y(n_1247)
);

AO22x2_ASAP7_75t_L g1248 ( 
.A1(n_1152),
.A2(n_1153),
.B1(n_1155),
.B2(n_1154),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1153),
.B(n_1155),
.Y(n_1249)
);

CKINVDCx6p67_ASAP7_75t_R g1250 ( 
.A(n_1192),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1191),
.A2(n_1172),
.B(n_1185),
.C(n_1200),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1202),
.Y(n_1252)
);

HB1xp67_ASAP7_75t_L g1253 ( 
.A(n_1206),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1230),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1222),
.Y(n_1255)
);

OR2x2_ASAP7_75t_L g1256 ( 
.A(n_1236),
.B(n_1154),
.Y(n_1256)
);

OR2x2_ASAP7_75t_L g1257 ( 
.A(n_1236),
.B(n_1169),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1244),
.B(n_1169),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1227),
.B(n_1173),
.Y(n_1259)
);

OR2x2_ASAP7_75t_L g1260 ( 
.A(n_1242),
.B(n_1173),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1243),
.B(n_1241),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1227),
.B(n_1173),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1249),
.B(n_1180),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1217),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1221),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1228),
.Y(n_1266)
);

BUFx6f_ASAP7_75t_L g1267 ( 
.A(n_1252),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1209),
.A2(n_1185),
.B1(n_1188),
.B2(n_1178),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1241),
.B(n_1180),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1222),
.B(n_1148),
.Y(n_1270)
);

INVx2_ASAP7_75t_SL g1271 ( 
.A(n_1208),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1237),
.B(n_1148),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1248),
.Y(n_1273)
);

NOR2x1_ASAP7_75t_SL g1274 ( 
.A(n_1220),
.B(n_1177),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1216),
.A2(n_1209),
.B1(n_1246),
.B2(n_1177),
.Y(n_1275)
);

AND2x2_ASAP7_75t_L g1276 ( 
.A(n_1237),
.B(n_1162),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1251),
.B(n_1175),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1248),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1248),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1207),
.Y(n_1280)
);

NOR2xp33_ASAP7_75t_SL g1281 ( 
.A(n_1268),
.B(n_1250),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1261),
.B(n_1212),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1256),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1260),
.B(n_1218),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1256),
.Y(n_1285)
);

AND2x4_ASAP7_75t_L g1286 ( 
.A(n_1280),
.B(n_1210),
.Y(n_1286)
);

AOI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1275),
.A2(n_1216),
.B1(n_1251),
.B2(n_1240),
.Y(n_1287)
);

AO21x2_ASAP7_75t_L g1288 ( 
.A1(n_1274),
.A2(n_1245),
.B(n_1162),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1253),
.Y(n_1289)
);

OAI221xp5_ASAP7_75t_L g1290 ( 
.A1(n_1277),
.A2(n_1240),
.B1(n_1213),
.B2(n_1220),
.C(n_1229),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1254),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1259),
.B(n_1247),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1271),
.Y(n_1293)
);

BUFx2_ASAP7_75t_SL g1294 ( 
.A(n_1271),
.Y(n_1294)
);

NOR3xp33_ASAP7_75t_L g1295 ( 
.A(n_1276),
.B(n_1172),
.C(n_1225),
.Y(n_1295)
);

INVxp67_ASAP7_75t_SL g1296 ( 
.A(n_1257),
.Y(n_1296)
);

OR2x6_ASAP7_75t_L g1297 ( 
.A(n_1280),
.B(n_1220),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1264),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1264),
.B(n_1162),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1261),
.B(n_1214),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1265),
.Y(n_1301)
);

AND2x2_ASAP7_75t_L g1302 ( 
.A(n_1294),
.B(n_1258),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1288),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1298),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1292),
.B(n_1247),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1289),
.B(n_1262),
.Y(n_1306)
);

NOR4xp25_ASAP7_75t_SL g1307 ( 
.A(n_1290),
.B(n_1273),
.C(n_1279),
.D(n_1255),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1288),
.Y(n_1308)
);

INVx1_ASAP7_75t_SL g1309 ( 
.A(n_1284),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1301),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1286),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1283),
.B(n_1263),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1291),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1302),
.B(n_1282),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1310),
.B(n_1309),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1304),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1306),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1312),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1303),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1303),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1311),
.B(n_1293),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1308),
.Y(n_1322)
);

NOR2xp33_ASAP7_75t_L g1323 ( 
.A(n_1305),
.B(n_1300),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1308),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1311),
.B(n_1287),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1313),
.Y(n_1326)
);

OR2x6_ASAP7_75t_L g1327 ( 
.A(n_1313),
.B(n_1297),
.Y(n_1327)
);

OAI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1305),
.A2(n_1281),
.B(n_1295),
.Y(n_1328)
);

NOR2xp33_ASAP7_75t_SL g1329 ( 
.A(n_1328),
.B(n_1281),
.Y(n_1329)
);

AOI31xp33_ASAP7_75t_L g1330 ( 
.A1(n_1328),
.A2(n_1290),
.A3(n_1239),
.B(n_1192),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1314),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1318),
.B(n_1296),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1323),
.B(n_1285),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1316),
.Y(n_1334)
);

OR2x2_ASAP7_75t_L g1335 ( 
.A(n_1315),
.B(n_1257),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1321),
.B(n_1272),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1325),
.B(n_1192),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1317),
.B(n_1286),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1329),
.A2(n_1295),
.B1(n_1326),
.B2(n_1327),
.Y(n_1339)
);

AOI22xp5_ASAP7_75t_SL g1340 ( 
.A1(n_1329),
.A2(n_1334),
.B1(n_1338),
.B2(n_1330),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1332),
.Y(n_1341)
);

OAI21xp33_ASAP7_75t_L g1342 ( 
.A1(n_1331),
.A2(n_1276),
.B(n_1269),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1335),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1333),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1336),
.B(n_1337),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1330),
.A2(n_1297),
.B1(n_1327),
.B2(n_1322),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1330),
.A2(n_1307),
.B1(n_1297),
.B2(n_1327),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1340),
.A2(n_1270),
.B1(n_1299),
.B2(n_1273),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1343),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1341),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_L g1351 ( 
.A(n_1344),
.B(n_1324),
.Y(n_1351)
);

AOI21xp33_ASAP7_75t_SL g1352 ( 
.A1(n_1347),
.A2(n_1192),
.B(n_1319),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1345),
.B(n_1299),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1342),
.B(n_1320),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1349),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1351),
.B(n_1339),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1350),
.Y(n_1357)
);

XNOR2x1_ASAP7_75t_L g1358 ( 
.A(n_1348),
.B(n_1347),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1354),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1352),
.Y(n_1360)
);

INVxp67_ASAP7_75t_L g1361 ( 
.A(n_1353),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1348),
.A2(n_1346),
.B(n_1274),
.Y(n_1362)
);

OAI211xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1350),
.A2(n_1232),
.B(n_1178),
.C(n_1233),
.Y(n_1363)
);

NOR3xp33_ASAP7_75t_L g1364 ( 
.A(n_1356),
.B(n_1179),
.C(n_1197),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1361),
.B(n_1272),
.Y(n_1365)
);

NAND2xp33_ASAP7_75t_SL g1366 ( 
.A(n_1355),
.B(n_1198),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1360),
.B(n_1198),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_1359),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1357),
.B(n_1258),
.Y(n_1369)
);

O2A1O1Ixp33_ASAP7_75t_L g1370 ( 
.A1(n_1363),
.A2(n_1232),
.B(n_1177),
.C(n_1197),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1358),
.B(n_1278),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1368),
.B(n_1362),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1370),
.A2(n_1367),
.B(n_1366),
.Y(n_1373)
);

NAND4xp25_ASAP7_75t_L g1374 ( 
.A(n_1365),
.B(n_1198),
.C(n_1239),
.D(n_1231),
.Y(n_1374)
);

AOI222xp33_ASAP7_75t_L g1375 ( 
.A1(n_1371),
.A2(n_1278),
.B1(n_1219),
.B2(n_1224),
.C1(n_1215),
.C2(n_1172),
.Y(n_1375)
);

NAND2xp33_ASAP7_75t_R g1376 ( 
.A(n_1369),
.B(n_1189),
.Y(n_1376)
);

AOI222xp33_ASAP7_75t_L g1377 ( 
.A1(n_1364),
.A2(n_1215),
.B1(n_1171),
.B2(n_1234),
.C1(n_1223),
.C2(n_1226),
.Y(n_1377)
);

AOI322xp5_ASAP7_75t_L g1378 ( 
.A1(n_1371),
.A2(n_1211),
.A3(n_1226),
.B1(n_1238),
.B2(n_1266),
.C1(n_1162),
.C2(n_1235),
.Y(n_1378)
);

AOI21xp33_ASAP7_75t_SL g1379 ( 
.A1(n_1372),
.A2(n_1183),
.B(n_1189),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1373),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_1374),
.Y(n_1381)
);

NAND4xp25_ASAP7_75t_SL g1382 ( 
.A(n_1378),
.B(n_1198),
.C(n_1193),
.D(n_1195),
.Y(n_1382)
);

XNOR2xp5_ASAP7_75t_L g1383 ( 
.A(n_1376),
.B(n_1205),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1377),
.A2(n_1375),
.B(n_1189),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1373),
.B(n_1260),
.Y(n_1385)
);

AOI222xp33_ASAP7_75t_L g1386 ( 
.A1(n_1372),
.A2(n_1171),
.B1(n_1211),
.B2(n_1235),
.C1(n_1202),
.C2(n_1161),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1372),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1373),
.B(n_1267),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1387),
.Y(n_1389)
);

AOI22xp5_ASAP7_75t_L g1390 ( 
.A1(n_1382),
.A2(n_1202),
.B1(n_1205),
.B2(n_1189),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1380),
.B(n_1267),
.Y(n_1391)
);

NAND4xp75_ASAP7_75t_L g1392 ( 
.A(n_1388),
.B(n_1235),
.C(n_1193),
.D(n_1195),
.Y(n_1392)
);

NAND4xp75_ASAP7_75t_L g1393 ( 
.A(n_1384),
.B(n_1235),
.C(n_1203),
.D(n_1186),
.Y(n_1393)
);

AO22x2_ASAP7_75t_L g1394 ( 
.A1(n_1385),
.A2(n_1203),
.B1(n_1186),
.B2(n_1175),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1383),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1381),
.B(n_1267),
.Y(n_1396)
);

NOR2xp33_ASAP7_75t_L g1397 ( 
.A(n_1381),
.B(n_1205),
.Y(n_1397)
);

A2O1A1Ixp33_ASAP7_75t_SL g1398 ( 
.A1(n_1386),
.A2(n_1186),
.B(n_1159),
.C(n_1203),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1379),
.Y(n_1399)
);

XOR2xp5_ASAP7_75t_L g1400 ( 
.A(n_1380),
.B(n_1267),
.Y(n_1400)
);

NOR3xp33_ASAP7_75t_L g1401 ( 
.A(n_1380),
.B(n_1183),
.C(n_1168),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1389),
.B(n_1267),
.Y(n_1402)
);

NOR2xp67_ASAP7_75t_SL g1403 ( 
.A(n_1395),
.B(n_1252),
.Y(n_1403)
);

NOR3xp33_ASAP7_75t_SL g1404 ( 
.A(n_1396),
.B(n_1203),
.C(n_1252),
.Y(n_1404)
);

AOI31xp33_ASAP7_75t_SL g1405 ( 
.A1(n_1391),
.A2(n_1397),
.A3(n_1400),
.B(n_1401),
.Y(n_1405)
);

AND2x4_ASAP7_75t_L g1406 ( 
.A(n_1399),
.B(n_1252),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1402),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1406),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1405),
.B(n_1390),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1407),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1408),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1410),
.A2(n_1409),
.B1(n_1411),
.B2(n_1394),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1410),
.Y(n_1413)
);

OR3x2_ASAP7_75t_L g1414 ( 
.A(n_1413),
.B(n_1403),
.C(n_1404),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1412),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1415),
.A2(n_1393),
.B1(n_1392),
.B2(n_1394),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1416),
.A2(n_1414),
.B1(n_1398),
.B2(n_1168),
.Y(n_1417)
);

AOI211xp5_ASAP7_75t_L g1418 ( 
.A1(n_1417),
.A2(n_1203),
.B(n_1159),
.C(n_1156),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1418),
.Y(n_1419)
);

OAI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1419),
.A2(n_1203),
.B1(n_1160),
.B2(n_1254),
.C(n_1161),
.Y(n_1420)
);

AOI211xp5_ASAP7_75t_L g1421 ( 
.A1(n_1420),
.A2(n_1156),
.B(n_1160),
.C(n_1164),
.Y(n_1421)
);


endmodule