module fake_jpeg_1559_n_659 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_659);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_659;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_378;
wire n_133;
wire n_132;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx8_ASAP7_75t_SL g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_15),
.B(n_17),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_60),
.Y(n_137)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_61),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g138 ( 
.A(n_63),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_66),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_9),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_67),
.B(n_72),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_68),
.Y(n_146)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_69),
.Y(n_174)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_10),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_74),
.B(n_86),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_33),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_75),
.B(n_85),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_79),
.Y(n_195)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_81),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_82),
.Y(n_184)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_20),
.B(n_10),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_87),
.Y(n_147)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_88),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_89),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_48),
.Y(n_90)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_90),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_10),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_91),
.B(n_121),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_92),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_93),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_95),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_43),
.B(n_8),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_96),
.B(n_113),
.Y(n_153)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_41),
.Y(n_97)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_97),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_98),
.Y(n_173)
);

BUFx8_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

CKINVDCx6p67_ASAP7_75t_R g134 ( 
.A(n_99),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_101),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_49),
.Y(n_102)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_102),
.Y(n_204)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_103),
.Y(n_135)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_104),
.Y(n_156)
);

BUFx24_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_105),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_49),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_106),
.Y(n_140)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_21),
.Y(n_107)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_41),
.Y(n_108)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_108),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_36),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_110),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_111),
.Y(n_171)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_19),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_57),
.Y(n_114)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_114),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_28),
.B(n_11),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_115),
.B(n_13),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_116),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_57),
.Y(n_117)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_21),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_21),
.Y(n_119)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_119),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_122),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_34),
.B(n_11),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_28),
.Y(n_122)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_21),
.Y(n_123)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_123),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_50),
.Y(n_125)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_50),
.Y(n_126)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_50),
.Y(n_127)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_44),
.Y(n_128)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_45),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_129),
.Y(n_193)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_50),
.Y(n_130)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_130),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_118),
.A2(n_28),
.B1(n_52),
.B2(n_55),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_144),
.A2(n_169),
.B1(n_175),
.B2(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_86),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_157),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_120),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_99),
.A2(n_52),
.B1(n_34),
.B2(n_55),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_94),
.A2(n_40),
.B1(n_35),
.B2(n_42),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_170),
.A2(n_194),
.B1(n_199),
.B2(n_25),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_63),
.A2(n_52),
.B1(n_40),
.B2(n_42),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_70),
.A2(n_52),
.B1(n_35),
.B2(n_27),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_92),
.A2(n_52),
.B1(n_27),
.B2(n_30),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_179),
.A2(n_187),
.B1(n_203),
.B2(n_105),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_108),
.B(n_30),
.C(n_29),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_180),
.B(n_19),
.Y(n_253)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_107),
.B(n_58),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_185),
.B(n_192),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_106),
.A2(n_29),
.B1(n_56),
.B2(n_51),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_119),
.B(n_58),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_95),
.A2(n_56),
.B1(n_51),
.B2(n_43),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_98),
.A2(n_25),
.B1(n_19),
.B2(n_3),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_125),
.B(n_12),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_201),
.B(n_202),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_100),
.B(n_12),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_93),
.A2(n_25),
.B1(n_19),
.B2(n_12),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_111),
.B(n_12),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_205),
.B(n_209),
.Y(n_285)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_69),
.Y(n_207)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_102),
.B(n_7),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_210),
.B(n_16),
.Y(n_289)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_77),
.Y(n_211)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_114),
.B(n_11),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_217),
.B(n_219),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_116),
.B(n_11),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_117),
.Y(n_220)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_129),
.B(n_15),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_0),
.Y(n_256)
);

AOI32xp33_ASAP7_75t_L g225 ( 
.A1(n_142),
.A2(n_145),
.A3(n_153),
.B1(n_133),
.B2(n_167),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_225),
.B(n_246),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_226),
.Y(n_352)
);

INVx11_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_227),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_177),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_228),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_231),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_174),
.A2(n_173),
.B1(n_182),
.B2(n_204),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_233),
.A2(n_261),
.B1(n_271),
.B2(n_241),
.Y(n_324)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_139),
.Y(n_234)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_234),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_235),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_236),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_159),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_237),
.Y(n_333)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_208),
.Y(n_240)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_240),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_222),
.A2(n_73),
.B1(n_90),
.B2(n_89),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_241),
.A2(n_278),
.B1(n_293),
.B2(n_297),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_151),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_243),
.B(n_250),
.Y(n_326)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_160),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_245),
.Y(n_331)
);

AOI32xp33_ASAP7_75t_L g246 ( 
.A1(n_135),
.A2(n_101),
.A3(n_19),
.B1(n_25),
.B2(n_82),
.Y(n_246)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_172),
.Y(n_247)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_247),
.Y(n_313)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_162),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_249),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_159),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_134),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_251),
.B(n_275),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_146),
.Y(n_252)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_252),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g353 ( 
.A(n_253),
.B(n_256),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_183),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_254),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_255),
.Y(n_305)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_141),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_257),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_193),
.B(n_65),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g349 ( 
.A(n_258),
.Y(n_349)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_158),
.Y(n_259)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_259),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_78),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_260),
.B(n_265),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_170),
.A2(n_76),
.B1(n_64),
.B2(n_62),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_168),
.Y(n_263)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_134),
.A2(n_25),
.B(n_19),
.C(n_16),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_161),
.Y(n_266)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_267),
.Y(n_311)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_137),
.Y(n_268)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_268),
.Y(n_325)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_213),
.Y(n_269)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_131),
.Y(n_270)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_270),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_194),
.A2(n_59),
.B1(n_25),
.B2(n_15),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_131),
.Y(n_272)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_272),
.Y(n_344)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_171),
.Y(n_273)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_273),
.Y(n_356)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_274),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_137),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_295),
.B1(n_204),
.B2(n_182),
.Y(n_314)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_218),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_277),
.B(n_279),
.Y(n_346)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_148),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_206),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_282),
.Y(n_354)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_176),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_281),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_163),
.B(n_6),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_200),
.B(n_6),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_283),
.B(n_284),
.Y(n_357)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_196),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_169),
.A2(n_15),
.B(n_17),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_286),
.A2(n_2),
.B(n_3),
.Y(n_362)
);

INVx4_ASAP7_75t_SL g287 ( 
.A(n_152),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_287),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_214),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_288),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_289),
.Y(n_335)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_143),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_290),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_291),
.Y(n_350)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_147),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_292),
.Y(n_359)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_198),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_199),
.A2(n_16),
.B1(n_18),
.B2(n_4),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_136),
.B(n_18),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_296),
.B(n_300),
.Y(n_364)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_136),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_174),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_299),
.Y(n_317)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_173),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_150),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_149),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_302),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_150),
.B(n_18),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_140),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_303),
.B(n_216),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_216),
.B(n_2),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_138),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_229),
.A2(n_203),
.B1(n_144),
.B2(n_187),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_308),
.A2(n_342),
.B1(n_298),
.B2(n_166),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_314),
.A2(n_347),
.B1(n_358),
.B2(n_363),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_253),
.B(n_140),
.C(n_156),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_315),
.B(n_328),
.C(n_338),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_304),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_256),
.A2(n_175),
.B(n_178),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_321),
.A2(n_291),
.B(n_268),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_324),
.A2(n_255),
.B1(n_252),
.B2(n_279),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_230),
.B(n_179),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g376 ( 
.A(n_332),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_248),
.B(n_138),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_285),
.B(n_223),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_340),
.B(n_265),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_229),
.A2(n_223),
.B1(n_221),
.B2(n_215),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_231),
.A2(n_221),
.B1(n_215),
.B2(n_191),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_294),
.A2(n_154),
.B1(n_184),
.B2(n_191),
.Y(n_358)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_362),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_237),
.A2(n_148),
.B1(n_166),
.B2(n_164),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_366),
.B(n_382),
.Y(n_417)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_317),
.Y(n_367)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_332),
.Y(n_369)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_322),
.A2(n_286),
.B(n_242),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_370),
.A2(n_401),
.B(n_411),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_322),
.A2(n_233),
.B1(n_258),
.B2(n_184),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_372),
.A2(n_377),
.B1(n_378),
.B2(n_396),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_232),
.C(n_234),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_373),
.B(n_381),
.C(n_386),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_318),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_374),
.B(n_404),
.Y(n_415)
);

OAI21xp33_ASAP7_75t_SL g436 ( 
.A1(n_375),
.A2(n_319),
.B(n_331),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_312),
.A2(n_132),
.B1(n_154),
.B2(n_176),
.Y(n_377)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_329),
.Y(n_379)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_379),
.Y(n_424)
);

OAI22xp33_ASAP7_75t_SL g380 ( 
.A1(n_327),
.A2(n_227),
.B1(n_264),
.B2(n_238),
.Y(n_380)
);

AOI22xp33_ASAP7_75t_L g439 ( 
.A1(n_380),
.A2(n_406),
.B1(n_413),
.B2(n_355),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_262),
.C(n_244),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_327),
.B(n_267),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_316),
.A2(n_284),
.B1(n_249),
.B2(n_273),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_383),
.A2(n_385),
.B1(n_391),
.B2(n_355),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_364),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_393),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_316),
.A2(n_280),
.B1(n_299),
.B2(n_239),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_353),
.B(n_240),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_387),
.A2(n_390),
.B(n_394),
.Y(n_430)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_329),
.Y(n_388)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_388),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_335),
.B(n_303),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_389),
.B(n_397),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g390 ( 
.A(n_362),
.B(n_300),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_315),
.B(n_266),
.C(n_275),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_402),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_281),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_321),
.A2(n_328),
.B(n_349),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_338),
.B(n_287),
.C(n_236),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_395),
.B(n_330),
.C(n_323),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_349),
.A2(n_308),
.B1(n_335),
.B2(n_333),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_326),
.B(n_354),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_320),
.B(n_269),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_400),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_333),
.A2(n_247),
.B(n_235),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_357),
.C(n_309),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_317),
.Y(n_403)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_403),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_345),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_350),
.B(n_254),
.C(n_272),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_405),
.B(n_339),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_347),
.A2(n_132),
.B1(n_278),
.B2(n_270),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_311),
.Y(n_407)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_407),
.Y(n_431)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_311),
.Y(n_408)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_408),
.Y(n_437)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_346),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_410),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_336),
.A2(n_2),
.B(n_3),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_412),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_337),
.A2(n_164),
.B1(n_4),
.B2(n_5),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_371),
.B(n_394),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_416),
.B(n_427),
.C(n_438),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_366),
.A2(n_342),
.B1(n_324),
.B2(n_306),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_420),
.A2(n_441),
.B1(n_445),
.B2(n_368),
.Y(n_455)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_372),
.A2(n_306),
.B1(n_330),
.B2(n_348),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_423),
.A2(n_439),
.B1(n_444),
.B2(n_447),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_384),
.B(n_359),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_426),
.B(n_376),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_371),
.B(n_358),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_428),
.B(n_448),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_313),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_432),
.B(n_434),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_381),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_410),
.Y(n_435)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_435),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_440),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_386),
.B(n_307),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_411),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_378),
.A2(n_336),
.B1(n_359),
.B2(n_344),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_399),
.A2(n_341),
.B1(n_344),
.B2(n_334),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_446),
.B(n_392),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_367),
.A2(n_341),
.B1(n_334),
.B2(n_343),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_375),
.B(n_307),
.Y(n_448)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_407),
.Y(n_452)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_452),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_SL g506 ( 
.A(n_454),
.B(n_438),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_455),
.A2(n_459),
.B1(n_427),
.B2(n_446),
.Y(n_500)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_430),
.A2(n_387),
.B(n_401),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_456),
.A2(n_462),
.B(n_473),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_442),
.Y(n_458)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_458),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_420),
.A2(n_396),
.B1(n_390),
.B2(n_403),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_450),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_460),
.B(n_465),
.Y(n_491)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_431),
.Y(n_461)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_461),
.Y(n_492)
);

A2O1A1O1Ixp25_ASAP7_75t_L g462 ( 
.A1(n_417),
.A2(n_375),
.B(n_382),
.C(n_400),
.D(n_393),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_430),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_466),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_313),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_467),
.B(n_468),
.Y(n_511)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_419),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_426),
.B(n_422),
.Y(n_469)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_469),
.Y(n_504)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_470),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_416),
.B(n_373),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_471),
.B(n_482),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_390),
.B(n_369),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_443),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_474),
.B(n_483),
.Y(n_514)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_437),
.Y(n_476)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_422),
.B(n_405),
.Y(n_478)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_478),
.Y(n_516)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_417),
.B(n_400),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_484),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_395),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_414),
.B(n_374),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_453),
.B(n_319),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_414),
.B(n_408),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_486),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_421),
.B(n_433),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_437),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_490),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_421),
.B(n_390),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_488),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_429),
.A2(n_385),
.B1(n_383),
.B2(n_377),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_489),
.A2(n_455),
.B1(n_477),
.B2(n_441),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_450),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_425),
.C(n_451),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_495),
.B(n_496),
.C(n_508),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_475),
.B(n_454),
.C(n_471),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_459),
.A2(n_429),
.B1(n_443),
.B2(n_418),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_497),
.A2(n_500),
.B1(n_513),
.B2(n_520),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_482),
.B(n_451),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_502),
.B(n_506),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_456),
.A2(n_444),
.B(n_445),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g555 ( 
.A1(n_505),
.A2(n_524),
.B(n_323),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_507),
.A2(n_466),
.B1(n_472),
.B2(n_483),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_479),
.B(n_428),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_479),
.B(n_428),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_510),
.B(n_515),
.C(n_517),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_474),
.A2(n_433),
.B1(n_452),
.B2(n_435),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_478),
.B(n_448),
.C(n_325),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_447),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_464),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_519),
.B(n_486),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_469),
.A2(n_449),
.B1(n_424),
.B2(n_442),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_463),
.B(n_325),
.C(n_339),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_525),
.C(n_472),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_488),
.A2(n_449),
.B1(n_424),
.B2(n_412),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_523),
.A2(n_470),
.B1(n_461),
.B2(n_457),
.Y(n_538)
);

AOI21x1_ASAP7_75t_SL g524 ( 
.A1(n_473),
.A2(n_424),
.B(n_398),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_467),
.B(n_309),
.C(n_305),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_490),
.Y(n_528)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_529),
.A2(n_543),
.B1(n_544),
.B2(n_545),
.Y(n_572)
);

OAI211xp5_ASAP7_75t_SL g530 ( 
.A1(n_493),
.A2(n_480),
.B(n_462),
.C(n_485),
.Y(n_530)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_530),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_521),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g568 ( 
.A(n_532),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_533),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_491),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g578 ( 
.A1(n_534),
.A2(n_536),
.B(n_539),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_504),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_521),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_537),
.B(n_552),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_538),
.A2(n_546),
.B1(n_548),
.B2(n_550),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_514),
.B(n_472),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_520),
.B(n_457),
.Y(n_540)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_540),
.Y(n_566)
);

CKINVDCx14_ASAP7_75t_R g541 ( 
.A(n_514),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_541),
.A2(n_555),
.B(n_539),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_504),
.B(n_476),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_542),
.B(n_547),
.Y(n_558)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_509),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_509),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_492),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_512),
.Y(n_546)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_511),
.Y(n_548)
);

BUFx24_ASAP7_75t_SL g549 ( 
.A(n_498),
.Y(n_549)
);

BUFx24_ASAP7_75t_SL g561 ( 
.A(n_549),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_507),
.A2(n_487),
.B1(n_489),
.B2(n_458),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_497),
.A2(n_505),
.B1(n_516),
.B2(n_503),
.Y(n_551)
);

XNOR2x1_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_513),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_511),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_523),
.B(n_379),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_554),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_493),
.A2(n_494),
.B1(n_524),
.B2(n_517),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_494),
.A2(n_412),
.B1(n_343),
.B2(n_388),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_556),
.B(n_508),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_526),
.B(n_496),
.C(n_495),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_559),
.B(n_560),
.C(n_562),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_526),
.B(n_502),
.C(n_501),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_535),
.B(n_501),
.C(n_522),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_535),
.B(n_506),
.C(n_515),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_563),
.B(n_575),
.C(n_532),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g585 ( 
.A(n_565),
.B(n_577),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g567 ( 
.A(n_531),
.B(n_510),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_SL g601 ( 
.A(n_567),
.B(n_543),
.Y(n_601)
);

XNOR2x1_ASAP7_75t_L g590 ( 
.A(n_569),
.B(n_573),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_536),
.B(n_525),
.Y(n_570)
);

NOR3xp33_ASAP7_75t_L g593 ( 
.A(n_570),
.B(n_533),
.C(n_537),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_531),
.B(n_305),
.C(n_518),
.Y(n_575)
);

FAx1_ASAP7_75t_SL g577 ( 
.A(n_530),
.B(n_518),
.CI(n_360),
.CON(n_577),
.SN(n_577)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_547),
.B(n_310),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_579),
.B(n_542),
.Y(n_583)
);

FAx1_ASAP7_75t_L g580 ( 
.A(n_554),
.B(n_348),
.CI(n_360),
.CON(n_580),
.SN(n_580)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_580),
.B(n_556),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g617 ( 
.A(n_583),
.B(n_586),
.Y(n_617)
);

OAI21xp5_ASAP7_75t_L g584 ( 
.A1(n_579),
.A2(n_528),
.B(n_551),
.Y(n_584)
);

NOR2xp67_ASAP7_75t_SL g605 ( 
.A(n_584),
.B(n_587),
.Y(n_605)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_558),
.B(n_527),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_575),
.B(n_527),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_588),
.Y(n_618)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_571),
.Y(n_589)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_589),
.Y(n_608)
);

BUFx24_ASAP7_75t_SL g591 ( 
.A(n_561),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_SL g614 ( 
.A(n_591),
.B(n_599),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_SL g592 ( 
.A1(n_571),
.A2(n_552),
.B1(n_548),
.B2(n_541),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_592),
.B(n_594),
.Y(n_602)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_593),
.Y(n_612)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_557),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_595),
.B(n_596),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g596 ( 
.A1(n_574),
.A2(n_538),
.B1(n_540),
.B2(n_553),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_572),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_600),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_576),
.A2(n_550),
.B1(n_529),
.B2(n_544),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_598),
.A2(n_580),
.B1(n_577),
.B2(n_569),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_558),
.B(n_545),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g600 ( 
.A(n_573),
.B(n_555),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_601),
.B(n_564),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_588),
.A2(n_578),
.B1(n_581),
.B2(n_568),
.Y(n_603)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_603),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g626 ( 
.A(n_604),
.B(n_365),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_559),
.C(n_560),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_606),
.B(n_609),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g607 ( 
.A1(n_585),
.A2(n_566),
.B1(n_580),
.B2(n_564),
.Y(n_607)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_607),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g611 ( 
.A(n_582),
.B(n_562),
.C(n_563),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_611),
.B(n_616),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_585),
.A2(n_577),
.B(n_546),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_SL g625 ( 
.A1(n_615),
.A2(n_331),
.B(n_356),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_587),
.B(n_583),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_612),
.B(n_586),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_620),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g620 ( 
.A(n_606),
.B(n_582),
.C(n_590),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_SL g622 ( 
.A1(n_615),
.A2(n_600),
.B(n_601),
.Y(n_622)
);

OAI21xp5_ASAP7_75t_SL g635 ( 
.A1(n_622),
.A2(n_630),
.B(n_618),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_611),
.B(n_590),
.C(n_567),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_623),
.B(n_624),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_614),
.B(n_310),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_625),
.B(n_631),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_626),
.B(n_628),
.Y(n_639)
);

AOI21xp5_ASAP7_75t_L g628 ( 
.A1(n_603),
.A2(n_356),
.B(n_365),
.Y(n_628)
);

OAI21xp5_ASAP7_75t_SL g630 ( 
.A1(n_602),
.A2(n_331),
.B(n_351),
.Y(n_630)
);

XNOR2xp5_ASAP7_75t_L g631 ( 
.A(n_617),
.B(n_616),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_631),
.B(n_610),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_633),
.B(n_635),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_629),
.B(n_608),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_636),
.A2(n_626),
.B(n_361),
.Y(n_647)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_622),
.B(n_617),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_637),
.B(n_641),
.Y(n_649)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_627),
.A2(n_618),
.B(n_613),
.C(n_604),
.Y(n_638)
);

A2O1A1Ixp33_ASAP7_75t_SL g646 ( 
.A1(n_638),
.A2(n_625),
.B(n_607),
.C(n_628),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_620),
.B(n_605),
.Y(n_641)
);

MAJIxp5_ASAP7_75t_L g643 ( 
.A(n_640),
.B(n_621),
.C(n_632),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_643),
.B(n_647),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_634),
.A2(n_638),
.B(n_637),
.Y(n_644)
);

AO21x1_ASAP7_75t_L g652 ( 
.A1(n_644),
.A2(n_646),
.B(n_639),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_SL g645 ( 
.A(n_642),
.B(n_623),
.Y(n_645)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_645),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_649),
.B(n_639),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_651),
.B(n_652),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g654 ( 
.A(n_653),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g656 ( 
.A1(n_654),
.A2(n_648),
.B(n_650),
.Y(n_656)
);

AO21x1_ASAP7_75t_L g657 ( 
.A1(n_656),
.A2(n_655),
.B(n_361),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_657),
.B(n_5),
.C(n_654),
.Y(n_658)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_658),
.B(n_5),
.Y(n_659)
);


endmodule