module fake_jpeg_3743_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx4f_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_33),
.Y(n_49)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_37),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_38),
.B(n_15),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_39),
.A2(n_17),
.B(n_25),
.C(n_24),
.Y(n_42)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_28),
.B1(n_15),
.B2(n_26),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_42),
.A2(n_60),
.B(n_20),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_28),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_47),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_45),
.Y(n_71)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_31),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_50),
.Y(n_87)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_22),
.B1(n_15),
.B2(n_17),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_52),
.A2(n_26),
.B1(n_39),
.B2(n_34),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_54),
.A2(n_59),
.B1(n_39),
.B2(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_34),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_63),
.A2(n_37),
.B1(n_41),
.B2(n_19),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_47),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_78),
.B1(n_83),
.B2(n_53),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_67),
.B(n_55),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_39),
.B(n_35),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_81),
.B1(n_85),
.B2(n_47),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_74),
.B1(n_51),
.B2(n_56),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_44),
.B1(n_43),
.B2(n_62),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_49),
.B(n_36),
.C(n_35),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_83),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_33),
.B1(n_32),
.B2(n_37),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_42),
.A2(n_34),
.B1(n_41),
.B2(n_32),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_36),
.B1(n_33),
.B2(n_37),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_19),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_88),
.A2(n_96),
.B1(n_83),
.B2(n_78),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_89),
.A2(n_95),
.B1(n_100),
.B2(n_104),
.Y(n_111)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_92),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_91),
.B(n_102),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_68),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_93),
.B(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_67),
.A2(n_79),
.B1(n_69),
.B2(n_85),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_78),
.A2(n_57),
.B1(n_61),
.B2(n_37),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_97),
.B(n_36),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_106),
.B(n_87),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_101),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_67),
.A2(n_79),
.B1(n_84),
.B2(n_81),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_72),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_49),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_75),
.A2(n_80),
.B1(n_78),
.B2(n_73),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_77),
.Y(n_107)
);

INVxp33_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_48),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_64),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_82),
.Y(n_121)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_115),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_122),
.B1(n_134),
.B2(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_75),
.B1(n_78),
.B2(n_83),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_88),
.B1(n_41),
.B2(n_53),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_98),
.A2(n_83),
.B(n_77),
.C(n_64),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_118),
.A2(n_106),
.B(n_103),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_70),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_70),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_123),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_96),
.Y(n_140)
);

AO22x1_ASAP7_75t_SL g122 ( 
.A1(n_97),
.A2(n_57),
.B1(n_36),
.B2(n_53),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_93),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_124),
.B(n_129),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_126),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_91),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_94),
.B(n_82),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_99),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_71),
.C(n_87),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_122),
.C(n_116),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_137),
.A2(n_161),
.B1(n_108),
.B2(n_105),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_141),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_95),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_143),
.A2(n_118),
.B(n_122),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_146),
.B(n_148),
.Y(n_176)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_149),
.B(n_157),
.C(n_132),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_113),
.B1(n_134),
.B2(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_153),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_152),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_123),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_136),
.B(n_107),
.Y(n_155)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_155),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_71),
.Y(n_156)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_156),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_105),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_129),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_114),
.B(n_48),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_160),
.A2(n_70),
.B(n_134),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_41),
.B1(n_90),
.B2(n_108),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_117),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_162),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_164),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_122),
.B(n_127),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_166),
.A2(n_170),
.B1(n_175),
.B2(n_179),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g199 ( 
.A1(n_167),
.A2(n_169),
.B(n_186),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_111),
.B(n_119),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_150),
.A2(n_111),
.B1(n_117),
.B2(n_105),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_147),
.A2(n_149),
.B1(n_140),
.B2(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_162),
.Y(n_190)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_142),
.Y(n_178)
);

INVxp33_ASAP7_75t_SL g194 ( 
.A(n_178),
.Y(n_194)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_45),
.B1(n_58),
.B2(n_46),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_181),
.C(n_157),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_45),
.C(n_58),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_184),
.A2(n_146),
.B1(n_155),
.B2(n_151),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_143),
.A2(n_160),
.B(n_153),
.Y(n_186)
);

NAND2xp33_ASAP7_75t_SL g187 ( 
.A(n_138),
.B(n_36),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_139),
.Y(n_208)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_137),
.B(n_36),
.CI(n_58),
.CON(n_188),
.SN(n_188)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_188),
.B(n_144),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_152),
.B(n_130),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_189),
.B(n_139),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_193),
.A2(n_195),
.B1(n_203),
.B2(n_212),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_145),
.B1(n_156),
.B2(n_137),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_157),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_197),
.B(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_198),
.B(n_200),
.Y(n_229)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_201),
.A2(n_174),
.B(n_177),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_171),
.A2(n_138),
.B1(n_144),
.B2(n_148),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_209),
.C(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_182),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_205),
.B(n_207),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_183),
.Y(n_206)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_206),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_166),
.A2(n_161),
.B1(n_154),
.B2(n_159),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_165),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_45),
.C(n_36),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_182),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_210),
.B(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_175),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_76),
.B1(n_131),
.B2(n_66),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_165),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_192),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_169),
.B(n_46),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_226),
.C(n_228),
.Y(n_242)
);

NOR2xp67_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_179),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_233),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_221),
.B(n_224),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_197),
.B(n_186),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_164),
.C(n_172),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_170),
.B1(n_183),
.B2(n_185),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_227),
.A2(n_199),
.B1(n_174),
.B2(n_208),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_163),
.C(n_188),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_230),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_188),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_235),
.C(n_168),
.Y(n_246)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_232),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_187),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_173),
.Y(n_235)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_236),
.Y(n_244)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_238),
.B(n_249),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_234),
.A2(n_195),
.B1(n_191),
.B2(n_203),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_243),
.B1(n_29),
.B2(n_23),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_142),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_199),
.B1(n_207),
.B2(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_245),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_252),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_194),
.C(n_168),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_253),
.C(n_254),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_178),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_23),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_131),
.B1(n_66),
.B2(n_19),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_251),
.A2(n_256),
.B1(n_217),
.B2(n_225),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_46),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_131),
.C(n_16),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_23),
.C(n_21),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_224),
.B(n_23),
.C(n_21),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_231),
.C(n_233),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_223),
.A2(n_29),
.B1(n_19),
.B2(n_21),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_257),
.B(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_229),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_254),
.Y(n_275)
);

AO221x1_ASAP7_75t_L g262 ( 
.A1(n_247),
.A2(n_223),
.B1(n_235),
.B2(n_232),
.C(n_221),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_268),
.B(n_269),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_263),
.B(n_272),
.C(n_1),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_29),
.B1(n_16),
.B2(n_14),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_266),
.A2(n_241),
.B1(n_250),
.B2(n_29),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_250),
.B(n_20),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_248),
.A2(n_20),
.B(n_18),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_0),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_271),
.A2(n_18),
.B(n_255),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_21),
.C(n_16),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_275),
.A2(n_281),
.B(n_282),
.Y(n_293)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

AOI322xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_261),
.A3(n_270),
.B1(n_272),
.B2(n_11),
.C1(n_6),
.C2(n_7),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_283),
.B(n_4),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_265),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_1),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_266),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_285),
.A2(n_287),
.B(n_3),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_264),
.B(n_1),
.Y(n_287)
);

AO21x1_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_267),
.B(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_294),
.Y(n_299)
);

AOI31xp67_ASAP7_75t_L g300 ( 
.A1(n_290),
.A2(n_283),
.A3(n_282),
.B(n_278),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_286),
.A2(n_261),
.B1(n_270),
.B2(n_4),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_292),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_296),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_298),
.C(n_7),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_5),
.B(n_7),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_303),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_289),
.A2(n_285),
.B1(n_280),
.B2(n_9),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_305),
.B(n_295),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_8),
.C(n_9),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_306),
.A2(n_304),
.B(n_301),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_299),
.A2(n_288),
.B1(n_292),
.B2(n_293),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_311),
.C(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

MAJx2_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_302),
.C(n_9),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_312),
.B(n_10),
.Y(n_316)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_9),
.B(n_10),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_315),
.Y(n_318)
);


endmodule