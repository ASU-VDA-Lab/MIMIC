module fake_jpeg_28828_n_157 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_157);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_157;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_46),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_15),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_23),
.B(n_20),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_3),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_1),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_74),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_2),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_75),
.B(n_77),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_2),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_66),
.B1(n_65),
.B2(n_67),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_81),
.A2(n_90),
.B1(n_54),
.B2(n_55),
.Y(n_105)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_62),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_67),
.B(n_59),
.Y(n_86)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_86),
.A2(n_65),
.B(n_49),
.C(n_59),
.D(n_64),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_87),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_62),
.B1(n_53),
.B2(n_48),
.Y(n_90)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_70),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_91),
.B(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_103),
.B(n_17),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_96),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_99),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_91),
.B(n_4),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_78),
.B(n_63),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_100),
.B(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_106),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_4),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_118)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_50),
.A3(n_27),
.B1(n_31),
.B2(n_47),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_5),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_87),
.B(n_6),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_80),
.C(n_83),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_116),
.C(n_117),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_26),
.C(n_44),
.Y(n_116)
);

AOI322xp5_ASAP7_75t_SL g117 ( 
.A1(n_103),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_12),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_42),
.B1(n_25),
.B2(n_32),
.Y(n_140)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_33),
.C(n_13),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_121),
.B(n_127),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_12),
.Y(n_122)
);

AOI21x1_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_125),
.B(n_128),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_123),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_45),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_18),
.C(n_21),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_96),
.B(n_22),
.Y(n_128)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_115),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_140),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_111),
.B1(n_119),
.B2(n_130),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_141),
.B(n_131),
.Y(n_147)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_142),
.B(n_143),
.Y(n_146)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_133),
.B(n_127),
.C(n_116),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_144),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_147),
.A2(n_141),
.B1(n_137),
.B2(n_132),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_150),
.B(n_151),
.Y(n_152)
);

OAI322xp33_ASAP7_75t_L g151 ( 
.A1(n_145),
.A2(n_135),
.A3(n_133),
.B1(n_136),
.B2(n_124),
.C1(n_117),
.C2(n_137),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_150),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_153),
.B(n_146),
.Y(n_154)
);

OAI221xp5_ASAP7_75t_L g155 ( 
.A1(n_154),
.A2(n_149),
.B1(n_148),
.B2(n_121),
.C(n_39),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_24),
.Y(n_156)
);

AOI221xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.C(n_41),
.Y(n_157)
);


endmodule