module fake_jpeg_14526_n_464 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_464);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_464;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_SL g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_4),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVxp33_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_33),
.B(n_9),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_49),
.B(n_50),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_9),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_9),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_59),
.B(n_73),
.Y(n_147)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_60),
.Y(n_145)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_63),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_67),
.Y(n_122)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_68),
.Y(n_139)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_70),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_7),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_74),
.Y(n_134)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_15),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_88),
.Y(n_116)
);

BUFx12f_ASAP7_75t_SL g77 ( 
.A(n_19),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_77),
.B(n_85),
.Y(n_99)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_78),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_16),
.B(n_7),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_90),
.Y(n_100)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_38),
.Y(n_83)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_87),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_23),
.Y(n_90)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_17),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_92),
.B(n_94),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_7),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_23),
.Y(n_95)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_95),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_96),
.Y(n_148)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_38),
.B1(n_45),
.B2(n_40),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_106),
.A2(n_118),
.B1(n_27),
.B2(n_45),
.Y(n_179)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_73),
.A2(n_18),
.B(n_37),
.C(n_32),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_117),
.B(n_35),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_95),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_59),
.A2(n_48),
.B(n_37),
.C(n_32),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_137),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_20),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_70),
.B(n_48),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_27),
.Y(n_186)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_149),
.Y(n_176)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_151),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVxp67_ASAP7_75t_SL g229 ( 
.A(n_153),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_154),
.B(n_158),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

AND2x2_ASAP7_75t_SL g158 ( 
.A(n_101),
.B(n_0),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_69),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_201),
.C(n_17),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_99),
.A2(n_40),
.B1(n_26),
.B2(n_78),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_161),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_163),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_164),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_103),
.B(n_24),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_117),
.B(n_127),
.Y(n_204)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_167),
.Y(n_215)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g235 ( 
.A(n_168),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_116),
.A2(n_80),
.B1(n_82),
.B2(n_72),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_172),
.B1(n_174),
.B2(n_179),
.Y(n_210)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_116),
.A2(n_71),
.B1(n_67),
.B2(n_65),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_118),
.A2(n_64),
.B1(n_58),
.B2(n_57),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_182),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_177),
.Y(n_240)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_178),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_56),
.B1(n_54),
.B2(n_51),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_181),
.A2(n_135),
.B1(n_109),
.B2(n_113),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_129),
.Y(n_182)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_111),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_183),
.Y(n_232)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_108),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_190),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_187),
.B(n_188),
.Y(n_236)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_189),
.B(n_192),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_145),
.A2(n_26),
.B1(n_47),
.B2(n_39),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g192 ( 
.A(n_105),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_193),
.B(n_194),
.Y(n_238)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_102),
.A2(n_47),
.B1(n_46),
.B2(n_39),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_105),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_110),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_197),
.B(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_200),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_144),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_147),
.B(n_24),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_204),
.B(n_212),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_158),
.B(n_132),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_206),
.B(n_214),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_208),
.B(n_11),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_185),
.A2(n_135),
.B1(n_115),
.B2(n_110),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_234),
.B1(n_189),
.B2(n_107),
.Y(n_248)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_154),
.A2(n_183),
.B(n_187),
.C(n_177),
.Y(n_212)
);

AOI32xp33_ASAP7_75t_L g213 ( 
.A1(n_201),
.A2(n_47),
.A3(n_22),
.B1(n_30),
.B2(n_35),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_213),
.A2(n_10),
.B(n_1),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_158),
.B(n_104),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_154),
.B(n_104),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_220),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_242),
.B1(n_192),
.B2(n_157),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_160),
.B(n_115),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_160),
.A2(n_139),
.B(n_140),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_15),
.B(n_1),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_169),
.B(n_47),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_241),
.C(n_196),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_165),
.A2(n_24),
.B(n_46),
.C(n_30),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_231),
.B(n_237),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_172),
.A2(n_113),
.B1(n_109),
.B2(n_121),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_165),
.B(n_121),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_165),
.B(n_139),
.C(n_22),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_174),
.A2(n_107),
.B1(n_20),
.B2(n_2),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_152),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_246),
.B(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_226),
.Y(n_247)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_247),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_248),
.A2(n_251),
.B1(n_256),
.B2(n_259),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_272),
.Y(n_291)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_235),
.Y(n_250)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_250),
.Y(n_296)
);

AO21x2_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_204),
.B(n_203),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_252),
.A2(n_254),
.B1(n_261),
.B2(n_263),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_210),
.A2(n_170),
.B1(n_171),
.B2(n_162),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_SL g255 ( 
.A1(n_218),
.A2(n_155),
.B(n_163),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_230),
.A2(n_180),
.B1(n_166),
.B2(n_151),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_208),
.B(n_159),
.C(n_176),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_274),
.C(n_282),
.Y(n_297)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_234),
.A2(n_193),
.B1(n_197),
.B2(n_168),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_210),
.A2(n_156),
.B1(n_199),
.B2(n_167),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_260),
.A2(n_278),
.B1(n_280),
.B2(n_232),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_206),
.A2(n_153),
.B1(n_184),
.B2(n_175),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_202),
.Y(n_262)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_262),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_219),
.A2(n_164),
.B1(n_0),
.B2(n_3),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_267),
.A2(n_212),
.B(n_223),
.Y(n_293)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_202),
.Y(n_268)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_203),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_269),
.B(n_270),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_217),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_224),
.B(n_10),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_271),
.B(n_233),
.Y(n_314)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_243),
.Y(n_273)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_216),
.B(n_11),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_243),
.Y(n_275)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_275),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_242),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_276),
.A2(n_279),
.B1(n_232),
.B2(n_240),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_238),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_277),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_209),
.A2(n_4),
.B1(n_6),
.B2(n_12),
.Y(n_278)
);

OAI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_240),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_216),
.A2(n_13),
.B1(n_14),
.B2(n_0),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_239),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_281),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_0),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_284),
.A2(n_273),
.B1(n_280),
.B2(n_235),
.Y(n_334)
);

BUFx24_ASAP7_75t_SL g285 ( 
.A(n_272),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_286),
.B(n_287),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_214),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_220),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_290),
.B(n_294),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_292),
.A2(n_316),
.B1(n_248),
.B2(n_260),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_265),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_253),
.B(n_231),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_241),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_301),
.A2(n_267),
.B(n_256),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_261),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_312),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_251),
.A2(n_225),
.B1(n_213),
.B2(n_233),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_308),
.A2(n_293),
.B1(n_306),
.B2(n_315),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_211),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_249),
.B(n_211),
.C(n_236),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_257),
.C(n_253),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_254),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_314),
.B(n_205),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_253),
.A2(n_235),
.B1(n_222),
.B2(n_227),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_317),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_321),
.C(n_335),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_264),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_308),
.A2(n_252),
.B1(n_264),
.B2(n_263),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_323),
.A2(n_325),
.B1(n_330),
.B2(n_334),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_326),
.A2(n_340),
.B1(n_343),
.B2(n_346),
.Y(n_349)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_309),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_327),
.B(n_336),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_286),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_332),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_276),
.B1(n_266),
.B2(n_275),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_287),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_316),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_291),
.B(n_282),
.C(n_274),
.Y(n_335)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_290),
.A2(n_278),
.B1(n_222),
.B2(n_227),
.Y(n_338)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_301),
.A2(n_215),
.B1(n_243),
.B2(n_205),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_244),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_311),
.C(n_297),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_342),
.B(n_345),
.Y(n_367)
);

AOI22x1_ASAP7_75t_L g343 ( 
.A1(n_294),
.A2(n_215),
.B1(n_221),
.B2(n_207),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_283),
.Y(n_344)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_344),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_298),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_SL g346 ( 
.A1(n_302),
.A2(n_229),
.B(n_215),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_300),
.B(n_244),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_347),
.B(n_289),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_359),
.C(n_363),
.Y(n_374)
);

OR2x2_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_310),
.Y(n_352)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_344),
.Y(n_353)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_353),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_355),
.B(n_318),
.Y(n_378)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_357),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_341),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_340),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_360),
.B(n_323),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_333),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_362),
.B(n_368),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_319),
.B(n_301),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_335),
.B(n_304),
.C(n_303),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_371),
.C(n_372),
.Y(n_384)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_337),
.Y(n_366)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_366),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_320),
.B(n_289),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_332),
.A2(n_312),
.B1(n_303),
.B2(n_304),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_369),
.A2(n_339),
.B1(n_288),
.B2(n_330),
.Y(n_394)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_322),
.Y(n_370)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_370),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_345),
.C(n_329),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_318),
.B(n_314),
.Y(n_372)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_373),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_361),
.A2(n_331),
.B1(n_324),
.B2(n_328),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_376),
.A2(n_389),
.B1(n_288),
.B2(n_292),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_367),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_377),
.B(n_388),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_378),
.B(n_365),
.Y(n_409)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_380),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_350),
.B(n_325),
.Y(n_381)
);

MAJx2_ASAP7_75t_L g408 ( 
.A(n_381),
.B(n_365),
.C(n_352),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_367),
.A2(n_328),
.B(n_343),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_382),
.B(n_349),
.Y(n_405)
);

FAx1_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_338),
.CI(n_343),
.CON(n_387),
.SN(n_387)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_387),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_358),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_360),
.A2(n_339),
.B1(n_284),
.B2(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_353),
.Y(n_391)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_391),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_394),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_299),
.C(n_283),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_359),
.C(n_364),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_398),
.B(n_404),
.C(n_406),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_395),
.B(n_351),
.C(n_363),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_399),
.B(n_400),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g400 ( 
.A(n_385),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_374),
.B(n_355),
.C(n_358),
.Y(n_404)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_405),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_374),
.B(n_369),
.C(n_372),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_310),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g423 ( 
.A(n_407),
.B(n_393),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_SL g414 ( 
.A(n_408),
.B(n_409),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_384),
.B(n_349),
.C(n_348),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_410),
.B(n_412),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_411),
.A2(n_394),
.B1(n_403),
.B2(n_401),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_295),
.C(n_357),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_401),
.A2(n_375),
.B(n_382),
.Y(n_416)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_416),
.B(n_387),
.C(n_409),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_417),
.A2(n_423),
.B1(n_426),
.B2(n_380),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_397),
.A2(n_386),
.B1(n_389),
.B2(n_376),
.Y(n_418)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_418),
.Y(n_431)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_420),
.B(n_421),
.Y(n_432)
);

BUFx24_ASAP7_75t_SL g421 ( 
.A(n_396),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_391),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_424),
.B(n_425),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_384),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_408),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_427),
.A2(n_354),
.B1(n_338),
.B2(n_299),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_424),
.B(n_422),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_429),
.B(n_433),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_417),
.B(n_406),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_430),
.B(n_435),
.C(n_436),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_413),
.A2(n_387),
.B1(n_383),
.B2(n_390),
.Y(n_433)
);

AO21x1_ASAP7_75t_L g439 ( 
.A1(n_434),
.A2(n_416),
.B(n_414),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_414),
.B(n_398),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_419),
.B(n_399),
.C(n_378),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_436),
.B(n_437),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_419),
.B(n_379),
.C(n_392),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_379),
.C(n_392),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_438),
.B(n_307),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_439),
.A2(n_446),
.B(n_447),
.Y(n_452)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_441),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_442),
.B(n_443),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_438),
.B(n_307),
.Y(n_444)
);

AOI21xp33_ASAP7_75t_L g449 ( 
.A1(n_444),
.A2(n_431),
.B(n_434),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_305),
.C(n_313),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_429),
.A2(n_305),
.B(n_296),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_440),
.B(n_437),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_448),
.B(n_453),
.Y(n_457)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_449),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_445),
.A2(n_428),
.B(n_435),
.Y(n_453)
);

INVx6_ASAP7_75t_L g455 ( 
.A(n_450),
.Y(n_455)
);

O2A1O1Ixp33_ASAP7_75t_SL g459 ( 
.A1(n_455),
.A2(n_456),
.B(n_452),
.C(n_444),
.Y(n_459)
);

NOR2x1_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_439),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_457),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_458),
.B(n_459),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g461 ( 
.A(n_460),
.B(n_454),
.C(n_432),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_461),
.B(n_456),
.C(n_296),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_221),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_463),
.B(n_207),
.Y(n_464)
);


endmodule