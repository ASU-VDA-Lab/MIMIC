module real_jpeg_10275_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx24_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_18),
.B1(n_19),
.B2(n_24),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_1),
.A2(n_24),
.B1(n_38),
.B2(n_39),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g68 ( 
.A(n_2),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_5),
.A2(n_18),
.B(n_51),
.C(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_5),
.B(n_18),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_5),
.A2(n_8),
.B(n_39),
.Y(n_88)
);

BUFx6f_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_8),
.A2(n_17),
.B(n_26),
.C(n_35),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_8),
.A2(n_29),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_8),
.A2(n_18),
.B1(n_19),
.B2(n_29),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_8),
.B(n_15),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_81),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_80),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_57),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_13),
.B(n_57),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_32),
.C(n_47),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_14),
.A2(n_47),
.B1(n_89),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_14),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_23),
.B(n_27),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_15),
.A2(n_23),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

A2O1A1Ixp33_ASAP7_75t_L g30 ( 
.A1(n_16),
.A2(n_17),
.B(n_26),
.C(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_19),
.B2(n_22),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_26),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g35 ( 
.A1(n_18),
.A2(n_22),
.B(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_19),
.A2(n_29),
.B(n_52),
.C(n_88),
.Y(n_87)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_29),
.B(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_29),
.B(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_32),
.A2(n_33),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_42),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_37),
.B(n_44),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_37),
.A2(n_44),
.B1(n_45),
.B2(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_38),
.B(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_70),
.B(n_72),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_47),
.A2(n_86),
.B1(n_87),
.B2(n_89),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_47),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_47),
.B(n_87),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_50),
.B(n_53),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_49),
.A2(n_51),
.B1(n_54),
.B2(n_55),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_75),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_62),
.B1(n_63),
.B2(n_74),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_69),
.B2(n_73),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_69),
.B(n_85),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_76),
.A2(n_78),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_96),
.C(n_104),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_77),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_108),
.B(n_114),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_99),
.B(n_107),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_90),
.B(n_98),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_94),
.B(n_97),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_96),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_95),
.B(n_96),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_96),
.A2(n_102),
.B1(n_103),
.B2(n_106),
.Y(n_101)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_100),
.B(n_101),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_109),
.B(n_110),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);


endmodule