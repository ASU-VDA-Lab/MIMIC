module fake_jpeg_21888_n_179 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_SL g16 ( 
.A(n_4),
.Y(n_16)
);

INVx11_ASAP7_75t_SL g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_22),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_35),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_17),
.B1(n_25),
.B2(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_15),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_48),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_18),
.B(n_30),
.C(n_27),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_46),
.B(n_49),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_59),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_31),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_26),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_32),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_19),
.B1(n_40),
.B2(n_2),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_27),
.B(n_30),
.C(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_58),
.B(n_48),
.Y(n_76)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_57),
.A2(n_24),
.B1(n_39),
.B2(n_34),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_60),
.Y(n_90)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_65),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_59),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_34),
.B1(n_38),
.B2(n_26),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_64),
.A2(n_69),
.B1(n_79),
.B2(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_28),
.B1(n_19),
.B2(n_38),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_53),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_50),
.B1(n_55),
.B2(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_15),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_78),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_76),
.Y(n_97)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_55),
.A2(n_40),
.B1(n_1),
.B2(n_3),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_0),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_1),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_83),
.A2(n_88),
.B1(n_66),
.B2(n_77),
.Y(n_115)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_62),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_51),
.C(n_53),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_88),
.C(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_8),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_94),
.B(n_5),
.Y(n_114)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_101),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_72),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_73),
.B(n_71),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_106),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_83),
.A2(n_66),
.B1(n_69),
.B2(n_73),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_103),
.B(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_87),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_82),
.B(n_72),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_67),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_74),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_111),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_101),
.B1(n_90),
.B2(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_119),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_95),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_77),
.Y(n_118)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_97),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_130),
.B(n_131),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_104),
.B(n_85),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_117),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_107),
.B1(n_105),
.B2(n_96),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_85),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_100),
.B(n_98),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_102),
.C(n_119),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_142),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_103),
.B1(n_112),
.B2(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_147),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_106),
.C(n_96),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_124),
.C(n_123),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_100),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_145),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_146),
.A2(n_5),
.B(n_6),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_145),
.A2(n_125),
.B1(n_120),
.B2(n_127),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_146),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_141),
.C(n_136),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_122),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_156),
.A2(n_139),
.B(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_143),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_151),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_160),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_162),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_142),
.C(n_11),
.Y(n_162)
);

NAND3xp33_ASAP7_75t_SL g163 ( 
.A(n_148),
.B(n_14),
.C(n_7),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_163),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_166),
.Y(n_169)
);

NOR4xp25_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_161),
.C(n_158),
.D(n_154),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_171),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_153),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_167),
.B(n_154),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_167),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g176 ( 
.A1(n_174),
.A2(n_7),
.B(n_13),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_169),
.B(n_168),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_173),
.C(n_13),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_177),
.Y(n_179)
);


endmodule