module fake_jpeg_9798_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_38),
.B(n_34),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_49),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_41),
.B(n_21),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_22),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_24),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_28),
.B1(n_22),
.B2(n_29),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_53),
.A2(n_40),
.B1(n_44),
.B2(n_30),
.Y(n_101)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_62),
.Y(n_105)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_63),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_22),
.B1(n_29),
.B2(n_24),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_58),
.A2(n_71),
.B1(n_75),
.B2(n_49),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_64),
.B(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_20),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_68),
.B(n_44),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_70),
.B(n_49),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_43),
.A2(n_29),
.B1(n_28),
.B2(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_25),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

AO22x2_ASAP7_75t_L g75 ( 
.A1(n_36),
.A2(n_32),
.B1(n_35),
.B2(n_17),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_77),
.B(n_21),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_56),
.A2(n_62),
.B1(n_75),
.B2(n_28),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_81),
.B(n_86),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_92),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_85),
.A2(n_87),
.B1(n_91),
.B2(n_101),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_46),
.B1(n_44),
.B2(n_41),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_63),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_89),
.B(n_90),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_41),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_100),
.B(n_16),
.Y(n_141)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_109),
.B1(n_112),
.B2(n_116),
.Y(n_130)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_69),
.B(n_40),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_78),
.C(n_31),
.Y(n_129)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_61),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_113),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

HB1xp67_ASAP7_75t_SL g142 ( 
.A(n_114),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_55),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_120),
.B(n_123),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_82),
.B(n_52),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_125),
.B(n_136),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_57),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_128),
.B(n_141),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_129),
.B(n_140),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_67),
.B1(n_68),
.B2(n_65),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_99),
.B1(n_97),
.B2(n_112),
.Y(n_154)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_85),
.A2(n_45),
.B1(n_42),
.B2(n_39),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_134),
.A2(n_146),
.B1(n_93),
.B2(n_109),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_107),
.A2(n_31),
.A3(n_30),
.B1(n_26),
.B2(n_16),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_80),
.A2(n_78),
.B1(n_45),
.B2(n_42),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_107),
.B(n_1),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_148),
.A2(n_129),
.B(n_128),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_121),
.B(n_84),
.Y(n_150)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_150),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_122),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_151),
.B(n_160),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_105),
.C(n_118),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_159),
.C(n_163),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_83),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_179),
.B1(n_133),
.B2(n_149),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_143),
.A2(n_114),
.B1(n_89),
.B2(n_103),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_161),
.B1(n_167),
.B2(n_169),
.Y(n_191)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_142),
.A2(n_111),
.B(n_32),
.C(n_39),
.D(n_42),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_156),
.B(n_17),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_83),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_130),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_170),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_119),
.C(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_124),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_143),
.A2(n_97),
.B1(n_93),
.B2(n_102),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_162),
.A2(n_138),
.B(n_17),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_42),
.C(n_45),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_39),
.C(n_59),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_163),
.C(n_154),
.Y(n_199)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_166),
.B(n_174),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_134),
.A2(n_26),
.B1(n_18),
.B2(n_19),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_34),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_172),
.B(n_176),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_34),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_175),
.Y(n_187)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_127),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_34),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_1),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_181),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_139),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_178),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_134),
.A2(n_98),
.B1(n_115),
.B2(n_18),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_141),
.B(n_1),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_135),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_182),
.B(n_183),
.Y(n_194)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_1),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_145),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_146),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_186),
.B(n_199),
.C(n_205),
.Y(n_222)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_216),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

MAJx2_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_137),
.C(n_145),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_198),
.B(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_211),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_158),
.A2(n_138),
.B1(n_133),
.B2(n_149),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_215),
.B1(n_4),
.B2(n_5),
.Y(n_243)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_156),
.B(n_147),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_212),
.B(n_214),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_165),
.B(n_147),
.C(n_104),
.Y(n_205)
);

XNOR2x1_ASAP7_75t_SL g206 ( 
.A(n_165),
.B(n_17),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_207),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_183),
.A2(n_124),
.B1(n_19),
.B2(n_27),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_208),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_88),
.C(n_96),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_213),
.C(n_182),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_176),
.A2(n_33),
.B1(n_27),
.B2(n_106),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_164),
.B(n_2),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_131),
.C(n_139),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_168),
.A2(n_17),
.B(n_33),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_169),
.A2(n_17),
.B1(n_131),
.B2(n_11),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_168),
.B1(n_173),
.B2(n_180),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_175),
.A2(n_2),
.B(n_3),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_3),
.B(n_4),
.Y(n_237)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_233),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_171),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_221),
.C(n_226),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_177),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_184),
.C(n_181),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_227),
.B(n_232),
.C(n_236),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_187),
.Y(n_229)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_202),
.B(n_172),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_242),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_160),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_193),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_174),
.C(n_178),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_217),
.B(n_189),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_201),
.B(n_178),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_238),
.B(n_5),
.C(n_6),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_187),
.B(n_4),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_241),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_185),
.A2(n_206),
.B1(n_203),
.B2(n_204),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_240),
.A2(n_243),
.B1(n_211),
.B2(n_196),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_190),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_209),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_200),
.B(n_11),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_SL g254 ( 
.A(n_245),
.B(n_214),
.C(n_212),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_204),
.B1(n_198),
.B2(n_199),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_247),
.A2(n_250),
.B1(n_259),
.B2(n_228),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_SL g270 ( 
.A(n_248),
.B(n_252),
.C(n_266),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_231),
.A2(n_195),
.B1(n_204),
.B2(n_208),
.Y(n_249)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_249),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_191),
.B1(n_205),
.B2(n_212),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_220),
.B(n_207),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_258),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_224),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_196),
.B1(n_6),
.B2(n_7),
.Y(n_255)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_235),
.B(n_11),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_257),
.B(n_234),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_12),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_12),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_267),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_243),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_265)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_265),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_222),
.B(n_226),
.C(n_232),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_246),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_277),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_229),
.Y(n_272)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_272),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_278),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_253),
.Y(n_275)
);

INVx13_ASAP7_75t_L g289 ( 
.A(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_218),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_239),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_279),
.B(n_283),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_260),
.A2(n_223),
.B1(n_224),
.B2(n_237),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_281),
.A2(n_257),
.B1(n_233),
.B2(n_234),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_256),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_256),
.C(n_264),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_248),
.B(n_254),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_247),
.A2(n_223),
.B(n_236),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_285),
.A2(n_264),
.B(n_227),
.Y(n_295)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_250),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_258),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_296),
.C(n_300),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_279),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g294 ( 
.A1(n_270),
.A2(n_249),
.B1(n_259),
.B2(n_266),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_294),
.A2(n_271),
.B(n_270),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_276),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_262),
.C(n_221),
.Y(n_296)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_297),
.Y(n_309)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_280),
.B(n_251),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_10),
.C(n_12),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_301),
.B(n_302),
.C(n_274),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_13),
.C(n_14),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_303),
.A2(n_315),
.B1(n_291),
.B2(n_301),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_286),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_294),
.Y(n_305)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_306),
.Y(n_322)
);

XNOR2x1_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_290),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_307),
.A2(n_298),
.B1(n_294),
.B2(n_290),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_296),
.C(n_288),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_313),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_272),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_314),
.B(n_13),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_273),
.B(n_278),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_317),
.B(n_320),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_319),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_311),
.B(n_291),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_321),
.A2(n_303),
.B(n_307),
.Y(n_326)
);

AOI211xp5_ASAP7_75t_L g334 ( 
.A1(n_326),
.A2(n_327),
.B(n_330),
.C(n_317),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_SL g327 ( 
.A(n_319),
.B(n_308),
.Y(n_327)
);

AND2x4_ASAP7_75t_SL g330 ( 
.A(n_322),
.B(n_313),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_329),
.A2(n_312),
.B1(n_318),
.B2(n_309),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_334),
.C(n_310),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g332 ( 
.A1(n_325),
.A2(n_323),
.B(n_324),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_332),
.B(n_333),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_328),
.B(n_316),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_332),
.Y(n_337)
);

OAI32xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_335),
.A3(n_310),
.B1(n_295),
.B2(n_276),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_300),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_283),
.B1(n_14),
.B2(n_15),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_14),
.Y(n_341)
);


endmodule