module fake_jpeg_7574_n_134 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_12),
.B1(n_21),
.B2(n_13),
.Y(n_38)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_18),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_19),
.B1(n_23),
.B2(n_20),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_40),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_12),
.B(n_21),
.C(n_22),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_15),
.Y(n_49)
);

CKINVDCx11_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_48),
.Y(n_66)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_44),
.B(n_53),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_13),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_45),
.A2(n_18),
.B(n_16),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_37),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_46),
.B(n_49),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_15),
.C(n_11),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_3),
.Y(n_77)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g54 ( 
.A1(n_32),
.A2(n_19),
.B1(n_11),
.B2(n_22),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_59),
.B1(n_36),
.B2(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_55),
.B(n_57),
.Y(n_79)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_0),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_60),
.B(n_7),
.C(n_8),
.Y(n_75)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_58),
.A2(n_18),
.B1(n_36),
.B2(n_4),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_32),
.A2(n_24),
.B1(n_23),
.B2(n_16),
.Y(n_59)
);

AND2x6_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_1),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_2),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_67),
.B(n_74),
.Y(n_90)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

OAI21xp33_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_5),
.B(n_50),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_2),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_44),
.B(n_47),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_76),
.B(n_78),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_7),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_4),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_80),
.B(n_82),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_81),
.A2(n_75),
.B1(n_69),
.B2(n_67),
.Y(n_102)
);

AOI222xp33_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_78),
.B1(n_74),
.B2(n_77),
.C1(n_87),
.C2(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_89),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_64),
.B(n_8),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_87),
.A2(n_88),
.B(n_76),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_65),
.A2(n_53),
.B(n_51),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_66),
.B(n_9),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_92),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_97),
.B(n_99),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_98),
.A2(n_100),
.B(n_63),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_102),
.B(n_103),
.Y(n_111)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_105),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_95),
.B(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_106),
.B(n_68),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_93),
.B1(n_83),
.B2(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_110),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_101),
.B1(n_87),
.B2(n_91),
.Y(n_112)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_113),
.A2(n_98),
.B(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_119),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_105),
.B(n_104),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_118),
.B(n_68),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_96),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_114),
.A2(n_117),
.B1(n_111),
.B2(n_108),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_124),
.B(n_85),
.C(n_77),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_116),
.A2(n_110),
.B(n_113),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_109),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_82),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_123),
.B(n_72),
.C(n_85),
.Y(n_125)
);

NOR2xp67_ASAP7_75t_SL g131 ( 
.A(n_125),
.B(n_127),
.Y(n_131)
);

A2O1A1Ixp33_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_128),
.B(n_124),
.C(n_123),
.Y(n_129)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_120),
.A2(n_109),
.B(n_71),
.C(n_51),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_128),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_130),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.Y(n_134)
);


endmodule