module fake_jpeg_2729_n_270 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_270);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_270;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_152;
wire n_73;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_8),
.B(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_12),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_40),
.B(n_45),
.Y(n_108)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_23),
.A2(n_8),
.B(n_13),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_42),
.B(n_49),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_52),
.Y(n_83)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_51),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_8),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_50),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_22),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_20),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_27),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_30),
.Y(n_60)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_40),
.B(n_19),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_52),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_66),
.B(n_75),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_43),
.A2(n_24),
.B1(n_28),
.B2(n_38),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_67),
.A2(n_74),
.B1(n_84),
.B2(n_86),
.Y(n_113)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_70),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_24),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g74 ( 
.A1(n_54),
.A2(n_28),
.B1(n_34),
.B2(n_33),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_35),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_41),
.A2(n_25),
.B1(n_15),
.B2(n_26),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_78),
.A2(n_79),
.B1(n_88),
.B2(n_101),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_41),
.A2(n_25),
.B1(n_15),
.B2(n_26),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_39),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_82),
.Y(n_118)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_16),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_39),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_87),
.B(n_105),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_27),
.B1(n_16),
.B2(n_32),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_31),
.B1(n_18),
.B2(n_32),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_90),
.A2(n_111),
.B1(n_58),
.B2(n_62),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_27),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_94),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_27),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_1),
.Y(n_140)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

CKINVDCx12_ASAP7_75t_R g98 ( 
.A(n_58),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_47),
.A2(n_31),
.B1(n_18),
.B2(n_36),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_102),
.Y(n_137)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_110),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_57),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_47),
.A2(n_36),
.B1(n_3),
.B2(n_4),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_123),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_83),
.B(n_63),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_120),
.B(n_125),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_140),
.Y(n_144)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_44),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_83),
.B(n_63),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_74),
.A2(n_44),
.B1(n_57),
.B2(n_61),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_126),
.A2(n_128),
.B1(n_132),
.B2(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_64),
.B(n_44),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_139),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_130),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_67),
.A2(n_36),
.B1(n_9),
.B2(n_10),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_91),
.B1(n_71),
.B2(n_89),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_36),
.B1(n_3),
.B2(n_4),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_7),
.C(n_13),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_107),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_1),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_77),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_3),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_70),
.A2(n_9),
.B1(n_11),
.B2(n_14),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_84),
.B1(n_99),
.B2(n_72),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_116),
.B(n_76),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_148),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_171),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_116),
.B(n_77),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_104),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_104),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_151),
.B(n_154),
.Y(n_183)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_152),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g154 ( 
.A(n_140),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_73),
.B(n_109),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_162),
.B(n_92),
.Y(n_195)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_95),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_113),
.A2(n_97),
.B1(n_103),
.B2(n_102),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_172),
.B1(n_136),
.B2(n_134),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_80),
.B1(n_100),
.B2(n_89),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_164),
.B1(n_165),
.B2(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_141),
.Y(n_175)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_114),
.A2(n_73),
.A3(n_92),
.B1(n_85),
.B2(n_107),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_114),
.A2(n_119),
.B1(n_113),
.B2(n_121),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_128),
.B1(n_140),
.B2(n_121),
.Y(n_169)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_120),
.A2(n_80),
.B1(n_100),
.B2(n_71),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_160),
.B1(n_167),
.B2(n_172),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_175),
.B(n_179),
.Y(n_203)
);

NOR2xp67_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_130),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_187),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_125),
.B1(n_139),
.B2(n_127),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_192),
.B1(n_153),
.B2(n_143),
.Y(n_206)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_144),
.A2(n_136),
.B1(n_142),
.B2(n_124),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_155),
.B(n_130),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_185),
.C(n_186),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_124),
.C(n_129),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_129),
.C(n_122),
.Y(n_186)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_112),
.C(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_188),
.B(n_190),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_138),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_137),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_191),
.B(n_153),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_159),
.A2(n_165),
.B1(n_167),
.B2(n_170),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_144),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_199),
.B1(n_205),
.B2(n_206),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_198),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_174),
.A2(n_144),
.B1(n_147),
.B2(n_156),
.Y(n_199)
);

AOI221xp5_ASAP7_75t_L g218 ( 
.A1(n_201),
.A2(n_211),
.B1(n_181),
.B2(n_192),
.C(n_195),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g202 ( 
.A(n_183),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_209),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_174),
.A2(n_168),
.B1(n_162),
.B2(n_143),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_207),
.Y(n_216)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_173),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_212),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_177),
.A2(n_91),
.B1(n_152),
.B2(n_166),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_193),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_188),
.C(n_180),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_213),
.B(n_215),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_180),
.C(n_182),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_186),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_224),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_218),
.A2(n_196),
.B1(n_211),
.B2(n_194),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_200),
.B(n_185),
.C(n_187),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_220),
.B(n_223),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_194),
.B(n_189),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_226),
.B(n_219),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_198),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_184),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_194),
.B(n_179),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_175),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_212),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_221),
.A2(n_210),
.B1(n_206),
.B2(n_197),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_219),
.A2(n_226),
.B1(n_205),
.B2(n_225),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_234),
.B1(n_235),
.B2(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_200),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_231),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_233),
.A2(n_229),
.B(n_232),
.Y(n_247)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_220),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_213),
.C(n_215),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_240),
.C(n_242),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_227),
.C(n_217),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_241),
.B(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_224),
.C(n_222),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_237),
.B(n_179),
.Y(n_243)
);

OAI21x1_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_228),
.B(n_209),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_214),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_250),
.Y(n_258)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_244),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_241),
.A2(n_237),
.B(n_233),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_239),
.B(n_231),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_253),
.B(n_246),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_254),
.Y(n_263)
);

NOR2xp67_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_242),
.Y(n_256)
);

OAI21x1_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_249),
.B(n_243),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_246),
.Y(n_259)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_259),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_260),
.A2(n_166),
.B(n_171),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_254),
.C(n_207),
.Y(n_261)
);

A2O1A1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_261),
.A2(n_258),
.B(n_190),
.C(n_255),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_263),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_9),
.C(n_4),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_262),
.C(n_85),
.Y(n_267)
);

AOI221xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_268),
.B1(n_264),
.B2(n_3),
.C(n_5),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_269),
.B(n_5),
.C(n_262),
.Y(n_270)
);


endmodule