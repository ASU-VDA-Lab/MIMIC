module fake_jpeg_4258_n_205 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx13_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_0),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_33),
.Y(n_52)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_35),
.B1(n_28),
.B2(n_24),
.Y(n_39)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx24_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_46),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_26),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_45),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_33),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_41),
.A2(n_43),
.B1(n_27),
.B2(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_28),
.B1(n_29),
.B2(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_15),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_49),
.B(n_15),
.Y(n_57)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_37),
.Y(n_75)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_53),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

OAI32xp33_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_45),
.A3(n_43),
.B1(n_41),
.B2(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_64),
.Y(n_86)
);

OR2x4_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_58),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_22),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_60),
.B(n_62),
.Y(n_95)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_36),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_19),
.C(n_23),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_67),
.A2(n_74),
.B1(n_15),
.B2(n_26),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_25),
.B(n_18),
.Y(n_97)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_29),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_71),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_23),
.B1(n_19),
.B2(n_21),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_42),
.B(n_34),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_66),
.B1(n_65),
.B2(n_60),
.Y(n_91)
);

AO21x2_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_51),
.B(n_34),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_78),
.A2(n_97),
.B(n_61),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_36),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_58),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_77),
.A2(n_48),
.B1(n_42),
.B2(n_23),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_82),
.B(n_84),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_21),
.B1(n_20),
.B2(n_27),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_27),
.B1(n_20),
.B2(n_17),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_56),
.A2(n_16),
.B1(n_17),
.B2(n_31),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_59),
.A2(n_16),
.B1(n_37),
.B2(n_32),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_91),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_36),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_70),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_58),
.A2(n_37),
.B1(n_36),
.B2(n_32),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_101),
.B(n_62),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_57),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_102),
.B(n_53),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_106),
.B(n_116),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_117),
.C(n_94),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_79),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_112),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_70),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_85),
.Y(n_132)
);

NOR4xp25_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_63),
.C(n_32),
.D(n_3),
.Y(n_114)
);

AOI21xp33_ASAP7_75t_SL g129 ( 
.A1(n_114),
.A2(n_93),
.B(n_84),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_115),
.B(n_118),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_25),
.B(n_73),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_78),
.A2(n_97),
.B(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_95),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_54),
.Y(n_119)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_78),
.A2(n_25),
.B(n_69),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_54),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_122),
.B(n_87),
.Y(n_125)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_125),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_138),
.C(n_117),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_131),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_108),
.A2(n_78),
.B1(n_101),
.B2(n_82),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_136),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_122),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_72),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_142),
.Y(n_159)
);

A2O1A1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_141),
.A2(n_103),
.B(n_114),
.C(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_83),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_124),
.B(n_143),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_126),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_106),
.C(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_148),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_116),
.C(n_115),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_110),
.C(n_102),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_150),
.B(n_154),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_151),
.B(n_152),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_110),
.C(n_108),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_107),
.B(n_105),
.C(n_120),
.D(n_98),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_156),
.B(n_142),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g180 ( 
.A1(n_160),
.A2(n_14),
.B(n_12),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_155),
.B(n_157),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_164),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_169),
.B(n_80),
.Y(n_179)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_170),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_149),
.A2(n_141),
.B1(n_126),
.B2(n_131),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_168),
.B1(n_153),
.B2(n_145),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_152),
.A2(n_137),
.B1(n_132),
.B2(n_141),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_158),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_144),
.B(n_11),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_160),
.A2(n_151),
.B1(n_156),
.B2(n_145),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_172),
.B(n_173),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g173 ( 
.A(n_167),
.B(n_163),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_145),
.C(n_128),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_176),
.B(n_178),
.C(n_172),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_80),
.C(n_98),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_166),
.Y(n_184)
);

OAI21x1_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_14),
.B(n_11),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_123),
.B1(n_92),
.B2(n_4),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_92),
.B1(n_2),
.B2(n_4),
.Y(n_185)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_170),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_176),
.B(n_175),
.C(n_6),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_187),
.B(n_188),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_185),
.B(n_175),
.Y(n_193)
);

OAI221xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.C(n_6),
.Y(n_191)
);

INVxp33_ASAP7_75t_SL g189 ( 
.A(n_178),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_189),
.A2(n_1),
.B(n_5),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_192),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_189),
.B1(n_182),
.B2(n_9),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_195),
.B(n_7),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_1),
.B(n_5),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_197),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_7),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_198),
.B(n_8),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_8),
.C(n_10),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_10),
.B(n_201),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_204),
.Y(n_205)
);


endmodule