module fake_ariane_2791_n_6325 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_6325);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_6325;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_5553;
wire n_6002;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_5717;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_5791;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_5712;
wire n_3954;
wire n_6297;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_6058;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_6293;
wire n_2482;
wire n_1682;
wire n_958;
wire n_6129;
wire n_2554;
wire n_4321;
wire n_5590;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_6313;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_6190;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_625;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_5896;
wire n_4567;
wire n_786;
wire n_5833;
wire n_6249;
wire n_6253;
wire n_6128;
wire n_3552;
wire n_2950;
wire n_6197;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_5744;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_3482;
wire n_6295;
wire n_5403;
wire n_823;
wire n_1900;
wire n_620;
wire n_6096;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_899;
wire n_3975;
wire n_5830;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_661;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_6161;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_6136;
wire n_1140;
wire n_3458;
wire n_5843;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_6156;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_5913;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5757;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_6236;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_5968;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_5586;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5971;
wire n_6319;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5984;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_619;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_5897;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_6261;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5778;
wire n_5179;
wire n_2435;
wire n_5680;
wire n_1932;
wire n_6210;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5974;
wire n_5723;
wire n_5922;
wire n_5549;
wire n_1087;
wire n_632;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_6044;
wire n_1841;
wire n_1680;
wire n_6206;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_5831;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_5708;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_646;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_6033;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_6060;
wire n_3108;
wire n_5788;
wire n_5983;
wire n_2632;
wire n_5557;
wire n_4314;
wire n_2980;
wire n_5951;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_6117;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_6009;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_670;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_6192;
wire n_5773;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_6263;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_6048;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_6234;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_6224;
wire n_5089;
wire n_5775;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_6142;
wire n_2617;
wire n_6119;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_6189;
wire n_1053;
wire n_5796;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_5960;
wire n_3007;
wire n_2267;
wire n_5858;
wire n_5985;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_6304;
wire n_4292;
wire n_2118;
wire n_688;
wire n_636;
wire n_1490;
wire n_5552;
wire n_6074;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_1104;
wire n_986;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5742;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_6229;
wire n_1863;
wire n_5933;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_616;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_5810;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_5818;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_5889;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_5450;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_6031;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_655;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_5719;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5904;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_6012;
wire n_704;
wire n_2958;
wire n_1714;
wire n_4429;
wire n_1044;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_608;
wire n_2457;
wire n_2992;
wire n_6124;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_5829;
wire n_2520;
wire n_811;
wire n_791;
wire n_5881;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_6201;
wire n_3450;
wire n_687;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_642;
wire n_5073;
wire n_1406;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_5894;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_6036;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_6102;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_6244;
wire n_4846;
wire n_1330;
wire n_906;
wire n_6204;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_5826;
wire n_4822;
wire n_5931;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_5532;
wire n_3740;
wire n_5441;
wire n_6179;
wire n_2417;
wire n_6059;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_5994;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_5772;
wire n_6188;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_5921;
wire n_6247;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_6104;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_6205;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_1593;
wire n_2610;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5884;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_5728;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_5679;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_5879;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_775;
wire n_667;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_5825;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_5629;
wire n_5759;
wire n_2411;
wire n_4631;
wire n_5999;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_6180;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_6004;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_6275;
wire n_3497;
wire n_4542;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_6141;
wire n_3595;
wire n_2068;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_6194;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5807;
wire n_5426;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_6318;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_1056;
wire n_5584;
wire n_674;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_6075;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_6068;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_6248;
wire n_848;
wire n_5125;
wire n_4922;
wire n_6066;
wire n_6080;
wire n_629;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_6150;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_5906;
wire n_2189;
wire n_5732;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_5780;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_6006;
wire n_3597;
wire n_5743;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_3786;
wire n_875;
wire n_6022;
wire n_2828;
wire n_1626;
wire n_5950;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_793;
wire n_5705;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_6116;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_5875;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_5848;
wire n_1679;
wire n_5834;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_5784;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_6209;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_6274;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_6237;
wire n_1525;
wire n_4628;
wire n_5982;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_6155;
wire n_2901;
wire n_3940;
wire n_6099;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5824;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_6203;
wire n_2138;
wire n_4230;
wire n_3040;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_5276;
wire n_2000;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_5763;
wire n_3633;
wire n_857;
wire n_6061;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_1064;
wire n_633;
wire n_1446;
wire n_1701;
wire n_6273;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_6174;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_5907;
wire n_784;
wire n_4339;
wire n_6013;
wire n_6182;
wire n_4690;
wire n_2987;
wire n_6279;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_5895;
wire n_2651;
wire n_753;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_3632;
wire n_2522;
wire n_1344;
wire n_4064;
wire n_6131;
wire n_3351;
wire n_5478;
wire n_6113;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_2324;
wire n_840;
wire n_5283;
wire n_3454;
wire n_5961;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_2740;
wire n_1991;
wire n_614;
wire n_4066;
wire n_6252;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_3445;
wire n_2105;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1148;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5949;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_6049;
wire n_5885;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_658;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_5856;
wire n_3872;
wire n_5760;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_5844;
wire n_6298;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_5938;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_6132;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_1168;
wire n_4663;
wire n_5840;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_656;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_3895;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_5917;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_6168;
wire n_5304;
wire n_5437;
wire n_1581;
wire n_3058;
wire n_946;
wire n_757;
wire n_5355;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_6284;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_5915;
wire n_1368;
wire n_963;
wire n_6306;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_1115;
wire n_4654;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5966;
wire n_5515;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_6046;
wire n_1233;
wire n_4493;
wire n_6055;
wire n_1808;
wire n_6091;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_6144;
wire n_1451;
wire n_1487;
wire n_675;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5753;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_6221;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_6285;
wire n_610;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_5901;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_6115;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_6272;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_5497;
wire n_5519;
wire n_6071;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_6178;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_6191;
wire n_2442;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_645;
wire n_5098;
wire n_721;
wire n_1084;
wire n_6000;
wire n_1276;
wire n_5145;
wire n_6072;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_5466;
wire n_1528;
wire n_3315;
wire n_6094;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_5738;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_5953;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_6098;
wire n_5995;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_612;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2685;
wire n_2061;
wire n_5987;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_6291;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_5873;
wire n_4498;
wire n_772;
wire n_1245;
wire n_5741;
wire n_2743;
wire n_1669;
wire n_3429;
wire n_2969;
wire n_1675;
wire n_2466;
wire n_676;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_6056;
wire n_5926;
wire n_5866;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_652;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_5877;
wire n_912;
wire n_4786;
wire n_6042;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_6315;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_6133;
wire n_2693;
wire n_5408;
wire n_5812;
wire n_5540;
wire n_5804;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_6241;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_5992;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_5981;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_5737;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_6083;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_6278;
wire n_2274;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_6101;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_5905;
wire n_6112;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_6271;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_926;
wire n_2296;
wire n_5735;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_6037;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_5787;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_5935;
wire n_4916;
wire n_5967;
wire n_6095;
wire n_4323;
wire n_5934;
wire n_1899;
wire n_6045;
wire n_5376;
wire n_3508;
wire n_6300;
wire n_4129;
wire n_5488;
wire n_1105;
wire n_5727;
wire n_3599;
wire n_5988;
wire n_5646;
wire n_4480;
wire n_5711;
wire n_3734;
wire n_5832;
wire n_6254;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_5891;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_6011;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_6176;
wire n_1963;
wire n_3868;
wire n_729;
wire n_6222;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_6308;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3568;
wire n_3216;
wire n_2708;
wire n_6187;
wire n_735;
wire n_4844;
wire n_6220;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_5650;
wire n_5729;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_6149;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_5762;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_5874;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_606;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_659;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_6034;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_5910;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_5941;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_6019;
wire n_4977;
wire n_2492;
wire n_3425;
wire n_2939;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_5936;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_5928;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_5785;
wire n_3411;
wire n_5222;
wire n_6165;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_6114;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_649;
wire n_1561;
wire n_5494;
wire n_5970;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_1557;
wire n_6166;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_4764;
wire n_2408;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_5800;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5766;
wire n_5293;
wire n_779;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_6047;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_6258;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_6026;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_5882;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_5606;
wire n_2310;
wire n_5911;
wire n_3600;
wire n_1023;
wire n_914;
wire n_689;
wire n_6139;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_638;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_5849;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_5841;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_685;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_617;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_918;
wire n_5645;
wire n_639;
wire n_5020;
wire n_673;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_6183;
wire n_6107;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_6003;
wire n_5443;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_5631;
wire n_3481;
wire n_5101;
wire n_6020;
wire n_2236;
wire n_6185;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_5608;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_622;
wire n_4584;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_5806;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_6213;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_5747;
wire n_1204;
wire n_2428;
wire n_994;
wire n_1360;
wire n_6063;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_6153;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_6202;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_5690;
wire n_1980;
wire n_5740;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_6082;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_679;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_6105;
wire n_826;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_5898;
wire n_607;
wire n_5923;
wire n_3687;
wire n_2787;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_5946;
wire n_1268;
wire n_2676;
wire n_4550;
wire n_2770;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_6163;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_5836;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_5739;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_6023;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_6196;
wire n_5425;
wire n_5273;
wire n_5839;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_5887;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_6321;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_5880;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_671;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_6064;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_684;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_6164;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_5730;
wire n_6292;
wire n_4165;
wire n_2056;
wire n_5754;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_5756;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_6015;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_662;
wire n_3461;
wire n_1410;
wire n_2297;
wire n_939;
wire n_4203;
wire n_5789;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_933;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_6073;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_4761;
wire n_2052;
wire n_4627;
wire n_4556;
wire n_6137;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_5751;
wire n_626;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_6120;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5997;
wire n_5375;
wire n_5438;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_6135;
wire n_1752;
wire n_2361;
wire n_3030;
wire n_4538;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_4730;
wire n_1296;
wire n_4421;
wire n_6230;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_5932;
wire n_6121;
wire n_3430;
wire n_1299;
wire n_5919;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_6001;
wire n_4971;
wire n_2095;
wire n_5664;
wire n_2738;
wire n_5890;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_5823;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5944;
wire n_6299;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_1069;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5725;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_4259;
wire n_5870;
wire n_2030;
wire n_6053;
wire n_850;
wire n_6233;
wire n_4299;
wire n_5625;
wire n_2407;
wire n_690;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_6010;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_5570;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_5265;
wire n_5955;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_6032;
wire n_1196;
wire n_5733;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_4575;
wire n_945;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_5978;
wire n_3220;
wire n_4581;
wire n_6008;
wire n_665;
wire n_4625;
wire n_6181;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_672;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_5290;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_6170;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_5845;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_5969;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_6005;
wire n_611;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_5736;
wire n_4929;
wire n_2874;
wire n_6029;
wire n_4117;
wire n_6025;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_6085;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_6062;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_5847;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_5718;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5546;
wire n_6294;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_6079;
wire n_6260;
wire n_680;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_5544;
wire n_5660;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_6314;
wire n_5610;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1468;
wire n_1253;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_6065;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_5808;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_5770;
wire n_5710;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_5799;
wire n_6265;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_6148;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_650;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_6087;
wire n_964;
wire n_2220;
wire n_6108;
wire n_6100;
wire n_4433;
wire n_2829;
wire n_5862;
wire n_1914;
wire n_2253;
wire n_5886;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_5802;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_6103;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_5883;
wire n_1095;
wire n_3078;
wire n_6078;
wire n_3971;
wire n_5630;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_6207;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5929;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_5975;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_5496;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_5991;
wire n_4952;
wire n_4426;
wire n_5956;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_6017;
wire n_3946;
wire n_5920;
wire n_2112;
wire n_2640;
wire n_6125;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_6097;
wire n_6057;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_6302;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_6223;
wire n_4039;
wire n_5793;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_5761;
wire n_677;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_5681;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_6195;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_627;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_5748;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_6200;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_5657;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5765;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_6106;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_6287;
wire n_2840;
wire n_6172;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_5957;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_666;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_6067;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_5867;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_6296;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_5822;
wire n_5786;
wire n_3586;
wire n_5817;
wire n_4160;
wire n_6109;
wire n_1668;
wire n_5798;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_5713;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_618;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_6309;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_5989;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_640;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_5908;
wire n_1352;
wire n_5431;
wire n_643;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_682;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_5752;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_5746;
wire n_686;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_4666;
wire n_4082;
wire n_3140;
wire n_2320;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_6016;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_5903;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_4721;
wire n_2170;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_5912;
wire n_5745;
wire n_6086;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5803;
wire n_5593;
wire n_5270;
wire n_5853;
wire n_6171;
wire n_3468;
wire n_5779;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_879;
wire n_5446;
wire n_4561;
wire n_1541;
wire n_3291;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_1185;
wire n_2475;
wire n_4715;
wire n_6157;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_1090;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_6162;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_6127;
wire n_1440;
wire n_6246;
wire n_1370;
wire n_5005;
wire n_6126;
wire n_1549;
wire n_6151;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_683;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_5755;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_4711;
wire n_2749;
wire n_5962;
wire n_660;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_6154;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_5801;
wire n_3904;
wire n_6054;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_613;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_5721;
wire n_2609;
wire n_6184;
wire n_1767;
wire n_4138;
wire n_3131;
wire n_1040;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_6312;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_6193;
wire n_3992;
wire n_6007;
wire n_621;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_6208;
wire n_2881;
wire n_6303;
wire n_3092;
wire n_6014;
wire n_4270;
wire n_697;
wire n_4620;
wire n_5397;
wire n_6255;
wire n_4924;
wire n_4044;
wire n_6270;
wire n_2305;
wire n_5996;
wire n_880;
wire n_5566;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_6276;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_5805;
wire n_932;
wire n_6266;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_5758;
wire n_5842;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_6147;
wire n_5692;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_6211;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_6093;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_5902;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_6215;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_969;
wire n_1663;
wire n_5952;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_5716;
wire n_3897;
wire n_1735;
wire n_5888;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_5980;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_5790;
wire n_4647;
wire n_3575;
wire n_6310;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_6259;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_6289;
wire n_4059;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_5948;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_648;
wire n_3273;
wire n_2918;
wire n_835;
wire n_6186;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_6035;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_5850;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_635;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_5940;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_6232;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_5860;
wire n_2422;
wire n_654;
wire n_2933;
wire n_3387;
wire n_6214;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_6143;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_6225;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_5859;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_6219;
wire n_723;
wire n_1393;
wire n_6175;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_6198;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1982;
wire n_641;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_6281;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_5878;
wire n_2674;
wire n_5820;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_954;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_5964;
wire n_2673;
wire n_6076;
wire n_4678;
wire n_664;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_5776;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_5909;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_5750;
wire n_1232;
wire n_1211;
wire n_996;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_5837;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_6226;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_6283;
wire n_4688;
wire n_4939;
wire n_5900;
wire n_1486;
wire n_3619;
wire n_6158;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_6122;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_5486;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_5851;
wire n_6317;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_6269;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_1214;
wire n_634;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_6088;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_5855;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_5861;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_5749;
wire n_6320;
wire n_6316;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_5998;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_6250;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_5827;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_5656;
wire n_1988;
wire n_5678;
wire n_5865;
wire n_6050;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_5815;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_5965;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_6024;
wire n_4768;
wire n_1889;
wire n_6090;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_6038;
wire n_2902;
wire n_6030;
wire n_6245;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_5871;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_6052;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_6280;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_5939;
wire n_1819;
wire n_3095;
wire n_947;
wire n_5792;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_4775;
wire n_696;
wire n_1442;
wire n_6256;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2549;
wire n_2499;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_5954;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_6324;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_669;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_6243;
wire n_5795;
wire n_5715;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_2155;
wire n_6231;
wire n_615;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_6041;
wire n_824;
wire n_5659;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_6323;
wire n_5720;
wire n_4267;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5854;
wire n_5958;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_5783;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_965;
wire n_5809;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_5993;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_836;
wire n_3464;
wire n_6290;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_5821;
wire n_713;
wire n_3179;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_6118;
wire n_706;
wire n_2120;
wire n_6028;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_6267;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_5943;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_6216;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_637;
wire n_5335;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_5771;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_6167;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_5698;
wire n_5731;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_6159;
wire n_2129;
wire n_5857;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_647;
wire n_2027;
wire n_2932;
wire n_6217;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_1467;
wire n_5209;
wire n_6307;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_5916;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_681;
wire n_3286;
wire n_5781;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_6140;
wire n_6111;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_6240;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_5673;
wire n_861;
wire n_5814;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_6069;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_6077;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_6040;
wire n_1890;
wire n_6305;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_657;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_5769;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_6239;
wire n_3208;
wire n_5768;
wire n_1342;
wire n_6199;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_5963;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_5972;
wire n_3400;
wire n_1466;
wire n_6177;
wire n_2581;
wire n_5937;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_6173;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_6218;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_624;
wire n_5577;
wire n_876;
wire n_5872;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_5976;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_5838;
wire n_3694;
wire n_771;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_5846;
wire n_2307;
wire n_3702;
wire n_5930;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_1324;
wire n_3543;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_6257;
wire n_4152;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_6039;
wire n_6286;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_5816;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_6018;
wire n_1286;
wire n_6021;
wire n_4617;
wire n_1685;
wire n_4611;
wire n_2477;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_5797;
wire n_1052;
wire n_4732;
wire n_2076;
wire n_2203;
wire n_5942;
wire n_5764;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_5777;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_6322;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_6130;
wire n_5868;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_644;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_5986;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_5794;
wire n_3141;
wire n_5272;
wire n_2053;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_6123;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_5722;
wire n_5811;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_623;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_628;
wire n_5863;
wire n_3790;
wire n_907;
wire n_6152;
wire n_5734;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_6169;
wire n_5774;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_609;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_5977;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_5959;
wire n_3563;
wire n_5945;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_6301;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_6282;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_5767;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_5973;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_5869;
wire n_5914;
wire n_2114;
wire n_3329;
wire n_3833;
wire n_2927;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_6043;
wire n_6268;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_6145;
wire n_2865;
wire n_5925;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_6311;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_6134;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_653;
wire n_6262;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5876;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_6160;
wire n_4667;
wire n_5813;
wire n_6235;
wire n_1471;
wire n_6212;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_5892;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_5714;
wire n_2169;
wire n_6089;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_5990;
wire n_2175;
wire n_1625;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_6138;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_6070;
wire n_5852;
wire n_5918;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_5947;
wire n_6242;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_5835;
wire n_668;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_5819;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_5893;
wire n_2710;
wire n_6092;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_6251;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_5726;
wire n_4371;
wire n_1902;
wire n_5828;
wire n_2784;
wire n_3898;
wire n_694;
wire n_6228;
wire n_4749;
wire n_5924;
wire n_1845;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_5899;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_6264;
wire n_5782;
wire n_630;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_5864;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_6084;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_6288;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_5709;
wire n_1764;
wire n_4807;
wire n_6277;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_5927;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_6051;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_6227;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_5696;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_6146;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_6081;
wire n_1249;
wire n_5724;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_5979;
wire n_6027;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_6110;
wire n_1762;
wire n_6238;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_231),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_389),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g608 ( 
.A(n_302),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_393),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_308),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_586),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_411),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_1),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_418),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_396),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_366),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_260),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_104),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_589),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_342),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_45),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_510),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_177),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_391),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_88),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_388),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_344),
.Y(n_627)
);

CKINVDCx20_ASAP7_75t_R g628 ( 
.A(n_74),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_180),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_364),
.Y(n_630)
);

CKINVDCx20_ASAP7_75t_R g631 ( 
.A(n_184),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_2),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_307),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_593),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_411),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_346),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_334),
.Y(n_637)
);

BUFx10_ASAP7_75t_L g638 ( 
.A(n_464),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_236),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_2),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_6),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_125),
.Y(n_642)
);

INVx1_ASAP7_75t_SL g643 ( 
.A(n_524),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_228),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_333),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_451),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_437),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_438),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_522),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_197),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_365),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_115),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_431),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_309),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_378),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_471),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_372),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_413),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_376),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_104),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_534),
.Y(n_661)
);

BUFx8_ASAP7_75t_SL g662 ( 
.A(n_348),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_540),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_151),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_492),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_332),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_360),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_28),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_519),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_386),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_513),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_386),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_418),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_159),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_452),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_602),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_285),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_393),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_224),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_486),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_40),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_355),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_521),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_329),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_536),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_423),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_495),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_4),
.Y(n_688)
);

BUFx10_ASAP7_75t_L g689 ( 
.A(n_327),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_164),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_554),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_140),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_112),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_179),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_116),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_125),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_472),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_444),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_234),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_526),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_37),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_394),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_82),
.Y(n_703)
);

CKINVDCx16_ASAP7_75t_R g704 ( 
.A(n_216),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_251),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_15),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_274),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_242),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_59),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_444),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_325),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_53),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_507),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_14),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_138),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_562),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_321),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_310),
.Y(n_718)
);

BUFx6f_ASAP7_75t_L g719 ( 
.A(n_39),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_58),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_546),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_548),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_103),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_247),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_398),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_384),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_445),
.Y(n_727)
);

BUFx5_ASAP7_75t_L g728 ( 
.A(n_2),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_253),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_473),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_461),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_590),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_417),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_261),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_226),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_126),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_27),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_525),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_487),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_43),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_335),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_204),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_103),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_80),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_178),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_381),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_40),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_345),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_441),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_304),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_467),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_402),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_308),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_541),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_422),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_349),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_533),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_453),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_501),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_447),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_452),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_140),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_299),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_458),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_374),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_603),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_15),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_379),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_230),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_340),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_516),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_501),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_232),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_525),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_101),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_436),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_185),
.Y(n_777)
);

CKINVDCx16_ASAP7_75t_R g778 ( 
.A(n_196),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_520),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_372),
.Y(n_780)
);

INVx1_ASAP7_75t_SL g781 ( 
.A(n_251),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_52),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_414),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_433),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_223),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_324),
.Y(n_786)
);

CKINVDCx5p33_ASAP7_75t_R g787 ( 
.A(n_514),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_497),
.Y(n_788)
);

BUFx10_ASAP7_75t_L g789 ( 
.A(n_119),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_120),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_87),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_548),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_194),
.Y(n_793)
);

CKINVDCx20_ASAP7_75t_R g794 ( 
.A(n_537),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_401),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_395),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_159),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_567),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_352),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_194),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_69),
.Y(n_801)
);

BUFx10_ASAP7_75t_L g802 ( 
.A(n_106),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_13),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_487),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_378),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_328),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_5),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_392),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_258),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_594),
.Y(n_810)
);

HB1xp67_ASAP7_75t_L g811 ( 
.A(n_399),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_371),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_459),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_388),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_245),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_221),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_84),
.Y(n_817)
);

BUFx6f_ASAP7_75t_L g818 ( 
.A(n_239),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_211),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_245),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_329),
.Y(n_821)
);

CKINVDCx20_ASAP7_75t_R g822 ( 
.A(n_23),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_575),
.Y(n_823)
);

INVx1_ASAP7_75t_SL g824 ( 
.A(n_423),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_534),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_79),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_250),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_558),
.Y(n_828)
);

INVx2_ASAP7_75t_L g829 ( 
.A(n_382),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_356),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_201),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_142),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_78),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_284),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_539),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_421),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_70),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_550),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_429),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_597),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_434),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_397),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_347),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_604),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_172),
.Y(n_845)
);

CKINVDCx20_ASAP7_75t_R g846 ( 
.A(n_415),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_480),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_102),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_289),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_21),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_567),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_81),
.Y(n_852)
);

CKINVDCx20_ASAP7_75t_R g853 ( 
.A(n_219),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_13),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_169),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_374),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_577),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_321),
.Y(n_858)
);

BUFx6f_ASAP7_75t_L g859 ( 
.A(n_463),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_280),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_58),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_201),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_332),
.Y(n_863)
);

BUFx6f_ASAP7_75t_L g864 ( 
.A(n_547),
.Y(n_864)
);

CKINVDCx20_ASAP7_75t_R g865 ( 
.A(n_542),
.Y(n_865)
);

CKINVDCx20_ASAP7_75t_R g866 ( 
.A(n_508),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_430),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_437),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_318),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_136),
.Y(n_870)
);

BUFx10_ASAP7_75t_L g871 ( 
.A(n_226),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_424),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_20),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_35),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_9),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_205),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_383),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_202),
.Y(n_878)
);

CKINVDCx5p33_ASAP7_75t_R g879 ( 
.A(n_577),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_479),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_249),
.Y(n_881)
);

CKINVDCx20_ASAP7_75t_R g882 ( 
.A(n_412),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_330),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_478),
.Y(n_884)
);

BUFx2_ASAP7_75t_L g885 ( 
.A(n_200),
.Y(n_885)
);

CKINVDCx20_ASAP7_75t_R g886 ( 
.A(n_410),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_432),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_214),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_375),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_603),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_407),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_170),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_139),
.Y(n_893)
);

BUFx10_ASAP7_75t_L g894 ( 
.A(n_574),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_442),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_362),
.Y(n_896)
);

CKINVDCx20_ASAP7_75t_R g897 ( 
.A(n_186),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_356),
.Y(n_898)
);

BUFx5_ASAP7_75t_L g899 ( 
.A(n_28),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_377),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_45),
.Y(n_901)
);

CKINVDCx5p33_ASAP7_75t_R g902 ( 
.A(n_278),
.Y(n_902)
);

BUFx10_ASAP7_75t_L g903 ( 
.A(n_274),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_263),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_563),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_293),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_17),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_48),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_10),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_1),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_275),
.Y(n_911)
);

CKINVDCx20_ASAP7_75t_R g912 ( 
.A(n_109),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_166),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_175),
.Y(n_914)
);

BUFx2_ASAP7_75t_SL g915 ( 
.A(n_561),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_457),
.Y(n_916)
);

CKINVDCx20_ASAP7_75t_R g917 ( 
.A(n_538),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_305),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_94),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_90),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_390),
.Y(n_921)
);

INVx2_ASAP7_75t_SL g922 ( 
.A(n_189),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_161),
.Y(n_923)
);

CKINVDCx20_ASAP7_75t_R g924 ( 
.A(n_41),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_171),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_489),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_336),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_481),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_443),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_500),
.Y(n_930)
);

CKINVDCx20_ASAP7_75t_R g931 ( 
.A(n_8),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_543),
.Y(n_932)
);

INVx1_ASAP7_75t_SL g933 ( 
.A(n_56),
.Y(n_933)
);

INVxp67_ASAP7_75t_SL g934 ( 
.A(n_202),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_493),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_174),
.Y(n_936)
);

INVx1_ASAP7_75t_SL g937 ( 
.A(n_60),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_56),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_87),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_570),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_134),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_340),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_562),
.Y(n_943)
);

BUFx5_ASAP7_75t_L g944 ( 
.A(n_70),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_258),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_210),
.Y(n_946)
);

BUFx5_ASAP7_75t_L g947 ( 
.A(n_366),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_168),
.Y(n_948)
);

BUFx10_ASAP7_75t_L g949 ( 
.A(n_126),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_529),
.Y(n_950)
);

CKINVDCx20_ASAP7_75t_R g951 ( 
.A(n_593),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_156),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_246),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_385),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_490),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_224),
.Y(n_956)
);

BUFx10_ASAP7_75t_L g957 ( 
.A(n_259),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_67),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_605),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_359),
.Y(n_960)
);

CKINVDCx14_ASAP7_75t_R g961 ( 
.A(n_574),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_215),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_601),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_571),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_545),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_373),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_27),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_605),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_602),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_540),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_572),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_173),
.Y(n_972)
);

CKINVDCx5p33_ASAP7_75t_R g973 ( 
.A(n_53),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_123),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_89),
.Y(n_975)
);

BUFx10_ASAP7_75t_L g976 ( 
.A(n_96),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_415),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_13),
.Y(n_978)
);

CKINVDCx20_ASAP7_75t_R g979 ( 
.A(n_23),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_282),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_464),
.Y(n_981)
);

CKINVDCx20_ASAP7_75t_R g982 ( 
.A(n_310),
.Y(n_982)
);

CKINVDCx16_ASAP7_75t_R g983 ( 
.A(n_435),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_334),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_531),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_441),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_280),
.Y(n_987)
);

BUFx8_ASAP7_75t_SL g988 ( 
.A(n_446),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_587),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_592),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_177),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_468),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_416),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_138),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_256),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_513),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_597),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_16),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_460),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_541),
.Y(n_1000)
);

BUFx10_ASAP7_75t_L g1001 ( 
.A(n_586),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_213),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_146),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_331),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_465),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_302),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_17),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_3),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_100),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_504),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_264),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_11),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_157),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_SL g1014 ( 
.A(n_428),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_331),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_400),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_72),
.Y(n_1017)
);

BUFx6f_ASAP7_75t_L g1018 ( 
.A(n_564),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_342),
.Y(n_1019)
);

BUFx3_ASAP7_75t_L g1020 ( 
.A(n_337),
.Y(n_1020)
);

CKINVDCx20_ASAP7_75t_R g1021 ( 
.A(n_532),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_493),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_130),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_403),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_514),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_582),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_180),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_39),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_262),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_214),
.Y(n_1030)
);

INVx1_ASAP7_75t_SL g1031 ( 
.A(n_322),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_287),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_3),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_200),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_324),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_229),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_435),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_554),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_448),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_400),
.Y(n_1040)
);

CKINVDCx5p33_ASAP7_75t_R g1041 ( 
.A(n_419),
.Y(n_1041)
);

CKINVDCx5p33_ASAP7_75t_R g1042 ( 
.A(n_338),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_523),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_79),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_523),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_449),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_127),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_490),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_113),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_491),
.Y(n_1050)
);

INVx1_ASAP7_75t_SL g1051 ( 
.A(n_106),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_419),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_266),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_494),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_243),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_511),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_31),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_425),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_375),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_16),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_494),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_551),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_477),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_585),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_36),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_284),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_466),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_561),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_195),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_368),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_107),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_462),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_83),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_262),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_51),
.Y(n_1075)
);

CKINVDCx14_ASAP7_75t_R g1076 ( 
.A(n_588),
.Y(n_1076)
);

BUFx2_ASAP7_75t_SL g1077 ( 
.A(n_1),
.Y(n_1077)
);

BUFx2_ASAP7_75t_SL g1078 ( 
.A(n_157),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_549),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_528),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_341),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_275),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_361),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_85),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_41),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_77),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_553),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_48),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_404),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_263),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_291),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_535),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_565),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_147),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_345),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_544),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_349),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_133),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_344),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_496),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_431),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_222),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_89),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_137),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_257),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_511),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_347),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_486),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_91),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_380),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_300),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_357),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_420),
.Y(n_1113)
);

CKINVDCx5p33_ASAP7_75t_R g1114 ( 
.A(n_502),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_537),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_387),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_32),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_500),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_575),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_481),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_521),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_466),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_961),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_694),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_688),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_728),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_688),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_961),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_688),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_728),
.Y(n_1130)
);

INVxp67_ASAP7_75t_SL g1131 ( 
.A(n_706),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_1014),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_738),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_738),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_728),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_713),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_738),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_728),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_608),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_738),
.Y(n_1140)
);

INVxp67_ASAP7_75t_SL g1141 ( 
.A(n_706),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_862),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_862),
.Y(n_1143)
);

NOR2xp67_ASAP7_75t_L g1144 ( 
.A(n_862),
.B(n_0),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_728),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1076),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_728),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_706),
.B(n_0),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_862),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_713),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_713),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_1076),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_728),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_717),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_717),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_728),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_717),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_718),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_694),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_662),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_662),
.Y(n_1161)
);

BUFx6f_ASAP7_75t_L g1162 ( 
.A(n_719),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_608),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_718),
.Y(n_1164)
);

CKINVDCx16_ASAP7_75t_R g1165 ( 
.A(n_704),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_718),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_731),
.Y(n_1167)
);

INVx1_ASAP7_75t_SL g1168 ( 
.A(n_1014),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_728),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_988),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_731),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_731),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_988),
.Y(n_1173)
);

XNOR2xp5_ASAP7_75t_L g1174 ( 
.A(n_640),
.B(n_767),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_704),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_797),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_797),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_797),
.Y(n_1178)
);

OR2x2_ASAP7_75t_L g1179 ( 
.A(n_672),
.B(n_0),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_898),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_898),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_778),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_898),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_999),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_778),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_999),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_616),
.Y(n_1187)
);

CKINVDCx16_ASAP7_75t_R g1188 ( 
.A(n_983),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_999),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_983),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_875),
.Y(n_1191)
);

BUFx6f_ASAP7_75t_L g1192 ( 
.A(n_719),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1020),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_1090),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1090),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1114),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1020),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_1119),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1121),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1020),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_616),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_672),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1024),
.Y(n_1203)
);

CKINVDCx14_ASAP7_75t_R g1204 ( 
.A(n_638),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_869),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1024),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1024),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_728),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_606),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_719),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_631),
.Y(n_1211)
);

BUFx2_ASAP7_75t_L g1212 ( 
.A(n_869),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1053),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_899),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1053),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_611),
.Y(n_1216)
);

NOR2xp67_ASAP7_75t_L g1217 ( 
.A(n_875),
.B(n_3),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1053),
.Y(n_1218)
);

HB1xp67_ASAP7_75t_SL g1219 ( 
.A(n_613),
.Y(n_1219)
);

INVxp67_ASAP7_75t_L g1220 ( 
.A(n_811),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1070),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1070),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1070),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_612),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_719),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_899),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_899),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_719),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_619),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_621),
.Y(n_1230)
);

NOR2xp67_ASAP7_75t_L g1231 ( 
.A(n_875),
.B(n_4),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_622),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_899),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_899),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_623),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_624),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_899),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_811),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_899),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_719),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_899),
.Y(n_1241)
);

CKINVDCx5p33_ASAP7_75t_R g1242 ( 
.A(n_626),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_627),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_899),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_899),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_641),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_641),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_629),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_944),
.B(n_4),
.Y(n_1249)
);

CKINVDCx14_ASAP7_75t_R g1250 ( 
.A(n_638),
.Y(n_1250)
);

INVx3_ASAP7_75t_L g1251 ( 
.A(n_727),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_641),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_630),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1057),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_695),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_633),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_635),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_1045),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1057),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_637),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1057),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_639),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_642),
.Y(n_1263)
);

BUFx5_ASAP7_75t_L g1264 ( 
.A(n_632),
.Y(n_1264)
);

INVxp67_ASAP7_75t_SL g1265 ( 
.A(n_632),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_670),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_670),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_628),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_628),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_670),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_645),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_647),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_648),
.Y(n_1273)
);

BUFx5_ASAP7_75t_L g1274 ( 
.A(n_807),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_709),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_649),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_724),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_709),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1045),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_727),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_709),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_650),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_814),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_814),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_652),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_814),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_922),
.Y(n_1287)
);

INVx2_ASAP7_75t_L g1288 ( 
.A(n_944),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_922),
.Y(n_1289)
);

CKINVDCx5p33_ASAP7_75t_R g1290 ( 
.A(n_653),
.Y(n_1290)
);

CKINVDCx20_ASAP7_75t_R g1291 ( 
.A(n_724),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_638),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_922),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_944),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_654),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_727),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_885),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_655),
.Y(n_1298)
);

BUFx6f_ASAP7_75t_L g1299 ( 
.A(n_727),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_966),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_966),
.Y(n_1301)
);

CKINVDCx16_ASAP7_75t_R g1302 ( 
.A(n_638),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_727),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_656),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_659),
.Y(n_1305)
);

CKINVDCx16_ASAP7_75t_R g1306 ( 
.A(n_689),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_820),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_660),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_661),
.Y(n_1309)
);

HB1xp67_ASAP7_75t_L g1310 ( 
.A(n_885),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_664),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_966),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_807),
.Y(n_1313)
);

INVxp67_ASAP7_75t_SL g1314 ( 
.A(n_910),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_944),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_667),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_910),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_671),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_689),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_677),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_678),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_682),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1008),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1008),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_820),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_665),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_665),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_665),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_684),
.Y(n_1329)
);

NOR2xp67_ASAP7_75t_L g1330 ( 
.A(n_651),
.B(n_5),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_666),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_944),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_666),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_666),
.Y(n_1334)
);

CKINVDCx5p33_ASAP7_75t_R g1335 ( 
.A(n_692),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_681),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_702),
.Y(n_1337)
);

BUFx8_ASAP7_75t_SL g1338 ( 
.A(n_951),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_681),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_681),
.Y(n_1340)
);

CKINVDCx16_ASAP7_75t_R g1341 ( 
.A(n_689),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_693),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_697),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_944),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_822),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_703),
.Y(n_1346)
);

CKINVDCx14_ASAP7_75t_R g1347 ( 
.A(n_689),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_749),
.Y(n_1348)
);

INVxp67_ASAP7_75t_L g1349 ( 
.A(n_1077),
.Y(n_1349)
);

BUFx3_ASAP7_75t_L g1350 ( 
.A(n_944),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_749),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_749),
.Y(n_1352)
);

BUFx3_ASAP7_75t_L g1353 ( 
.A(n_944),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_705),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_651),
.B(n_5),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_777),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_944),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_777),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_SL g1359 ( 
.A(n_668),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_777),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_707),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_710),
.Y(n_1362)
);

CKINVDCx16_ASAP7_75t_R g1363 ( 
.A(n_789),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_785),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_712),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_785),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_716),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_722),
.Y(n_1368)
);

CKINVDCx16_ASAP7_75t_R g1369 ( 
.A(n_789),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_785),
.Y(n_1370)
);

BUFx8_ASAP7_75t_SL g1371 ( 
.A(n_951),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_789),
.Y(n_1372)
);

OR2x2_ASAP7_75t_L g1373 ( 
.A(n_791),
.B(n_6),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_944),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_873),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_791),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_791),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_723),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_725),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_726),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_753),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_947),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_729),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_829),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_829),
.Y(n_1385)
);

INVx1_ASAP7_75t_SL g1386 ( 
.A(n_780),
.Y(n_1386)
);

CKINVDCx20_ASAP7_75t_R g1387 ( 
.A(n_794),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_846),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_829),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_1077),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_730),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_853),
.Y(n_1392)
);

CKINVDCx20_ASAP7_75t_R g1393 ( 
.A(n_865),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_947),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_839),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_732),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_839),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_839),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_947),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_868),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_733),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_739),
.Y(n_1402)
);

BUFx5_ASAP7_75t_L g1403 ( 
.A(n_607),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_740),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_868),
.Y(n_1405)
);

BUFx6f_ASAP7_75t_L g1406 ( 
.A(n_727),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_868),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1006),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_947),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1006),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1006),
.Y(n_1411)
);

INVx1_ASAP7_75t_SL g1412 ( 
.A(n_866),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1025),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1025),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_880),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1025),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1036),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1036),
.Y(n_1418)
);

CKINVDCx16_ASAP7_75t_R g1419 ( 
.A(n_789),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_741),
.Y(n_1420)
);

NOR2xp67_ASAP7_75t_L g1421 ( 
.A(n_1086),
.B(n_6),
.Y(n_1421)
);

BUFx10_ASAP7_75t_L g1422 ( 
.A(n_736),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1086),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1086),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_882),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1102),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1102),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1102),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_714),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_607),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1122),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_742),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_609),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_744),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1122),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_745),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_886),
.Y(n_1437)
);

BUFx3_ASAP7_75t_L g1438 ( 
.A(n_947),
.Y(n_1438)
);

BUFx3_ASAP7_75t_L g1439 ( 
.A(n_947),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_746),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_747),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_750),
.Y(n_1442)
);

BUFx10_ASAP7_75t_L g1443 ( 
.A(n_736),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_609),
.Y(n_1444)
);

BUFx8_ASAP7_75t_SL g1445 ( 
.A(n_931),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_897),
.Y(n_1446)
);

INVx1_ASAP7_75t_SL g1447 ( 
.A(n_900),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_912),
.Y(n_1448)
);

BUFx2_ASAP7_75t_L g1449 ( 
.A(n_737),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_917),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_751),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_803),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_757),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_758),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_610),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_947),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_610),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_850),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_760),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_761),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_762),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_919),
.Y(n_1462)
);

BUFx10_ASAP7_75t_L g1463 ( 
.A(n_736),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_924),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_736),
.Y(n_1465)
);

BUFx2_ASAP7_75t_L g1466 ( 
.A(n_979),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_763),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_615),
.Y(n_1468)
);

INVxp67_ASAP7_75t_L g1469 ( 
.A(n_934),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_764),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_947),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_615),
.Y(n_1472)
);

CKINVDCx5p33_ASAP7_75t_R g1473 ( 
.A(n_765),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_947),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_617),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_766),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_768),
.Y(n_1477)
);

INVxp67_ASAP7_75t_L g1478 ( 
.A(n_934),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_617),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_620),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_770),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_947),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_736),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_736),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_620),
.B(n_7),
.Y(n_1485)
);

INVxp67_ASAP7_75t_L g1486 ( 
.A(n_1109),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1109),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_625),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_625),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_634),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_634),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_771),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_636),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_773),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_774),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_636),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_646),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_775),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_759),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_646),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_657),
.Y(n_1501)
);

BUFx6f_ASAP7_75t_L g1502 ( 
.A(n_759),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_776),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_915),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_657),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_658),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_779),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_658),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_663),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_782),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_759),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_663),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_783),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_759),
.Y(n_1514)
);

BUFx2_ASAP7_75t_L g1515 ( 
.A(n_854),
.Y(n_1515)
);

BUFx6f_ASAP7_75t_L g1516 ( 
.A(n_759),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_786),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_787),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_669),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_669),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_673),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_788),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_673),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_674),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_674),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_675),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_675),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_676),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_804),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_676),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_790),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_679),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_679),
.Y(n_1533)
);

INVxp67_ASAP7_75t_SL g1534 ( 
.A(n_804),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_680),
.Y(n_1535)
);

CKINVDCx20_ASAP7_75t_R g1536 ( 
.A(n_982),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_680),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_798),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1016),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_683),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_683),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_804),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_799),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_804),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_685),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_685),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_802),
.B(n_851),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_800),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_805),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_815),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_686),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_816),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_804),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_817),
.Y(n_1554)
);

CKINVDCx20_ASAP7_75t_R g1555 ( 
.A(n_1021),
.Y(n_1555)
);

CKINVDCx20_ASAP7_75t_R g1556 ( 
.A(n_1055),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_686),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_687),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_687),
.Y(n_1559)
);

INVxp67_ASAP7_75t_L g1560 ( 
.A(n_915),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_690),
.Y(n_1561)
);

BUFx6f_ASAP7_75t_L g1562 ( 
.A(n_804),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_690),
.Y(n_1563)
);

XOR2xp5_ASAP7_75t_L g1564 ( 
.A(n_907),
.B(n_7),
.Y(n_1564)
);

NOR2xp67_ASAP7_75t_L g1565 ( 
.A(n_691),
.B(n_7),
.Y(n_1565)
);

CKINVDCx5p33_ASAP7_75t_R g1566 ( 
.A(n_825),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_691),
.Y(n_1567)
);

NOR2xp67_ASAP7_75t_L g1568 ( 
.A(n_696),
.B(n_8),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_827),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_828),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_696),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_818),
.Y(n_1572)
);

INVxp67_ASAP7_75t_L g1573 ( 
.A(n_1078),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_698),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_698),
.Y(n_1575)
);

INVxp67_ASAP7_75t_L g1576 ( 
.A(n_1219),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1133),
.Y(n_1577)
);

BUFx2_ASAP7_75t_L g1578 ( 
.A(n_1175),
.Y(n_1578)
);

INVxp33_ASAP7_75t_L g1579 ( 
.A(n_1174),
.Y(n_1579)
);

INVxp33_ASAP7_75t_SL g1580 ( 
.A(n_1160),
.Y(n_1580)
);

BUFx6f_ASAP7_75t_L g1581 ( 
.A(n_1162),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1359),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1132),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1134),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_1168),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_1160),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1137),
.Y(n_1587)
);

CKINVDCx20_ASAP7_75t_R g1588 ( 
.A(n_1187),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1130),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1140),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1165),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1142),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1143),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1149),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1266),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1188),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1267),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1130),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1270),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_1161),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1201),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1349),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_1161),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1275),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1278),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1281),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1283),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1284),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1286),
.Y(n_1609)
);

CKINVDCx20_ASAP7_75t_R g1610 ( 
.A(n_1268),
.Y(n_1610)
);

CKINVDCx20_ASAP7_75t_R g1611 ( 
.A(n_1269),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1170),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1251),
.Y(n_1613)
);

CKINVDCx20_ASAP7_75t_R g1614 ( 
.A(n_1277),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1287),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1289),
.Y(n_1616)
);

INVxp33_ASAP7_75t_L g1617 ( 
.A(n_1174),
.Y(n_1617)
);

INVxp33_ASAP7_75t_SL g1618 ( 
.A(n_1170),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1293),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1291),
.Y(n_1620)
);

INVxp67_ASAP7_75t_SL g1621 ( 
.A(n_1390),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1300),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1301),
.Y(n_1623)
);

BUFx2_ASAP7_75t_SL g1624 ( 
.A(n_1547),
.Y(n_1624)
);

INVxp67_ASAP7_75t_SL g1625 ( 
.A(n_1135),
.Y(n_1625)
);

INVxp67_ASAP7_75t_SL g1626 ( 
.A(n_1135),
.Y(n_1626)
);

CKINVDCx5p33_ASAP7_75t_R g1627 ( 
.A(n_1173),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1312),
.Y(n_1628)
);

CKINVDCx16_ASAP7_75t_R g1629 ( 
.A(n_1302),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1150),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_1307),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1151),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1154),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1173),
.Y(n_1634)
);

CKINVDCx14_ASAP7_75t_R g1635 ( 
.A(n_1204),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1250),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1347),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1155),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1157),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1158),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1169),
.Y(n_1641)
);

INVxp67_ASAP7_75t_L g1642 ( 
.A(n_1449),
.Y(n_1642)
);

CKINVDCx5p33_ASAP7_75t_R g1643 ( 
.A(n_1338),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1164),
.Y(n_1644)
);

INVxp33_ASAP7_75t_L g1645 ( 
.A(n_1345),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1166),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1371),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1445),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1167),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_1211),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1171),
.Y(n_1651)
);

INVxp33_ASAP7_75t_L g1652 ( 
.A(n_1375),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1169),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1172),
.Y(n_1654)
);

BUFx2_ASAP7_75t_L g1655 ( 
.A(n_1175),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1176),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1177),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1178),
.Y(n_1658)
);

BUFx6f_ASAP7_75t_L g1659 ( 
.A(n_1162),
.Y(n_1659)
);

INVxp33_ASAP7_75t_L g1660 ( 
.A(n_1466),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1180),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1181),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1325),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1183),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1184),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1186),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1189),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1193),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1182),
.Y(n_1669)
);

CKINVDCx20_ASAP7_75t_R g1670 ( 
.A(n_1381),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_1255),
.Y(n_1671)
);

CKINVDCx5p33_ASAP7_75t_R g1672 ( 
.A(n_1337),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1197),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1346),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1200),
.Y(n_1675)
);

CKINVDCx16_ASAP7_75t_R g1676 ( 
.A(n_1306),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1203),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1182),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1206),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1207),
.Y(n_1680)
);

CKINVDCx16_ASAP7_75t_R g1681 ( 
.A(n_1341),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1213),
.Y(n_1682)
);

INVxp33_ASAP7_75t_L g1683 ( 
.A(n_1429),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1215),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1218),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1221),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1222),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1223),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1129),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1249),
.Y(n_1690)
);

INVxp33_ASAP7_75t_L g1691 ( 
.A(n_1458),
.Y(n_1691)
);

CKINVDCx20_ASAP7_75t_R g1692 ( 
.A(n_1387),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1265),
.Y(n_1693)
);

INVxp67_ASAP7_75t_SL g1694 ( 
.A(n_1208),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1386),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1314),
.Y(n_1696)
);

INVxp33_ASAP7_75t_SL g1697 ( 
.A(n_1123),
.Y(n_1697)
);

CKINVDCx5p33_ASAP7_75t_R g1698 ( 
.A(n_1392),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1125),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1127),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1534),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1542),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1412),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1430),
.Y(n_1704)
);

INVxp67_ASAP7_75t_SL g1705 ( 
.A(n_1208),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1431),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1251),
.Y(n_1707)
);

CKINVDCx20_ASAP7_75t_R g1708 ( 
.A(n_1388),
.Y(n_1708)
);

CKINVDCx5p33_ASAP7_75t_R g1709 ( 
.A(n_1447),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1433),
.Y(n_1710)
);

INVxp67_ASAP7_75t_SL g1711 ( 
.A(n_1504),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1435),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_1393),
.Y(n_1713)
);

INVxp33_ASAP7_75t_SL g1714 ( 
.A(n_1123),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1128),
.Y(n_1715)
);

CKINVDCx5p33_ASAP7_75t_R g1716 ( 
.A(n_1128),
.Y(n_1716)
);

INVxp33_ASAP7_75t_SL g1717 ( 
.A(n_1146),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1444),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_1415),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1455),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1425),
.Y(n_1721)
);

INVxp67_ASAP7_75t_L g1722 ( 
.A(n_1449),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1437),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1446),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1457),
.Y(n_1725)
);

BUFx2_ASAP7_75t_SL g1726 ( 
.A(n_1547),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1468),
.Y(n_1727)
);

CKINVDCx16_ASAP7_75t_R g1728 ( 
.A(n_1363),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1472),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1475),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1479),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1480),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1488),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1489),
.Y(n_1734)
);

CKINVDCx20_ASAP7_75t_R g1735 ( 
.A(n_1448),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1490),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1450),
.Y(n_1737)
);

INVxp67_ASAP7_75t_SL g1738 ( 
.A(n_1560),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1491),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1462),
.Y(n_1740)
);

INVxp67_ASAP7_75t_SL g1741 ( 
.A(n_1573),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1493),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1496),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1497),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1464),
.Y(n_1745)
);

INVxp33_ASAP7_75t_SL g1746 ( 
.A(n_1146),
.Y(n_1746)
);

BUFx3_ASAP7_75t_L g1747 ( 
.A(n_1228),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1185),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1500),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1501),
.Y(n_1750)
);

BUFx2_ASAP7_75t_L g1751 ( 
.A(n_1185),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1505),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1452),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1506),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1508),
.Y(n_1755)
);

BUFx2_ASAP7_75t_L g1756 ( 
.A(n_1190),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1509),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1512),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1152),
.Y(n_1759)
);

CKINVDCx5p33_ASAP7_75t_R g1760 ( 
.A(n_1152),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1519),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1520),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1521),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1523),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1524),
.Y(n_1765)
);

INVxp67_ASAP7_75t_SL g1766 ( 
.A(n_1350),
.Y(n_1766)
);

INVxp33_ASAP7_75t_SL g1767 ( 
.A(n_1196),
.Y(n_1767)
);

INVxp67_ASAP7_75t_SL g1768 ( 
.A(n_1353),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1525),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1526),
.Y(n_1770)
);

CKINVDCx5p33_ASAP7_75t_R g1771 ( 
.A(n_1196),
.Y(n_1771)
);

CKINVDCx5p33_ASAP7_75t_R g1772 ( 
.A(n_1198),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1527),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1528),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1530),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1532),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1533),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1535),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1537),
.Y(n_1779)
);

INVxp33_ASAP7_75t_SL g1780 ( 
.A(n_1198),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1251),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1162),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1199),
.Y(n_1783)
);

INVxp33_ASAP7_75t_SL g1784 ( 
.A(n_1199),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1209),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1540),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1541),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1209),
.Y(n_1788)
);

BUFx2_ASAP7_75t_L g1789 ( 
.A(n_1190),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1545),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_1216),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1228),
.Y(n_1792)
);

INVxp67_ASAP7_75t_SL g1793 ( 
.A(n_1357),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1546),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1452),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1216),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_1536),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1511),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1551),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1557),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1162),
.Y(n_1801)
);

CKINVDCx14_ASAP7_75t_R g1802 ( 
.A(n_1194),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1558),
.Y(n_1803)
);

CKINVDCx20_ASAP7_75t_R g1804 ( 
.A(n_1539),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1511),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1559),
.Y(n_1806)
);

CKINVDCx5p33_ASAP7_75t_R g1807 ( 
.A(n_1224),
.Y(n_1807)
);

CKINVDCx5p33_ASAP7_75t_R g1808 ( 
.A(n_1224),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1511),
.Y(n_1809)
);

INVx1_ASAP7_75t_SL g1810 ( 
.A(n_1555),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1515),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1229),
.Y(n_1812)
);

INVxp33_ASAP7_75t_L g1813 ( 
.A(n_1297),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1561),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1194),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1563),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1567),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1571),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1574),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1575),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1229),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1313),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1230),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1195),
.Y(n_1824)
);

CKINVDCx5p33_ASAP7_75t_R g1825 ( 
.A(n_1230),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1317),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1323),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1324),
.Y(n_1828)
);

CKINVDCx5p33_ASAP7_75t_R g1829 ( 
.A(n_1232),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1136),
.Y(n_1830)
);

CKINVDCx20_ASAP7_75t_R g1831 ( 
.A(n_1556),
.Y(n_1831)
);

INVxp33_ASAP7_75t_SL g1832 ( 
.A(n_1232),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1136),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1227),
.Y(n_1834)
);

CKINVDCx20_ASAP7_75t_R g1835 ( 
.A(n_1369),
.Y(n_1835)
);

CKINVDCx20_ASAP7_75t_R g1836 ( 
.A(n_1419),
.Y(n_1836)
);

BUFx6f_ASAP7_75t_L g1837 ( 
.A(n_1162),
.Y(n_1837)
);

CKINVDCx5p33_ASAP7_75t_R g1838 ( 
.A(n_1235),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1233),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1234),
.Y(n_1840)
);

INVxp67_ASAP7_75t_L g1841 ( 
.A(n_1124),
.Y(n_1841)
);

BUFx2_ASAP7_75t_SL g1842 ( 
.A(n_1292),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1237),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1357),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1239),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1241),
.Y(n_1846)
);

INVxp33_ASAP7_75t_SL g1847 ( 
.A(n_1235),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1244),
.Y(n_1848)
);

INVxp33_ASAP7_75t_L g1849 ( 
.A(n_1310),
.Y(n_1849)
);

CKINVDCx16_ASAP7_75t_R g1850 ( 
.A(n_1212),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1245),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1236),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1264),
.Y(n_1853)
);

CKINVDCx20_ASAP7_75t_R g1854 ( 
.A(n_1195),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1264),
.Y(n_1855)
);

INVxp67_ASAP7_75t_SL g1856 ( 
.A(n_1438),
.Y(n_1856)
);

INVxp33_ASAP7_75t_SL g1857 ( 
.A(n_1236),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1242),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1242),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1264),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1243),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1243),
.Y(n_1862)
);

CKINVDCx20_ASAP7_75t_R g1863 ( 
.A(n_1248),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1264),
.Y(n_1864)
);

INVxp33_ASAP7_75t_SL g1865 ( 
.A(n_1248),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1228),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1253),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1264),
.Y(n_1868)
);

CKINVDCx20_ASAP7_75t_R g1869 ( 
.A(n_1253),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1264),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1256),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1264),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1264),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1439),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1274),
.Y(n_1875)
);

INVxp67_ASAP7_75t_L g1876 ( 
.A(n_1159),
.Y(n_1876)
);

INVxp67_ASAP7_75t_SL g1877 ( 
.A(n_1439),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1256),
.Y(n_1878)
);

CKINVDCx5p33_ASAP7_75t_R g1879 ( 
.A(n_1257),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1274),
.Y(n_1880)
);

CKINVDCx20_ASAP7_75t_R g1881 ( 
.A(n_1257),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1274),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_1260),
.Y(n_1883)
);

INVxp67_ASAP7_75t_SL g1884 ( 
.A(n_1456),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1274),
.Y(n_1885)
);

INVxp67_ASAP7_75t_L g1886 ( 
.A(n_1205),
.Y(n_1886)
);

CKINVDCx20_ASAP7_75t_R g1887 ( 
.A(n_1260),
.Y(n_1887)
);

INVxp33_ASAP7_75t_SL g1888 ( 
.A(n_1262),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1192),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1212),
.Y(n_1890)
);

INVxp67_ASAP7_75t_SL g1891 ( 
.A(n_1456),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1274),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1274),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1274),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1262),
.Y(n_1895)
);

INVxp33_ASAP7_75t_SL g1896 ( 
.A(n_1263),
.Y(n_1896)
);

CKINVDCx20_ASAP7_75t_R g1897 ( 
.A(n_1263),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1271),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1271),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1272),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1246),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1247),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1252),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1292),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1254),
.Y(n_1905)
);

CKINVDCx20_ASAP7_75t_R g1906 ( 
.A(n_1272),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1259),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1261),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1192),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1326),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1327),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1273),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1192),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1328),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1331),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1333),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1273),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_1276),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1334),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1192),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1276),
.Y(n_1921)
);

INVxp33_ASAP7_75t_SL g1922 ( 
.A(n_1282),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1282),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1336),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1339),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_1285),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1340),
.Y(n_1927)
);

CKINVDCx16_ASAP7_75t_R g1928 ( 
.A(n_1319),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1348),
.Y(n_1929)
);

INVxp33_ASAP7_75t_SL g1930 ( 
.A(n_1285),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1351),
.Y(n_1931)
);

CKINVDCx16_ASAP7_75t_R g1932 ( 
.A(n_1319),
.Y(n_1932)
);

CKINVDCx20_ASAP7_75t_R g1933 ( 
.A(n_1290),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1192),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1290),
.Y(n_1935)
);

CKINVDCx5p33_ASAP7_75t_R g1936 ( 
.A(n_1295),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1352),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1372),
.Y(n_1938)
);

INVxp33_ASAP7_75t_SL g1939 ( 
.A(n_1295),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1356),
.Y(n_1940)
);

CKINVDCx20_ASAP7_75t_R g1941 ( 
.A(n_1298),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1298),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1358),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1360),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1613),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1613),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1928),
.B(n_1304),
.Y(n_1947)
);

OAI22x1_ASAP7_75t_L g1948 ( 
.A1(n_1890),
.A2(n_1564),
.B1(n_1220),
.B2(n_1238),
.Y(n_1948)
);

AND2x4_ASAP7_75t_L g1949 ( 
.A(n_1693),
.B(n_1372),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1707),
.Y(n_1950)
);

AND2x2_ASAP7_75t_SL g1951 ( 
.A(n_1932),
.B(n_1148),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1707),
.Y(n_1952)
);

AND2x4_ASAP7_75t_L g1953 ( 
.A(n_1696),
.B(n_1131),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1690),
.B(n_1141),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1624),
.B(n_1191),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1701),
.B(n_1148),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1702),
.B(n_1148),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1781),
.Y(n_1958)
);

OA21x2_ASAP7_75t_L g1959 ( 
.A1(n_1889),
.A2(n_1138),
.B(n_1126),
.Y(n_1959)
);

BUFx2_ASAP7_75t_L g1960 ( 
.A(n_1850),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1781),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1841),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1798),
.Y(n_1963)
);

NOR2x1_ASAP7_75t_L g1964 ( 
.A(n_1726),
.B(n_1179),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_L g1965 ( 
.A(n_1842),
.B(n_1179),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1602),
.B(n_1403),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1589),
.Y(n_1967)
);

OA21x2_ASAP7_75t_L g1968 ( 
.A1(n_1889),
.A2(n_1138),
.B(n_1126),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1621),
.B(n_1711),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1798),
.Y(n_1970)
);

XNOR2x2_ASAP7_75t_L g1971 ( 
.A(n_1723),
.B(n_1485),
.Y(n_1971)
);

BUFx3_ASAP7_75t_L g1972 ( 
.A(n_1589),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1738),
.B(n_1403),
.Y(n_1973)
);

INVx6_ASAP7_75t_L g1974 ( 
.A(n_1598),
.Y(n_1974)
);

INVx2_ASAP7_75t_L g1975 ( 
.A(n_1805),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1805),
.Y(n_1976)
);

HB1xp67_ASAP7_75t_L g1977 ( 
.A(n_1591),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1809),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1809),
.Y(n_1979)
);

BUFx6f_ASAP7_75t_L g1980 ( 
.A(n_1598),
.Y(n_1980)
);

BUFx6f_ASAP7_75t_L g1981 ( 
.A(n_1581),
.Y(n_1981)
);

BUFx12f_ASAP7_75t_L g1982 ( 
.A(n_1582),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1577),
.Y(n_1983)
);

BUFx3_ASAP7_75t_L g1984 ( 
.A(n_1747),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1581),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1581),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1584),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1587),
.Y(n_1988)
);

BUFx6f_ASAP7_75t_L g1989 ( 
.A(n_1581),
.Y(n_1989)
);

BUFx3_ASAP7_75t_L g1990 ( 
.A(n_1747),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_L g1991 ( 
.A(n_1715),
.B(n_1403),
.Y(n_1991)
);

INVx3_ASAP7_75t_L g1992 ( 
.A(n_1659),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1590),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1592),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1741),
.B(n_1403),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1834),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1593),
.Y(n_1997)
);

BUFx3_ASAP7_75t_L g1998 ( 
.A(n_1792),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1904),
.B(n_1403),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1659),
.Y(n_2000)
);

AND2x6_ASAP7_75t_L g2001 ( 
.A(n_1689),
.B(n_1355),
.Y(n_2001)
);

INVx5_ASAP7_75t_L g2002 ( 
.A(n_1659),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1839),
.Y(n_2003)
);

NOR2xp33_ASAP7_75t_L g2004 ( 
.A(n_1938),
.B(n_1304),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1594),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1840),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1843),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1901),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1845),
.Y(n_2009)
);

INVx3_ASAP7_75t_L g2010 ( 
.A(n_1782),
.Y(n_2010)
);

BUFx2_ASAP7_75t_L g2011 ( 
.A(n_1876),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1902),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1846),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1848),
.Y(n_2014)
);

AND2x6_ASAP7_75t_L g2015 ( 
.A(n_1699),
.B(n_699),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1697),
.B(n_1305),
.Y(n_2016)
);

AOI22x1_ASAP7_75t_SL g2017 ( 
.A1(n_1643),
.A2(n_967),
.B1(n_978),
.B2(n_909),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1596),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1642),
.A2(n_1478),
.B1(n_1486),
.B2(n_1469),
.Y(n_2019)
);

INVx6_ASAP7_75t_L g2020 ( 
.A(n_1866),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1851),
.Y(n_2021)
);

INVx2_ASAP7_75t_L g2022 ( 
.A(n_1909),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1903),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1905),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1704),
.B(n_1487),
.Y(n_2025)
);

AND2x4_ASAP7_75t_L g2026 ( 
.A(n_1830),
.B(n_1485),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1833),
.B(n_1373),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1907),
.Y(n_2028)
);

INVx3_ASAP7_75t_L g2029 ( 
.A(n_1782),
.Y(n_2029)
);

NOR2x1_ASAP7_75t_L g2030 ( 
.A(n_1900),
.B(n_1217),
.Y(n_2030)
);

INVxp33_ASAP7_75t_SL g2031 ( 
.A(n_1771),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1909),
.Y(n_2032)
);

CKINVDCx11_ASAP7_75t_R g2033 ( 
.A(n_1863),
.Y(n_2033)
);

INVx6_ASAP7_75t_L g2034 ( 
.A(n_1801),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1722),
.A2(n_1305),
.B1(n_1309),
.B2(n_1308),
.Y(n_2035)
);

OA21x2_ASAP7_75t_L g2036 ( 
.A1(n_1913),
.A2(n_1147),
.B(n_1145),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1697),
.B(n_1714),
.Y(n_2037)
);

BUFx12f_ASAP7_75t_L g2038 ( 
.A(n_1582),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1913),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1714),
.B(n_1308),
.Y(n_2040)
);

INVx4_ASAP7_75t_L g2041 ( 
.A(n_1801),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1908),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1910),
.Y(n_2043)
);

INVx3_ASAP7_75t_L g2044 ( 
.A(n_1801),
.Y(n_2044)
);

BUFx8_ASAP7_75t_SL g2045 ( 
.A(n_1670),
.Y(n_2045)
);

OAI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1753),
.A2(n_1231),
.B1(n_1258),
.B2(n_1139),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1944),
.Y(n_2047)
);

HB1xp67_ASAP7_75t_L g2048 ( 
.A(n_1886),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1943),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1920),
.Y(n_2050)
);

BUFx3_ASAP7_75t_L g2051 ( 
.A(n_1700),
.Y(n_2051)
);

AND2x6_ASAP7_75t_L g2052 ( 
.A(n_1630),
.B(n_699),
.Y(n_2052)
);

BUFx6f_ASAP7_75t_L g2053 ( 
.A(n_1837),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1911),
.Y(n_2054)
);

BUFx6f_ASAP7_75t_L g2055 ( 
.A(n_1837),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1795),
.Y(n_2056)
);

BUFx3_ASAP7_75t_L g2057 ( 
.A(n_1632),
.Y(n_2057)
);

AND2x6_ASAP7_75t_L g2058 ( 
.A(n_1633),
.B(n_700),
.Y(n_2058)
);

BUFx6f_ASAP7_75t_L g2059 ( 
.A(n_1920),
.Y(n_2059)
);

OAI22x1_ASAP7_75t_R g2060 ( 
.A1(n_1863),
.A2(n_1311),
.B1(n_1316),
.B2(n_1309),
.Y(n_2060)
);

BUFx3_ASAP7_75t_L g2061 ( 
.A(n_1638),
.Y(n_2061)
);

INVx3_ASAP7_75t_L g2062 ( 
.A(n_1934),
.Y(n_2062)
);

HB1xp67_ASAP7_75t_L g2063 ( 
.A(n_1811),
.Y(n_2063)
);

INVx3_ASAP7_75t_L g2064 ( 
.A(n_1934),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1914),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1853),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_1855),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1915),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1916),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_1919),
.Y(n_2070)
);

BUFx6f_ASAP7_75t_L g2071 ( 
.A(n_1860),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1924),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_SL g2073 ( 
.A(n_1862),
.B(n_1942),
.Y(n_2073)
);

INVx2_ASAP7_75t_L g2074 ( 
.A(n_1864),
.Y(n_2074)
);

AND2x6_ASAP7_75t_L g2075 ( 
.A(n_1639),
.B(n_700),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1640),
.B(n_1373),
.Y(n_2076)
);

INVx3_ASAP7_75t_L g2077 ( 
.A(n_1868),
.Y(n_2077)
);

BUFx6f_ASAP7_75t_L g2078 ( 
.A(n_1870),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1925),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1706),
.B(n_1364),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1710),
.B(n_1366),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_1578),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1927),
.Y(n_2083)
);

NOR2xp33_ASAP7_75t_L g2084 ( 
.A(n_1717),
.B(n_1311),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_1929),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1872),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1873),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_1875),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1880),
.Y(n_2089)
);

CKINVDCx11_ASAP7_75t_R g2090 ( 
.A(n_1869),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_1712),
.B(n_1370),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1882),
.Y(n_2092)
);

BUFx2_ASAP7_75t_L g2093 ( 
.A(n_1655),
.Y(n_2093)
);

AND2x6_ASAP7_75t_L g2094 ( 
.A(n_1644),
.B(n_701),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_1931),
.Y(n_2095)
);

OAI22x1_ASAP7_75t_SL g2096 ( 
.A1(n_1643),
.A2(n_998),
.B1(n_1012),
.B2(n_1007),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_1678),
.Y(n_2097)
);

BUFx6f_ASAP7_75t_L g2098 ( 
.A(n_1885),
.Y(n_2098)
);

INVx5_ASAP7_75t_L g2099 ( 
.A(n_1625),
.Y(n_2099)
);

BUFx6f_ASAP7_75t_L g2100 ( 
.A(n_1892),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_1767),
.A2(n_1318),
.B1(n_1320),
.B2(n_1316),
.Y(n_2101)
);

INVx5_ASAP7_75t_L g2102 ( 
.A(n_1626),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1893),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1937),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1940),
.Y(n_2105)
);

INVx2_ASAP7_75t_L g2106 ( 
.A(n_1894),
.Y(n_2106)
);

HB1xp67_ASAP7_75t_L g2107 ( 
.A(n_1650),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1646),
.Y(n_2108)
);

BUFx6f_ASAP7_75t_L g2109 ( 
.A(n_1649),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_1751),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1651),
.Y(n_2111)
);

INVx3_ASAP7_75t_L g2112 ( 
.A(n_1654),
.Y(n_2112)
);

INVx3_ASAP7_75t_L g2113 ( 
.A(n_1656),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1766),
.B(n_1318),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1647),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1657),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1715),
.B(n_1320),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1658),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1661),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_1662),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1664),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_1717),
.B(n_1321),
.Y(n_2122)
);

BUFx6f_ASAP7_75t_L g2123 ( 
.A(n_1665),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1666),
.Y(n_2124)
);

CKINVDCx5p33_ASAP7_75t_R g2125 ( 
.A(n_1647),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1667),
.Y(n_2126)
);

BUFx3_ASAP7_75t_L g2127 ( 
.A(n_1668),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1673),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1675),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1677),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1679),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_1680),
.Y(n_2132)
);

OAI21x1_ASAP7_75t_L g2133 ( 
.A1(n_1682),
.A2(n_1147),
.B(n_1145),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_SL g2134 ( 
.A(n_1716),
.B(n_1321),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1684),
.Y(n_2135)
);

AND2x6_ASAP7_75t_L g2136 ( 
.A(n_1685),
.B(n_1686),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1687),
.Y(n_2137)
);

OAI22xp5_ASAP7_75t_L g2138 ( 
.A1(n_1802),
.A2(n_1279),
.B1(n_1330),
.B2(n_1060),
.Y(n_2138)
);

CKINVDCx16_ASAP7_75t_R g2139 ( 
.A(n_1629),
.Y(n_2139)
);

BUFx3_ASAP7_75t_L g2140 ( 
.A(n_1688),
.Y(n_2140)
);

BUFx2_ASAP7_75t_L g2141 ( 
.A(n_1756),
.Y(n_2141)
);

OAI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_1716),
.A2(n_1117),
.B1(n_1033),
.B2(n_618),
.Y(n_2142)
);

AND2x6_ASAP7_75t_L g2143 ( 
.A(n_1718),
.B(n_701),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1595),
.Y(n_2144)
);

BUFx6f_ASAP7_75t_L g2145 ( 
.A(n_1822),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1720),
.B(n_1565),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1597),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1768),
.B(n_1322),
.Y(n_2148)
);

BUFx6f_ASAP7_75t_L g2149 ( 
.A(n_1826),
.Y(n_2149)
);

BUFx6f_ASAP7_75t_L g2150 ( 
.A(n_1827),
.Y(n_2150)
);

OA21x2_ASAP7_75t_L g2151 ( 
.A1(n_1828),
.A2(n_1156),
.B(n_1153),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1599),
.Y(n_2152)
);

INVx5_ASAP7_75t_L g2153 ( 
.A(n_1641),
.Y(n_2153)
);

BUFx6f_ASAP7_75t_L g2154 ( 
.A(n_1725),
.Y(n_2154)
);

NAND2xp33_ASAP7_75t_L g2155 ( 
.A(n_1759),
.B(n_818),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1604),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_1727),
.Y(n_2157)
);

AND2x2_ASAP7_75t_L g2158 ( 
.A(n_1729),
.B(n_1376),
.Y(n_2158)
);

INVxp67_ASAP7_75t_L g2159 ( 
.A(n_1650),
.Y(n_2159)
);

INVx2_ASAP7_75t_L g2160 ( 
.A(n_1605),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_1606),
.Y(n_2161)
);

OA21x2_ASAP7_75t_L g2162 ( 
.A1(n_1607),
.A2(n_1156),
.B(n_1153),
.Y(n_2162)
);

INVx3_ASAP7_75t_L g2163 ( 
.A(n_1608),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_1609),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1648),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_1746),
.B(n_1322),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1615),
.Y(n_2167)
);

INVx2_ASAP7_75t_SL g2168 ( 
.A(n_1583),
.Y(n_2168)
);

OA21x2_ASAP7_75t_L g2169 ( 
.A1(n_1616),
.A2(n_1226),
.B(n_1214),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1730),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1619),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1622),
.Y(n_2172)
);

INVx3_ASAP7_75t_L g2173 ( 
.A(n_1623),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_1671),
.Y(n_2174)
);

AND2x4_ASAP7_75t_L g2175 ( 
.A(n_1731),
.B(n_1568),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_1789),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1628),
.Y(n_2177)
);

AOI22xp5_ASAP7_75t_L g2178 ( 
.A1(n_1767),
.A2(n_1335),
.B1(n_1342),
.B2(n_1329),
.Y(n_2178)
);

AND2x2_ASAP7_75t_L g2179 ( 
.A(n_1732),
.B(n_1377),
.Y(n_2179)
);

INVx4_ASAP7_75t_L g2180 ( 
.A(n_1636),
.Y(n_2180)
);

AND2x4_ASAP7_75t_L g2181 ( 
.A(n_1733),
.B(n_1421),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1734),
.Y(n_2182)
);

OAI22x1_ASAP7_75t_L g2183 ( 
.A1(n_1771),
.A2(n_1202),
.B1(n_1163),
.B2(n_618),
.Y(n_2183)
);

AND2x6_ASAP7_75t_L g2184 ( 
.A(n_1736),
.B(n_708),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_1739),
.Y(n_2185)
);

OAI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_1759),
.A2(n_643),
.B1(n_644),
.B2(n_614),
.Y(n_2186)
);

INVx2_ASAP7_75t_L g2187 ( 
.A(n_1742),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1743),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1744),
.Y(n_2189)
);

NAND2xp5_ASAP7_75t_L g2190 ( 
.A(n_1793),
.B(n_1329),
.Y(n_2190)
);

BUFx6f_ASAP7_75t_L g2191 ( 
.A(n_1749),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1750),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_1752),
.Y(n_2193)
);

CKINVDCx5p33_ASAP7_75t_R g2194 ( 
.A(n_1648),
.Y(n_2194)
);

BUFx8_ASAP7_75t_L g2195 ( 
.A(n_1676),
.Y(n_2195)
);

NAND2xp33_ASAP7_75t_L g2196 ( 
.A(n_1760),
.B(n_818),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1671),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1754),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1755),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1844),
.B(n_1335),
.Y(n_2200)
);

INVx2_ASAP7_75t_L g2201 ( 
.A(n_1757),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1758),
.B(n_1384),
.Y(n_2202)
);

INVx2_ASAP7_75t_L g2203 ( 
.A(n_1761),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1762),
.Y(n_2204)
);

AND2x2_ASAP7_75t_SL g2205 ( 
.A(n_1681),
.B(n_708),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1763),
.Y(n_2206)
);

BUFx3_ASAP7_75t_L g2207 ( 
.A(n_1764),
.Y(n_2207)
);

AOI22xp5_ASAP7_75t_L g2208 ( 
.A1(n_1780),
.A2(n_1343),
.B1(n_1354),
.B2(n_1342),
.Y(n_2208)
);

INVxp33_ASAP7_75t_SL g2209 ( 
.A(n_1772),
.Y(n_2209)
);

AND2x4_ASAP7_75t_L g2210 ( 
.A(n_1765),
.B(n_1144),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1769),
.B(n_1770),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_1773),
.B(n_1385),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_1780),
.A2(n_1354),
.B1(n_1361),
.B2(n_1343),
.Y(n_2213)
);

OAI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_1760),
.A2(n_643),
.B1(n_644),
.B2(n_614),
.Y(n_2214)
);

AND2x2_ASAP7_75t_L g2215 ( 
.A(n_1774),
.B(n_1389),
.Y(n_2215)
);

AND2x6_ASAP7_75t_L g2216 ( 
.A(n_1775),
.B(n_711),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_1856),
.B(n_1361),
.Y(n_2217)
);

CKINVDCx11_ASAP7_75t_R g2218 ( 
.A(n_1869),
.Y(n_2218)
);

AND2x6_ASAP7_75t_L g2219 ( 
.A(n_1776),
.B(n_711),
.Y(n_2219)
);

INVx2_ASAP7_75t_SL g2220 ( 
.A(n_1583),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1777),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1874),
.B(n_1362),
.Y(n_2222)
);

INVx2_ASAP7_75t_L g2223 ( 
.A(n_1778),
.Y(n_2223)
);

BUFx6f_ASAP7_75t_L g2224 ( 
.A(n_1779),
.Y(n_2224)
);

NAND2xp5_ASAP7_75t_L g2225 ( 
.A(n_1877),
.B(n_1362),
.Y(n_2225)
);

INVx5_ASAP7_75t_L g2226 ( 
.A(n_1653),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1786),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_1787),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_1790),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1794),
.Y(n_2230)
);

INVx2_ASAP7_75t_L g2231 ( 
.A(n_1799),
.Y(n_2231)
);

INVx3_ASAP7_75t_L g2232 ( 
.A(n_1800),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_1884),
.B(n_1365),
.Y(n_2233)
);

BUFx6f_ASAP7_75t_L g2234 ( 
.A(n_1803),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1806),
.Y(n_2235)
);

CKINVDCx14_ASAP7_75t_R g2236 ( 
.A(n_1635),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_1814),
.Y(n_2237)
);

BUFx2_ASAP7_75t_L g2238 ( 
.A(n_1854),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1816),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_L g2240 ( 
.A(n_1746),
.B(n_1365),
.Y(n_2240)
);

OA21x2_ASAP7_75t_L g2241 ( 
.A1(n_1817),
.A2(n_1226),
.B(n_1214),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1818),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1724),
.Y(n_2243)
);

AND2x6_ASAP7_75t_L g2244 ( 
.A(n_1819),
.B(n_715),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1820),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1891),
.Y(n_2246)
);

AND2x4_ASAP7_75t_L g2247 ( 
.A(n_1576),
.B(n_1395),
.Y(n_2247)
);

BUFx6f_ASAP7_75t_L g2248 ( 
.A(n_1867),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_1694),
.B(n_1367),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_1871),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_1705),
.Y(n_2251)
);

OAI22x1_ASAP7_75t_R g2252 ( 
.A1(n_1881),
.A2(n_1368),
.B1(n_1378),
.B2(n_1367),
.Y(n_2252)
);

OAI21x1_ASAP7_75t_L g2253 ( 
.A1(n_1861),
.A2(n_1294),
.B(n_1288),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1585),
.Y(n_2254)
);

HB1xp67_ASAP7_75t_L g2255 ( 
.A(n_1695),
.Y(n_2255)
);

BUFx6f_ASAP7_75t_L g2256 ( 
.A(n_1878),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1585),
.B(n_1368),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1895),
.Y(n_2258)
);

AND2x4_ASAP7_75t_L g2259 ( 
.A(n_1669),
.B(n_1397),
.Y(n_2259)
);

INVx3_ASAP7_75t_L g2260 ( 
.A(n_1879),
.Y(n_2260)
);

BUFx2_ASAP7_75t_L g2261 ( 
.A(n_1854),
.Y(n_2261)
);

OAI22xp5_ASAP7_75t_SL g2262 ( 
.A1(n_1588),
.A2(n_1379),
.B1(n_1380),
.B2(n_1378),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1748),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1898),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_1918),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1815),
.Y(n_2266)
);

BUFx6f_ASAP7_75t_L g2267 ( 
.A(n_1921),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1824),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_1772),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1783),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1783),
.Y(n_2271)
);

BUFx6f_ASAP7_75t_L g2272 ( 
.A(n_1785),
.Y(n_2272)
);

OAI22xp5_ASAP7_75t_L g2273 ( 
.A1(n_1784),
.A2(n_752),
.B1(n_756),
.B2(n_748),
.Y(n_2273)
);

AND2x4_ASAP7_75t_L g2274 ( 
.A(n_1637),
.B(n_1398),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_1785),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1788),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_1683),
.B(n_1380),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_1637),
.B(n_1383),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_1788),
.Y(n_2279)
);

AND2x4_ASAP7_75t_L g2280 ( 
.A(n_1791),
.B(n_1400),
.Y(n_2280)
);

INVx2_ASAP7_75t_L g2281 ( 
.A(n_1791),
.Y(n_2281)
);

AND2x2_ASAP7_75t_SL g2282 ( 
.A(n_1728),
.B(n_818),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_1784),
.B(n_1383),
.Y(n_2283)
);

BUFx12f_ASAP7_75t_L g2284 ( 
.A(n_1586),
.Y(n_2284)
);

INVx3_ASAP7_75t_L g2285 ( 
.A(n_1796),
.Y(n_2285)
);

INVx2_ASAP7_75t_SL g2286 ( 
.A(n_1796),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1807),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_1807),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_1808),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_1808),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_1812),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_1812),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_1821),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1691),
.B(n_1405),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_1821),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1823),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_1823),
.Y(n_2297)
);

INVx2_ASAP7_75t_L g2298 ( 
.A(n_1825),
.Y(n_2298)
);

OA21x2_ASAP7_75t_L g2299 ( 
.A1(n_1825),
.A2(n_1294),
.B(n_1288),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_1829),
.Y(n_2300)
);

INVx4_ASAP7_75t_L g2301 ( 
.A(n_1829),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_1813),
.B(n_1407),
.Y(n_2302)
);

CKINVDCx6p67_ASAP7_75t_R g2303 ( 
.A(n_1835),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_1838),
.Y(n_2304)
);

AND2x2_ASAP7_75t_SL g2305 ( 
.A(n_1832),
.B(n_818),
.Y(n_2305)
);

BUFx6f_ASAP7_75t_L g2306 ( 
.A(n_1838),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1852),
.Y(n_2307)
);

AND2x6_ASAP7_75t_L g2308 ( 
.A(n_1810),
.B(n_715),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1852),
.Y(n_2309)
);

CKINVDCx5p33_ASAP7_75t_R g2310 ( 
.A(n_1737),
.Y(n_2310)
);

AOI22xp5_ASAP7_75t_SL g2311 ( 
.A1(n_1881),
.A2(n_1548),
.B1(n_1549),
.B2(n_1543),
.Y(n_2311)
);

NAND2xp5_ASAP7_75t_L g2312 ( 
.A(n_1832),
.B(n_1391),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1858),
.Y(n_2313)
);

CKINVDCx11_ASAP7_75t_R g2314 ( 
.A(n_1887),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_1858),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_1695),
.Y(n_2316)
);

BUFx6f_ASAP7_75t_L g2317 ( 
.A(n_1859),
.Y(n_2317)
);

NOR2xp33_ASAP7_75t_L g2318 ( 
.A(n_1847),
.B(n_1391),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1859),
.Y(n_2319)
);

NAND2xp5_ASAP7_75t_L g2320 ( 
.A(n_1847),
.B(n_1396),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1883),
.Y(n_2321)
);

BUFx8_ASAP7_75t_L g2322 ( 
.A(n_1580),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_1883),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_1899),
.Y(n_2324)
);

INVx2_ASAP7_75t_L g2325 ( 
.A(n_1899),
.Y(n_2325)
);

BUFx12f_ASAP7_75t_L g2326 ( 
.A(n_1600),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1857),
.B(n_1396),
.Y(n_2327)
);

CKINVDCx5p33_ASAP7_75t_R g2328 ( 
.A(n_1740),
.Y(n_2328)
);

BUFx6f_ASAP7_75t_L g2329 ( 
.A(n_1912),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1912),
.Y(n_2330)
);

INVx2_ASAP7_75t_L g2331 ( 
.A(n_1923),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1857),
.B(n_1401),
.Y(n_2332)
);

AND2x2_ASAP7_75t_L g2333 ( 
.A(n_1849),
.B(n_1408),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1923),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1865),
.B(n_1401),
.Y(n_2335)
);

INVx3_ASAP7_75t_L g2336 ( 
.A(n_1936),
.Y(n_2336)
);

INVx4_ASAP7_75t_L g2337 ( 
.A(n_1936),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_1672),
.B(n_1410),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_1865),
.B(n_1402),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_SL g2340 ( 
.A(n_1888),
.B(n_1402),
.Y(n_2340)
);

OA21x2_ASAP7_75t_L g2341 ( 
.A1(n_1698),
.A2(n_1332),
.B(n_1315),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_1674),
.Y(n_2342)
);

INVx2_ASAP7_75t_L g2343 ( 
.A(n_1698),
.Y(n_2343)
);

NOR2x1_ASAP7_75t_L g2344 ( 
.A(n_1887),
.B(n_1411),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_1888),
.B(n_1404),
.Y(n_2345)
);

AOI22xp5_ASAP7_75t_L g2346 ( 
.A1(n_1896),
.A2(n_1420),
.B1(n_1432),
.B2(n_1404),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_1896),
.B(n_1420),
.Y(n_2347)
);

BUFx2_ASAP7_75t_L g2348 ( 
.A(n_1897),
.Y(n_2348)
);

BUFx3_ASAP7_75t_L g2349 ( 
.A(n_1922),
.Y(n_2349)
);

NAND2xp5_ASAP7_75t_L g2350 ( 
.A(n_1922),
.B(n_1432),
.Y(n_2350)
);

NAND2xp33_ASAP7_75t_L g2351 ( 
.A(n_1600),
.B(n_818),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1930),
.Y(n_2352)
);

AND2x4_ASAP7_75t_L g2353 ( 
.A(n_1941),
.B(n_1413),
.Y(n_2353)
);

NAND2xp33_ASAP7_75t_L g2354 ( 
.A(n_1603),
.B(n_859),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_1930),
.Y(n_2355)
);

OA21x2_ASAP7_75t_L g2356 ( 
.A1(n_1703),
.A2(n_1332),
.B(n_1315),
.Y(n_2356)
);

OA22x2_ASAP7_75t_SL g2357 ( 
.A1(n_1939),
.A2(n_721),
.B1(n_734),
.B2(n_720),
.Y(n_2357)
);

BUFx2_ASAP7_75t_L g2358 ( 
.A(n_1897),
.Y(n_2358)
);

BUFx8_ASAP7_75t_L g2359 ( 
.A(n_1580),
.Y(n_2359)
);

OAI22x1_ASAP7_75t_L g2360 ( 
.A1(n_1703),
.A2(n_752),
.B1(n_756),
.B2(n_748),
.Y(n_2360)
);

INVx2_ASAP7_75t_L g2361 ( 
.A(n_1709),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_1709),
.Y(n_2362)
);

OAI22xp5_ASAP7_75t_L g2363 ( 
.A1(n_1939),
.A2(n_813),
.B1(n_824),
.B2(n_781),
.Y(n_2363)
);

AND2x2_ASAP7_75t_L g2364 ( 
.A(n_1645),
.B(n_1414),
.Y(n_2364)
);

BUFx3_ASAP7_75t_L g2365 ( 
.A(n_1618),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1618),
.B(n_1434),
.Y(n_2366)
);

AND2x2_ASAP7_75t_L g2367 ( 
.A(n_1652),
.B(n_1416),
.Y(n_2367)
);

CKINVDCx5p33_ASAP7_75t_R g2368 ( 
.A(n_2045),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_1946),
.Y(n_2369)
);

INVx2_ASAP7_75t_L g2370 ( 
.A(n_1945),
.Y(n_2370)
);

CKINVDCx5p33_ASAP7_75t_R g2371 ( 
.A(n_2165),
.Y(n_2371)
);

HB1xp67_ASAP7_75t_L g2372 ( 
.A(n_1960),
.Y(n_2372)
);

CKINVDCx5p33_ASAP7_75t_R g2373 ( 
.A(n_2165),
.Y(n_2373)
);

CKINVDCx5p33_ASAP7_75t_R g2374 ( 
.A(n_2194),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1955),
.B(n_1434),
.Y(n_2375)
);

INVxp67_ASAP7_75t_L g2376 ( 
.A(n_1962),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_1946),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_1963),
.Y(n_2378)
);

CKINVDCx5p33_ASAP7_75t_R g2379 ( 
.A(n_2194),
.Y(n_2379)
);

NOR2xp33_ASAP7_75t_L g2380 ( 
.A(n_2257),
.B(n_1660),
.Y(n_2380)
);

INVx2_ASAP7_75t_L g2381 ( 
.A(n_1945),
.Y(n_2381)
);

BUFx8_ASAP7_75t_L g2382 ( 
.A(n_1960),
.Y(n_2382)
);

NAND2xp5_ASAP7_75t_L g2383 ( 
.A(n_1955),
.B(n_1436),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_1963),
.Y(n_2384)
);

AOI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2305),
.A2(n_1440),
.B1(n_1441),
.B2(n_1436),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1950),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_2272),
.B(n_2275),
.Y(n_2387)
);

INVx2_ASAP7_75t_L g2388 ( 
.A(n_1950),
.Y(n_2388)
);

CKINVDCx5p33_ASAP7_75t_R g2389 ( 
.A(n_2115),
.Y(n_2389)
);

CKINVDCx20_ASAP7_75t_R g2390 ( 
.A(n_2033),
.Y(n_2390)
);

BUFx6f_ASAP7_75t_L g2391 ( 
.A(n_1967),
.Y(n_2391)
);

CKINVDCx5p33_ASAP7_75t_R g2392 ( 
.A(n_2115),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2168),
.B(n_1440),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1978),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2168),
.B(n_1441),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1978),
.Y(n_2396)
);

INVx3_ASAP7_75t_L g2397 ( 
.A(n_2162),
.Y(n_2397)
);

INVx1_ASAP7_75t_L g2398 ( 
.A(n_2144),
.Y(n_2398)
);

AND2x4_ASAP7_75t_L g2399 ( 
.A(n_2272),
.B(n_1906),
.Y(n_2399)
);

CKINVDCx5p33_ASAP7_75t_R g2400 ( 
.A(n_2125),
.Y(n_2400)
);

CKINVDCx5p33_ASAP7_75t_R g2401 ( 
.A(n_2125),
.Y(n_2401)
);

BUFx6f_ASAP7_75t_L g2402 ( 
.A(n_1967),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_1954),
.B(n_1442),
.Y(n_2403)
);

CKINVDCx5p33_ASAP7_75t_R g2404 ( 
.A(n_2243),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_1952),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2144),
.Y(n_2406)
);

INVx2_ASAP7_75t_L g2407 ( 
.A(n_1952),
.Y(n_2407)
);

BUFx6f_ASAP7_75t_L g2408 ( 
.A(n_1967),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2156),
.Y(n_2409)
);

CKINVDCx20_ASAP7_75t_R g2410 ( 
.A(n_2090),
.Y(n_2410)
);

CKINVDCx5p33_ASAP7_75t_R g2411 ( 
.A(n_2243),
.Y(n_2411)
);

OAI21x1_ASAP7_75t_L g2412 ( 
.A1(n_2133),
.A2(n_1374),
.B(n_1344),
.Y(n_2412)
);

HB1xp67_ASAP7_75t_L g2413 ( 
.A(n_2011),
.Y(n_2413)
);

CKINVDCx5p33_ASAP7_75t_R g2414 ( 
.A(n_2310),
.Y(n_2414)
);

CKINVDCx5p33_ASAP7_75t_R g2415 ( 
.A(n_2310),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2156),
.Y(n_2416)
);

CKINVDCx5p33_ASAP7_75t_R g2417 ( 
.A(n_2328),
.Y(n_2417)
);

INVx3_ASAP7_75t_L g2418 ( 
.A(n_2162),
.Y(n_2418)
);

INVx2_ASAP7_75t_L g2419 ( 
.A(n_1958),
.Y(n_2419)
);

CKINVDCx5p33_ASAP7_75t_R g2420 ( 
.A(n_2328),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_2164),
.Y(n_2421)
);

HB1xp67_ASAP7_75t_L g2422 ( 
.A(n_2011),
.Y(n_2422)
);

CKINVDCx20_ASAP7_75t_R g2423 ( 
.A(n_2218),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2254),
.B(n_1835),
.Y(n_2424)
);

INVx1_ASAP7_75t_L g2425 ( 
.A(n_2172),
.Y(n_2425)
);

INVx3_ASAP7_75t_L g2426 ( 
.A(n_2162),
.Y(n_2426)
);

NOR2xp33_ASAP7_75t_R g2427 ( 
.A(n_2236),
.B(n_1906),
.Y(n_2427)
);

CKINVDCx5p33_ASAP7_75t_R g2428 ( 
.A(n_2284),
.Y(n_2428)
);

HB1xp67_ASAP7_75t_L g2429 ( 
.A(n_2082),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1953),
.B(n_1442),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2177),
.Y(n_2431)
);

CKINVDCx20_ASAP7_75t_R g2432 ( 
.A(n_2314),
.Y(n_2432)
);

BUFx6f_ASAP7_75t_L g2433 ( 
.A(n_1967),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2111),
.Y(n_2434)
);

INVx2_ASAP7_75t_L g2435 ( 
.A(n_1958),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_1961),
.Y(n_2436)
);

NAND2xp5_ASAP7_75t_L g2437 ( 
.A(n_1953),
.B(n_1451),
.Y(n_2437)
);

NOR2xp33_ASAP7_75t_L g2438 ( 
.A(n_2254),
.B(n_1836),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2111),
.Y(n_2439)
);

CKINVDCx5p33_ASAP7_75t_R g2440 ( 
.A(n_2284),
.Y(n_2440)
);

BUFx3_ASAP7_75t_L g2441 ( 
.A(n_1974),
.Y(n_2441)
);

INVx3_ASAP7_75t_L g2442 ( 
.A(n_2162),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2119),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2119),
.Y(n_2444)
);

CKINVDCx5p33_ASAP7_75t_R g2445 ( 
.A(n_1982),
.Y(n_2445)
);

NOR2xp33_ASAP7_75t_R g2446 ( 
.A(n_2139),
.B(n_1917),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_1967),
.Y(n_2447)
);

BUFx3_ASAP7_75t_L g2448 ( 
.A(n_1974),
.Y(n_2448)
);

INVx3_ASAP7_75t_L g2449 ( 
.A(n_2169),
.Y(n_2449)
);

INVx2_ASAP7_75t_L g2450 ( 
.A(n_1961),
.Y(n_2450)
);

CKINVDCx5p33_ASAP7_75t_R g2451 ( 
.A(n_1982),
.Y(n_2451)
);

CKINVDCx20_ASAP7_75t_R g2452 ( 
.A(n_2139),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_2272),
.B(n_1917),
.Y(n_2453)
);

NOR2xp33_ASAP7_75t_L g2454 ( 
.A(n_2220),
.B(n_1836),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2082),
.Y(n_2455)
);

NAND2xp33_ASAP7_75t_R g2456 ( 
.A(n_2031),
.B(n_1745),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2220),
.B(n_1451),
.Y(n_2457)
);

CKINVDCx5p33_ASAP7_75t_R g2458 ( 
.A(n_2038),
.Y(n_2458)
);

CKINVDCx5p33_ASAP7_75t_R g2459 ( 
.A(n_2038),
.Y(n_2459)
);

CKINVDCx20_ASAP7_75t_R g2460 ( 
.A(n_2060),
.Y(n_2460)
);

AND2x6_ASAP7_75t_L g2461 ( 
.A(n_1965),
.B(n_720),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2121),
.Y(n_2462)
);

INVx2_ASAP7_75t_SL g2463 ( 
.A(n_2020),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2121),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2124),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2277),
.B(n_1453),
.Y(n_2466)
);

CKINVDCx20_ASAP7_75t_R g2467 ( 
.A(n_2060),
.Y(n_2467)
);

INVx2_ASAP7_75t_L g2468 ( 
.A(n_1970),
.Y(n_2468)
);

CKINVDCx20_ASAP7_75t_R g2469 ( 
.A(n_2252),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2124),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_1970),
.Y(n_2471)
);

CKINVDCx5p33_ASAP7_75t_R g2472 ( 
.A(n_2031),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_L g2473 ( 
.A(n_1953),
.B(n_1453),
.Y(n_2473)
);

BUFx2_ASAP7_75t_L g2474 ( 
.A(n_2093),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2126),
.Y(n_2475)
);

CKINVDCx20_ASAP7_75t_R g2476 ( 
.A(n_2252),
.Y(n_2476)
);

BUFx6f_ASAP7_75t_L g2477 ( 
.A(n_1980),
.Y(n_2477)
);

CKINVDCx5p33_ASAP7_75t_R g2478 ( 
.A(n_2209),
.Y(n_2478)
);

CKINVDCx5p33_ASAP7_75t_R g2479 ( 
.A(n_2209),
.Y(n_2479)
);

CKINVDCx5p33_ASAP7_75t_R g2480 ( 
.A(n_2326),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_1975),
.Y(n_2481)
);

INVx3_ASAP7_75t_L g2482 ( 
.A(n_2169),
.Y(n_2482)
);

NAND2xp5_ASAP7_75t_L g2483 ( 
.A(n_2232),
.B(n_1454),
.Y(n_2483)
);

CKINVDCx5p33_ASAP7_75t_R g2484 ( 
.A(n_2326),
.Y(n_2484)
);

INVx3_ASAP7_75t_L g2485 ( 
.A(n_2169),
.Y(n_2485)
);

XOR2xp5_ASAP7_75t_L g2486 ( 
.A(n_2311),
.B(n_1670),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2126),
.Y(n_2487)
);

OA21x2_ASAP7_75t_L g2488 ( 
.A1(n_2133),
.A2(n_1374),
.B(n_1344),
.Y(n_2488)
);

INVx2_ASAP7_75t_L g2489 ( 
.A(n_1975),
.Y(n_2489)
);

BUFx2_ASAP7_75t_L g2490 ( 
.A(n_2093),
.Y(n_2490)
);

CKINVDCx20_ASAP7_75t_R g2491 ( 
.A(n_2303),
.Y(n_2491)
);

CKINVDCx20_ASAP7_75t_R g2492 ( 
.A(n_2303),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_1976),
.Y(n_2493)
);

INVxp67_ASAP7_75t_L g2494 ( 
.A(n_2107),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_1976),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_1979),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_L g2497 ( 
.A(n_2232),
.B(n_1454),
.Y(n_2497)
);

INVx1_ASAP7_75t_L g2498 ( 
.A(n_2130),
.Y(n_2498)
);

CKINVDCx20_ASAP7_75t_R g2499 ( 
.A(n_2262),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2130),
.Y(n_2500)
);

INVx1_ASAP7_75t_SL g2501 ( 
.A(n_2097),
.Y(n_2501)
);

INVx3_ASAP7_75t_L g2502 ( 
.A(n_2169),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2135),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_SL g2504 ( 
.A(n_1951),
.B(n_1603),
.Y(n_2504)
);

BUFx6f_ASAP7_75t_L g2505 ( 
.A(n_1980),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2232),
.B(n_1459),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_1959),
.Y(n_2507)
);

CKINVDCx5p33_ASAP7_75t_R g2508 ( 
.A(n_2322),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_2137),
.Y(n_2509)
);

NAND2xp5_ASAP7_75t_L g2510 ( 
.A(n_2246),
.B(n_1459),
.Y(n_2510)
);

INVx3_ASAP7_75t_L g2511 ( 
.A(n_1980),
.Y(n_2511)
);

BUFx3_ASAP7_75t_L g2512 ( 
.A(n_1974),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_1959),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_1959),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_1980),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_1951),
.B(n_1460),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2137),
.Y(n_2517)
);

CKINVDCx20_ASAP7_75t_R g2518 ( 
.A(n_2348),
.Y(n_2518)
);

CKINVDCx5p33_ASAP7_75t_R g2519 ( 
.A(n_2322),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_2322),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2246),
.B(n_1460),
.Y(n_2521)
);

BUFx6f_ASAP7_75t_L g2522 ( 
.A(n_1980),
.Y(n_2522)
);

BUFx6f_ASAP7_75t_L g2523 ( 
.A(n_2066),
.Y(n_2523)
);

CKINVDCx5p33_ASAP7_75t_R g2524 ( 
.A(n_2359),
.Y(n_2524)
);

CKINVDCx5p33_ASAP7_75t_R g2525 ( 
.A(n_2359),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_1959),
.Y(n_2526)
);

CKINVDCx5p33_ASAP7_75t_R g2527 ( 
.A(n_2359),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2182),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2182),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2188),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2189),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2174),
.B(n_1461),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2189),
.Y(n_2533)
);

INVx3_ASAP7_75t_L g2534 ( 
.A(n_2151),
.Y(n_2534)
);

INVx3_ASAP7_75t_L g2535 ( 
.A(n_2151),
.Y(n_2535)
);

CKINVDCx5p33_ASAP7_75t_R g2536 ( 
.A(n_2195),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_1968),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_L g2538 ( 
.A(n_2066),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2192),
.Y(n_2539)
);

CKINVDCx5p33_ASAP7_75t_R g2540 ( 
.A(n_2195),
.Y(n_2540)
);

CKINVDCx5p33_ASAP7_75t_R g2541 ( 
.A(n_2349),
.Y(n_2541)
);

INVx3_ASAP7_75t_L g2542 ( 
.A(n_2151),
.Y(n_2542)
);

INVx1_ASAP7_75t_L g2543 ( 
.A(n_2192),
.Y(n_2543)
);

BUFx2_ASAP7_75t_L g2544 ( 
.A(n_2097),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_2349),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2199),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2365),
.Y(n_2547)
);

CKINVDCx5p33_ASAP7_75t_R g2548 ( 
.A(n_2365),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2197),
.B(n_1461),
.Y(n_2549)
);

CKINVDCx5p33_ASAP7_75t_R g2550 ( 
.A(n_2301),
.Y(n_2550)
);

INVx1_ASAP7_75t_SL g2551 ( 
.A(n_2110),
.Y(n_2551)
);

HB1xp67_ASAP7_75t_L g2552 ( 
.A(n_2110),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_1969),
.B(n_1467),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2199),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2318),
.B(n_1612),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2204),
.Y(n_2556)
);

CKINVDCx20_ASAP7_75t_R g2557 ( 
.A(n_2348),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2255),
.B(n_1467),
.Y(n_2558)
);

BUFx6f_ASAP7_75t_L g2559 ( 
.A(n_2066),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_L g2560 ( 
.A(n_2339),
.B(n_1612),
.Y(n_2560)
);

HB1xp67_ASAP7_75t_L g2561 ( 
.A(n_2141),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2204),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2347),
.B(n_1627),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2221),
.Y(n_2564)
);

CKINVDCx5p33_ASAP7_75t_R g2565 ( 
.A(n_2301),
.Y(n_2565)
);

BUFx2_ASAP7_75t_L g2566 ( 
.A(n_2141),
.Y(n_2566)
);

XNOR2xp5_ASAP7_75t_L g2567 ( 
.A(n_2282),
.B(n_1692),
.Y(n_2567)
);

NOR2xp33_ASAP7_75t_L g2568 ( 
.A(n_2016),
.B(n_1627),
.Y(n_2568)
);

NAND2xp5_ASAP7_75t_SL g2569 ( 
.A(n_1951),
.B(n_1634),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2221),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_2040),
.B(n_1634),
.Y(n_2571)
);

CKINVDCx5p33_ASAP7_75t_R g2572 ( 
.A(n_2301),
.Y(n_2572)
);

CKINVDCx5p33_ASAP7_75t_R g2573 ( 
.A(n_2337),
.Y(n_2573)
);

BUFx2_ASAP7_75t_L g2574 ( 
.A(n_2176),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2228),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_2251),
.B(n_1470),
.Y(n_2576)
);

INVx3_ASAP7_75t_L g2577 ( 
.A(n_2151),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_1968),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2337),
.Y(n_2579)
);

CKINVDCx5p33_ASAP7_75t_R g2580 ( 
.A(n_2337),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2228),
.Y(n_2581)
);

HB1xp67_ASAP7_75t_L g2582 ( 
.A(n_2176),
.Y(n_2582)
);

CKINVDCx5p33_ASAP7_75t_R g2583 ( 
.A(n_2316),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_1983),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2305),
.B(n_1481),
.Y(n_2585)
);

CKINVDCx5p33_ASAP7_75t_R g2586 ( 
.A(n_2272),
.Y(n_2586)
);

NOR2xp67_ASAP7_75t_L g2587 ( 
.A(n_2180),
.B(n_2159),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_1983),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2251),
.B(n_1470),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_1987),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_2251),
.B(n_1473),
.Y(n_2591)
);

OA21x2_ASAP7_75t_L g2592 ( 
.A1(n_2253),
.A2(n_1394),
.B(n_1382),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_SL g2593 ( 
.A(n_2305),
.B(n_1518),
.Y(n_2593)
);

HB1xp67_ASAP7_75t_L g2594 ( 
.A(n_1977),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_1968),
.Y(n_2595)
);

AND2x4_ASAP7_75t_L g2596 ( 
.A(n_2272),
.B(n_1933),
.Y(n_2596)
);

CKINVDCx5p33_ASAP7_75t_R g2597 ( 
.A(n_2275),
.Y(n_2597)
);

CKINVDCx5p33_ASAP7_75t_R g2598 ( 
.A(n_2275),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_1968),
.Y(n_2599)
);

AND2x2_ASAP7_75t_L g2600 ( 
.A(n_2343),
.B(n_2361),
.Y(n_2600)
);

OA21x2_ASAP7_75t_L g2601 ( 
.A1(n_2253),
.A2(n_1394),
.B(n_1382),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2343),
.B(n_2361),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_1988),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2362),
.B(n_1473),
.Y(n_2604)
);

BUFx6f_ASAP7_75t_L g2605 ( 
.A(n_2066),
.Y(n_2605)
);

CKINVDCx20_ASAP7_75t_R g2606 ( 
.A(n_2358),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2362),
.B(n_1476),
.Y(n_2607)
);

INVx2_ASAP7_75t_L g2608 ( 
.A(n_2036),
.Y(n_2608)
);

BUFx6f_ASAP7_75t_L g2609 ( 
.A(n_2066),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_1949),
.B(n_1476),
.Y(n_2610)
);

AND2x2_ASAP7_75t_SL g2611 ( 
.A(n_2282),
.B(n_721),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_1949),
.B(n_1477),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_1949),
.B(n_1477),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_1988),
.Y(n_2614)
);

CKINVDCx5p33_ASAP7_75t_R g2615 ( 
.A(n_2275),
.Y(n_2615)
);

INVxp67_ASAP7_75t_L g2616 ( 
.A(n_2063),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_L g2617 ( 
.A(n_2001),
.B(n_1481),
.Y(n_2617)
);

CKINVDCx20_ASAP7_75t_R g2618 ( 
.A(n_2358),
.Y(n_2618)
);

CKINVDCx5p33_ASAP7_75t_R g2619 ( 
.A(n_2289),
.Y(n_2619)
);

NOR2xp33_ASAP7_75t_R g2620 ( 
.A(n_2279),
.B(n_1926),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2001),
.B(n_2147),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2036),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2036),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2289),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2036),
.Y(n_2625)
);

CKINVDCx8_ASAP7_75t_R g2626 ( 
.A(n_2238),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_1993),
.Y(n_2627)
);

INVx1_ASAP7_75t_SL g2628 ( 
.A(n_2018),
.Y(n_2628)
);

INVxp67_ASAP7_75t_L g2629 ( 
.A(n_2048),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_1993),
.Y(n_2630)
);

INVx2_ASAP7_75t_L g2631 ( 
.A(n_2241),
.Y(n_2631)
);

AND2x6_ASAP7_75t_L g2632 ( 
.A(n_1964),
.B(n_734),
.Y(n_2632)
);

BUFx2_ASAP7_75t_L g2633 ( 
.A(n_2238),
.Y(n_2633)
);

CKINVDCx20_ASAP7_75t_R g2634 ( 
.A(n_2261),
.Y(n_2634)
);

INVx6_ASAP7_75t_L g2635 ( 
.A(n_2180),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2071),
.Y(n_2636)
);

BUFx6f_ASAP7_75t_L g2637 ( 
.A(n_2071),
.Y(n_2637)
);

BUFx2_ASAP7_75t_L g2638 ( 
.A(n_2261),
.Y(n_2638)
);

CKINVDCx20_ASAP7_75t_R g2639 ( 
.A(n_2101),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_1994),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2241),
.Y(n_2641)
);

CKINVDCx20_ASAP7_75t_R g2642 ( 
.A(n_2178),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_2289),
.Y(n_2643)
);

BUFx2_ASAP7_75t_SL g2644 ( 
.A(n_2286),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_SL g2645 ( 
.A(n_2289),
.B(n_1518),
.Y(n_2645)
);

CKINVDCx5p33_ASAP7_75t_R g2646 ( 
.A(n_2289),
.Y(n_2646)
);

NAND2xp5_ASAP7_75t_L g2647 ( 
.A(n_2001),
.B(n_1492),
.Y(n_2647)
);

BUFx6f_ASAP7_75t_L g2648 ( 
.A(n_2071),
.Y(n_2648)
);

CKINVDCx5p33_ASAP7_75t_R g2649 ( 
.A(n_2291),
.Y(n_2649)
);

CKINVDCx5p33_ASAP7_75t_R g2650 ( 
.A(n_2291),
.Y(n_2650)
);

AND2x4_ASAP7_75t_L g2651 ( 
.A(n_2291),
.B(n_2306),
.Y(n_2651)
);

CKINVDCx20_ASAP7_75t_R g2652 ( 
.A(n_2208),
.Y(n_2652)
);

AND2x4_ASAP7_75t_L g2653 ( 
.A(n_2291),
.B(n_1926),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_1994),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_1997),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2241),
.Y(n_2656)
);

INVx3_ASAP7_75t_L g2657 ( 
.A(n_2241),
.Y(n_2657)
);

CKINVDCx5p33_ASAP7_75t_R g2658 ( 
.A(n_2291),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_L g2659 ( 
.A(n_2001),
.B(n_1494),
.Y(n_2659)
);

CKINVDCx5p33_ASAP7_75t_R g2660 ( 
.A(n_2306),
.Y(n_2660)
);

BUFx6f_ASAP7_75t_L g2661 ( 
.A(n_2071),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_2306),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2067),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_1997),
.Y(n_2664)
);

INVx3_ASAP7_75t_L g2665 ( 
.A(n_2059),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2005),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2005),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_L g2668 ( 
.A(n_2001),
.B(n_1494),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_2059),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2067),
.Y(n_2670)
);

INVx2_ASAP7_75t_L g2671 ( 
.A(n_2074),
.Y(n_2671)
);

CKINVDCx20_ASAP7_75t_R g2672 ( 
.A(n_2213),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2364),
.B(n_1495),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_1996),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_1996),
.Y(n_2675)
);

BUFx2_ASAP7_75t_SL g2676 ( 
.A(n_2286),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_2071),
.Y(n_2677)
);

BUFx8_ASAP7_75t_L g2678 ( 
.A(n_2248),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2003),
.Y(n_2679)
);

CKINVDCx5p33_ASAP7_75t_R g2680 ( 
.A(n_2306),
.Y(n_2680)
);

CKINVDCx5p33_ASAP7_75t_R g2681 ( 
.A(n_2306),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_L g2682 ( 
.A(n_2001),
.B(n_1495),
.Y(n_2682)
);

NOR2xp33_ASAP7_75t_L g2683 ( 
.A(n_2084),
.B(n_1933),
.Y(n_2683)
);

CKINVDCx20_ASAP7_75t_R g2684 ( 
.A(n_2346),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2003),
.Y(n_2685)
);

CKINVDCx16_ASAP7_75t_R g2686 ( 
.A(n_2180),
.Y(n_2686)
);

CKINVDCx5p33_ASAP7_75t_R g2687 ( 
.A(n_2317),
.Y(n_2687)
);

CKINVDCx20_ASAP7_75t_R g2688 ( 
.A(n_2037),
.Y(n_2688)
);

INVx3_ASAP7_75t_L g2689 ( 
.A(n_2059),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2006),
.Y(n_2690)
);

HB1xp67_ASAP7_75t_L g2691 ( 
.A(n_2353),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2006),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2317),
.Y(n_2693)
);

INVx3_ASAP7_75t_L g2694 ( 
.A(n_2059),
.Y(n_2694)
);

CKINVDCx5p33_ASAP7_75t_R g2695 ( 
.A(n_2317),
.Y(n_2695)
);

CKINVDCx5p33_ASAP7_75t_R g2696 ( 
.A(n_2317),
.Y(n_2696)
);

CKINVDCx20_ASAP7_75t_R g2697 ( 
.A(n_2317),
.Y(n_2697)
);

INVx3_ASAP7_75t_L g2698 ( 
.A(n_2059),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2074),
.Y(n_2699)
);

CKINVDCx20_ASAP7_75t_R g2700 ( 
.A(n_2329),
.Y(n_2700)
);

INVx1_ASAP7_75t_L g2701 ( 
.A(n_2007),
.Y(n_2701)
);

CKINVDCx5p33_ASAP7_75t_R g2702 ( 
.A(n_2329),
.Y(n_2702)
);

HB1xp67_ASAP7_75t_L g2703 ( 
.A(n_2353),
.Y(n_2703)
);

AND2x2_ASAP7_75t_L g2704 ( 
.A(n_2364),
.B(n_1498),
.Y(n_2704)
);

INVxp67_ASAP7_75t_SL g2705 ( 
.A(n_1972),
.Y(n_2705)
);

CKINVDCx5p33_ASAP7_75t_R g2706 ( 
.A(n_2329),
.Y(n_2706)
);

CKINVDCx5p33_ASAP7_75t_R g2707 ( 
.A(n_2329),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2007),
.Y(n_2708)
);

NOR2xp67_ASAP7_75t_L g2709 ( 
.A(n_2122),
.B(n_1498),
.Y(n_2709)
);

BUFx3_ASAP7_75t_L g2710 ( 
.A(n_1974),
.Y(n_2710)
);

AND2x6_ASAP7_75t_L g2711 ( 
.A(n_2280),
.B(n_735),
.Y(n_2711)
);

BUFx3_ASAP7_75t_L g2712 ( 
.A(n_1972),
.Y(n_2712)
);

BUFx10_ASAP7_75t_L g2713 ( 
.A(n_2166),
.Y(n_2713)
);

CKINVDCx20_ASAP7_75t_R g2714 ( 
.A(n_2329),
.Y(n_2714)
);

BUFx2_ASAP7_75t_L g2715 ( 
.A(n_2282),
.Y(n_2715)
);

BUFx6f_ASAP7_75t_L g2716 ( 
.A(n_2078),
.Y(n_2716)
);

CKINVDCx5p33_ASAP7_75t_R g2717 ( 
.A(n_2248),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2009),
.Y(n_2718)
);

HB1xp67_ASAP7_75t_L g2719 ( 
.A(n_2353),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2009),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2013),
.Y(n_2721)
);

CKINVDCx5p33_ASAP7_75t_R g2722 ( 
.A(n_2248),
.Y(n_2722)
);

BUFx6f_ASAP7_75t_L g2723 ( 
.A(n_2078),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2086),
.Y(n_2724)
);

CKINVDCx20_ASAP7_75t_R g2725 ( 
.A(n_2035),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2013),
.Y(n_2726)
);

INVx5_ASAP7_75t_L g2727 ( 
.A(n_2136),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_SL g2728 ( 
.A(n_2248),
.B(n_1513),
.Y(n_2728)
);

CKINVDCx20_ASAP7_75t_R g2729 ( 
.A(n_2240),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2014),
.Y(n_2730)
);

INVx2_ASAP7_75t_L g2731 ( 
.A(n_2086),
.Y(n_2731)
);

INVx3_ASAP7_75t_L g2732 ( 
.A(n_2041),
.Y(n_2732)
);

CKINVDCx5p33_ASAP7_75t_R g2733 ( 
.A(n_2250),
.Y(n_2733)
);

CKINVDCx20_ASAP7_75t_R g2734 ( 
.A(n_2073),
.Y(n_2734)
);

CKINVDCx20_ASAP7_75t_R g2735 ( 
.A(n_2283),
.Y(n_2735)
);

INVx3_ASAP7_75t_L g2736 ( 
.A(n_2041),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2014),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2021),
.Y(n_2738)
);

BUFx6f_ASAP7_75t_L g2739 ( 
.A(n_2078),
.Y(n_2739)
);

INVx1_ASAP7_75t_SL g2740 ( 
.A(n_2338),
.Y(n_2740)
);

AND2x4_ASAP7_75t_L g2741 ( 
.A(n_2250),
.B(n_1935),
.Y(n_2741)
);

CKINVDCx20_ASAP7_75t_R g2742 ( 
.A(n_2312),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2001),
.B(n_1503),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2021),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2008),
.Y(n_2745)
);

CKINVDCx5p33_ASAP7_75t_R g2746 ( 
.A(n_2250),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2147),
.B(n_1503),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2087),
.Y(n_2748)
);

CKINVDCx5p33_ASAP7_75t_R g2749 ( 
.A(n_2250),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2250),
.Y(n_2750)
);

BUFx6f_ASAP7_75t_L g2751 ( 
.A(n_2078),
.Y(n_2751)
);

CKINVDCx5p33_ASAP7_75t_R g2752 ( 
.A(n_2256),
.Y(n_2752)
);

CKINVDCx5p33_ASAP7_75t_R g2753 ( 
.A(n_2256),
.Y(n_2753)
);

CKINVDCx20_ASAP7_75t_R g2754 ( 
.A(n_2320),
.Y(n_2754)
);

CKINVDCx20_ASAP7_75t_R g2755 ( 
.A(n_2327),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2147),
.B(n_1507),
.Y(n_2756)
);

CKINVDCx5p33_ASAP7_75t_R g2757 ( 
.A(n_2256),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2008),
.Y(n_2758)
);

AND2x2_ASAP7_75t_L g2759 ( 
.A(n_2367),
.B(n_1507),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2012),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2012),
.Y(n_2761)
);

CKINVDCx20_ASAP7_75t_R g2762 ( 
.A(n_2332),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2087),
.Y(n_2763)
);

AND2x2_ASAP7_75t_L g2764 ( 
.A(n_2367),
.B(n_1510),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_2256),
.Y(n_2765)
);

INVx2_ASAP7_75t_L g2766 ( 
.A(n_2088),
.Y(n_2766)
);

AND2x4_ASAP7_75t_L g2767 ( 
.A(n_2256),
.B(n_1941),
.Y(n_2767)
);

BUFx6f_ASAP7_75t_L g2768 ( 
.A(n_2078),
.Y(n_2768)
);

CKINVDCx20_ASAP7_75t_R g2769 ( 
.A(n_2335),
.Y(n_2769)
);

BUFx6f_ASAP7_75t_L g2770 ( 
.A(n_2092),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2023),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_L g2772 ( 
.A(n_2163),
.B(n_1510),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2023),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2088),
.Y(n_2774)
);

INVx3_ASAP7_75t_L g2775 ( 
.A(n_2041),
.Y(n_2775)
);

NOR2xp33_ASAP7_75t_R g2776 ( 
.A(n_2285),
.B(n_1692),
.Y(n_2776)
);

CKINVDCx20_ASAP7_75t_R g2777 ( 
.A(n_2345),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2024),
.Y(n_2778)
);

BUFx6f_ASAP7_75t_L g2779 ( 
.A(n_2092),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2294),
.B(n_1513),
.Y(n_2780)
);

INVx6_ASAP7_75t_L g2781 ( 
.A(n_2145),
.Y(n_2781)
);

CKINVDCx20_ASAP7_75t_R g2782 ( 
.A(n_2350),
.Y(n_2782)
);

INVxp67_ASAP7_75t_L g2783 ( 
.A(n_2056),
.Y(n_2783)
);

INVx1_ASAP7_75t_L g2784 ( 
.A(n_2024),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2028),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2076),
.B(n_1522),
.Y(n_2786)
);

INVx2_ASAP7_75t_L g2787 ( 
.A(n_2089),
.Y(n_2787)
);

INVx1_ASAP7_75t_L g2788 ( 
.A(n_2028),
.Y(n_2788)
);

CKINVDCx5p33_ASAP7_75t_R g2789 ( 
.A(n_2265),
.Y(n_2789)
);

OAI21x1_ASAP7_75t_L g2790 ( 
.A1(n_2077),
.A2(n_1409),
.B(n_1399),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2042),
.Y(n_2791)
);

CKINVDCx5p33_ASAP7_75t_R g2792 ( 
.A(n_2265),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2042),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2043),
.Y(n_2794)
);

INVx3_ASAP7_75t_L g2795 ( 
.A(n_1992),
.Y(n_2795)
);

AND3x2_ASAP7_75t_L g2796 ( 
.A(n_2352),
.B(n_1713),
.C(n_1708),
.Y(n_2796)
);

INVx2_ASAP7_75t_L g2797 ( 
.A(n_2089),
.Y(n_2797)
);

OAI21x1_ASAP7_75t_L g2798 ( 
.A1(n_2077),
.A2(n_1409),
.B(n_1399),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2103),
.Y(n_2799)
);

BUFx6f_ASAP7_75t_L g2800 ( 
.A(n_2092),
.Y(n_2800)
);

INVx2_ASAP7_75t_L g2801 ( 
.A(n_2103),
.Y(n_2801)
);

CKINVDCx5p33_ASAP7_75t_R g2802 ( 
.A(n_2265),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2043),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2163),
.B(n_1517),
.Y(n_2804)
);

CKINVDCx5p33_ASAP7_75t_R g2805 ( 
.A(n_2265),
.Y(n_2805)
);

BUFx8_ASAP7_75t_L g2806 ( 
.A(n_2265),
.Y(n_2806)
);

BUFx6f_ASAP7_75t_L g2807 ( 
.A(n_2092),
.Y(n_2807)
);

BUFx6f_ASAP7_75t_L g2808 ( 
.A(n_2092),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2047),
.Y(n_2809)
);

INVx3_ASAP7_75t_L g2810 ( 
.A(n_1992),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2047),
.Y(n_2811)
);

AOI22xp5_ASAP7_75t_L g2812 ( 
.A1(n_2585),
.A2(n_2290),
.B1(n_2292),
.B2(n_2281),
.Y(n_2812)
);

AOI22xp33_ASAP7_75t_L g2813 ( 
.A1(n_2611),
.A2(n_1971),
.B1(n_2308),
.B2(n_2205),
.Y(n_2813)
);

INVx3_ASAP7_75t_L g2814 ( 
.A(n_2727),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_SL g2815 ( 
.A(n_2717),
.B(n_2267),
.Y(n_2815)
);

INVx2_ASAP7_75t_L g2816 ( 
.A(n_2663),
.Y(n_2816)
);

BUFx3_ASAP7_75t_L g2817 ( 
.A(n_2678),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2670),
.Y(n_2818)
);

BUFx2_ASAP7_75t_L g2819 ( 
.A(n_2474),
.Y(n_2819)
);

OR2x6_ASAP7_75t_L g2820 ( 
.A(n_2715),
.B(n_2267),
.Y(n_2820)
);

INVx3_ASAP7_75t_L g2821 ( 
.A(n_2727),
.Y(n_2821)
);

AOI22xp33_ASAP7_75t_SL g2822 ( 
.A1(n_2611),
.A2(n_1971),
.B1(n_2205),
.B2(n_2308),
.Y(n_2822)
);

AND2x4_ASAP7_75t_L g2823 ( 
.A(n_2387),
.B(n_2207),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_SL g2824 ( 
.A(n_2717),
.B(n_2267),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2670),
.Y(n_2825)
);

AOI22xp33_ASAP7_75t_SL g2826 ( 
.A1(n_2460),
.A2(n_2308),
.B1(n_2363),
.B2(n_2273),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2671),
.Y(n_2827)
);

INVx2_ASAP7_75t_SL g2828 ( 
.A(n_2781),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2600),
.B(n_2285),
.Y(n_2829)
);

NAND2xp5_ASAP7_75t_SL g2830 ( 
.A(n_2722),
.B(n_2267),
.Y(n_2830)
);

AND2x6_ASAP7_75t_L g2831 ( 
.A(n_2621),
.B(n_2267),
.Y(n_2831)
);

BUFx2_ASAP7_75t_L g2832 ( 
.A(n_2490),
.Y(n_2832)
);

BUFx3_ASAP7_75t_L g2833 ( 
.A(n_2678),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2671),
.Y(n_2834)
);

INVx4_ASAP7_75t_L g2835 ( 
.A(n_2727),
.Y(n_2835)
);

INVx2_ASAP7_75t_SL g2836 ( 
.A(n_2781),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2699),
.Y(n_2837)
);

CKINVDCx5p33_ASAP7_75t_R g2838 ( 
.A(n_2456),
.Y(n_2838)
);

INVx2_ASAP7_75t_SL g2839 ( 
.A(n_2781),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2699),
.Y(n_2840)
);

BUFx6f_ASAP7_75t_L g2841 ( 
.A(n_2523),
.Y(n_2841)
);

OR2x6_ASAP7_75t_L g2842 ( 
.A(n_2387),
.B(n_2207),
.Y(n_2842)
);

INVx2_ASAP7_75t_SL g2843 ( 
.A(n_2441),
.Y(n_2843)
);

INVx3_ASAP7_75t_L g2844 ( 
.A(n_2727),
.Y(n_2844)
);

AND2x2_ASAP7_75t_L g2845 ( 
.A(n_2740),
.B(n_2076),
.Y(n_2845)
);

CKINVDCx20_ASAP7_75t_R g2846 ( 
.A(n_2390),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2724),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2724),
.Y(n_2848)
);

INVx1_ASAP7_75t_SL g2849 ( 
.A(n_2501),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2731),
.Y(n_2850)
);

INVx3_ASAP7_75t_L g2851 ( 
.A(n_2727),
.Y(n_2851)
);

INVx3_ASAP7_75t_L g2852 ( 
.A(n_2523),
.Y(n_2852)
);

NOR2xp33_ASAP7_75t_L g2853 ( 
.A(n_2555),
.B(n_2352),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2602),
.B(n_2336),
.Y(n_2854)
);

INVx4_ASAP7_75t_L g2855 ( 
.A(n_2523),
.Y(n_2855)
);

INVx3_ASAP7_75t_L g2856 ( 
.A(n_2523),
.Y(n_2856)
);

NAND3xp33_ASAP7_75t_L g2857 ( 
.A(n_2683),
.B(n_2004),
.C(n_2355),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2560),
.B(n_2338),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2748),
.Y(n_2859)
);

INVx2_ASAP7_75t_L g2860 ( 
.A(n_2748),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2763),
.Y(n_2861)
);

BUFx8_ASAP7_75t_SL g2862 ( 
.A(n_2390),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_2763),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_2563),
.B(n_2355),
.Y(n_2864)
);

INVxp67_ASAP7_75t_SL g2865 ( 
.A(n_2538),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2766),
.Y(n_2866)
);

INVx2_ASAP7_75t_SL g2867 ( 
.A(n_2441),
.Y(n_2867)
);

BUFx3_ASAP7_75t_L g2868 ( 
.A(n_2678),
.Y(n_2868)
);

OR2x6_ASAP7_75t_L g2869 ( 
.A(n_2387),
.B(n_2281),
.Y(n_2869)
);

NAND2xp5_ASAP7_75t_L g2870 ( 
.A(n_2568),
.B(n_2571),
.Y(n_2870)
);

BUFx6f_ASAP7_75t_L g2871 ( 
.A(n_2538),
.Y(n_2871)
);

NAND2xp33_ASAP7_75t_L g2872 ( 
.A(n_2550),
.B(n_2260),
.Y(n_2872)
);

NOR2xp33_ASAP7_75t_L g2873 ( 
.A(n_2729),
.B(n_2380),
.Y(n_2873)
);

CKINVDCx20_ASAP7_75t_R g2874 ( 
.A(n_2410),
.Y(n_2874)
);

INVx3_ASAP7_75t_L g2875 ( 
.A(n_2538),
.Y(n_2875)
);

INVx2_ASAP7_75t_L g2876 ( 
.A(n_2774),
.Y(n_2876)
);

INVx3_ASAP7_75t_L g2877 ( 
.A(n_2538),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2774),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2787),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2787),
.Y(n_2880)
);

OR2x6_ASAP7_75t_L g2881 ( 
.A(n_2651),
.B(n_2290),
.Y(n_2881)
);

AOI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2585),
.A2(n_2295),
.B1(n_2296),
.B2(n_2292),
.Y(n_2882)
);

HB1xp67_ASAP7_75t_L g2883 ( 
.A(n_2551),
.Y(n_2883)
);

INVx8_ASAP7_75t_L g2884 ( 
.A(n_2711),
.Y(n_2884)
);

INVx4_ASAP7_75t_L g2885 ( 
.A(n_2559),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2375),
.B(n_2295),
.Y(n_2886)
);

INVxp33_ASAP7_75t_SL g2887 ( 
.A(n_2427),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2797),
.Y(n_2888)
);

AO22x2_ASAP7_75t_L g2889 ( 
.A1(n_2516),
.A2(n_2186),
.B1(n_2214),
.B2(n_2046),
.Y(n_2889)
);

INVx2_ASAP7_75t_SL g2890 ( 
.A(n_2448),
.Y(n_2890)
);

INVx3_ASAP7_75t_L g2891 ( 
.A(n_2559),
.Y(n_2891)
);

INVx2_ASAP7_75t_L g2892 ( 
.A(n_2797),
.Y(n_2892)
);

NAND2xp33_ASAP7_75t_L g2893 ( 
.A(n_2550),
.B(n_2260),
.Y(n_2893)
);

INVx3_ASAP7_75t_L g2894 ( 
.A(n_2559),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2799),
.Y(n_2895)
);

INVx2_ASAP7_75t_L g2896 ( 
.A(n_2799),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2801),
.Y(n_2897)
);

INVx1_ASAP7_75t_L g2898 ( 
.A(n_2801),
.Y(n_2898)
);

NAND2xp33_ASAP7_75t_SL g2899 ( 
.A(n_2565),
.B(n_2260),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2369),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2370),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2377),
.Y(n_2902)
);

INVx4_ASAP7_75t_L g2903 ( 
.A(n_2559),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2383),
.B(n_2296),
.Y(n_2904)
);

NAND2xp33_ASAP7_75t_L g2905 ( 
.A(n_2565),
.B(n_2298),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2576),
.B(n_2298),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2729),
.B(n_2269),
.Y(n_2907)
);

NOR2xp33_ASAP7_75t_L g2908 ( 
.A(n_2688),
.B(n_2269),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2378),
.Y(n_2909)
);

AOI22xp33_ASAP7_75t_SL g2910 ( 
.A1(n_2460),
.A2(n_2308),
.B1(n_2142),
.B2(n_1713),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2384),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2370),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2381),
.Y(n_2913)
);

INVx2_ASAP7_75t_SL g2914 ( 
.A(n_2448),
.Y(n_2914)
);

CKINVDCx20_ASAP7_75t_R g2915 ( 
.A(n_2410),
.Y(n_2915)
);

INVx2_ASAP7_75t_L g2916 ( 
.A(n_2381),
.Y(n_2916)
);

INVx2_ASAP7_75t_L g2917 ( 
.A(n_2386),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2386),
.Y(n_2918)
);

INVx3_ASAP7_75t_L g2919 ( 
.A(n_2605),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2388),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2589),
.B(n_2304),
.Y(n_2921)
);

INVx3_ASAP7_75t_L g2922 ( 
.A(n_2605),
.Y(n_2922)
);

BUFx2_ASAP7_75t_L g2923 ( 
.A(n_2544),
.Y(n_2923)
);

INVx2_ASAP7_75t_SL g2924 ( 
.A(n_2512),
.Y(n_2924)
);

INVx3_ASAP7_75t_L g2925 ( 
.A(n_2605),
.Y(n_2925)
);

INVx1_ASAP7_75t_SL g2926 ( 
.A(n_2566),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2388),
.Y(n_2927)
);

INVxp33_ASAP7_75t_SL g2928 ( 
.A(n_2404),
.Y(n_2928)
);

INVx4_ASAP7_75t_L g2929 ( 
.A(n_2605),
.Y(n_2929)
);

NAND2xp33_ASAP7_75t_L g2930 ( 
.A(n_2572),
.B(n_2304),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2591),
.B(n_2325),
.Y(n_2931)
);

INVx2_ASAP7_75t_SL g2932 ( 
.A(n_2512),
.Y(n_2932)
);

INVx4_ASAP7_75t_L g2933 ( 
.A(n_2609),
.Y(n_2933)
);

OR2x6_ASAP7_75t_L g2934 ( 
.A(n_2651),
.B(n_2325),
.Y(n_2934)
);

INVxp67_ASAP7_75t_SL g2935 ( 
.A(n_2609),
.Y(n_2935)
);

INVx1_ASAP7_75t_L g2936 ( 
.A(n_2394),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2553),
.B(n_2330),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2396),
.Y(n_2938)
);

INVx2_ASAP7_75t_SL g2939 ( 
.A(n_2710),
.Y(n_2939)
);

INVx5_ASAP7_75t_L g2940 ( 
.A(n_2609),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2405),
.Y(n_2941)
);

BUFx6f_ASAP7_75t_L g2942 ( 
.A(n_2609),
.Y(n_2942)
);

BUFx6f_ASAP7_75t_L g2943 ( 
.A(n_2636),
.Y(n_2943)
);

NOR2xp33_ASAP7_75t_L g2944 ( 
.A(n_2688),
.B(n_2270),
.Y(n_2944)
);

OAI22x1_ASAP7_75t_L g2945 ( 
.A1(n_2486),
.A2(n_2331),
.B1(n_2330),
.B2(n_2271),
.Y(n_2945)
);

INVx2_ASAP7_75t_L g2946 ( 
.A(n_2405),
.Y(n_2946)
);

BUFx3_ASAP7_75t_L g2947 ( 
.A(n_2806),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2398),
.Y(n_2948)
);

INVx4_ASAP7_75t_L g2949 ( 
.A(n_2636),
.Y(n_2949)
);

INVx2_ASAP7_75t_L g2950 ( 
.A(n_2407),
.Y(n_2950)
);

OAI22xp33_ASAP7_75t_SL g2951 ( 
.A1(n_2691),
.A2(n_2323),
.B1(n_2271),
.B2(n_2276),
.Y(n_2951)
);

NAND3xp33_ASAP7_75t_L g2952 ( 
.A(n_2376),
.B(n_2276),
.C(n_2270),
.Y(n_2952)
);

AND3x2_ASAP7_75t_L g2953 ( 
.A(n_2454),
.B(n_2767),
.C(n_2741),
.Y(n_2953)
);

NOR2xp33_ASAP7_75t_L g2954 ( 
.A(n_2466),
.B(n_2287),
.Y(n_2954)
);

NAND2xp5_ASAP7_75t_SL g2955 ( 
.A(n_2733),
.B(n_2331),
.Y(n_2955)
);

INVx1_ASAP7_75t_L g2956 ( 
.A(n_2406),
.Y(n_2956)
);

AND2x4_ASAP7_75t_L g2957 ( 
.A(n_2651),
.B(n_2051),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2407),
.Y(n_2958)
);

INVx3_ASAP7_75t_L g2959 ( 
.A(n_2636),
.Y(n_2959)
);

BUFx6f_ASAP7_75t_L g2960 ( 
.A(n_2636),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2419),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2419),
.Y(n_2962)
);

INVx3_ASAP7_75t_L g2963 ( 
.A(n_2637),
.Y(n_2963)
);

OAI22xp33_ASAP7_75t_L g2964 ( 
.A1(n_2385),
.A2(n_2288),
.B1(n_2293),
.B2(n_2287),
.Y(n_2964)
);

INVx3_ASAP7_75t_L g2965 ( 
.A(n_2637),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2435),
.Y(n_2966)
);

CKINVDCx6p67_ASAP7_75t_R g2967 ( 
.A(n_2452),
.Y(n_2967)
);

INVx1_ASAP7_75t_L g2968 ( 
.A(n_2435),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2436),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2436),
.Y(n_2970)
);

INVx3_ASAP7_75t_L g2971 ( 
.A(n_2637),
.Y(n_2971)
);

BUFx2_ASAP7_75t_L g2972 ( 
.A(n_2574),
.Y(n_2972)
);

NOR2xp33_ASAP7_75t_L g2973 ( 
.A(n_2628),
.B(n_2288),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2450),
.Y(n_2974)
);

BUFx10_ASAP7_75t_L g2975 ( 
.A(n_2411),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2450),
.Y(n_2976)
);

INVx2_ASAP7_75t_L g2977 ( 
.A(n_2468),
.Y(n_2977)
);

INVx2_ASAP7_75t_SL g2978 ( 
.A(n_2710),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2713),
.B(n_2293),
.Y(n_2979)
);

BUFx6f_ASAP7_75t_L g2980 ( 
.A(n_2637),
.Y(n_2980)
);

INVx2_ASAP7_75t_L g2981 ( 
.A(n_2468),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2471),
.Y(n_2982)
);

AOI22xp33_ASAP7_75t_L g2983 ( 
.A1(n_2711),
.A2(n_2308),
.B1(n_2247),
.B2(n_2146),
.Y(n_2983)
);

CKINVDCx16_ASAP7_75t_R g2984 ( 
.A(n_2446),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2471),
.Y(n_2985)
);

NOR2xp33_ASAP7_75t_L g2986 ( 
.A(n_2713),
.B(n_2297),
.Y(n_2986)
);

NAND3xp33_ASAP7_75t_L g2987 ( 
.A(n_2616),
.B(n_2323),
.C(n_2321),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2481),
.Y(n_2988)
);

INVx1_ASAP7_75t_L g2989 ( 
.A(n_2481),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2489),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_SL g2991 ( 
.A(n_2733),
.B(n_2746),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2489),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2711),
.A2(n_2308),
.B1(n_2247),
.B2(n_2146),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_SL g2994 ( 
.A(n_2746),
.B(n_2264),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2493),
.Y(n_2995)
);

AOI22xp5_ASAP7_75t_L g2996 ( 
.A1(n_2586),
.A2(n_2597),
.B1(n_2615),
.B2(n_2598),
.Y(n_2996)
);

NAND2xp5_ASAP7_75t_SL g2997 ( 
.A(n_2749),
.B(n_2264),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2493),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2495),
.Y(n_2999)
);

INVx1_ASAP7_75t_L g3000 ( 
.A(n_2495),
.Y(n_3000)
);

NOR2xp33_ASAP7_75t_L g3001 ( 
.A(n_2713),
.B(n_2297),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2496),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2507),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2403),
.B(n_2114),
.Y(n_3004)
);

INVx2_ASAP7_75t_L g3005 ( 
.A(n_2507),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2513),
.Y(n_3006)
);

BUFx3_ASAP7_75t_L g3007 ( 
.A(n_2806),
.Y(n_3007)
);

BUFx3_ASAP7_75t_L g3008 ( 
.A(n_2806),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2709),
.B(n_2148),
.Y(n_3009)
);

OR2x6_ASAP7_75t_L g3010 ( 
.A(n_2399),
.B(n_2185),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2409),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2513),
.Y(n_3012)
);

CKINVDCx20_ASAP7_75t_R g3013 ( 
.A(n_2423),
.Y(n_3013)
);

OAI22xp5_ASAP7_75t_L g3014 ( 
.A1(n_2586),
.A2(n_2307),
.B1(n_2309),
.B2(n_2300),
.Y(n_3014)
);

BUFx6f_ASAP7_75t_L g3015 ( 
.A(n_2648),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2514),
.Y(n_3016)
);

AO22x2_ASAP7_75t_L g3017 ( 
.A1(n_2516),
.A2(n_2280),
.B1(n_2308),
.B2(n_2342),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_SL g3018 ( 
.A(n_2749),
.B(n_2300),
.Y(n_3018)
);

BUFx10_ASAP7_75t_L g3019 ( 
.A(n_2411),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2514),
.Y(n_3020)
);

NAND2xp5_ASAP7_75t_SL g3021 ( 
.A(n_2750),
.B(n_2307),
.Y(n_3021)
);

CKINVDCx6p67_ASAP7_75t_R g3022 ( 
.A(n_2452),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2780),
.B(n_2190),
.Y(n_3023)
);

INVx2_ASAP7_75t_SL g3024 ( 
.A(n_2635),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2526),
.Y(n_3025)
);

INVx3_ASAP7_75t_L g3026 ( 
.A(n_2648),
.Y(n_3026)
);

BUFx10_ASAP7_75t_L g3027 ( 
.A(n_2414),
.Y(n_3027)
);

INVx1_ASAP7_75t_L g3028 ( 
.A(n_2416),
.Y(n_3028)
);

NAND3xp33_ASAP7_75t_L g3029 ( 
.A(n_2629),
.B(n_2313),
.C(n_2309),
.Y(n_3029)
);

NAND2xp33_ASAP7_75t_L g3030 ( 
.A(n_2572),
.B(n_2324),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2421),
.Y(n_3031)
);

BUFx3_ASAP7_75t_L g3032 ( 
.A(n_2382),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_SL g3033 ( 
.A(n_2750),
.B(n_2752),
.Y(n_3033)
);

BUFx2_ASAP7_75t_L g3034 ( 
.A(n_2429),
.Y(n_3034)
);

BUFx2_ASAP7_75t_L g3035 ( 
.A(n_2455),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_L g3036 ( 
.A(n_2472),
.B(n_2313),
.Y(n_3036)
);

BUFx6f_ASAP7_75t_L g3037 ( 
.A(n_2648),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2425),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2673),
.B(n_2200),
.Y(n_3039)
);

INVx2_ASAP7_75t_L g3040 ( 
.A(n_2526),
.Y(n_3040)
);

INVx3_ASAP7_75t_L g3041 ( 
.A(n_2661),
.Y(n_3041)
);

INVx2_ASAP7_75t_L g3042 ( 
.A(n_2537),
.Y(n_3042)
);

INVx2_ASAP7_75t_L g3043 ( 
.A(n_2537),
.Y(n_3043)
);

AND2x4_ASAP7_75t_L g3044 ( 
.A(n_2697),
.B(n_2051),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2578),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2578),
.Y(n_3046)
);

INVx3_ASAP7_75t_L g3047 ( 
.A(n_2661),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2595),
.Y(n_3048)
);

NAND3xp33_ASAP7_75t_L g3049 ( 
.A(n_2783),
.B(n_2319),
.C(n_2315),
.Y(n_3049)
);

NOR2xp33_ASAP7_75t_L g3050 ( 
.A(n_2472),
.B(n_2315),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2704),
.B(n_2217),
.Y(n_3051)
);

INVx2_ASAP7_75t_L g3052 ( 
.A(n_2595),
.Y(n_3052)
);

CKINVDCx5p33_ASAP7_75t_R g3053 ( 
.A(n_2414),
.Y(n_3053)
);

INVx2_ASAP7_75t_SL g3054 ( 
.A(n_2635),
.Y(n_3054)
);

AND2x2_ASAP7_75t_L g3055 ( 
.A(n_2759),
.B(n_2076),
.Y(n_3055)
);

INVx2_ASAP7_75t_SL g3056 ( 
.A(n_2635),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2431),
.Y(n_3057)
);

INVx4_ASAP7_75t_L g3058 ( 
.A(n_2661),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_SL g3059 ( 
.A(n_2752),
.B(n_2319),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2599),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2599),
.Y(n_3061)
);

AND2x2_ASAP7_75t_L g3062 ( 
.A(n_2764),
.B(n_2294),
.Y(n_3062)
);

OR2x6_ASAP7_75t_L g3063 ( 
.A(n_2399),
.B(n_2185),
.Y(n_3063)
);

INVx2_ASAP7_75t_L g3064 ( 
.A(n_2608),
.Y(n_3064)
);

OAI22xp33_ASAP7_75t_L g3065 ( 
.A1(n_2430),
.A2(n_2321),
.B1(n_2334),
.B2(n_2324),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2434),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2439),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_SL g3068 ( 
.A(n_2753),
.B(n_2334),
.Y(n_3068)
);

INVx3_ASAP7_75t_L g3069 ( 
.A(n_2661),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2608),
.Y(n_3070)
);

INVx2_ASAP7_75t_SL g3071 ( 
.A(n_2597),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_SL g3072 ( 
.A(n_2753),
.B(n_2222),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2622),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2478),
.B(n_2366),
.Y(n_3074)
);

BUFx4f_ASAP7_75t_L g3075 ( 
.A(n_2711),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2443),
.Y(n_3076)
);

NOR2xp33_ASAP7_75t_L g3077 ( 
.A(n_2478),
.B(n_2479),
.Y(n_3077)
);

AND2x2_ASAP7_75t_L g3078 ( 
.A(n_2786),
.B(n_2027),
.Y(n_3078)
);

AOI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2598),
.A2(n_2280),
.B1(n_2258),
.B2(n_2233),
.Y(n_3079)
);

AOI22xp33_ASAP7_75t_L g3080 ( 
.A1(n_2711),
.A2(n_2703),
.B1(n_2719),
.B2(n_2247),
.Y(n_3080)
);

AOI22xp5_ASAP7_75t_L g3081 ( 
.A1(n_2615),
.A2(n_2258),
.B1(n_2249),
.B2(n_2225),
.Y(n_3081)
);

AND2x2_ASAP7_75t_L g3082 ( 
.A(n_2786),
.B(n_2027),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2444),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2483),
.B(n_2497),
.Y(n_3084)
);

INVx2_ASAP7_75t_SL g3085 ( 
.A(n_2619),
.Y(n_3085)
);

NOR2xp33_ASAP7_75t_L g3086 ( 
.A(n_2479),
.B(n_1719),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_SL g3087 ( 
.A(n_2757),
.B(n_1984),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2622),
.Y(n_3088)
);

NAND3xp33_ASAP7_75t_L g3089 ( 
.A(n_2415),
.B(n_1522),
.C(n_1517),
.Y(n_3089)
);

NAND2xp33_ASAP7_75t_L g3090 ( 
.A(n_2573),
.B(n_2136),
.Y(n_3090)
);

INVx4_ASAP7_75t_L g3091 ( 
.A(n_2677),
.Y(n_3091)
);

INVx1_ASAP7_75t_L g3092 ( 
.A(n_2462),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2464),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2677),
.Y(n_3094)
);

INVx1_ASAP7_75t_L g3095 ( 
.A(n_2465),
.Y(n_3095)
);

BUFx2_ASAP7_75t_L g3096 ( 
.A(n_2552),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2470),
.Y(n_3097)
);

BUFx10_ASAP7_75t_L g3098 ( 
.A(n_2415),
.Y(n_3098)
);

NAND3xp33_ASAP7_75t_L g3099 ( 
.A(n_2417),
.B(n_1538),
.C(n_1531),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_SL g3100 ( 
.A(n_2765),
.B(n_1990),
.Y(n_3100)
);

NAND2xp5_ASAP7_75t_L g3101 ( 
.A(n_2506),
.B(n_2027),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2747),
.B(n_2342),
.Y(n_3102)
);

OAI22xp33_ASAP7_75t_L g3103 ( 
.A1(n_2437),
.A2(n_2266),
.B1(n_2268),
.B2(n_2263),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2475),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2623),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2487),
.Y(n_3106)
);

INVx4_ASAP7_75t_L g3107 ( 
.A(n_2677),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2623),
.Y(n_3108)
);

AO21x2_ASAP7_75t_L g3109 ( 
.A1(n_2617),
.A2(n_2106),
.B(n_2054),
.Y(n_3109)
);

INVx4_ASAP7_75t_L g3110 ( 
.A(n_2677),
.Y(n_3110)
);

INVx2_ASAP7_75t_L g3111 ( 
.A(n_2625),
.Y(n_3111)
);

INVx3_ASAP7_75t_L g3112 ( 
.A(n_2716),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2789),
.B(n_1998),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2498),
.Y(n_3114)
);

BUFx2_ASAP7_75t_L g3115 ( 
.A(n_2561),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_2619),
.Y(n_3116)
);

INVx4_ASAP7_75t_L g3117 ( 
.A(n_2716),
.Y(n_3117)
);

AOI22xp33_ASAP7_75t_L g3118 ( 
.A1(n_2711),
.A2(n_2146),
.B1(n_2175),
.B2(n_2210),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2382),
.Y(n_3119)
);

NAND2xp5_ASAP7_75t_SL g3120 ( 
.A(n_2789),
.B(n_1998),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2625),
.Y(n_3121)
);

INVx2_ASAP7_75t_SL g3122 ( 
.A(n_2624),
.Y(n_3122)
);

BUFx8_ASAP7_75t_SL g3123 ( 
.A(n_2432),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2494),
.B(n_1719),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2631),
.Y(n_3125)
);

INVx4_ASAP7_75t_L g3126 ( 
.A(n_2716),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_SL g3127 ( 
.A(n_2792),
.B(n_2263),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2500),
.Y(n_3128)
);

CKINVDCx6p67_ASAP7_75t_R g3129 ( 
.A(n_2432),
.Y(n_3129)
);

INVx2_ASAP7_75t_SL g3130 ( 
.A(n_2624),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_SL g3131 ( 
.A(n_2792),
.B(n_2266),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2503),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2509),
.Y(n_3133)
);

INVx2_ASAP7_75t_L g3134 ( 
.A(n_2631),
.Y(n_3134)
);

AND2x6_ASAP7_75t_L g3135 ( 
.A(n_2716),
.B(n_2210),
.Y(n_3135)
);

AOI22xp33_ASAP7_75t_L g3136 ( 
.A1(n_2725),
.A2(n_2175),
.B1(n_2210),
.B2(n_2181),
.Y(n_3136)
);

BUFx2_ASAP7_75t_L g3137 ( 
.A(n_2582),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2517),
.Y(n_3138)
);

NAND2xp33_ASAP7_75t_R g3139 ( 
.A(n_2620),
.B(n_2278),
.Y(n_3139)
);

INVx2_ASAP7_75t_L g3140 ( 
.A(n_2641),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2528),
.B(n_2302),
.Y(n_3141)
);

INVxp33_ASAP7_75t_L g3142 ( 
.A(n_2372),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2529),
.Y(n_3143)
);

BUFx6f_ASAP7_75t_L g3144 ( 
.A(n_2723),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2530),
.Y(n_3145)
);

OAI22x1_ASAP7_75t_L g3146 ( 
.A1(n_2567),
.A2(n_2268),
.B1(n_2344),
.B2(n_2274),
.Y(n_3146)
);

AND2x4_ASAP7_75t_L g3147 ( 
.A(n_2697),
.B(n_2057),
.Y(n_3147)
);

INVx2_ASAP7_75t_L g3148 ( 
.A(n_2641),
.Y(n_3148)
);

INVx2_ASAP7_75t_SL g3149 ( 
.A(n_2643),
.Y(n_3149)
);

NOR2xp33_ASAP7_75t_L g3150 ( 
.A(n_2413),
.B(n_1721),
.Y(n_3150)
);

AOI22xp33_ASAP7_75t_L g3151 ( 
.A1(n_2725),
.A2(n_2175),
.B1(n_2181),
.B2(n_2143),
.Y(n_3151)
);

AND2x6_ASAP7_75t_L g3152 ( 
.A(n_2723),
.B(n_2181),
.Y(n_3152)
);

CKINVDCx5p33_ASAP7_75t_R g3153 ( 
.A(n_2417),
.Y(n_3153)
);

INVx3_ASAP7_75t_L g3154 ( 
.A(n_2723),
.Y(n_3154)
);

INVx2_ASAP7_75t_L g3155 ( 
.A(n_2656),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2531),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2533),
.Y(n_3157)
);

OAI21xp33_ASAP7_75t_L g3158 ( 
.A1(n_2610),
.A2(n_1538),
.B(n_1531),
.Y(n_3158)
);

INVx1_ASAP7_75t_L g3159 ( 
.A(n_2539),
.Y(n_3159)
);

INVx2_ASAP7_75t_SL g3160 ( 
.A(n_2643),
.Y(n_3160)
);

AO22x2_ASAP7_75t_L g3161 ( 
.A1(n_2674),
.A2(n_2357),
.B1(n_2259),
.B2(n_2138),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_2723),
.Y(n_3162)
);

INVx1_ASAP7_75t_L g3163 ( 
.A(n_2543),
.Y(n_3163)
);

INVx2_ASAP7_75t_L g3164 ( 
.A(n_2397),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2397),
.Y(n_3165)
);

INVx2_ASAP7_75t_L g3166 ( 
.A(n_2397),
.Y(n_3166)
);

BUFx6f_ASAP7_75t_L g3167 ( 
.A(n_2739),
.Y(n_3167)
);

CKINVDCx6p67_ASAP7_75t_R g3168 ( 
.A(n_2686),
.Y(n_3168)
);

AOI22xp5_ASAP7_75t_L g3169 ( 
.A1(n_2646),
.A2(n_2340),
.B1(n_1991),
.B2(n_2134),
.Y(n_3169)
);

NOR2x1p5_ASAP7_75t_L g3170 ( 
.A(n_2508),
.B(n_2274),
.Y(n_3170)
);

NOR2xp33_ASAP7_75t_L g3171 ( 
.A(n_2422),
.B(n_1721),
.Y(n_3171)
);

INVx2_ASAP7_75t_L g3172 ( 
.A(n_2418),
.Y(n_3172)
);

INVx3_ASAP7_75t_L g3173 ( 
.A(n_2739),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2756),
.B(n_2026),
.Y(n_3174)
);

AOI22xp33_ASAP7_75t_L g3175 ( 
.A1(n_2639),
.A2(n_2184),
.B1(n_2216),
.B2(n_2143),
.Y(n_3175)
);

BUFx6f_ASAP7_75t_L g3176 ( 
.A(n_2739),
.Y(n_3176)
);

INVx5_ASAP7_75t_L g3177 ( 
.A(n_2739),
.Y(n_3177)
);

BUFx3_ASAP7_75t_L g3178 ( 
.A(n_2382),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2418),
.Y(n_3179)
);

BUFx2_ASAP7_75t_L g3180 ( 
.A(n_2633),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2546),
.Y(n_3181)
);

INVx2_ASAP7_75t_L g3182 ( 
.A(n_2418),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_2772),
.B(n_2026),
.Y(n_3183)
);

INVx1_ASAP7_75t_L g3184 ( 
.A(n_2554),
.Y(n_3184)
);

INVx2_ASAP7_75t_L g3185 ( 
.A(n_2426),
.Y(n_3185)
);

INVx1_ASAP7_75t_L g3186 ( 
.A(n_2556),
.Y(n_3186)
);

INVx2_ASAP7_75t_L g3187 ( 
.A(n_2426),
.Y(n_3187)
);

OAI22xp33_ASAP7_75t_L g3188 ( 
.A1(n_2473),
.A2(n_2117),
.B1(n_1947),
.B2(n_1548),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2804),
.B(n_2026),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2562),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2426),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2442),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_2564),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2442),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2442),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2570),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2449),
.Y(n_3197)
);

AOI22xp5_ASAP7_75t_L g3198 ( 
.A1(n_2646),
.A2(n_2030),
.B1(n_2274),
.B2(n_2136),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2575),
.Y(n_3199)
);

INVx2_ASAP7_75t_L g3200 ( 
.A(n_2449),
.Y(n_3200)
);

INVx2_ASAP7_75t_SL g3201 ( 
.A(n_2649),
.Y(n_3201)
);

NAND2xp5_ASAP7_75t_L g3202 ( 
.A(n_2604),
.B(n_2607),
.Y(n_3202)
);

OAI22xp33_ASAP7_75t_L g3203 ( 
.A1(n_2639),
.A2(n_1549),
.B1(n_1550),
.B2(n_1543),
.Y(n_3203)
);

NOR3xp33_ASAP7_75t_L g3204 ( 
.A(n_2504),
.B(n_2019),
.C(n_1552),
.Y(n_3204)
);

BUFx3_ASAP7_75t_L g3205 ( 
.A(n_2700),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2581),
.Y(n_3206)
);

NOR2xp33_ASAP7_75t_L g3207 ( 
.A(n_2541),
.B(n_1735),
.Y(n_3207)
);

INVx2_ASAP7_75t_L g3208 ( 
.A(n_2449),
.Y(n_3208)
);

NAND3xp33_ASAP7_75t_L g3209 ( 
.A(n_2420),
.B(n_1552),
.C(n_1550),
.Y(n_3209)
);

NAND2xp5_ASAP7_75t_L g3210 ( 
.A(n_2584),
.B(n_2025),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_2588),
.B(n_2302),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_2590),
.Y(n_3212)
);

INVx8_ASAP7_75t_L g3213 ( 
.A(n_2649),
.Y(n_3213)
);

INVx3_ASAP7_75t_L g3214 ( 
.A(n_2751),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2482),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_2482),
.Y(n_3216)
);

INVx2_ASAP7_75t_L g3217 ( 
.A(n_2482),
.Y(n_3217)
);

INVx1_ASAP7_75t_SL g3218 ( 
.A(n_2638),
.Y(n_3218)
);

NAND3xp33_ASAP7_75t_L g3219 ( 
.A(n_2420),
.B(n_1566),
.C(n_1554),
.Y(n_3219)
);

BUFx6f_ASAP7_75t_L g3220 ( 
.A(n_2751),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2603),
.Y(n_3221)
);

CKINVDCx5p33_ASAP7_75t_R g3222 ( 
.A(n_2371),
.Y(n_3222)
);

HB1xp67_ASAP7_75t_L g3223 ( 
.A(n_2594),
.Y(n_3223)
);

INVx2_ASAP7_75t_L g3224 ( 
.A(n_2485),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2614),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_2627),
.Y(n_3226)
);

AO21x2_ASAP7_75t_L g3227 ( 
.A1(n_2647),
.A2(n_2106),
.B(n_2054),
.Y(n_3227)
);

HB1xp67_ASAP7_75t_L g3228 ( 
.A(n_2583),
.Y(n_3228)
);

INVx3_ASAP7_75t_L g3229 ( 
.A(n_2751),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_2630),
.B(n_2025),
.Y(n_3230)
);

INVx1_ASAP7_75t_L g3231 ( 
.A(n_2640),
.Y(n_3231)
);

INVx2_ASAP7_75t_SL g3232 ( 
.A(n_2650),
.Y(n_3232)
);

NAND2xp5_ASAP7_75t_L g3233 ( 
.A(n_2654),
.B(n_2333),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2655),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2664),
.Y(n_3235)
);

INVx2_ASAP7_75t_L g3236 ( 
.A(n_2485),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_SL g3237 ( 
.A(n_2802),
.B(n_2805),
.Y(n_3237)
);

NOR2xp33_ASAP7_75t_L g3238 ( 
.A(n_2545),
.B(n_1797),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2666),
.B(n_2333),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2485),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2667),
.Y(n_3241)
);

INVx2_ASAP7_75t_L g3242 ( 
.A(n_2502),
.Y(n_3242)
);

INVx1_ASAP7_75t_L g3243 ( 
.A(n_2745),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_2758),
.Y(n_3244)
);

INVxp67_ASAP7_75t_L g3245 ( 
.A(n_2393),
.Y(n_3245)
);

AND2x2_ASAP7_75t_L g3246 ( 
.A(n_2760),
.B(n_2211),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_2761),
.Y(n_3247)
);

AOI22xp5_ASAP7_75t_L g3248 ( 
.A1(n_2650),
.A2(n_2136),
.B1(n_2259),
.B2(n_2351),
.Y(n_3248)
);

OR2x2_ASAP7_75t_L g3249 ( 
.A(n_2612),
.B(n_1579),
.Y(n_3249)
);

INVxp33_ASAP7_75t_L g3250 ( 
.A(n_2776),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_2771),
.B(n_2163),
.Y(n_3251)
);

AND2x6_ASAP7_75t_L g3252 ( 
.A(n_2751),
.B(n_2768),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2773),
.B(n_2173),
.Y(n_3253)
);

NAND2xp33_ASAP7_75t_R g3254 ( 
.A(n_2445),
.B(n_2341),
.Y(n_3254)
);

OAI21xp33_ASAP7_75t_SL g3255 ( 
.A1(n_2778),
.A2(n_2065),
.B(n_2049),
.Y(n_3255)
);

INVx2_ASAP7_75t_L g3256 ( 
.A(n_2502),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_2784),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3011),
.Y(n_3258)
);

INVxp33_ASAP7_75t_L g3259 ( 
.A(n_3150),
.Y(n_3259)
);

INVx2_ASAP7_75t_SL g3260 ( 
.A(n_3032),
.Y(n_3260)
);

OR2x6_ASAP7_75t_L g3261 ( 
.A(n_2884),
.B(n_2741),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3028),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_3031),
.Y(n_3263)
);

NAND2xp33_ASAP7_75t_R g3264 ( 
.A(n_2838),
.B(n_2658),
.Y(n_3264)
);

OR2x2_ASAP7_75t_SL g3265 ( 
.A(n_2984),
.B(n_2467),
.Y(n_3265)
);

NOR2xp33_ASAP7_75t_L g3266 ( 
.A(n_2870),
.B(n_2735),
.Y(n_3266)
);

AOI21xp5_ASAP7_75t_L g3267 ( 
.A1(n_3084),
.A2(n_2668),
.B(n_2659),
.Y(n_3267)
);

OAI21xp5_ASAP7_75t_L g3268 ( 
.A1(n_3255),
.A2(n_2798),
.B(n_2790),
.Y(n_3268)
);

AND2x2_ASAP7_75t_L g3269 ( 
.A(n_3055),
.B(n_2399),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3055),
.B(n_2453),
.Y(n_3270)
);

NAND2xp5_ASAP7_75t_L g3271 ( 
.A(n_2853),
.B(n_2785),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3038),
.Y(n_3272)
);

XNOR2x2_ASAP7_75t_SL g3273 ( 
.A(n_2822),
.B(n_2360),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3038),
.Y(n_3274)
);

INVxp33_ASAP7_75t_L g3275 ( 
.A(n_3171),
.Y(n_3275)
);

INVx2_ASAP7_75t_SL g3276 ( 
.A(n_3032),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2816),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2864),
.B(n_2788),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3057),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_3066),
.Y(n_3280)
);

INVx1_ASAP7_75t_L g3281 ( 
.A(n_3066),
.Y(n_3281)
);

INVxp67_ASAP7_75t_SL g3282 ( 
.A(n_3125),
.Y(n_3282)
);

AND2x2_ASAP7_75t_L g3283 ( 
.A(n_2845),
.B(n_2453),
.Y(n_3283)
);

XOR2xp5_ASAP7_75t_L g3284 ( 
.A(n_2846),
.B(n_1804),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_3067),
.Y(n_3285)
);

INVx2_ASAP7_75t_L g3286 ( 
.A(n_2847),
.Y(n_3286)
);

NOR2xp33_ASAP7_75t_L g3287 ( 
.A(n_2858),
.B(n_2873),
.Y(n_3287)
);

CKINVDCx5p33_ASAP7_75t_R g3288 ( 
.A(n_2862),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3076),
.Y(n_3289)
);

AND2x2_ASAP7_75t_L g3290 ( 
.A(n_2845),
.B(n_2453),
.Y(n_3290)
);

INVx1_ASAP7_75t_L g3291 ( 
.A(n_3083),
.Y(n_3291)
);

CKINVDCx20_ASAP7_75t_R g3292 ( 
.A(n_3123),
.Y(n_3292)
);

INVx1_ASAP7_75t_L g3293 ( 
.A(n_3083),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3092),
.Y(n_3294)
);

INVxp67_ASAP7_75t_SL g3295 ( 
.A(n_3125),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2954),
.B(n_3004),
.Y(n_3296)
);

BUFx3_ASAP7_75t_L g3297 ( 
.A(n_2819),
.Y(n_3297)
);

NAND2xp33_ASAP7_75t_R g3298 ( 
.A(n_2838),
.B(n_2658),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3092),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3246),
.B(n_2791),
.Y(n_3300)
);

INVxp67_ASAP7_75t_SL g3301 ( 
.A(n_3134),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3246),
.B(n_2793),
.Y(n_3302)
);

AND2x2_ASAP7_75t_L g3303 ( 
.A(n_3078),
.B(n_2596),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3093),
.Y(n_3304)
);

NAND2xp5_ASAP7_75t_L g3305 ( 
.A(n_3141),
.B(n_2803),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_3095),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3095),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3097),
.Y(n_3308)
);

INVx2_ASAP7_75t_L g3309 ( 
.A(n_2847),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_2908),
.B(n_2735),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3097),
.Y(n_3311)
);

XNOR2x2_ASAP7_75t_L g3312 ( 
.A(n_2889),
.B(n_2360),
.Y(n_3312)
);

INVxp33_ASAP7_75t_L g3313 ( 
.A(n_2883),
.Y(n_3313)
);

XNOR2x2_ASAP7_75t_L g3314 ( 
.A(n_2889),
.B(n_2183),
.Y(n_3314)
);

BUFx6f_ASAP7_75t_L g3315 ( 
.A(n_2817),
.Y(n_3315)
);

AND2x2_ASAP7_75t_L g3316 ( 
.A(n_3082),
.B(n_2596),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3104),
.Y(n_3317)
);

NOR2xp33_ASAP7_75t_L g3318 ( 
.A(n_2944),
.B(n_2742),
.Y(n_3318)
);

CKINVDCx5p33_ASAP7_75t_R g3319 ( 
.A(n_2846),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3106),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3114),
.Y(n_3321)
);

CKINVDCx16_ASAP7_75t_R g3322 ( 
.A(n_2874),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_3114),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_3128),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_2926),
.B(n_1617),
.Y(n_3325)
);

NOR2xp33_ASAP7_75t_L g3326 ( 
.A(n_3074),
.B(n_2907),
.Y(n_3326)
);

INVx2_ASAP7_75t_L g3327 ( 
.A(n_2860),
.Y(n_3327)
);

BUFx6f_ASAP7_75t_SL g3328 ( 
.A(n_3119),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3132),
.Y(n_3329)
);

OAI21xp5_ASAP7_75t_L g3330 ( 
.A1(n_3164),
.A2(n_2412),
.B(n_2682),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_3132),
.Y(n_3331)
);

AND2x6_ASAP7_75t_L g3332 ( 
.A(n_2814),
.B(n_2653),
.Y(n_3332)
);

AND2x6_ASAP7_75t_L g3333 ( 
.A(n_2814),
.B(n_2653),
.Y(n_3333)
);

NOR2xp67_ASAP7_75t_L g3334 ( 
.A(n_3222),
.B(n_2508),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3133),
.Y(n_3335)
);

NAND2x1p5_ASAP7_75t_L g3336 ( 
.A(n_3075),
.B(n_2712),
.Y(n_3336)
);

NOR2xp33_ASAP7_75t_L g3337 ( 
.A(n_2857),
.B(n_2742),
.Y(n_3337)
);

CKINVDCx5p33_ASAP7_75t_R g3338 ( 
.A(n_2874),
.Y(n_3338)
);

XNOR2x2_ASAP7_75t_L g3339 ( 
.A(n_2889),
.B(n_2183),
.Y(n_3339)
);

CKINVDCx20_ASAP7_75t_R g3340 ( 
.A(n_2915),
.Y(n_3340)
);

NOR2xp33_ASAP7_75t_L g3341 ( 
.A(n_3023),
.B(n_2754),
.Y(n_3341)
);

INVx2_ASAP7_75t_L g3342 ( 
.A(n_2860),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3138),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_3143),
.Y(n_3344)
);

INVxp67_ASAP7_75t_L g3345 ( 
.A(n_3034),
.Y(n_3345)
);

NOR2xp33_ASAP7_75t_L g3346 ( 
.A(n_3039),
.B(n_2754),
.Y(n_3346)
);

INVxp33_ASAP7_75t_L g3347 ( 
.A(n_3124),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3143),
.Y(n_3348)
);

XOR2xp5_ASAP7_75t_L g3349 ( 
.A(n_2915),
.B(n_1831),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_3145),
.Y(n_3350)
);

INVx2_ASAP7_75t_L g3351 ( 
.A(n_2861),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3145),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_3141),
.B(n_2794),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_2861),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3156),
.Y(n_3355)
);

INVx1_ASAP7_75t_L g3356 ( 
.A(n_3156),
.Y(n_3356)
);

INVx1_ASAP7_75t_L g3357 ( 
.A(n_3157),
.Y(n_3357)
);

NAND2xp5_ASAP7_75t_SL g3358 ( 
.A(n_3075),
.B(n_2660),
.Y(n_3358)
);

OAI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_3164),
.A2(n_2743),
.B(n_2809),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3211),
.B(n_2811),
.Y(n_3360)
);

NOR2xp33_ASAP7_75t_L g3361 ( 
.A(n_3051),
.B(n_3202),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3159),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3159),
.Y(n_3363)
);

NAND2xp33_ASAP7_75t_SL g3364 ( 
.A(n_3071),
.B(n_2579),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3163),
.Y(n_3365)
);

NAND2xp33_ASAP7_75t_R g3366 ( 
.A(n_2887),
.B(n_2660),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3163),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_2817),
.Y(n_3368)
);

XNOR2x2_ASAP7_75t_L g3369 ( 
.A(n_2889),
.B(n_1948),
.Y(n_3369)
);

NAND2xp5_ASAP7_75t_L g3370 ( 
.A(n_3211),
.B(n_2675),
.Y(n_3370)
);

NOR2xp33_ASAP7_75t_L g3371 ( 
.A(n_3249),
.B(n_2755),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3181),
.Y(n_3372)
);

INVx2_ASAP7_75t_L g3373 ( 
.A(n_2863),
.Y(n_3373)
);

CKINVDCx20_ASAP7_75t_R g3374 ( 
.A(n_3013),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_3181),
.Y(n_3375)
);

INVx3_ASAP7_75t_L g3376 ( 
.A(n_3252),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3184),
.Y(n_3377)
);

CKINVDCx20_ASAP7_75t_R g3378 ( 
.A(n_3013),
.Y(n_3378)
);

NAND2x1p5_ASAP7_75t_L g3379 ( 
.A(n_3075),
.B(n_2940),
.Y(n_3379)
);

XNOR2xp5_ASAP7_75t_L g3380 ( 
.A(n_3053),
.B(n_2467),
.Y(n_3380)
);

BUFx3_ASAP7_75t_L g3381 ( 
.A(n_2819),
.Y(n_3381)
);

AND2x2_ASAP7_75t_L g3382 ( 
.A(n_3082),
.B(n_2653),
.Y(n_3382)
);

INVx2_ASAP7_75t_SL g3383 ( 
.A(n_3178),
.Y(n_3383)
);

BUFx2_ASAP7_75t_L g3384 ( 
.A(n_2832),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3062),
.B(n_2395),
.Y(n_3385)
);

NOR2xp33_ASAP7_75t_L g3386 ( 
.A(n_3249),
.B(n_2755),
.Y(n_3386)
);

INVx1_ASAP7_75t_L g3387 ( 
.A(n_3184),
.Y(n_3387)
);

XNOR2x2_ASAP7_75t_L g3388 ( 
.A(n_3161),
.B(n_1948),
.Y(n_3388)
);

NOR2xp33_ASAP7_75t_SL g3389 ( 
.A(n_3086),
.B(n_2428),
.Y(n_3389)
);

AOI21xp5_ASAP7_75t_L g3390 ( 
.A1(n_3090),
.A2(n_2681),
.B(n_2662),
.Y(n_3390)
);

NOR2xp33_ASAP7_75t_L g3391 ( 
.A(n_2973),
.B(n_2762),
.Y(n_3391)
);

INVx1_ASAP7_75t_L g3392 ( 
.A(n_3186),
.Y(n_3392)
);

INVx2_ASAP7_75t_L g3393 ( 
.A(n_2863),
.Y(n_3393)
);

INVx2_ASAP7_75t_L g3394 ( 
.A(n_2866),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3190),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3190),
.Y(n_3396)
);

XNOR2x2_ASAP7_75t_L g3397 ( 
.A(n_3161),
.B(n_2424),
.Y(n_3397)
);

INVx4_ASAP7_75t_SL g3398 ( 
.A(n_3135),
.Y(n_3398)
);

AND2x2_ASAP7_75t_L g3399 ( 
.A(n_3062),
.B(n_2457),
.Y(n_3399)
);

INVx1_ASAP7_75t_L g3400 ( 
.A(n_3193),
.Y(n_3400)
);

BUFx3_ASAP7_75t_L g3401 ( 
.A(n_2832),
.Y(n_3401)
);

NOR2xp33_ASAP7_75t_L g3402 ( 
.A(n_3036),
.B(n_2762),
.Y(n_3402)
);

NOR2xp33_ASAP7_75t_L g3403 ( 
.A(n_3050),
.B(n_2769),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3193),
.Y(n_3404)
);

OR2x6_ASAP7_75t_L g3405 ( 
.A(n_2884),
.B(n_2741),
.Y(n_3405)
);

NOR2xp33_ASAP7_75t_L g3406 ( 
.A(n_3245),
.B(n_2769),
.Y(n_3406)
);

INVx2_ASAP7_75t_L g3407 ( 
.A(n_2866),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_2937),
.B(n_2777),
.Y(n_3408)
);

INVx1_ASAP7_75t_L g3409 ( 
.A(n_3196),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_3196),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3199),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3199),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3206),
.Y(n_3413)
);

INVxp67_ASAP7_75t_SL g3414 ( 
.A(n_3134),
.Y(n_3414)
);

INVx2_ASAP7_75t_SL g3415 ( 
.A(n_2923),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3174),
.B(n_2777),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3212),
.Y(n_3417)
);

NOR2xp33_ASAP7_75t_L g3418 ( 
.A(n_3183),
.B(n_2782),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3212),
.B(n_2679),
.Y(n_3419)
);

CKINVDCx20_ASAP7_75t_R g3420 ( 
.A(n_3129),
.Y(n_3420)
);

OAI21xp5_ASAP7_75t_L g3421 ( 
.A1(n_3165),
.A2(n_3172),
.B(n_3166),
.Y(n_3421)
);

INVx1_ASAP7_75t_L g3422 ( 
.A(n_3221),
.Y(n_3422)
);

INVx1_ASAP7_75t_L g3423 ( 
.A(n_3221),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_3225),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3226),
.Y(n_3425)
);

CKINVDCx20_ASAP7_75t_R g3426 ( 
.A(n_3053),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_2996),
.B(n_2662),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_3226),
.Y(n_3428)
);

AND2x4_ASAP7_75t_L g3429 ( 
.A(n_2833),
.B(n_2712),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_3231),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_3231),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_L g3432 ( 
.A(n_3234),
.B(n_3235),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3235),
.Y(n_3433)
);

INVx1_ASAP7_75t_L g3434 ( 
.A(n_3241),
.Y(n_3434)
);

BUFx6f_ASAP7_75t_L g3435 ( 
.A(n_2833),
.Y(n_3435)
);

INVx1_ASAP7_75t_L g3436 ( 
.A(n_3241),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_3243),
.Y(n_3437)
);

CKINVDCx16_ASAP7_75t_R g3438 ( 
.A(n_2975),
.Y(n_3438)
);

INVx1_ASAP7_75t_L g3439 ( 
.A(n_3243),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_2876),
.Y(n_3440)
);

NOR2xp33_ASAP7_75t_L g3441 ( 
.A(n_3189),
.B(n_2782),
.Y(n_3441)
);

INVx2_ASAP7_75t_L g3442 ( 
.A(n_2876),
.Y(n_3442)
);

AND2x2_ASAP7_75t_L g3443 ( 
.A(n_2923),
.B(n_2767),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3244),
.Y(n_3444)
);

NOR2xp33_ASAP7_75t_L g3445 ( 
.A(n_3101),
.B(n_2642),
.Y(n_3445)
);

AND2x6_ASAP7_75t_L g3446 ( 
.A(n_2814),
.B(n_2502),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_L g3447 ( 
.A(n_2886),
.B(n_2642),
.Y(n_3447)
);

INVxp33_ASAP7_75t_L g3448 ( 
.A(n_3207),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3244),
.Y(n_3449)
);

AND2x4_ASAP7_75t_L g3450 ( 
.A(n_2868),
.B(n_2700),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_2904),
.B(n_2652),
.Y(n_3451)
);

AND2x2_ASAP7_75t_L g3452 ( 
.A(n_2972),
.B(n_2767),
.Y(n_3452)
);

NAND2xp33_ASAP7_75t_R g3453 ( 
.A(n_2887),
.B(n_2680),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3247),
.Y(n_3454)
);

XOR2xp5_ASAP7_75t_L g3455 ( 
.A(n_3153),
.B(n_1588),
.Y(n_3455)
);

NAND2xp5_ASAP7_75t_L g3456 ( 
.A(n_3247),
.B(n_2685),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3257),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3257),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_2900),
.B(n_2690),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_2948),
.Y(n_3460)
);

XOR2xp5_ASAP7_75t_L g3461 ( 
.A(n_3153),
.B(n_1601),
.Y(n_3461)
);

OR2x2_ASAP7_75t_L g3462 ( 
.A(n_2849),
.B(n_3218),
.Y(n_3462)
);

INVx1_ASAP7_75t_L g3463 ( 
.A(n_2956),
.Y(n_3463)
);

NOR2xp33_ASAP7_75t_L g3464 ( 
.A(n_3102),
.B(n_2652),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2900),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_2902),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_2902),
.Y(n_3467)
);

INVx2_ASAP7_75t_L g3468 ( 
.A(n_2892),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_2972),
.B(n_2532),
.Y(n_3469)
);

INVx1_ASAP7_75t_L g3470 ( 
.A(n_2909),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_2909),
.Y(n_3471)
);

AOI21xp5_ASAP7_75t_L g3472 ( 
.A1(n_3090),
.A2(n_2687),
.B(n_2680),
.Y(n_3472)
);

NAND2x1p5_ASAP7_75t_L g3473 ( 
.A(n_2940),
.B(n_2768),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_2911),
.Y(n_3474)
);

BUFx6f_ASAP7_75t_SL g3475 ( 
.A(n_2975),
.Y(n_3475)
);

INVx1_ASAP7_75t_L g3476 ( 
.A(n_2911),
.Y(n_3476)
);

INVx2_ASAP7_75t_L g3477 ( 
.A(n_2892),
.Y(n_3477)
);

INVx1_ASAP7_75t_L g3478 ( 
.A(n_2936),
.Y(n_3478)
);

AND2x4_ASAP7_75t_L g3479 ( 
.A(n_2868),
.B(n_2714),
.Y(n_3479)
);

INVx2_ASAP7_75t_SL g3480 ( 
.A(n_2975),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_2936),
.Y(n_3481)
);

INVx1_ASAP7_75t_SL g3482 ( 
.A(n_3180),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_2938),
.Y(n_3483)
);

INVx2_ASAP7_75t_L g3484 ( 
.A(n_2895),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_2938),
.Y(n_3485)
);

OAI21xp5_ASAP7_75t_L g3486 ( 
.A1(n_3165),
.A2(n_2593),
.B(n_2488),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_2818),
.Y(n_3487)
);

XOR2xp5_ASAP7_75t_L g3488 ( 
.A(n_2928),
.B(n_1601),
.Y(n_3488)
);

OR2x2_ASAP7_75t_SL g3489 ( 
.A(n_3228),
.B(n_2469),
.Y(n_3489)
);

NOR2xp33_ASAP7_75t_L g3490 ( 
.A(n_3034),
.B(n_2672),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_2825),
.Y(n_3491)
);

OAI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_3166),
.A2(n_3179),
.B(n_3172),
.Y(n_3492)
);

CKINVDCx14_ASAP7_75t_R g3493 ( 
.A(n_2967),
.Y(n_3493)
);

INVx1_ASAP7_75t_SL g3494 ( 
.A(n_3180),
.Y(n_3494)
);

INVx1_ASAP7_75t_L g3495 ( 
.A(n_2825),
.Y(n_3495)
);

XOR2x2_ASAP7_75t_L g3496 ( 
.A(n_3238),
.B(n_2796),
.Y(n_3496)
);

INVx1_ASAP7_75t_L g3497 ( 
.A(n_2827),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_2827),
.Y(n_3498)
);

CKINVDCx20_ASAP7_75t_R g3499 ( 
.A(n_3168),
.Y(n_3499)
);

INVx1_ASAP7_75t_L g3500 ( 
.A(n_2834),
.Y(n_3500)
);

XOR2xp5_ASAP7_75t_L g3501 ( 
.A(n_2928),
.B(n_1610),
.Y(n_3501)
);

INVx1_ASAP7_75t_L g3502 ( 
.A(n_2834),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_2837),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_2837),
.Y(n_3504)
);

AND2x4_ASAP7_75t_L g3505 ( 
.A(n_2947),
.B(n_2714),
.Y(n_3505)
);

INVx1_ASAP7_75t_L g3506 ( 
.A(n_2840),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_2840),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_2848),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_2848),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_2850),
.Y(n_3510)
);

AND2x2_ASAP7_75t_L g3511 ( 
.A(n_3035),
.B(n_2549),
.Y(n_3511)
);

CKINVDCx5p33_ASAP7_75t_R g3512 ( 
.A(n_3168),
.Y(n_3512)
);

CKINVDCx5p33_ASAP7_75t_R g3513 ( 
.A(n_3139),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_2850),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3035),
.B(n_2672),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3096),
.B(n_2558),
.Y(n_3516)
);

INVxp67_ASAP7_75t_SL g3517 ( 
.A(n_3140),
.Y(n_3517)
);

INVx4_ASAP7_75t_SL g3518 ( 
.A(n_3135),
.Y(n_3518)
);

NOR2xp33_ASAP7_75t_L g3519 ( 
.A(n_3096),
.B(n_2684),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_2859),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_2878),
.Y(n_3521)
);

INVxp67_ASAP7_75t_SL g3522 ( 
.A(n_3140),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_3115),
.B(n_2684),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3115),
.B(n_2438),
.Y(n_3524)
);

NAND2x1p5_ASAP7_75t_L g3525 ( 
.A(n_2940),
.B(n_2768),
.Y(n_3525)
);

INVx1_ASAP7_75t_L g3526 ( 
.A(n_2878),
.Y(n_3526)
);

NAND2x1p5_ASAP7_75t_L g3527 ( 
.A(n_2940),
.B(n_2768),
.Y(n_3527)
);

NAND2xp33_ASAP7_75t_R g3528 ( 
.A(n_2953),
.B(n_2681),
.Y(n_3528)
);

INVx2_ASAP7_75t_L g3529 ( 
.A(n_2896),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_2879),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_2879),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_2880),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_2880),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_2888),
.Y(n_3534)
);

INVx1_ASAP7_75t_L g3535 ( 
.A(n_2888),
.Y(n_3535)
);

AOI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3009),
.A2(n_2693),
.B(n_2687),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_2979),
.B(n_2693),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_2898),
.Y(n_3538)
);

NAND2xp33_ASAP7_75t_R g3539 ( 
.A(n_3044),
.B(n_2695),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_2898),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3210),
.Y(n_3541)
);

BUFx5_ASAP7_75t_L g3542 ( 
.A(n_3252),
.Y(n_3542)
);

CKINVDCx20_ASAP7_75t_R g3543 ( 
.A(n_3022),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3230),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3233),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3239),
.Y(n_3546)
);

INVxp67_ASAP7_75t_SL g3547 ( 
.A(n_3148),
.Y(n_3547)
);

INVx1_ASAP7_75t_L g3548 ( 
.A(n_2961),
.Y(n_3548)
);

NAND2x1_ASAP7_75t_L g3549 ( 
.A(n_3252),
.B(n_2835),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_2897),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_2961),
.Y(n_3551)
);

XOR2xp5_ASAP7_75t_L g3552 ( 
.A(n_3250),
.B(n_1610),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_2966),
.Y(n_3553)
);

INVxp33_ASAP7_75t_L g3554 ( 
.A(n_3223),
.Y(n_3554)
);

AND2x4_ASAP7_75t_L g3555 ( 
.A(n_2947),
.B(n_2587),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_2966),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_2968),
.Y(n_3557)
);

BUFx3_ASAP7_75t_L g3558 ( 
.A(n_3137),
.Y(n_3558)
);

INVx1_ASAP7_75t_L g3559 ( 
.A(n_2968),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_2970),
.Y(n_3560)
);

BUFx3_ASAP7_75t_L g3561 ( 
.A(n_3137),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_2970),
.Y(n_3562)
);

AND2x2_ASAP7_75t_L g3563 ( 
.A(n_3044),
.B(n_2259),
.Y(n_3563)
);

INVxp33_ASAP7_75t_L g3564 ( 
.A(n_3142),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_2976),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_2897),
.Y(n_3566)
);

XOR2xp5_ASAP7_75t_L g3567 ( 
.A(n_2910),
.B(n_1611),
.Y(n_3567)
);

INVx1_ASAP7_75t_L g3568 ( 
.A(n_2976),
.Y(n_3568)
);

XOR2xp5_ASAP7_75t_L g3569 ( 
.A(n_3203),
.B(n_1611),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_2985),
.Y(n_3570)
);

CKINVDCx5p33_ASAP7_75t_R g3571 ( 
.A(n_3022),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_2985),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_2988),
.Y(n_3573)
);

AND2x2_ASAP7_75t_SL g3574 ( 
.A(n_2813),
.B(n_2354),
.Y(n_3574)
);

INVx1_ASAP7_75t_L g3575 ( 
.A(n_2988),
.Y(n_3575)
);

INVx2_ASAP7_75t_SL g3576 ( 
.A(n_3019),
.Y(n_3576)
);

INVx2_ASAP7_75t_L g3577 ( 
.A(n_2901),
.Y(n_3577)
);

AND2x2_ASAP7_75t_L g3578 ( 
.A(n_3044),
.B(n_2583),
.Y(n_3578)
);

XNOR2xp5_ASAP7_75t_L g3579 ( 
.A(n_3170),
.B(n_2469),
.Y(n_3579)
);

NOR2xp33_ASAP7_75t_L g3580 ( 
.A(n_2906),
.B(n_2547),
.Y(n_3580)
);

INVx1_ASAP7_75t_L g3581 ( 
.A(n_2989),
.Y(n_3581)
);

XOR2xp5_ASAP7_75t_L g3582 ( 
.A(n_3089),
.B(n_1614),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_2989),
.Y(n_3583)
);

AND2x2_ASAP7_75t_SL g3584 ( 
.A(n_2983),
.B(n_2155),
.Y(n_3584)
);

CKINVDCx5p33_ASAP7_75t_R g3585 ( 
.A(n_3019),
.Y(n_3585)
);

INVx2_ASAP7_75t_L g3586 ( 
.A(n_2901),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_2990),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_2995),
.Y(n_3588)
);

INVx1_ASAP7_75t_L g3589 ( 
.A(n_2995),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_2998),
.Y(n_3590)
);

CKINVDCx20_ASAP7_75t_R g3591 ( 
.A(n_3019),
.Y(n_3591)
);

INVx1_ASAP7_75t_L g3592 ( 
.A(n_2998),
.Y(n_3592)
);

INVx1_ASAP7_75t_L g3593 ( 
.A(n_3000),
.Y(n_3593)
);

CKINVDCx5p33_ASAP7_75t_R g3594 ( 
.A(n_3027),
.Y(n_3594)
);

INVx1_ASAP7_75t_L g3595 ( 
.A(n_3000),
.Y(n_3595)
);

INVx1_ASAP7_75t_L g3596 ( 
.A(n_3002),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3002),
.Y(n_3597)
);

INVx1_ASAP7_75t_SL g3598 ( 
.A(n_3205),
.Y(n_3598)
);

INVx1_ASAP7_75t_L g3599 ( 
.A(n_2912),
.Y(n_3599)
);

INVx1_ASAP7_75t_L g3600 ( 
.A(n_2912),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_2913),
.Y(n_3601)
);

INVxp67_ASAP7_75t_L g3602 ( 
.A(n_3462),
.Y(n_3602)
);

INVx1_ASAP7_75t_L g3603 ( 
.A(n_3460),
.Y(n_3603)
);

NAND2xp5_ASAP7_75t_L g3604 ( 
.A(n_3296),
.B(n_2548),
.Y(n_3604)
);

O2A1O1Ixp5_ASAP7_75t_L g3605 ( 
.A1(n_3267),
.A2(n_2824),
.B(n_2830),
.C(n_2815),
.Y(n_3605)
);

INVxp67_ASAP7_75t_L g3606 ( 
.A(n_3384),
.Y(n_3606)
);

INVx2_ASAP7_75t_L g3607 ( 
.A(n_3277),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3463),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_L g3609 ( 
.A(n_3296),
.B(n_3326),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3287),
.B(n_3361),
.Y(n_3610)
);

INVxp67_ASAP7_75t_SL g3611 ( 
.A(n_3282),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_3271),
.B(n_2695),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3287),
.B(n_2548),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3361),
.B(n_2986),
.Y(n_3614)
);

INVx2_ASAP7_75t_SL g3615 ( 
.A(n_3315),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3258),
.Y(n_3616)
);

INVxp67_ASAP7_75t_SL g3617 ( 
.A(n_3282),
.Y(n_3617)
);

INVxp67_ASAP7_75t_L g3618 ( 
.A(n_3469),
.Y(n_3618)
);

INVx2_ASAP7_75t_L g3619 ( 
.A(n_3286),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3271),
.B(n_3001),
.Y(n_3620)
);

OR2x6_ASAP7_75t_L g3621 ( 
.A(n_3261),
.B(n_2884),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_3278),
.B(n_3077),
.Y(n_3622)
);

NAND2xp5_ASAP7_75t_L g3623 ( 
.A(n_3278),
.B(n_2371),
.Y(n_3623)
);

INVx3_ASAP7_75t_L g3624 ( 
.A(n_3376),
.Y(n_3624)
);

NOR2xp33_ASAP7_75t_R g3625 ( 
.A(n_3366),
.B(n_2440),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_SL g3626 ( 
.A(n_3580),
.B(n_2696),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_SL g3627 ( 
.A(n_3580),
.B(n_2696),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3266),
.B(n_2373),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_3391),
.B(n_2374),
.Y(n_3629)
);

NOR2xp33_ASAP7_75t_L g3630 ( 
.A(n_3391),
.B(n_3347),
.Y(n_3630)
);

AND2x2_ASAP7_75t_L g3631 ( 
.A(n_3445),
.B(n_2826),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_L g3632 ( 
.A1(n_3397),
.A2(n_3369),
.B1(n_3339),
.B2(n_3314),
.Y(n_3632)
);

AND2x6_ASAP7_75t_SL g3633 ( 
.A(n_3371),
.B(n_2476),
.Y(n_3633)
);

INVx1_ASAP7_75t_L g3634 ( 
.A(n_3262),
.Y(n_3634)
);

NOR2x1p5_ASAP7_75t_L g3635 ( 
.A(n_3288),
.B(n_2519),
.Y(n_3635)
);

NAND2xp5_ASAP7_75t_L g3636 ( 
.A(n_3447),
.B(n_2374),
.Y(n_3636)
);

AOI22xp33_ASAP7_75t_L g3637 ( 
.A1(n_3312),
.A2(n_2945),
.B1(n_3017),
.B2(n_3146),
.Y(n_3637)
);

NOR2xp33_ASAP7_75t_L g3638 ( 
.A(n_3445),
.B(n_3447),
.Y(n_3638)
);

INVx2_ASAP7_75t_L g3639 ( 
.A(n_3309),
.Y(n_3639)
);

INVx8_ASAP7_75t_L g3640 ( 
.A(n_3328),
.Y(n_3640)
);

INVx1_ASAP7_75t_L g3641 ( 
.A(n_3263),
.Y(n_3641)
);

INVxp67_ASAP7_75t_L g3642 ( 
.A(n_3511),
.Y(n_3642)
);

AND2x2_ASAP7_75t_L g3643 ( 
.A(n_3451),
.B(n_3147),
.Y(n_3643)
);

INVxp67_ASAP7_75t_SL g3644 ( 
.A(n_3295),
.Y(n_3644)
);

NAND2xp5_ASAP7_75t_L g3645 ( 
.A(n_3451),
.B(n_2379),
.Y(n_3645)
);

INVx3_ASAP7_75t_L g3646 ( 
.A(n_3376),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_SL g3647 ( 
.A(n_3402),
.B(n_2702),
.Y(n_3647)
);

AOI22xp5_ASAP7_75t_L g3648 ( 
.A1(n_3402),
.A2(n_3403),
.B1(n_3318),
.B2(n_3310),
.Y(n_3648)
);

AOI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3388),
.A2(n_2945),
.B1(n_3017),
.B2(n_3146),
.Y(n_3649)
);

O2A1O1Ixp33_ASAP7_75t_L g3650 ( 
.A1(n_3403),
.A2(n_2964),
.B(n_3065),
.C(n_3030),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_SL g3651 ( 
.A(n_3310),
.B(n_2702),
.Y(n_3651)
);

AND2x2_ASAP7_75t_L g3652 ( 
.A(n_3464),
.B(n_3147),
.Y(n_3652)
);

AOI22xp5_ASAP7_75t_L g3653 ( 
.A1(n_3318),
.A2(n_2499),
.B1(n_2476),
.B2(n_2389),
.Y(n_3653)
);

AND2x4_ASAP7_75t_L g3654 ( 
.A(n_3261),
.B(n_3007),
.Y(n_3654)
);

AND2x2_ASAP7_75t_L g3655 ( 
.A(n_3464),
.B(n_3147),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_SL g3656 ( 
.A(n_3416),
.B(n_2706),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_SL g3657 ( 
.A(n_3416),
.B(n_2706),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3341),
.B(n_2379),
.Y(n_3658)
);

INVx2_ASAP7_75t_SL g3659 ( 
.A(n_3315),
.Y(n_3659)
);

AOI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3341),
.A2(n_2499),
.B1(n_2392),
.B2(n_2400),
.Y(n_3660)
);

NAND2xp5_ASAP7_75t_L g3661 ( 
.A(n_3346),
.B(n_3408),
.Y(n_3661)
);

AND2x2_ASAP7_75t_L g3662 ( 
.A(n_3524),
.B(n_2392),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3418),
.B(n_2401),
.Y(n_3663)
);

INVx2_ASAP7_75t_L g3664 ( 
.A(n_3327),
.Y(n_3664)
);

OAI22xp33_ASAP7_75t_L g3665 ( 
.A1(n_3305),
.A2(n_3079),
.B1(n_2812),
.B2(n_2882),
.Y(n_3665)
);

OAI221xp5_ASAP7_75t_L g3666 ( 
.A1(n_3337),
.A2(n_2626),
.B1(n_3204),
.B2(n_2613),
.C(n_3158),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3342),
.Y(n_3667)
);

HB1xp67_ASAP7_75t_L g3668 ( 
.A(n_3345),
.Y(n_3668)
);

AND2x6_ASAP7_75t_SL g3669 ( 
.A(n_3371),
.B(n_2368),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3351),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3354),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3418),
.B(n_2644),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3272),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3441),
.B(n_2676),
.Y(n_3674)
);

NOR2xp33_ASAP7_75t_L g3675 ( 
.A(n_3441),
.B(n_2626),
.Y(n_3675)
);

NAND2xp33_ASAP7_75t_L g3676 ( 
.A(n_3542),
.B(n_2580),
.Y(n_3676)
);

INVx2_ASAP7_75t_L g3677 ( 
.A(n_3373),
.Y(n_3677)
);

NAND2xp5_ASAP7_75t_L g3678 ( 
.A(n_3541),
.B(n_3103),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3544),
.B(n_3081),
.Y(n_3679)
);

AO22x1_ASAP7_75t_L g3680 ( 
.A1(n_3513),
.A2(n_2524),
.B1(n_2525),
.B2(n_2520),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_3315),
.Y(n_3681)
);

INVx2_ASAP7_75t_L g3682 ( 
.A(n_3393),
.Y(n_3682)
);

BUFx2_ASAP7_75t_SL g3683 ( 
.A(n_3426),
.Y(n_3683)
);

AOI221xp5_ASAP7_75t_L g3684 ( 
.A1(n_3337),
.A2(n_3161),
.B1(n_3188),
.B2(n_824),
.C(n_830),
.Y(n_3684)
);

OR2x2_ASAP7_75t_L g3685 ( 
.A(n_3490),
.B(n_3515),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3385),
.B(n_2921),
.Y(n_3686)
);

OAI22xp33_ASAP7_75t_L g3687 ( 
.A1(n_3305),
.A2(n_2707),
.B1(n_3063),
.B2(n_3010),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3394),
.Y(n_3688)
);

O2A1O1Ixp33_ASAP7_75t_L g3689 ( 
.A1(n_3353),
.A2(n_3030),
.B(n_3014),
.C(n_2931),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_3515),
.B(n_3071),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_L g3691 ( 
.A(n_3399),
.B(n_2580),
.Y(n_3691)
);

INVx2_ASAP7_75t_L g3692 ( 
.A(n_3407),
.Y(n_3692)
);

AOI22xp5_ASAP7_75t_L g3693 ( 
.A1(n_3386),
.A2(n_2557),
.B1(n_2606),
.B2(n_2518),
.Y(n_3693)
);

NOR2xp67_ASAP7_75t_L g3694 ( 
.A(n_3512),
.B(n_2536),
.Y(n_3694)
);

BUFx6f_ASAP7_75t_L g3695 ( 
.A(n_3368),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3448),
.B(n_1614),
.Y(n_3696)
);

AOI22xp5_ASAP7_75t_L g3697 ( 
.A1(n_3386),
.A2(n_3406),
.B1(n_3569),
.B2(n_3389),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3574),
.A2(n_3017),
.B1(n_3161),
.B2(n_2993),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3274),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_L g3700 ( 
.A(n_3545),
.B(n_3546),
.Y(n_3700)
);

AND2x6_ASAP7_75t_L g3701 ( 
.A(n_3398),
.B(n_3007),
.Y(n_3701)
);

INVx2_ASAP7_75t_L g3702 ( 
.A(n_3440),
.Y(n_3702)
);

NOR2xp33_ASAP7_75t_L g3703 ( 
.A(n_3259),
.B(n_1620),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3516),
.B(n_3300),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_L g3705 ( 
.A(n_3300),
.B(n_3136),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3442),
.Y(n_3706)
);

INVx2_ASAP7_75t_L g3707 ( 
.A(n_3468),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_L g3708 ( 
.A(n_3302),
.B(n_2829),
.Y(n_3708)
);

OAI22xp5_ASAP7_75t_L g3709 ( 
.A1(n_3275),
.A2(n_3169),
.B1(n_2952),
.B2(n_3029),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_L g3710 ( 
.A(n_3302),
.B(n_2854),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_SL g3711 ( 
.A(n_3519),
.B(n_3085),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3353),
.B(n_2510),
.Y(n_3712)
);

AND2x2_ASAP7_75t_L g3713 ( 
.A(n_3523),
.B(n_3010),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3523),
.B(n_3010),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3360),
.B(n_2521),
.Y(n_3715)
);

AO221x1_ASAP7_75t_L g3716 ( 
.A1(n_3273),
.A2(n_3017),
.B1(n_2942),
.B2(n_2943),
.C(n_2871),
.Y(n_3716)
);

NOR3xp33_ASAP7_75t_L g3717 ( 
.A(n_3406),
.B(n_2569),
.C(n_2951),
.Y(n_3717)
);

NOR2xp33_ASAP7_75t_L g3718 ( 
.A(n_3455),
.B(n_1631),
.Y(n_3718)
);

NAND2xp5_ASAP7_75t_SL g3719 ( 
.A(n_3537),
.B(n_3116),
.Y(n_3719)
);

AND2x2_ASAP7_75t_L g3720 ( 
.A(n_3443),
.B(n_3452),
.Y(n_3720)
);

AOI22xp33_ASAP7_75t_L g3721 ( 
.A1(n_3574),
.A2(n_3567),
.B1(n_3273),
.B2(n_3290),
.Y(n_3721)
);

AOI22xp5_ASAP7_75t_L g3722 ( 
.A1(n_3264),
.A2(n_2518),
.B1(n_2606),
.B2(n_2557),
.Y(n_3722)
);

INVx1_ASAP7_75t_L g3723 ( 
.A(n_3279),
.Y(n_3723)
);

NAND2xp5_ASAP7_75t_SL g3724 ( 
.A(n_3482),
.B(n_3116),
.Y(n_3724)
);

INVx2_ASAP7_75t_L g3725 ( 
.A(n_3477),
.Y(n_3725)
);

INVx1_ASAP7_75t_L g3726 ( 
.A(n_3280),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3360),
.B(n_3122),
.Y(n_3727)
);

AND2x2_ASAP7_75t_L g3728 ( 
.A(n_3578),
.B(n_3563),
.Y(n_3728)
);

AOI21xp5_ASAP7_75t_L g3729 ( 
.A1(n_3267),
.A2(n_2930),
.B(n_2905),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3281),
.Y(n_3730)
);

INVx2_ASAP7_75t_L g3731 ( 
.A(n_3484),
.Y(n_3731)
);

NOR2xp33_ASAP7_75t_L g3732 ( 
.A(n_3461),
.B(n_1663),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_L g3733 ( 
.A(n_3283),
.B(n_3494),
.Y(n_3733)
);

NOR2xp33_ASAP7_75t_L g3734 ( 
.A(n_3284),
.B(n_1663),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_3370),
.B(n_3122),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3370),
.B(n_3130),
.Y(n_3736)
);

NAND2xp5_ASAP7_75t_L g3737 ( 
.A(n_3415),
.B(n_3432),
.Y(n_3737)
);

INVx3_ASAP7_75t_L g3738 ( 
.A(n_3379),
.Y(n_3738)
);

NOR2xp33_ASAP7_75t_L g3739 ( 
.A(n_3349),
.B(n_2618),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_L g3740 ( 
.A(n_3432),
.B(n_3130),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3269),
.B(n_3149),
.Y(n_3741)
);

AOI21xp5_ASAP7_75t_L g3742 ( 
.A1(n_3268),
.A2(n_2930),
.B(n_2905),
.Y(n_3742)
);

INVxp67_ASAP7_75t_L g3743 ( 
.A(n_3558),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_SL g3744 ( 
.A(n_3561),
.B(n_3149),
.Y(n_3744)
);

OAI22xp33_ASAP7_75t_L g3745 ( 
.A1(n_3539),
.A2(n_3063),
.B1(n_3010),
.B2(n_2869),
.Y(n_3745)
);

AOI22xp5_ASAP7_75t_L g3746 ( 
.A1(n_3264),
.A2(n_2634),
.B1(n_2524),
.B2(n_2525),
.Y(n_3746)
);

AO221x1_ASAP7_75t_L g3747 ( 
.A1(n_3368),
.A2(n_2942),
.B1(n_2943),
.B2(n_2871),
.C(n_2841),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3285),
.Y(n_3748)
);

OAI221xp5_ASAP7_75t_L g3749 ( 
.A1(n_3582),
.A2(n_3049),
.B1(n_2987),
.B2(n_3118),
.C(n_3151),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3289),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_3270),
.B(n_3160),
.Y(n_3751)
);

AOI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3584),
.A2(n_3063),
.B1(n_2701),
.B2(n_2708),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_3488),
.B(n_2634),
.Y(n_3753)
);

OAI22xp5_ASAP7_75t_SL g3754 ( 
.A1(n_3501),
.A2(n_2491),
.B1(n_2492),
.B2(n_2520),
.Y(n_3754)
);

AND2x6_ASAP7_75t_SL g3755 ( 
.A(n_3450),
.B(n_2368),
.Y(n_3755)
);

NOR2x1p5_ASAP7_75t_L g3756 ( 
.A(n_3319),
.B(n_2527),
.Y(n_3756)
);

INVx2_ASAP7_75t_L g3757 ( 
.A(n_3529),
.Y(n_3757)
);

OR2x2_ASAP7_75t_L g3758 ( 
.A(n_3297),
.B(n_3063),
.Y(n_3758)
);

AOI22xp5_ASAP7_75t_L g3759 ( 
.A1(n_3298),
.A2(n_2527),
.B1(n_2484),
.B2(n_2480),
.Y(n_3759)
);

OR2x2_ASAP7_75t_L g3760 ( 
.A(n_3381),
.B(n_2869),
.Y(n_3760)
);

NAND2xp5_ASAP7_75t_L g3761 ( 
.A(n_3303),
.B(n_3160),
.Y(n_3761)
);

NOR2xp33_ASAP7_75t_L g3762 ( 
.A(n_3325),
.B(n_3099),
.Y(n_3762)
);

NAND2xp5_ASAP7_75t_L g3763 ( 
.A(n_3316),
.B(n_3201),
.Y(n_3763)
);

NOR2xp33_ASAP7_75t_L g3764 ( 
.A(n_3564),
.B(n_3209),
.Y(n_3764)
);

AND2x2_ASAP7_75t_L g3765 ( 
.A(n_3382),
.B(n_3027),
.Y(n_3765)
);

BUFx6f_ASAP7_75t_L g3766 ( 
.A(n_3435),
.Y(n_3766)
);

NOR2xp33_ASAP7_75t_L g3767 ( 
.A(n_3554),
.B(n_3201),
.Y(n_3767)
);

CKINVDCx5p33_ASAP7_75t_R g3768 ( 
.A(n_3292),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3291),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3293),
.Y(n_3770)
);

INVx3_ASAP7_75t_L g3771 ( 
.A(n_3379),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_3401),
.B(n_3294),
.Y(n_3772)
);

AOI22xp33_ASAP7_75t_L g3773 ( 
.A1(n_3584),
.A2(n_2718),
.B1(n_2720),
.B2(n_2692),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3299),
.Y(n_3774)
);

INVx1_ASAP7_75t_L g3775 ( 
.A(n_3304),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_3390),
.B(n_3232),
.Y(n_3776)
);

AOI22xp5_ASAP7_75t_L g3777 ( 
.A1(n_3366),
.A2(n_2492),
.B1(n_2451),
.B2(n_2458),
.Y(n_3777)
);

NOR2xp33_ASAP7_75t_L g3778 ( 
.A(n_3313),
.B(n_3219),
.Y(n_3778)
);

NOR2xp33_ASAP7_75t_L g3779 ( 
.A(n_3552),
.B(n_3127),
.Y(n_3779)
);

AOI21xp5_ASAP7_75t_L g3780 ( 
.A1(n_3268),
.A2(n_2893),
.B(n_2872),
.Y(n_3780)
);

NAND2xp5_ASAP7_75t_SL g3781 ( 
.A(n_3390),
.B(n_3213),
.Y(n_3781)
);

INVx1_ASAP7_75t_L g3782 ( 
.A(n_3306),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3307),
.Y(n_3783)
);

A2O1A1Ixp33_ASAP7_75t_L g3784 ( 
.A1(n_3536),
.A2(n_3198),
.B(n_3175),
.C(n_3248),
.Y(n_3784)
);

NAND2xp5_ASAP7_75t_SL g3785 ( 
.A(n_3472),
.B(n_3213),
.Y(n_3785)
);

AOI22xp33_ASAP7_75t_L g3786 ( 
.A1(n_3496),
.A2(n_2726),
.B1(n_2730),
.B2(n_2721),
.Y(n_3786)
);

NAND2xp5_ASAP7_75t_L g3787 ( 
.A(n_3308),
.B(n_2734),
.Y(n_3787)
);

NAND2xp5_ASAP7_75t_SL g3788 ( 
.A(n_3472),
.B(n_3213),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3311),
.B(n_2734),
.Y(n_3789)
);

NAND2xp5_ASAP7_75t_SL g3790 ( 
.A(n_3322),
.B(n_3213),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_L g3791 ( 
.A(n_3317),
.B(n_2823),
.Y(n_3791)
);

NOR2xp33_ASAP7_75t_L g3792 ( 
.A(n_3479),
.B(n_3131),
.Y(n_3792)
);

AOI22xp5_ASAP7_75t_L g3793 ( 
.A1(n_3453),
.A2(n_2451),
.B1(n_2458),
.B2(n_2445),
.Y(n_3793)
);

NOR2xp33_ASAP7_75t_L g3794 ( 
.A(n_3479),
.B(n_3018),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3320),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_L g3796 ( 
.A(n_3321),
.B(n_2823),
.Y(n_3796)
);

BUFx6f_ASAP7_75t_SL g3797 ( 
.A(n_3505),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3550),
.Y(n_3798)
);

OR2x2_ASAP7_75t_L g3799 ( 
.A(n_3505),
.B(n_2869),
.Y(n_3799)
);

INVx2_ASAP7_75t_SL g3800 ( 
.A(n_3435),
.Y(n_3800)
);

OR2x2_ASAP7_75t_L g3801 ( 
.A(n_3598),
.B(n_2869),
.Y(n_3801)
);

INVx1_ASAP7_75t_L g3802 ( 
.A(n_3323),
.Y(n_3802)
);

NOR2xp33_ASAP7_75t_L g3803 ( 
.A(n_3340),
.B(n_2459),
.Y(n_3803)
);

NOR2x1p5_ASAP7_75t_L g3804 ( 
.A(n_3338),
.B(n_3008),
.Y(n_3804)
);

NAND2xp5_ASAP7_75t_L g3805 ( 
.A(n_3324),
.B(n_2823),
.Y(n_3805)
);

INVx1_ASAP7_75t_L g3806 ( 
.A(n_3329),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3331),
.Y(n_3807)
);

AND2x2_ASAP7_75t_SL g3808 ( 
.A(n_3398),
.B(n_2872),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_L g3809 ( 
.A(n_3374),
.B(n_3098),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3335),
.B(n_2957),
.Y(n_3810)
);

AOI22xp33_ASAP7_75t_L g3811 ( 
.A1(n_3332),
.A2(n_2738),
.B1(n_2744),
.B2(n_2737),
.Y(n_3811)
);

INVx4_ASAP7_75t_L g3812 ( 
.A(n_3398),
.Y(n_3812)
);

AOI22xp33_ASAP7_75t_L g3813 ( 
.A1(n_3332),
.A2(n_2632),
.B1(n_3080),
.B2(n_2461),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3343),
.Y(n_3814)
);

INVx1_ASAP7_75t_L g3815 ( 
.A(n_3344),
.Y(n_3815)
);

NOR2xp67_ASAP7_75t_L g3816 ( 
.A(n_3480),
.B(n_2536),
.Y(n_3816)
);

AND2x6_ASAP7_75t_SL g3817 ( 
.A(n_3380),
.B(n_2540),
.Y(n_3817)
);

NOR2xp33_ASAP7_75t_L g3818 ( 
.A(n_3378),
.B(n_3098),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3429),
.B(n_3098),
.Y(n_3819)
);

AOI21xp5_ASAP7_75t_L g3820 ( 
.A1(n_3330),
.A2(n_2893),
.B(n_3251),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3348),
.Y(n_3821)
);

AOI21xp5_ASAP7_75t_L g3822 ( 
.A1(n_3330),
.A2(n_3253),
.B(n_3182),
.Y(n_3822)
);

OR2x6_ASAP7_75t_L g3823 ( 
.A(n_3261),
.B(n_2884),
.Y(n_3823)
);

AOI21xp5_ASAP7_75t_L g3824 ( 
.A1(n_3419),
.A2(n_3182),
.B(n_3179),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3579),
.B(n_802),
.Y(n_3825)
);

BUFx3_ASAP7_75t_L g3826 ( 
.A(n_3499),
.Y(n_3826)
);

NOR2xp33_ASAP7_75t_L g3827 ( 
.A(n_3438),
.B(n_2645),
.Y(n_3827)
);

NOR2xp33_ASAP7_75t_L g3828 ( 
.A(n_3555),
.B(n_3021),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3350),
.B(n_2957),
.Y(n_3829)
);

OR2x6_ASAP7_75t_L g3830 ( 
.A(n_3405),
.B(n_2842),
.Y(n_3830)
);

NAND2xp5_ASAP7_75t_SL g3831 ( 
.A(n_3518),
.B(n_2957),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3352),
.Y(n_3832)
);

INVxp67_ASAP7_75t_SL g3833 ( 
.A(n_3295),
.Y(n_3833)
);

AND2x2_ASAP7_75t_L g3834 ( 
.A(n_3334),
.B(n_802),
.Y(n_3834)
);

CKINVDCx5p33_ASAP7_75t_R g3835 ( 
.A(n_3328),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3566),
.Y(n_3836)
);

NOR2xp33_ASAP7_75t_L g3837 ( 
.A(n_3555),
.B(n_3059),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_SL g3838 ( 
.A(n_3518),
.B(n_2899),
.Y(n_3838)
);

INVx2_ASAP7_75t_L g3839 ( 
.A(n_3577),
.Y(n_3839)
);

NOR2xp33_ASAP7_75t_L g3840 ( 
.A(n_3489),
.B(n_3068),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_SL g3841 ( 
.A(n_3427),
.B(n_2991),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3364),
.B(n_3033),
.Y(n_3842)
);

OR2x6_ASAP7_75t_L g3843 ( 
.A(n_3405),
.B(n_2842),
.Y(n_3843)
);

INVx2_ASAP7_75t_SL g3844 ( 
.A(n_3260),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_SL g3845 ( 
.A(n_3542),
.B(n_3237),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3421),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_L g3847 ( 
.A(n_3405),
.B(n_3072),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3355),
.B(n_1566),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_3586),
.Y(n_3849)
);

INVxp67_ASAP7_75t_L g3850 ( 
.A(n_3332),
.Y(n_3850)
);

OAI221xp5_ASAP7_75t_L g3851 ( 
.A1(n_3356),
.A2(n_830),
.B1(n_838),
.B2(n_813),
.C(n_781),
.Y(n_3851)
);

OR2x6_ASAP7_75t_L g3852 ( 
.A(n_3276),
.B(n_2842),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3357),
.Y(n_3853)
);

INVx2_ASAP7_75t_L g3854 ( 
.A(n_3487),
.Y(n_3854)
);

NAND2xp5_ASAP7_75t_SL g3855 ( 
.A(n_3542),
.B(n_2940),
.Y(n_3855)
);

BUFx5_ASAP7_75t_L g3856 ( 
.A(n_3446),
.Y(n_3856)
);

NOR2xp33_ASAP7_75t_L g3857 ( 
.A(n_3585),
.B(n_2728),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_L g3858 ( 
.A(n_3362),
.B(n_3363),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3365),
.B(n_1569),
.Y(n_3859)
);

AND2x4_ASAP7_75t_SL g3860 ( 
.A(n_3420),
.B(n_2881),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3367),
.B(n_1570),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_3372),
.B(n_1570),
.Y(n_3862)
);

NOR2xp33_ASAP7_75t_L g3863 ( 
.A(n_3594),
.B(n_2540),
.Y(n_3863)
);

NAND2xp33_ASAP7_75t_L g3864 ( 
.A(n_3542),
.B(n_3252),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_SL g3865 ( 
.A(n_3542),
.B(n_3177),
.Y(n_3865)
);

NAND2xp33_ASAP7_75t_SL g3866 ( 
.A(n_3475),
.B(n_3024),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_SL g3867 ( 
.A(n_3542),
.B(n_3177),
.Y(n_3867)
);

AOI22xp33_ASAP7_75t_SL g3868 ( 
.A1(n_3332),
.A2(n_2017),
.B1(n_3333),
.B2(n_2632),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3375),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_SL g3870 ( 
.A(n_3536),
.B(n_3177),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3576),
.B(n_3177),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3377),
.Y(n_3872)
);

INVxp67_ASAP7_75t_L g3873 ( 
.A(n_3333),
.Y(n_3873)
);

NAND2xp5_ASAP7_75t_L g3874 ( 
.A(n_3387),
.B(n_2632),
.Y(n_3874)
);

CKINVDCx5p33_ASAP7_75t_R g3875 ( 
.A(n_3475),
.Y(n_3875)
);

NAND2xp33_ASAP7_75t_L g3876 ( 
.A(n_3571),
.B(n_3252),
.Y(n_3876)
);

INVx8_ASAP7_75t_L g3877 ( 
.A(n_3333),
.Y(n_3877)
);

NAND3xp33_ASAP7_75t_L g3878 ( 
.A(n_3419),
.B(n_2196),
.C(n_2955),
.Y(n_3878)
);

BUFx6f_ASAP7_75t_L g3879 ( 
.A(n_3473),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3392),
.B(n_2632),
.Y(n_3880)
);

BUFx5_ASAP7_75t_L g3881 ( 
.A(n_3446),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_3491),
.Y(n_3882)
);

NOR2xp33_ASAP7_75t_L g3883 ( 
.A(n_3265),
.B(n_2994),
.Y(n_3883)
);

OAI22xp5_ASAP7_75t_L g3884 ( 
.A1(n_3456),
.A2(n_3459),
.B1(n_2934),
.B2(n_2881),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_3395),
.B(n_2632),
.Y(n_3885)
);

NOR2xp33_ASAP7_75t_L g3886 ( 
.A(n_3591),
.B(n_2997),
.Y(n_3886)
);

NOR2xp33_ASAP7_75t_L g3887 ( 
.A(n_3493),
.B(n_3008),
.Y(n_3887)
);

OR2x6_ASAP7_75t_L g3888 ( 
.A(n_3383),
.B(n_2842),
.Y(n_3888)
);

AOI22xp5_ASAP7_75t_L g3889 ( 
.A1(n_3333),
.A2(n_2881),
.B1(n_2934),
.B2(n_3135),
.Y(n_3889)
);

AND2x2_ASAP7_75t_SL g3890 ( 
.A(n_3528),
.B(n_2835),
.Y(n_3890)
);

NAND2x1_ASAP7_75t_L g3891 ( 
.A(n_3446),
.B(n_3252),
.Y(n_3891)
);

INVx2_ASAP7_75t_L g3892 ( 
.A(n_3495),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3336),
.B(n_3177),
.Y(n_3893)
);

CKINVDCx5p33_ASAP7_75t_R g3894 ( 
.A(n_3543),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3396),
.B(n_2461),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_3400),
.B(n_2461),
.Y(n_3896)
);

NOR2xp33_ASAP7_75t_L g3897 ( 
.A(n_3404),
.B(n_2934),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_L g3898 ( 
.A(n_3409),
.B(n_2461),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_SL g3899 ( 
.A(n_3336),
.B(n_2841),
.Y(n_3899)
);

INVx2_ASAP7_75t_L g3900 ( 
.A(n_3497),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3410),
.B(n_2461),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_L g3902 ( 
.A(n_3411),
.B(n_2461),
.Y(n_3902)
);

AOI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_3528),
.A2(n_3135),
.B1(n_3152),
.B2(n_2820),
.Y(n_3903)
);

AND2x2_ASAP7_75t_L g3904 ( 
.A(n_3412),
.B(n_802),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_3358),
.B(n_2841),
.Y(n_3905)
);

NOR2xp33_ASAP7_75t_L g3906 ( 
.A(n_3413),
.B(n_2096),
.Y(n_3906)
);

NOR2xp33_ASAP7_75t_L g3907 ( 
.A(n_3417),
.B(n_2017),
.Y(n_3907)
);

NAND2xp5_ASAP7_75t_SL g3908 ( 
.A(n_3358),
.B(n_2841),
.Y(n_3908)
);

NAND2xp5_ASAP7_75t_L g3909 ( 
.A(n_3422),
.B(n_2080),
.Y(n_3909)
);

OR2x2_ASAP7_75t_L g3910 ( 
.A(n_3423),
.B(n_2820),
.Y(n_3910)
);

AOI21xp5_ASAP7_75t_L g3911 ( 
.A1(n_3459),
.A2(n_3187),
.B(n_3185),
.Y(n_3911)
);

AND2x2_ASAP7_75t_L g3912 ( 
.A(n_3424),
.B(n_851),
.Y(n_3912)
);

NAND3xp33_ASAP7_75t_L g3913 ( 
.A(n_3425),
.B(n_3100),
.C(n_3087),
.Y(n_3913)
);

NOR2xp33_ASAP7_75t_L g3914 ( 
.A(n_3428),
.B(n_2820),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3620),
.B(n_3430),
.Y(n_3915)
);

BUFx3_ASAP7_75t_L g3916 ( 
.A(n_3640),
.Y(n_3916)
);

AO22x1_ASAP7_75t_L g3917 ( 
.A1(n_3638),
.A2(n_3152),
.B1(n_3135),
.B2(n_2831),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3610),
.B(n_3431),
.Y(n_3918)
);

INVx1_ASAP7_75t_L g3919 ( 
.A(n_3603),
.Y(n_3919)
);

INVx3_ASAP7_75t_L g3920 ( 
.A(n_3812),
.Y(n_3920)
);

NOR2xp33_ASAP7_75t_L g3921 ( 
.A(n_3609),
.B(n_838),
.Y(n_3921)
);

INVx3_ASAP7_75t_L g3922 ( 
.A(n_3812),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3608),
.Y(n_3923)
);

AOI21xp5_ASAP7_75t_L g3924 ( 
.A1(n_3676),
.A2(n_3549),
.B(n_3359),
.Y(n_3924)
);

AOI22xp33_ASAP7_75t_L g3925 ( 
.A1(n_3716),
.A2(n_2820),
.B1(n_3152),
.B2(n_2198),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3616),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3854),
.Y(n_3927)
);

INVx4_ASAP7_75t_L g3928 ( 
.A(n_3640),
.Y(n_3928)
);

OAI22xp5_ASAP7_75t_SL g3929 ( 
.A1(n_3648),
.A2(n_887),
.B1(n_933),
.B2(n_861),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3611),
.B(n_3617),
.Y(n_3930)
);

INVx4_ASAP7_75t_L g3931 ( 
.A(n_3768),
.Y(n_3931)
);

BUFx6f_ASAP7_75t_L g3932 ( 
.A(n_3695),
.Y(n_3932)
);

BUFx12f_ASAP7_75t_L g3933 ( 
.A(n_3894),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_SL g3934 ( 
.A(n_3614),
.B(n_2871),
.Y(n_3934)
);

AOI22xp5_ASAP7_75t_L g3935 ( 
.A1(n_3638),
.A2(n_3135),
.B1(n_3152),
.B2(n_3254),
.Y(n_3935)
);

AND2x2_ASAP7_75t_L g3936 ( 
.A(n_3720),
.B(n_861),
.Y(n_3936)
);

INVx2_ASAP7_75t_SL g3937 ( 
.A(n_3804),
.Y(n_3937)
);

A2O1A1Ixp33_ASAP7_75t_L g3938 ( 
.A1(n_3650),
.A2(n_3434),
.B(n_3436),
.C(n_3433),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3634),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_SL g3940 ( 
.A(n_3622),
.B(n_2871),
.Y(n_3940)
);

OAI22xp33_ASAP7_75t_L g3941 ( 
.A1(n_3684),
.A2(n_933),
.B1(n_937),
.B2(n_887),
.Y(n_3941)
);

AOI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3684),
.A2(n_3152),
.B1(n_2198),
.B2(n_2201),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_L g3943 ( 
.A(n_3611),
.B(n_3437),
.Y(n_3943)
);

NOR2xp33_ASAP7_75t_L g3944 ( 
.A(n_3604),
.B(n_937),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_L g3945 ( 
.A(n_3617),
.B(n_3439),
.Y(n_3945)
);

INVx6_ASAP7_75t_L g3946 ( 
.A(n_3695),
.Y(n_3946)
);

AOI22xp5_ASAP7_75t_L g3947 ( 
.A1(n_3631),
.A2(n_3135),
.B1(n_3152),
.B2(n_2831),
.Y(n_3947)
);

INVx5_ASAP7_75t_L g3948 ( 
.A(n_3877),
.Y(n_3948)
);

INVx2_ASAP7_75t_SL g3949 ( 
.A(n_3695),
.Y(n_3949)
);

NAND2x1p5_ASAP7_75t_L g3950 ( 
.A(n_3891),
.B(n_2855),
.Y(n_3950)
);

AND2x6_ASAP7_75t_L g3951 ( 
.A(n_3903),
.B(n_3498),
.Y(n_3951)
);

INVx2_ASAP7_75t_L g3952 ( 
.A(n_3882),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_L g3953 ( 
.A(n_3644),
.B(n_3833),
.Y(n_3953)
);

HB1xp67_ASAP7_75t_L g3954 ( 
.A(n_3668),
.Y(n_3954)
);

INVx2_ASAP7_75t_L g3955 ( 
.A(n_3892),
.Y(n_3955)
);

OR2x4_ASAP7_75t_L g3956 ( 
.A(n_3840),
.B(n_3444),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3641),
.Y(n_3957)
);

INVx2_ASAP7_75t_L g3958 ( 
.A(n_3900),
.Y(n_3958)
);

INVx2_ASAP7_75t_L g3959 ( 
.A(n_3607),
.Y(n_3959)
);

OAI22xp5_ASAP7_75t_L g3960 ( 
.A1(n_3698),
.A2(n_3449),
.B1(n_3457),
.B2(n_3454),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3644),
.B(n_3458),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3650),
.B(n_2942),
.Y(n_3962)
);

BUFx3_ASAP7_75t_L g3963 ( 
.A(n_3826),
.Y(n_3963)
);

INVx8_ASAP7_75t_L g3964 ( 
.A(n_3877),
.Y(n_3964)
);

OAI22xp5_ASAP7_75t_L g3965 ( 
.A1(n_3698),
.A2(n_3465),
.B1(n_3467),
.B2(n_3466),
.Y(n_3965)
);

AND3x2_ASAP7_75t_SL g3966 ( 
.A(n_3755),
.B(n_3669),
.C(n_3633),
.Y(n_3966)
);

AND2x4_ASAP7_75t_L g3967 ( 
.A(n_3830),
.B(n_3470),
.Y(n_3967)
);

AND2x2_ASAP7_75t_SL g3968 ( 
.A(n_3721),
.B(n_3471),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3833),
.B(n_3474),
.Y(n_3969)
);

INVx2_ASAP7_75t_SL g3970 ( 
.A(n_3766),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3704),
.B(n_3476),
.Y(n_3971)
);

NOR2xp33_ASAP7_75t_L g3972 ( 
.A(n_3613),
.B(n_1005),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3686),
.B(n_3478),
.Y(n_3973)
);

NAND2xp33_ASAP7_75t_SL g3974 ( 
.A(n_3625),
.B(n_3024),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3623),
.B(n_3481),
.Y(n_3975)
);

BUFx6f_ASAP7_75t_L g3976 ( 
.A(n_3766),
.Y(n_3976)
);

HB1xp67_ASAP7_75t_L g3977 ( 
.A(n_3606),
.Y(n_3977)
);

INVx1_ASAP7_75t_SL g3978 ( 
.A(n_3801),
.Y(n_3978)
);

A2O1A1Ixp33_ASAP7_75t_L g3979 ( 
.A1(n_3689),
.A2(n_3483),
.B(n_3485),
.C(n_3120),
.Y(n_3979)
);

NOR2xp67_ASAP7_75t_L g3980 ( 
.A(n_3759),
.B(n_2855),
.Y(n_3980)
);

NAND2xp5_ASAP7_75t_L g3981 ( 
.A(n_3708),
.B(n_3500),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3673),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3710),
.B(n_3502),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3619),
.Y(n_3984)
);

AOI22xp5_ASAP7_75t_SL g3985 ( 
.A1(n_3675),
.A2(n_1049),
.B1(n_1051),
.B2(n_1031),
.Y(n_3985)
);

BUFx2_ASAP7_75t_L g3986 ( 
.A(n_3743),
.Y(n_3986)
);

BUFx2_ASAP7_75t_L g3987 ( 
.A(n_3743),
.Y(n_3987)
);

INVx3_ASAP7_75t_L g3988 ( 
.A(n_3701),
.Y(n_3988)
);

AOI22xp33_ASAP7_75t_L g3989 ( 
.A1(n_3721),
.A2(n_3152),
.B1(n_2201),
.B2(n_2203),
.Y(n_3989)
);

INVx1_ASAP7_75t_L g3990 ( 
.A(n_3699),
.Y(n_3990)
);

BUFx6f_ASAP7_75t_L g3991 ( 
.A(n_3766),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_3672),
.B(n_3674),
.Y(n_3992)
);

BUFx4f_ASAP7_75t_L g3993 ( 
.A(n_3701),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_3697),
.B(n_2942),
.Y(n_3994)
);

HB1xp67_ASAP7_75t_L g3995 ( 
.A(n_3606),
.Y(n_3995)
);

INVxp67_ASAP7_75t_SL g3996 ( 
.A(n_3737),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_L g3997 ( 
.A(n_3740),
.B(n_3712),
.Y(n_3997)
);

INVx5_ASAP7_75t_L g3998 ( 
.A(n_3877),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3715),
.B(n_3503),
.Y(n_3999)
);

BUFx6f_ASAP7_75t_L g4000 ( 
.A(n_3701),
.Y(n_4000)
);

INVx1_ASAP7_75t_SL g4001 ( 
.A(n_3760),
.Y(n_4001)
);

INVx4_ASAP7_75t_L g4002 ( 
.A(n_3875),
.Y(n_4002)
);

BUFx6f_ASAP7_75t_L g4003 ( 
.A(n_3701),
.Y(n_4003)
);

BUFx10_ASAP7_75t_L g4004 ( 
.A(n_3803),
.Y(n_4004)
);

BUFx2_ASAP7_75t_L g4005 ( 
.A(n_3618),
.Y(n_4005)
);

INVx1_ASAP7_75t_L g4006 ( 
.A(n_3723),
.Y(n_4006)
);

INVx1_ASAP7_75t_L g4007 ( 
.A(n_3726),
.Y(n_4007)
);

INVx3_ASAP7_75t_L g4008 ( 
.A(n_3701),
.Y(n_4008)
);

BUFx3_ASAP7_75t_L g4009 ( 
.A(n_3835),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3639),
.Y(n_4010)
);

CKINVDCx5p33_ASAP7_75t_R g4011 ( 
.A(n_3817),
.Y(n_4011)
);

CKINVDCx5p33_ASAP7_75t_R g4012 ( 
.A(n_3683),
.Y(n_4012)
);

INVxp67_ASAP7_75t_SL g4013 ( 
.A(n_3772),
.Y(n_4013)
);

INVxp67_ASAP7_75t_L g4014 ( 
.A(n_3662),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3884),
.B(n_3504),
.Y(n_4015)
);

NAND2x1_ASAP7_75t_L g4016 ( 
.A(n_3747),
.B(n_3252),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_L g4017 ( 
.A(n_3661),
.B(n_3700),
.Y(n_4017)
);

OAI22xp5_ASAP7_75t_L g4018 ( 
.A1(n_3685),
.A2(n_1078),
.B1(n_1049),
.B2(n_1051),
.Y(n_4018)
);

AOI22xp33_ASAP7_75t_L g4019 ( 
.A1(n_3632),
.A2(n_2203),
.B1(n_2206),
.B2(n_2187),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3664),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3730),
.Y(n_4021)
);

NAND2x1p5_ASAP7_75t_L g4022 ( 
.A(n_3890),
.B(n_2855),
.Y(n_4022)
);

NOR2x1_ASAP7_75t_L g4023 ( 
.A(n_3842),
.B(n_3113),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_L g4024 ( 
.A(n_3602),
.B(n_3506),
.Y(n_4024)
);

BUFx3_ASAP7_75t_L g4025 ( 
.A(n_3819),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_SL g4026 ( 
.A(n_3687),
.B(n_2942),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3748),
.Y(n_4027)
);

INVx3_ASAP7_75t_L g4028 ( 
.A(n_3879),
.Y(n_4028)
);

A2O1A1Ixp33_ASAP7_75t_L g4029 ( 
.A1(n_3689),
.A2(n_3666),
.B(n_3742),
.C(n_3675),
.Y(n_4029)
);

INVx2_ASAP7_75t_L g4030 ( 
.A(n_3667),
.Y(n_4030)
);

OR2x6_ASAP7_75t_L g4031 ( 
.A(n_3621),
.B(n_3823),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3602),
.B(n_3507),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3750),
.B(n_3508),
.Y(n_4033)
);

INVx2_ASAP7_75t_L g4034 ( 
.A(n_3670),
.Y(n_4034)
);

AND2x4_ASAP7_75t_L g4035 ( 
.A(n_3830),
.B(n_3593),
.Y(n_4035)
);

OAI21xp5_ASAP7_75t_L g4036 ( 
.A1(n_3729),
.A2(n_3486),
.B(n_2831),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3769),
.B(n_3509),
.Y(n_4037)
);

AOI22xp5_ASAP7_75t_L g4038 ( 
.A1(n_3703),
.A2(n_2831),
.B1(n_2705),
.B2(n_2143),
.Y(n_4038)
);

AND2x2_ASAP7_75t_L g4039 ( 
.A(n_3728),
.B(n_1031),
.Y(n_4039)
);

INVx2_ASAP7_75t_SL g4040 ( 
.A(n_3635),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3770),
.B(n_3510),
.Y(n_4041)
);

NAND2xp5_ASAP7_75t_SL g4042 ( 
.A(n_3687),
.B(n_2943),
.Y(n_4042)
);

BUFx6f_ASAP7_75t_L g4043 ( 
.A(n_3654),
.Y(n_4043)
);

AOI22xp5_ASAP7_75t_L g4044 ( 
.A1(n_3762),
.A2(n_2831),
.B1(n_2143),
.B2(n_2216),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_SL g4045 ( 
.A(n_3665),
.B(n_2943),
.Y(n_4045)
);

OR2x6_ASAP7_75t_L g4046 ( 
.A(n_3621),
.B(n_3421),
.Y(n_4046)
);

O2A1O1Ixp33_ASAP7_75t_L g4047 ( 
.A1(n_3709),
.A2(n_743),
.B(n_754),
.C(n_735),
.Y(n_4047)
);

NAND2xp5_ASAP7_75t_L g4048 ( 
.A(n_3774),
.B(n_3775),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_3782),
.Y(n_4049)
);

INVxp67_ASAP7_75t_L g4050 ( 
.A(n_3696),
.Y(n_4050)
);

NOR2xp33_ASAP7_75t_L g4051 ( 
.A(n_3734),
.B(n_3629),
.Y(n_4051)
);

NOR2xp33_ASAP7_75t_L g4052 ( 
.A(n_3718),
.B(n_831),
.Y(n_4052)
);

NOR2xp33_ASAP7_75t_L g4053 ( 
.A(n_3732),
.B(n_832),
.Y(n_4053)
);

BUFx6f_ASAP7_75t_L g4054 ( 
.A(n_3654),
.Y(n_4054)
);

NAND3xp33_ASAP7_75t_SL g4055 ( 
.A(n_3660),
.B(n_836),
.C(n_833),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_L g4056 ( 
.A(n_3783),
.B(n_3514),
.Y(n_4056)
);

INVx6_ASAP7_75t_L g4057 ( 
.A(n_3756),
.Y(n_4057)
);

INVx2_ASAP7_75t_SL g4058 ( 
.A(n_3615),
.Y(n_4058)
);

INVx1_ASAP7_75t_L g4059 ( 
.A(n_3795),
.Y(n_4059)
);

BUFx6f_ASAP7_75t_L g4060 ( 
.A(n_3879),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_SL g4061 ( 
.A(n_3665),
.B(n_3678),
.Y(n_4061)
);

AND2x2_ASAP7_75t_L g4062 ( 
.A(n_3618),
.B(n_851),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_SL g4063 ( 
.A(n_3679),
.B(n_2943),
.Y(n_4063)
);

BUFx2_ASAP7_75t_L g4064 ( 
.A(n_3642),
.Y(n_4064)
);

NOR2xp33_ASAP7_75t_L g4065 ( 
.A(n_3628),
.B(n_840),
.Y(n_4065)
);

AOI22xp5_ASAP7_75t_L g4066 ( 
.A1(n_3749),
.A2(n_2831),
.B1(n_2143),
.B2(n_2216),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3802),
.B(n_3520),
.Y(n_4067)
);

NAND2xp33_ASAP7_75t_L g4068 ( 
.A(n_3636),
.B(n_2831),
.Y(n_4068)
);

BUFx3_ASAP7_75t_L g4069 ( 
.A(n_3887),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3806),
.B(n_3521),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_3807),
.Y(n_4071)
);

INVx3_ASAP7_75t_L g4072 ( 
.A(n_3879),
.Y(n_4072)
);

AOI22xp5_ASAP7_75t_L g4073 ( 
.A1(n_3749),
.A2(n_2143),
.B1(n_2216),
.B2(n_2184),
.Y(n_4073)
);

INVx1_ASAP7_75t_L g4074 ( 
.A(n_3814),
.Y(n_4074)
);

INVx2_ASAP7_75t_SL g4075 ( 
.A(n_3659),
.Y(n_4075)
);

AOI22xp33_ASAP7_75t_L g4076 ( 
.A1(n_3632),
.A2(n_2206),
.B1(n_2223),
.B2(n_2187),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3815),
.Y(n_4077)
);

INVx2_ASAP7_75t_L g4078 ( 
.A(n_3671),
.Y(n_4078)
);

AND2x2_ASAP7_75t_L g4079 ( 
.A(n_3642),
.B(n_851),
.Y(n_4079)
);

OAI22xp5_ASAP7_75t_SL g4080 ( 
.A1(n_3653),
.A2(n_801),
.B1(n_823),
.B2(n_755),
.Y(n_4080)
);

AOI22xp33_ASAP7_75t_L g4081 ( 
.A1(n_3637),
.A2(n_2227),
.B1(n_2230),
.B2(n_2223),
.Y(n_4081)
);

AOI22xp5_ASAP7_75t_L g4082 ( 
.A1(n_3630),
.A2(n_2143),
.B1(n_2216),
.B2(n_2184),
.Y(n_4082)
);

INVx3_ASAP7_75t_L g4083 ( 
.A(n_3621),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3821),
.B(n_3526),
.Y(n_4084)
);

INVx3_ASAP7_75t_L g4085 ( 
.A(n_3823),
.Y(n_4085)
);

INVx2_ASAP7_75t_L g4086 ( 
.A(n_3677),
.Y(n_4086)
);

CKINVDCx5p33_ASAP7_75t_R g4087 ( 
.A(n_3754),
.Y(n_4087)
);

INVx2_ASAP7_75t_L g4088 ( 
.A(n_3682),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3832),
.Y(n_4089)
);

INVx2_ASAP7_75t_SL g4090 ( 
.A(n_3681),
.Y(n_4090)
);

BUFx4f_ASAP7_75t_L g4091 ( 
.A(n_3823),
.Y(n_4091)
);

AND2x4_ASAP7_75t_L g4092 ( 
.A(n_3830),
.B(n_3583),
.Y(n_4092)
);

AOI22xp33_ASAP7_75t_SL g4093 ( 
.A1(n_3851),
.A2(n_2219),
.B1(n_2244),
.B2(n_2184),
.Y(n_4093)
);

INVx3_ASAP7_75t_L g4094 ( 
.A(n_3624),
.Y(n_4094)
);

BUFx6f_ASAP7_75t_L g4095 ( 
.A(n_3843),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3688),
.Y(n_4096)
);

INVx3_ASAP7_75t_L g4097 ( 
.A(n_3624),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3692),
.Y(n_4098)
);

INVx1_ASAP7_75t_SL g4099 ( 
.A(n_3713),
.Y(n_4099)
);

NAND2xp5_ASAP7_75t_L g4100 ( 
.A(n_3853),
.B(n_3530),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3869),
.Y(n_4101)
);

INVx4_ASAP7_75t_L g4102 ( 
.A(n_3860),
.Y(n_4102)
);

BUFx6f_ASAP7_75t_L g4103 ( 
.A(n_3843),
.Y(n_4103)
);

INVx1_ASAP7_75t_L g4104 ( 
.A(n_3872),
.Y(n_4104)
);

BUFx6f_ASAP7_75t_L g4105 ( 
.A(n_3843),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_SL g4106 ( 
.A(n_3626),
.B(n_2960),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_SL g4107 ( 
.A(n_3627),
.B(n_2960),
.Y(n_4107)
);

NAND3xp33_ASAP7_75t_SL g4108 ( 
.A(n_3666),
.B(n_843),
.C(n_842),
.Y(n_4108)
);

OR2x6_ASAP7_75t_L g4109 ( 
.A(n_3850),
.B(n_3492),
.Y(n_4109)
);

OAI22xp33_ASAP7_75t_L g4110 ( 
.A1(n_3851),
.A2(n_801),
.B1(n_823),
.B2(n_755),
.Y(n_4110)
);

OR2x4_ASAP7_75t_L g4111 ( 
.A(n_3827),
.B(n_2145),
.Y(n_4111)
);

AND2x6_ASAP7_75t_L g4112 ( 
.A(n_3889),
.B(n_3531),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_SL g4113 ( 
.A(n_3645),
.B(n_3808),
.Y(n_4113)
);

AOI22xp33_ASAP7_75t_L g4114 ( 
.A1(n_3637),
.A2(n_2230),
.B1(n_2231),
.B2(n_2227),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_3705),
.B(n_3532),
.Y(n_4115)
);

BUFx6f_ASAP7_75t_L g4116 ( 
.A(n_3852),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_3858),
.B(n_3533),
.Y(n_4117)
);

AOI22xp33_ASAP7_75t_L g4118 ( 
.A1(n_3649),
.A2(n_2235),
.B1(n_2237),
.B2(n_2231),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_3808),
.B(n_2960),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_L g4120 ( 
.A(n_3727),
.B(n_3534),
.Y(n_4120)
);

NAND2x1p5_ASAP7_75t_L g4121 ( 
.A(n_3890),
.B(n_2885),
.Y(n_4121)
);

AND2x2_ASAP7_75t_L g4122 ( 
.A(n_3643),
.B(n_871),
.Y(n_4122)
);

AOI21xp5_ASAP7_75t_L g4123 ( 
.A1(n_3864),
.A2(n_3414),
.B(n_3301),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_SL g4124 ( 
.A(n_3868),
.B(n_2960),
.Y(n_4124)
);

INVx2_ASAP7_75t_SL g4125 ( 
.A(n_3800),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_3702),
.Y(n_4126)
);

BUFx2_ASAP7_75t_L g4127 ( 
.A(n_3652),
.Y(n_4127)
);

INVx1_ASAP7_75t_L g4128 ( 
.A(n_3706),
.Y(n_4128)
);

OR2x2_ASAP7_75t_L g4129 ( 
.A(n_3733),
.B(n_3535),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_SL g4130 ( 
.A(n_3868),
.B(n_2960),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_3735),
.B(n_3538),
.Y(n_4131)
);

NAND2xp5_ASAP7_75t_L g4132 ( 
.A(n_3736),
.B(n_3540),
.Y(n_4132)
);

BUFx3_ASAP7_75t_L g4133 ( 
.A(n_3844),
.Y(n_4133)
);

AND2x6_ASAP7_75t_L g4134 ( 
.A(n_3738),
.B(n_3548),
.Y(n_4134)
);

INVx1_ASAP7_75t_SL g4135 ( 
.A(n_3714),
.Y(n_4135)
);

O2A1O1Ixp33_ASAP7_75t_L g4136 ( 
.A1(n_3612),
.A2(n_754),
.B(n_769),
.C(n_743),
.Y(n_4136)
);

INVx1_ASAP7_75t_L g4137 ( 
.A(n_3707),
.Y(n_4137)
);

BUFx6f_ASAP7_75t_L g4138 ( 
.A(n_3852),
.Y(n_4138)
);

INVxp67_ASAP7_75t_L g4139 ( 
.A(n_3778),
.Y(n_4139)
);

INVxp67_ASAP7_75t_L g4140 ( 
.A(n_3778),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_3725),
.Y(n_4141)
);

BUFx2_ASAP7_75t_L g4142 ( 
.A(n_3655),
.Y(n_4142)
);

NOR2xp33_ASAP7_75t_L g4143 ( 
.A(n_3658),
.B(n_848),
.Y(n_4143)
);

AOI22xp33_ASAP7_75t_L g4144 ( 
.A1(n_3649),
.A2(n_2237),
.B1(n_2239),
.B2(n_2235),
.Y(n_4144)
);

INVx5_ASAP7_75t_L g4145 ( 
.A(n_3852),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_3731),
.Y(n_4146)
);

A2O1A1Ixp33_ASAP7_75t_L g4147 ( 
.A1(n_3742),
.A2(n_2057),
.B(n_2127),
.C(n_2061),
.Y(n_4147)
);

NAND2xp5_ASAP7_75t_L g4148 ( 
.A(n_3914),
.B(n_3551),
.Y(n_4148)
);

INVxp67_ASAP7_75t_L g4149 ( 
.A(n_3767),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3757),
.Y(n_4150)
);

BUFx6f_ASAP7_75t_L g4151 ( 
.A(n_3888),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_3914),
.B(n_3553),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3752),
.B(n_3556),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_3798),
.Y(n_4154)
);

INVx2_ASAP7_75t_L g4155 ( 
.A(n_3836),
.Y(n_4155)
);

INVx1_ASAP7_75t_L g4156 ( 
.A(n_3839),
.Y(n_4156)
);

INVx2_ASAP7_75t_L g4157 ( 
.A(n_3849),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3752),
.B(n_3557),
.Y(n_4158)
);

INVxp67_ASAP7_75t_L g4159 ( 
.A(n_3767),
.Y(n_4159)
);

NOR3xp33_ASAP7_75t_SL g4160 ( 
.A(n_3790),
.B(n_860),
.C(n_858),
.Y(n_4160)
);

BUFx6f_ASAP7_75t_L g4161 ( 
.A(n_3888),
.Y(n_4161)
);

AND2x2_ASAP7_75t_L g4162 ( 
.A(n_3904),
.B(n_871),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_3773),
.B(n_3559),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3791),
.Y(n_4164)
);

NOR2x2_ASAP7_75t_L g4165 ( 
.A(n_3888),
.B(n_2239),
.Y(n_4165)
);

BUFx4f_ASAP7_75t_SL g4166 ( 
.A(n_3744),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3773),
.B(n_3846),
.Y(n_4167)
);

INVx1_ASAP7_75t_L g4168 ( 
.A(n_3796),
.Y(n_4168)
);

AOI22xp33_ASAP7_75t_L g4169 ( 
.A1(n_3786),
.A2(n_2245),
.B1(n_2116),
.B2(n_2118),
.Y(n_4169)
);

AND2x6_ASAP7_75t_SL g4170 ( 
.A(n_3739),
.B(n_769),
.Y(n_4170)
);

INVx2_ASAP7_75t_L g4171 ( 
.A(n_3805),
.Y(n_4171)
);

NOR3xp33_ASAP7_75t_SL g4172 ( 
.A(n_3809),
.B(n_870),
.C(n_867),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_3810),
.Y(n_4173)
);

AO22x1_ASAP7_75t_L g4174 ( 
.A1(n_3907),
.A2(n_784),
.B1(n_792),
.B2(n_772),
.Y(n_4174)
);

NAND2xp33_ASAP7_75t_L g4175 ( 
.A(n_3663),
.B(n_3054),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3846),
.B(n_3560),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_3897),
.B(n_3562),
.Y(n_4177)
);

AOI22xp5_ASAP7_75t_SL g4178 ( 
.A1(n_3753),
.A2(n_812),
.B1(n_844),
.B2(n_792),
.Y(n_4178)
);

INVx1_ASAP7_75t_L g4179 ( 
.A(n_3829),
.Y(n_4179)
);

INVx3_ASAP7_75t_L g4180 ( 
.A(n_3646),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3910),
.Y(n_4181)
);

CKINVDCx5p33_ASAP7_75t_R g4182 ( 
.A(n_3863),
.Y(n_4182)
);

NAND2xp5_ASAP7_75t_SL g4183 ( 
.A(n_3647),
.B(n_2980),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_SL g4184 ( 
.A(n_3717),
.B(n_2980),
.Y(n_4184)
);

OR2x6_ASAP7_75t_L g4185 ( 
.A(n_3850),
.B(n_3492),
.Y(n_4185)
);

INVx1_ASAP7_75t_L g4186 ( 
.A(n_3909),
.Y(n_4186)
);

HB1xp67_ASAP7_75t_L g4187 ( 
.A(n_3758),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_3787),
.B(n_3565),
.Y(n_4188)
);

BUFx6f_ASAP7_75t_L g4189 ( 
.A(n_3799),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_3913),
.Y(n_4190)
);

BUFx3_ASAP7_75t_L g4191 ( 
.A(n_3818),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_3789),
.B(n_3568),
.Y(n_4192)
);

CKINVDCx5p33_ASAP7_75t_R g4193 ( 
.A(n_3680),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3874),
.Y(n_4194)
);

NOR2xp33_ASAP7_75t_L g4195 ( 
.A(n_3722),
.B(n_3693),
.Y(n_4195)
);

NOR2xp33_ASAP7_75t_L g4196 ( 
.A(n_3764),
.B(n_876),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3745),
.B(n_3570),
.Y(n_4197)
);

OR2x6_ASAP7_75t_L g4198 ( 
.A(n_3873),
.B(n_3572),
.Y(n_4198)
);

NAND2xp5_ASAP7_75t_L g4199 ( 
.A(n_3745),
.B(n_3573),
.Y(n_4199)
);

INVx2_ASAP7_75t_L g4200 ( 
.A(n_3741),
.Y(n_4200)
);

NAND2xp5_ASAP7_75t_L g4201 ( 
.A(n_3824),
.B(n_3575),
.Y(n_4201)
);

INVx2_ASAP7_75t_L g4202 ( 
.A(n_3751),
.Y(n_4202)
);

OR2x2_ASAP7_75t_L g4203 ( 
.A(n_3690),
.B(n_3581),
.Y(n_4203)
);

AOI22xp5_ASAP7_75t_L g4204 ( 
.A1(n_3717),
.A2(n_2184),
.B1(n_2219),
.B2(n_2216),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_L g4205 ( 
.A(n_3824),
.B(n_3587),
.Y(n_4205)
);

NAND2xp5_ASAP7_75t_L g4206 ( 
.A(n_3911),
.B(n_3588),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3880),
.Y(n_4207)
);

INVx3_ASAP7_75t_L g4208 ( 
.A(n_3646),
.Y(n_4208)
);

NOR2xp33_ASAP7_75t_L g4209 ( 
.A(n_3746),
.B(n_879),
.Y(n_4209)
);

BUFx12f_ASAP7_75t_L g4210 ( 
.A(n_3834),
.Y(n_4210)
);

NAND2xp5_ASAP7_75t_L g4211 ( 
.A(n_3911),
.B(n_3589),
.Y(n_4211)
);

NAND2xp5_ASAP7_75t_SL g4212 ( 
.A(n_3873),
.B(n_2980),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_3885),
.Y(n_4213)
);

INVx4_ASAP7_75t_L g4214 ( 
.A(n_3797),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3776),
.B(n_3590),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_3847),
.B(n_3592),
.Y(n_4216)
);

INVx3_ASAP7_75t_L g4217 ( 
.A(n_3738),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3895),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_L g4219 ( 
.A(n_3847),
.B(n_3595),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_SL g4220 ( 
.A(n_3651),
.B(n_2980),
.Y(n_4220)
);

NOR2xp33_ASAP7_75t_L g4221 ( 
.A(n_3779),
.B(n_884),
.Y(n_4221)
);

NOR2xp33_ASAP7_75t_L g4222 ( 
.A(n_3779),
.B(n_3906),
.Y(n_4222)
);

BUFx6f_ASAP7_75t_L g4223 ( 
.A(n_3831),
.Y(n_4223)
);

NAND2xp5_ASAP7_75t_L g4224 ( 
.A(n_3896),
.B(n_3596),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_3761),
.Y(n_4225)
);

OR2x6_ASAP7_75t_L g4226 ( 
.A(n_3781),
.B(n_3597),
.Y(n_4226)
);

NOR2xp33_ASAP7_75t_L g4227 ( 
.A(n_3711),
.B(n_888),
.Y(n_4227)
);

NAND2x1p5_ASAP7_75t_L g4228 ( 
.A(n_3771),
.B(n_2885),
.Y(n_4228)
);

NOR2xp33_ASAP7_75t_L g4229 ( 
.A(n_3777),
.B(n_889),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_3763),
.Y(n_4230)
);

INVx1_ASAP7_75t_L g4231 ( 
.A(n_3898),
.Y(n_4231)
);

AOI22xp5_ASAP7_75t_L g4232 ( 
.A1(n_3792),
.A2(n_2184),
.B1(n_2219),
.B2(n_2216),
.Y(n_4232)
);

BUFx6f_ASAP7_75t_L g4233 ( 
.A(n_3765),
.Y(n_4233)
);

BUFx3_ASAP7_75t_L g4234 ( 
.A(n_3793),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_3901),
.Y(n_4235)
);

OAI22xp33_ASAP7_75t_L g4236 ( 
.A1(n_3691),
.A2(n_819),
.B1(n_845),
.B2(n_793),
.Y(n_4236)
);

INVx2_ASAP7_75t_L g4237 ( 
.A(n_3902),
.Y(n_4237)
);

OAI22xp5_ASAP7_75t_SL g4238 ( 
.A1(n_3857),
.A2(n_819),
.B1(n_845),
.B2(n_793),
.Y(n_4238)
);

NAND2xp5_ASAP7_75t_L g4239 ( 
.A(n_3841),
.B(n_3547),
.Y(n_4239)
);

HB1xp67_ASAP7_75t_L g4240 ( 
.A(n_3792),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_3794),
.Y(n_4241)
);

INVx1_ASAP7_75t_L g4242 ( 
.A(n_3794),
.Y(n_4242)
);

AOI21xp5_ASAP7_75t_L g4243 ( 
.A1(n_3780),
.A2(n_3820),
.B(n_3876),
.Y(n_4243)
);

A2O1A1Ixp33_ASAP7_75t_L g4244 ( 
.A1(n_3784),
.A2(n_2061),
.B(n_2140),
.C(n_2127),
.Y(n_4244)
);

CKINVDCx5p33_ASAP7_75t_R g4245 ( 
.A(n_3797),
.Y(n_4245)
);

AND2x2_ASAP7_75t_L g4246 ( 
.A(n_3912),
.B(n_871),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_3719),
.Y(n_4247)
);

HB1xp67_ASAP7_75t_L g4248 ( 
.A(n_3724),
.Y(n_4248)
);

BUFx2_ASAP7_75t_L g4249 ( 
.A(n_3866),
.Y(n_4249)
);

NAND2xp5_ASAP7_75t_L g4250 ( 
.A(n_3780),
.B(n_3547),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_SL g4251 ( 
.A(n_3811),
.B(n_3015),
.Y(n_4251)
);

BUFx2_ASAP7_75t_L g4252 ( 
.A(n_3828),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_3785),
.B(n_3301),
.Y(n_4253)
);

NOR2xp33_ASAP7_75t_L g4254 ( 
.A(n_3886),
.B(n_890),
.Y(n_4254)
);

INVx4_ASAP7_75t_L g4255 ( 
.A(n_3928),
.Y(n_4255)
);

AND2x2_ASAP7_75t_L g4256 ( 
.A(n_4127),
.B(n_3883),
.Y(n_4256)
);

BUFx6f_ASAP7_75t_L g4257 ( 
.A(n_4043),
.Y(n_4257)
);

INVx4_ASAP7_75t_L g4258 ( 
.A(n_3928),
.Y(n_4258)
);

INVx1_ASAP7_75t_SL g4259 ( 
.A(n_4249),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_3996),
.B(n_3822),
.Y(n_4260)
);

AOI22xp33_ASAP7_75t_L g4261 ( 
.A1(n_3929),
.A2(n_3825),
.B1(n_3813),
.B2(n_3657),
.Y(n_4261)
);

INVx3_ASAP7_75t_SL g4262 ( 
.A(n_4245),
.Y(n_4262)
);

AND2x4_ASAP7_75t_L g4263 ( 
.A(n_4031),
.B(n_3816),
.Y(n_4263)
);

AND2x4_ASAP7_75t_L g4264 ( 
.A(n_4031),
.B(n_3788),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_3997),
.B(n_3822),
.Y(n_4265)
);

INVx1_ASAP7_75t_L g4266 ( 
.A(n_4048),
.Y(n_4266)
);

NAND2xp5_ASAP7_75t_L g4267 ( 
.A(n_3997),
.B(n_3820),
.Y(n_4267)
);

INVxp67_ASAP7_75t_L g4268 ( 
.A(n_3954),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3943),
.B(n_3656),
.Y(n_4269)
);

BUFx2_ASAP7_75t_L g4270 ( 
.A(n_3986),
.Y(n_4270)
);

INVx5_ASAP7_75t_L g4271 ( 
.A(n_4134),
.Y(n_4271)
);

CKINVDCx5p33_ASAP7_75t_R g4272 ( 
.A(n_3933),
.Y(n_4272)
);

NAND2xp5_ASAP7_75t_L g4273 ( 
.A(n_3943),
.B(n_3870),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4142),
.B(n_3837),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_3945),
.B(n_3856),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_3927),
.Y(n_4276)
);

INVx2_ASAP7_75t_L g4277 ( 
.A(n_3952),
.Y(n_4277)
);

INVx3_ASAP7_75t_L g4278 ( 
.A(n_4198),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_3945),
.B(n_3856),
.Y(n_4279)
);

NAND2xp5_ASAP7_75t_L g4280 ( 
.A(n_3961),
.B(n_3856),
.Y(n_4280)
);

OR2x4_ASAP7_75t_L g4281 ( 
.A(n_4195),
.B(n_3848),
.Y(n_4281)
);

INVx5_ASAP7_75t_L g4282 ( 
.A(n_4134),
.Y(n_4282)
);

AO21x2_ASAP7_75t_L g4283 ( 
.A1(n_4123),
.A2(n_3908),
.B(n_3905),
.Y(n_4283)
);

AND2x6_ASAP7_75t_L g4284 ( 
.A(n_4000),
.B(n_3771),
.Y(n_4284)
);

BUFx6f_ASAP7_75t_L g4285 ( 
.A(n_4043),
.Y(n_4285)
);

INVx1_ASAP7_75t_L g4286 ( 
.A(n_3926),
.Y(n_4286)
);

NOR2xp33_ASAP7_75t_R g4287 ( 
.A(n_4182),
.B(n_3859),
.Y(n_4287)
);

NAND2xp5_ASAP7_75t_L g4288 ( 
.A(n_3961),
.B(n_3856),
.Y(n_4288)
);

BUFx3_ASAP7_75t_L g4289 ( 
.A(n_4069),
.Y(n_4289)
);

BUFx6f_ASAP7_75t_L g4290 ( 
.A(n_4043),
.Y(n_4290)
);

INVx3_ASAP7_75t_L g4291 ( 
.A(n_4198),
.Y(n_4291)
);

NAND3xp33_ASAP7_75t_SL g4292 ( 
.A(n_4047),
.B(n_3813),
.C(n_3861),
.Y(n_4292)
);

BUFx2_ASAP7_75t_L g4293 ( 
.A(n_3987),
.Y(n_4293)
);

AOI22xp33_ASAP7_75t_L g4294 ( 
.A1(n_3968),
.A2(n_3599),
.B1(n_3601),
.B2(n_3600),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_3939),
.Y(n_4295)
);

BUFx2_ASAP7_75t_L g4296 ( 
.A(n_4005),
.Y(n_4296)
);

AND2x2_ASAP7_75t_L g4297 ( 
.A(n_4240),
.B(n_4064),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_3957),
.Y(n_4298)
);

OR2x6_ASAP7_75t_L g4299 ( 
.A(n_4031),
.B(n_3838),
.Y(n_4299)
);

NOR2xp33_ASAP7_75t_R g4300 ( 
.A(n_4193),
.B(n_3862),
.Y(n_4300)
);

NAND2xp5_ASAP7_75t_L g4301 ( 
.A(n_3969),
.B(n_3856),
.Y(n_4301)
);

NAND2xp5_ASAP7_75t_SL g4302 ( 
.A(n_4017),
.B(n_3980),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_3969),
.B(n_3856),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_3955),
.Y(n_4304)
);

INVx2_ASAP7_75t_L g4305 ( 
.A(n_3958),
.Y(n_4305)
);

BUFx6f_ASAP7_75t_L g4306 ( 
.A(n_4054),
.Y(n_4306)
);

INVx3_ASAP7_75t_L g4307 ( 
.A(n_4198),
.Y(n_4307)
);

AND2x4_ASAP7_75t_L g4308 ( 
.A(n_4099),
.B(n_3871),
.Y(n_4308)
);

NOR2xp33_ASAP7_75t_L g4309 ( 
.A(n_4051),
.B(n_3694),
.Y(n_4309)
);

AND2x6_ASAP7_75t_SL g4310 ( 
.A(n_4222),
.B(n_772),
.Y(n_4310)
);

INVx2_ASAP7_75t_SL g4311 ( 
.A(n_3916),
.Y(n_4311)
);

INVx1_ASAP7_75t_SL g4312 ( 
.A(n_4165),
.Y(n_4312)
);

AO21x2_ASAP7_75t_L g4313 ( 
.A1(n_3935),
.A2(n_3845),
.B(n_3227),
.Y(n_4313)
);

AND2x4_ASAP7_75t_L g4314 ( 
.A(n_4099),
.B(n_3899),
.Y(n_4314)
);

INVx1_ASAP7_75t_L g4315 ( 
.A(n_3982),
.Y(n_4315)
);

AND2x2_ASAP7_75t_L g4316 ( 
.A(n_4241),
.B(n_784),
.Y(n_4316)
);

INVx3_ASAP7_75t_L g4317 ( 
.A(n_3967),
.Y(n_4317)
);

INVx2_ASAP7_75t_L g4318 ( 
.A(n_3959),
.Y(n_4318)
);

OR2x2_ASAP7_75t_L g4319 ( 
.A(n_4135),
.B(n_1417),
.Y(n_4319)
);

AOI22xp33_ASAP7_75t_L g4320 ( 
.A1(n_3941),
.A2(n_2245),
.B1(n_2116),
.B2(n_2118),
.Y(n_4320)
);

INVx1_ASAP7_75t_L g4321 ( 
.A(n_3990),
.Y(n_4321)
);

BUFx10_ASAP7_75t_L g4322 ( 
.A(n_4057),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_SL g4323 ( 
.A(n_4139),
.B(n_3881),
.Y(n_4323)
);

CKINVDCx5p33_ASAP7_75t_R g4324 ( 
.A(n_4012),
.Y(n_4324)
);

INVx3_ASAP7_75t_L g4325 ( 
.A(n_3967),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_4061),
.B(n_3881),
.Y(n_4326)
);

BUFx6f_ASAP7_75t_L g4327 ( 
.A(n_4054),
.Y(n_4327)
);

A2O1A1Ixp33_ASAP7_75t_L g4328 ( 
.A1(n_3921),
.A2(n_3878),
.B(n_3605),
.C(n_796),
.Y(n_4328)
);

AOI22xp33_ASAP7_75t_L g4329 ( 
.A1(n_3989),
.A2(n_4108),
.B1(n_4080),
.B2(n_4110),
.Y(n_4329)
);

NAND2xp5_ASAP7_75t_SL g4330 ( 
.A(n_4140),
.B(n_3881),
.Y(n_4330)
);

INVx2_ASAP7_75t_SL g4331 ( 
.A(n_4057),
.Y(n_4331)
);

INVx2_ASAP7_75t_L g4332 ( 
.A(n_3984),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4010),
.Y(n_4333)
);

INVxp67_ASAP7_75t_L g4334 ( 
.A(n_4190),
.Y(n_4334)
);

INVx2_ASAP7_75t_SL g4335 ( 
.A(n_3963),
.Y(n_4335)
);

BUFx6f_ASAP7_75t_L g4336 ( 
.A(n_4054),
.Y(n_4336)
);

AND2x4_ASAP7_75t_SL g4337 ( 
.A(n_4102),
.B(n_2885),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_4013),
.B(n_3881),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_L g4339 ( 
.A(n_4176),
.B(n_3881),
.Y(n_4339)
);

INVx4_ASAP7_75t_L g4340 ( 
.A(n_3932),
.Y(n_4340)
);

AOI21xp5_ASAP7_75t_L g4341 ( 
.A1(n_4243),
.A2(n_3517),
.B(n_3414),
.Y(n_4341)
);

INVx3_ASAP7_75t_L g4342 ( 
.A(n_4233),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4006),
.Y(n_4343)
);

INVx2_ASAP7_75t_L g4344 ( 
.A(n_4020),
.Y(n_4344)
);

AND2x4_ASAP7_75t_L g4345 ( 
.A(n_4135),
.B(n_3893),
.Y(n_4345)
);

INVx3_ASAP7_75t_L g4346 ( 
.A(n_4233),
.Y(n_4346)
);

INVx5_ASAP7_75t_L g4347 ( 
.A(n_4134),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_3978),
.B(n_3855),
.Y(n_4348)
);

INVx2_ASAP7_75t_L g4349 ( 
.A(n_4030),
.Y(n_4349)
);

AOI22xp5_ASAP7_75t_L g4350 ( 
.A1(n_4238),
.A2(n_2219),
.B1(n_2244),
.B2(n_2184),
.Y(n_4350)
);

AND2x4_ASAP7_75t_L g4351 ( 
.A(n_3978),
.B(n_4001),
.Y(n_4351)
);

INVx2_ASAP7_75t_L g4352 ( 
.A(n_4034),
.Y(n_4352)
);

INVx1_ASAP7_75t_L g4353 ( 
.A(n_4007),
.Y(n_4353)
);

NAND2xp33_ASAP7_75t_SL g4354 ( 
.A(n_3937),
.B(n_3015),
.Y(n_4354)
);

BUFx6f_ASAP7_75t_L g4355 ( 
.A(n_4000),
.Y(n_4355)
);

AOI22xp5_ASAP7_75t_L g4356 ( 
.A1(n_4196),
.A2(n_2244),
.B1(n_2219),
.B2(n_894),
.Y(n_4356)
);

AOI22xp5_ASAP7_75t_L g4357 ( 
.A1(n_4221),
.A2(n_2244),
.B1(n_2219),
.B2(n_894),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_4176),
.B(n_3517),
.Y(n_4358)
);

INVx4_ASAP7_75t_L g4359 ( 
.A(n_3932),
.Y(n_4359)
);

INVx5_ASAP7_75t_L g4360 ( 
.A(n_4134),
.Y(n_4360)
);

INVx1_ASAP7_75t_SL g4361 ( 
.A(n_4252),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4021),
.Y(n_4362)
);

BUFx6f_ASAP7_75t_L g4363 ( 
.A(n_4000),
.Y(n_4363)
);

BUFx6f_ASAP7_75t_L g4364 ( 
.A(n_4003),
.Y(n_4364)
);

BUFx6f_ASAP7_75t_L g4365 ( 
.A(n_4003),
.Y(n_4365)
);

NOR2xp33_ASAP7_75t_L g4366 ( 
.A(n_4052),
.B(n_891),
.Y(n_4366)
);

HB1xp67_ASAP7_75t_L g4367 ( 
.A(n_3977),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_4078),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_3930),
.B(n_3522),
.Y(n_4369)
);

NOR3xp33_ASAP7_75t_SL g4370 ( 
.A(n_4055),
.B(n_4011),
.C(n_4065),
.Y(n_4370)
);

INVx2_ASAP7_75t_L g4371 ( 
.A(n_4086),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_4088),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4027),
.Y(n_4373)
);

BUFx4f_ASAP7_75t_L g4374 ( 
.A(n_4003),
.Y(n_4374)
);

NAND2xp5_ASAP7_75t_L g4375 ( 
.A(n_3930),
.B(n_3522),
.Y(n_4375)
);

HB1xp67_ASAP7_75t_L g4376 ( 
.A(n_3995),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_3953),
.B(n_4115),
.Y(n_4377)
);

INVx2_ASAP7_75t_L g4378 ( 
.A(n_4096),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4049),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_SL g4380 ( 
.A(n_4191),
.B(n_3605),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_4098),
.Y(n_4381)
);

AOI22xp5_ASAP7_75t_L g4382 ( 
.A1(n_4174),
.A2(n_2244),
.B1(n_894),
.B2(n_903),
.Y(n_4382)
);

OAI21xp5_ASAP7_75t_L g4383 ( 
.A1(n_4029),
.A2(n_3867),
.B(n_3865),
.Y(n_4383)
);

BUFx2_ASAP7_75t_L g4384 ( 
.A(n_4025),
.Y(n_4384)
);

BUFx12f_ASAP7_75t_SL g4385 ( 
.A(n_3931),
.Y(n_4385)
);

NAND2xp33_ASAP7_75t_SL g4386 ( 
.A(n_4160),
.B(n_3015),
.Y(n_4386)
);

INVx1_ASAP7_75t_L g4387 ( 
.A(n_4059),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_L g4388 ( 
.A(n_3953),
.B(n_3109),
.Y(n_4388)
);

OAI22xp5_ASAP7_75t_L g4389 ( 
.A1(n_3942),
.A2(n_806),
.B1(n_808),
.B2(n_795),
.Y(n_4389)
);

NOR2xp33_ASAP7_75t_R g4390 ( 
.A(n_3974),
.B(n_3229),
.Y(n_4390)
);

BUFx3_ASAP7_75t_L g4391 ( 
.A(n_4133),
.Y(n_4391)
);

BUFx2_ASAP7_75t_L g4392 ( 
.A(n_3956),
.Y(n_4392)
);

HB1xp67_ASAP7_75t_L g4393 ( 
.A(n_4216),
.Y(n_4393)
);

INVx3_ASAP7_75t_L g4394 ( 
.A(n_4233),
.Y(n_4394)
);

INVx4_ASAP7_75t_L g4395 ( 
.A(n_3932),
.Y(n_4395)
);

OR2x6_ASAP7_75t_L g4396 ( 
.A(n_4046),
.B(n_3473),
.Y(n_4396)
);

CKINVDCx5p33_ASAP7_75t_R g4397 ( 
.A(n_4009),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4071),
.Y(n_4398)
);

INVx1_ASAP7_75t_L g4399 ( 
.A(n_4074),
.Y(n_4399)
);

AND2x2_ASAP7_75t_L g4400 ( 
.A(n_4242),
.B(n_4200),
.Y(n_4400)
);

INVx3_ASAP7_75t_L g4401 ( 
.A(n_3976),
.Y(n_4401)
);

OAI21xp5_ASAP7_75t_L g4402 ( 
.A1(n_4244),
.A2(n_2935),
.B(n_2865),
.Y(n_4402)
);

NOR2x1_ASAP7_75t_L g4403 ( 
.A(n_3992),
.B(n_2903),
.Y(n_4403)
);

NOR2xp33_ASAP7_75t_R g4404 ( 
.A(n_4087),
.B(n_3229),
.Y(n_4404)
);

NOR3xp33_ASAP7_75t_SL g4405 ( 
.A(n_4143),
.B(n_893),
.C(n_892),
.Y(n_4405)
);

INVx3_ASAP7_75t_L g4406 ( 
.A(n_3976),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_4115),
.B(n_3109),
.Y(n_4407)
);

NOR2xp33_ASAP7_75t_L g4408 ( 
.A(n_4053),
.B(n_896),
.Y(n_4408)
);

NOR2xp33_ASAP7_75t_R g4409 ( 
.A(n_4166),
.B(n_3229),
.Y(n_4409)
);

INVx3_ASAP7_75t_L g4410 ( 
.A(n_3976),
.Y(n_4410)
);

O2A1O1Ixp33_ASAP7_75t_L g4411 ( 
.A1(n_4018),
.A2(n_809),
.B(n_810),
.C(n_808),
.Y(n_4411)
);

AND2x4_ASAP7_75t_L g4412 ( 
.A(n_4001),
.B(n_2903),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_4155),
.Y(n_4413)
);

INVx2_ASAP7_75t_L g4414 ( 
.A(n_4157),
.Y(n_4414)
);

CKINVDCx11_ASAP7_75t_R g4415 ( 
.A(n_4004),
.Y(n_4415)
);

NAND2xp5_ASAP7_75t_SL g4416 ( 
.A(n_4234),
.B(n_3015),
.Y(n_4416)
);

BUFx4f_ASAP7_75t_SL g4417 ( 
.A(n_4210),
.Y(n_4417)
);

INVx2_ASAP7_75t_L g4418 ( 
.A(n_4126),
.Y(n_4418)
);

NAND2xp5_ASAP7_75t_SL g4419 ( 
.A(n_4023),
.B(n_3037),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_SL g4420 ( 
.A(n_3991),
.B(n_3037),
.Y(n_4420)
);

BUFx6f_ASAP7_75t_L g4421 ( 
.A(n_3991),
.Y(n_4421)
);

BUFx2_ASAP7_75t_L g4422 ( 
.A(n_3956),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4077),
.Y(n_4423)
);

AND2x2_ASAP7_75t_L g4424 ( 
.A(n_4202),
.B(n_809),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4120),
.B(n_3227),
.Y(n_4425)
);

AND2x4_ASAP7_75t_SL g4426 ( 
.A(n_4102),
.B(n_2929),
.Y(n_4426)
);

AND3x1_ASAP7_75t_L g4427 ( 
.A(n_4172),
.B(n_812),
.C(n_810),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4089),
.Y(n_4428)
);

AOI211xp5_ASAP7_75t_L g4429 ( 
.A1(n_4018),
.A2(n_826),
.B(n_834),
.C(n_821),
.Y(n_4429)
);

INVx5_ASAP7_75t_L g4430 ( 
.A(n_4046),
.Y(n_4430)
);

INVx2_ASAP7_75t_L g4431 ( 
.A(n_4128),
.Y(n_4431)
);

OR2x6_ASAP7_75t_L g4432 ( 
.A(n_4046),
.B(n_3525),
.Y(n_4432)
);

HB1xp67_ASAP7_75t_L g4433 ( 
.A(n_4216),
.Y(n_4433)
);

AND2x2_ASAP7_75t_L g4434 ( 
.A(n_4225),
.B(n_821),
.Y(n_4434)
);

OR2x6_ASAP7_75t_L g4435 ( 
.A(n_4109),
.B(n_3525),
.Y(n_4435)
);

XNOR2xp5_ASAP7_75t_L g4436 ( 
.A(n_3985),
.B(n_8),
.Y(n_4436)
);

NAND2xp5_ASAP7_75t_L g4437 ( 
.A(n_4120),
.B(n_2080),
.Y(n_4437)
);

AND2x2_ASAP7_75t_L g4438 ( 
.A(n_4230),
.B(n_826),
.Y(n_4438)
);

OAI22xp5_ASAP7_75t_L g4439 ( 
.A1(n_4073),
.A2(n_835),
.B1(n_837),
.B2(n_834),
.Y(n_4439)
);

NAND2xp5_ASAP7_75t_SL g4440 ( 
.A(n_4149),
.B(n_3037),
.Y(n_4440)
);

AND2x2_ASAP7_75t_L g4441 ( 
.A(n_4159),
.B(n_835),
.Y(n_4441)
);

INVx2_ASAP7_75t_L g4442 ( 
.A(n_4137),
.Y(n_4442)
);

AND2x4_ASAP7_75t_L g4443 ( 
.A(n_4083),
.B(n_2929),
.Y(n_4443)
);

INVx1_ASAP7_75t_L g4444 ( 
.A(n_4101),
.Y(n_4444)
);

INVx2_ASAP7_75t_L g4445 ( 
.A(n_4141),
.Y(n_4445)
);

BUFx6f_ASAP7_75t_L g4446 ( 
.A(n_4091),
.Y(n_4446)
);

NOR2xp33_ASAP7_75t_R g4447 ( 
.A(n_4040),
.B(n_2852),
.Y(n_4447)
);

NAND2xp5_ASAP7_75t_L g4448 ( 
.A(n_4131),
.B(n_2081),
.Y(n_4448)
);

NAND2xp5_ASAP7_75t_L g4449 ( 
.A(n_4131),
.B(n_2081),
.Y(n_4449)
);

INVx2_ASAP7_75t_SL g4450 ( 
.A(n_3946),
.Y(n_4450)
);

AOI22xp5_ASAP7_75t_L g4451 ( 
.A1(n_4254),
.A2(n_2244),
.B1(n_903),
.B2(n_957),
.Y(n_4451)
);

NAND2xp5_ASAP7_75t_L g4452 ( 
.A(n_4132),
.B(n_2091),
.Y(n_4452)
);

HB1xp67_ASAP7_75t_L g4453 ( 
.A(n_4219),
.Y(n_4453)
);

AO22x1_ASAP7_75t_L g4454 ( 
.A1(n_4214),
.A2(n_841),
.B1(n_844),
.B2(n_837),
.Y(n_4454)
);

INVx2_ASAP7_75t_L g4455 ( 
.A(n_4146),
.Y(n_4455)
);

INVx2_ASAP7_75t_SL g4456 ( 
.A(n_3946),
.Y(n_4456)
);

HB1xp67_ASAP7_75t_L g4457 ( 
.A(n_4219),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4104),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_4132),
.B(n_2091),
.Y(n_4459)
);

INVx1_ASAP7_75t_L g4460 ( 
.A(n_3919),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_SL g4461 ( 
.A(n_4223),
.B(n_3037),
.Y(n_4461)
);

INVx1_ASAP7_75t_L g4462 ( 
.A(n_3923),
.Y(n_4462)
);

AND2x4_ASAP7_75t_L g4463 ( 
.A(n_4083),
.B(n_2929),
.Y(n_4463)
);

NAND2xp5_ASAP7_75t_L g4464 ( 
.A(n_3915),
.B(n_2158),
.Y(n_4464)
);

INVxp67_ASAP7_75t_L g4465 ( 
.A(n_4184),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_SL g4466 ( 
.A(n_4223),
.B(n_3144),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_3915),
.B(n_2158),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4150),
.Y(n_4468)
);

HB1xp67_ASAP7_75t_L g4469 ( 
.A(n_4203),
.Y(n_4469)
);

NOR3xp33_ASAP7_75t_SL g4470 ( 
.A(n_4229),
.B(n_904),
.C(n_902),
.Y(n_4470)
);

OR2x6_ASAP7_75t_L g4471 ( 
.A(n_4109),
.B(n_3527),
.Y(n_4471)
);

NAND2xp5_ASAP7_75t_L g4472 ( 
.A(n_3918),
.B(n_2179),
.Y(n_4472)
);

NOR3xp33_ASAP7_75t_SL g4473 ( 
.A(n_4209),
.B(n_906),
.C(n_905),
.Y(n_4473)
);

OAI22xp33_ASAP7_75t_L g4474 ( 
.A1(n_4066),
.A2(n_874),
.B1(n_921),
.B2(n_855),
.Y(n_4474)
);

CKINVDCx5p33_ASAP7_75t_R g4475 ( 
.A(n_4002),
.Y(n_4475)
);

HB1xp67_ASAP7_75t_L g4476 ( 
.A(n_4239),
.Y(n_4476)
);

INVx2_ASAP7_75t_L g4477 ( 
.A(n_4154),
.Y(n_4477)
);

NOR2xp33_ASAP7_75t_L g4478 ( 
.A(n_4050),
.B(n_908),
.Y(n_4478)
);

BUFx2_ASAP7_75t_L g4479 ( 
.A(n_4248),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4033),
.Y(n_4480)
);

AND2x4_ASAP7_75t_L g4481 ( 
.A(n_4085),
.B(n_2933),
.Y(n_4481)
);

NAND2xp5_ASAP7_75t_L g4482 ( 
.A(n_3918),
.B(n_2179),
.Y(n_4482)
);

OR2x6_ASAP7_75t_L g4483 ( 
.A(n_4109),
.B(n_3527),
.Y(n_4483)
);

OR2x6_ASAP7_75t_SL g4484 ( 
.A(n_3966),
.B(n_913),
.Y(n_4484)
);

INVx5_ASAP7_75t_L g4485 ( 
.A(n_3988),
.Y(n_4485)
);

NAND2xp5_ASAP7_75t_SL g4486 ( 
.A(n_4223),
.B(n_3144),
.Y(n_4486)
);

NAND2xp5_ASAP7_75t_L g4487 ( 
.A(n_3981),
.B(n_2202),
.Y(n_4487)
);

CKINVDCx5p33_ASAP7_75t_R g4488 ( 
.A(n_4002),
.Y(n_4488)
);

NAND2xp5_ASAP7_75t_SL g4489 ( 
.A(n_4015),
.B(n_3144),
.Y(n_4489)
);

AOI21xp5_ASAP7_75t_L g4490 ( 
.A1(n_4250),
.A2(n_4016),
.B(n_4036),
.Y(n_4490)
);

INVx3_ASAP7_75t_L g4491 ( 
.A(n_4226),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_3981),
.B(n_2202),
.Y(n_4492)
);

NOR2xp33_ASAP7_75t_R g4493 ( 
.A(n_3964),
.B(n_2852),
.Y(n_4493)
);

INVx6_ASAP7_75t_L g4494 ( 
.A(n_3948),
.Y(n_4494)
);

BUFx2_ASAP7_75t_L g4495 ( 
.A(n_4111),
.Y(n_4495)
);

NAND2xp5_ASAP7_75t_L g4496 ( 
.A(n_3983),
.B(n_2212),
.Y(n_4496)
);

BUFx2_ASAP7_75t_L g4497 ( 
.A(n_4111),
.Y(n_4497)
);

INVx2_ASAP7_75t_L g4498 ( 
.A(n_4156),
.Y(n_4498)
);

NAND2xp5_ASAP7_75t_L g4499 ( 
.A(n_3983),
.B(n_3999),
.Y(n_4499)
);

NAND2xp5_ASAP7_75t_L g4500 ( 
.A(n_3999),
.B(n_2212),
.Y(n_4500)
);

BUFx12f_ASAP7_75t_L g4501 ( 
.A(n_4170),
.Y(n_4501)
);

INVx5_ASAP7_75t_L g4502 ( 
.A(n_3988),
.Y(n_4502)
);

INVx2_ASAP7_75t_SL g4503 ( 
.A(n_4214),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_4117),
.B(n_2215),
.Y(n_4504)
);

INVx2_ASAP7_75t_L g4505 ( 
.A(n_4181),
.Y(n_4505)
);

CKINVDCx16_ASAP7_75t_R g4506 ( 
.A(n_4039),
.Y(n_4506)
);

NAND2xp5_ASAP7_75t_L g4507 ( 
.A(n_4117),
.B(n_2215),
.Y(n_4507)
);

AOI22xp5_ASAP7_75t_L g4508 ( 
.A1(n_4113),
.A2(n_2244),
.B1(n_894),
.B2(n_949),
.Y(n_4508)
);

NOR2xp33_ASAP7_75t_R g4509 ( 
.A(n_3964),
.B(n_4175),
.Y(n_4509)
);

AND2x2_ASAP7_75t_L g4510 ( 
.A(n_4014),
.B(n_847),
.Y(n_4510)
);

INVx2_ASAP7_75t_L g4511 ( 
.A(n_4033),
.Y(n_4511)
);

BUFx2_ASAP7_75t_L g4512 ( 
.A(n_4247),
.Y(n_4512)
);

HB1xp67_ASAP7_75t_L g4513 ( 
.A(n_4239),
.Y(n_4513)
);

INVxp67_ASAP7_75t_L g4514 ( 
.A(n_4215),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_4148),
.B(n_3185),
.Y(n_4515)
);

INVx2_ASAP7_75t_SL g4516 ( 
.A(n_4058),
.Y(n_4516)
);

BUFx6f_ASAP7_75t_L g4517 ( 
.A(n_4091),
.Y(n_4517)
);

CKINVDCx5p33_ASAP7_75t_R g4518 ( 
.A(n_3936),
.Y(n_4518)
);

INVx1_ASAP7_75t_L g4519 ( 
.A(n_4037),
.Y(n_4519)
);

INVx2_ASAP7_75t_L g4520 ( 
.A(n_4041),
.Y(n_4520)
);

INVx4_ASAP7_75t_L g4521 ( 
.A(n_3964),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_4148),
.B(n_3187),
.Y(n_4522)
);

AOI22xp33_ASAP7_75t_L g4523 ( 
.A1(n_4093),
.A2(n_2120),
.B1(n_2128),
.B2(n_2108),
.Y(n_4523)
);

AND2x4_ASAP7_75t_L g4524 ( 
.A(n_4085),
.B(n_2933),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_L g4525 ( 
.A(n_4152),
.B(n_4015),
.Y(n_4525)
);

INVx1_ASAP7_75t_L g4526 ( 
.A(n_4041),
.Y(n_4526)
);

NAND2xp5_ASAP7_75t_L g4527 ( 
.A(n_4152),
.B(n_3191),
.Y(n_4527)
);

AO21x2_ASAP7_75t_L g4528 ( 
.A1(n_4251),
.A2(n_3005),
.B(n_3003),
.Y(n_4528)
);

OAI22xp5_ASAP7_75t_L g4529 ( 
.A1(n_4204),
.A2(n_852),
.B1(n_855),
.B2(n_849),
.Y(n_4529)
);

BUFx2_ASAP7_75t_L g4530 ( 
.A(n_4226),
.Y(n_4530)
);

INVx2_ASAP7_75t_L g4531 ( 
.A(n_4056),
.Y(n_4531)
);

INVx1_ASAP7_75t_SL g4532 ( 
.A(n_4129),
.Y(n_4532)
);

INVx3_ASAP7_75t_L g4533 ( 
.A(n_4226),
.Y(n_4533)
);

AND2x4_ASAP7_75t_L g4534 ( 
.A(n_4035),
.B(n_2933),
.Y(n_4534)
);

AND2x4_ASAP7_75t_L g4535 ( 
.A(n_4035),
.B(n_2949),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_L g4536 ( 
.A(n_4168),
.B(n_3191),
.Y(n_4536)
);

BUFx10_ASAP7_75t_L g4537 ( 
.A(n_4227),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_4056),
.Y(n_4538)
);

AND2x4_ASAP7_75t_L g4539 ( 
.A(n_4092),
.B(n_4187),
.Y(n_4539)
);

NAND2xp5_ASAP7_75t_L g4540 ( 
.A(n_4173),
.B(n_3192),
.Y(n_4540)
);

NAND2xp5_ASAP7_75t_SL g4541 ( 
.A(n_4060),
.B(n_3144),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_4067),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_SL g4543 ( 
.A(n_3920),
.B(n_3162),
.Y(n_4543)
);

NOR2xp33_ASAP7_75t_R g4544 ( 
.A(n_3949),
.B(n_2852),
.Y(n_4544)
);

BUFx3_ASAP7_75t_L g4545 ( 
.A(n_4075),
.Y(n_4545)
);

BUFx6f_ASAP7_75t_L g4546 ( 
.A(n_3993),
.Y(n_4546)
);

INVx3_ASAP7_75t_L g4547 ( 
.A(n_4092),
.Y(n_4547)
);

INVx3_ASAP7_75t_L g4548 ( 
.A(n_4022),
.Y(n_4548)
);

NAND2xp5_ASAP7_75t_SL g4549 ( 
.A(n_3920),
.B(n_3162),
.Y(n_4549)
);

AOI22xp33_ASAP7_75t_L g4550 ( 
.A1(n_3951),
.A2(n_2131),
.B1(n_2149),
.B2(n_2145),
.Y(n_4550)
);

INVx1_ASAP7_75t_L g4551 ( 
.A(n_4070),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_L g4552 ( 
.A(n_4179),
.B(n_3192),
.Y(n_4552)
);

AND2x4_ASAP7_75t_L g4553 ( 
.A(n_4145),
.B(n_2949),
.Y(n_4553)
);

INVx1_ASAP7_75t_L g4554 ( 
.A(n_4070),
.Y(n_4554)
);

NAND2xp5_ASAP7_75t_L g4555 ( 
.A(n_3971),
.B(n_3194),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_4084),
.Y(n_4556)
);

INVx1_ASAP7_75t_L g4557 ( 
.A(n_4084),
.Y(n_4557)
);

NOR2xp33_ASAP7_75t_L g4558 ( 
.A(n_3944),
.B(n_914),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4100),
.Y(n_4559)
);

OR2x2_ASAP7_75t_L g4560 ( 
.A(n_4024),
.B(n_4032),
.Y(n_4560)
);

NAND2xp5_ASAP7_75t_L g4561 ( 
.A(n_4167),
.B(n_3194),
.Y(n_4561)
);

HB1xp67_ASAP7_75t_L g4562 ( 
.A(n_4177),
.Y(n_4562)
);

NAND2xp5_ASAP7_75t_L g4563 ( 
.A(n_4167),
.B(n_3195),
.Y(n_4563)
);

BUFx2_ASAP7_75t_L g4564 ( 
.A(n_4022),
.Y(n_4564)
);

INVx4_ASAP7_75t_L g4565 ( 
.A(n_3922),
.Y(n_4565)
);

INVx4_ASAP7_75t_L g4566 ( 
.A(n_3922),
.Y(n_4566)
);

AND2x4_ASAP7_75t_L g4567 ( 
.A(n_4145),
.B(n_2949),
.Y(n_4567)
);

NAND2xp5_ASAP7_75t_L g4568 ( 
.A(n_4177),
.B(n_3951),
.Y(n_4568)
);

AND2x4_ASAP7_75t_L g4569 ( 
.A(n_4145),
.B(n_3058),
.Y(n_4569)
);

BUFx2_ASAP7_75t_L g4570 ( 
.A(n_4121),
.Y(n_4570)
);

NAND2xp5_ASAP7_75t_L g4571 ( 
.A(n_3951),
.B(n_3195),
.Y(n_4571)
);

HB1xp67_ASAP7_75t_L g4572 ( 
.A(n_4100),
.Y(n_4572)
);

INVx1_ASAP7_75t_L g4573 ( 
.A(n_4215),
.Y(n_4573)
);

INVx3_ASAP7_75t_L g4574 ( 
.A(n_4121),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_3951),
.B(n_3197),
.Y(n_4575)
);

NAND2xp5_ASAP7_75t_L g4576 ( 
.A(n_3973),
.B(n_3197),
.Y(n_4576)
);

AND2x4_ASAP7_75t_L g4577 ( 
.A(n_4145),
.B(n_3058),
.Y(n_4577)
);

INVxp67_ASAP7_75t_SL g4578 ( 
.A(n_4201),
.Y(n_4578)
);

BUFx6f_ASAP7_75t_L g4579 ( 
.A(n_4116),
.Y(n_4579)
);

NOR2xp33_ASAP7_75t_R g4580 ( 
.A(n_3970),
.B(n_3214),
.Y(n_4580)
);

NAND2xp5_ASAP7_75t_L g4581 ( 
.A(n_4164),
.B(n_3200),
.Y(n_4581)
);

NAND3xp33_ASAP7_75t_L g4582 ( 
.A(n_3972),
.B(n_4178),
.C(n_3938),
.Y(n_4582)
);

AOI21xp5_ASAP7_75t_L g4583 ( 
.A1(n_4036),
.A2(n_3167),
.B(n_3162),
.Y(n_4583)
);

NOR2xp33_ASAP7_75t_L g4584 ( 
.A(n_3975),
.B(n_916),
.Y(n_4584)
);

NAND2xp5_ASAP7_75t_L g4585 ( 
.A(n_4171),
.B(n_3200),
.Y(n_4585)
);

AOI22xp5_ASAP7_75t_L g4586 ( 
.A1(n_4112),
.A2(n_903),
.B1(n_957),
.B2(n_871),
.Y(n_4586)
);

BUFx5_ASAP7_75t_L g4587 ( 
.A(n_4112),
.Y(n_4587)
);

INVx1_ASAP7_75t_L g4588 ( 
.A(n_4224),
.Y(n_4588)
);

AND2x4_ASAP7_75t_L g4589 ( 
.A(n_4116),
.B(n_3058),
.Y(n_4589)
);

HB1xp67_ASAP7_75t_L g4590 ( 
.A(n_4235),
.Y(n_4590)
);

INVx3_ASAP7_75t_L g4591 ( 
.A(n_4217),
.Y(n_4591)
);

BUFx6f_ASAP7_75t_L g4592 ( 
.A(n_4116),
.Y(n_4592)
);

INVx1_ASAP7_75t_L g4593 ( 
.A(n_4224),
.Y(n_4593)
);

NAND2xp5_ASAP7_75t_L g4594 ( 
.A(n_4153),
.B(n_4158),
.Y(n_4594)
);

NAND2xp5_ASAP7_75t_L g4595 ( 
.A(n_4153),
.B(n_3208),
.Y(n_4595)
);

INVx2_ASAP7_75t_SL g4596 ( 
.A(n_4090),
.Y(n_4596)
);

AND2x4_ASAP7_75t_L g4597 ( 
.A(n_4138),
.B(n_3091),
.Y(n_4597)
);

INVx1_ASAP7_75t_L g4598 ( 
.A(n_4197),
.Y(n_4598)
);

NAND3xp33_ASAP7_75t_SL g4599 ( 
.A(n_4044),
.B(n_852),
.C(n_849),
.Y(n_4599)
);

INVx2_ASAP7_75t_SL g4600 ( 
.A(n_4125),
.Y(n_4600)
);

NAND2xp33_ASAP7_75t_L g4601 ( 
.A(n_3979),
.B(n_3162),
.Y(n_4601)
);

NOR2xp33_ASAP7_75t_L g4602 ( 
.A(n_4186),
.B(n_920),
.Y(n_4602)
);

INVx1_ASAP7_75t_L g4603 ( 
.A(n_4197),
.Y(n_4603)
);

NAND2xp5_ASAP7_75t_L g4604 ( 
.A(n_4158),
.B(n_3208),
.Y(n_4604)
);

INVx5_ASAP7_75t_L g4605 ( 
.A(n_4271),
.Y(n_4605)
);

OAI22xp5_ASAP7_75t_L g4606 ( 
.A1(n_4582),
.A2(n_3947),
.B1(n_4082),
.B2(n_4232),
.Y(n_4606)
);

A2O1A1Ixp33_ASAP7_75t_L g4607 ( 
.A1(n_4411),
.A2(n_4162),
.B(n_4246),
.C(n_4038),
.Y(n_4607)
);

OR2x6_ASAP7_75t_L g4608 ( 
.A(n_4435),
.B(n_3917),
.Y(n_4608)
);

AND2x2_ASAP7_75t_L g4609 ( 
.A(n_4297),
.B(n_4062),
.Y(n_4609)
);

A2O1A1Ixp33_ASAP7_75t_SL g4610 ( 
.A1(n_4309),
.A2(n_4136),
.B(n_857),
.C(n_863),
.Y(n_4610)
);

NAND2xp5_ASAP7_75t_L g4611 ( 
.A(n_4393),
.B(n_4207),
.Y(n_4611)
);

A2O1A1Ixp33_ASAP7_75t_L g4612 ( 
.A1(n_4411),
.A2(n_4124),
.B(n_4130),
.C(n_4122),
.Y(n_4612)
);

BUFx6f_ASAP7_75t_L g4613 ( 
.A(n_4446),
.Y(n_4613)
);

NOR2xp33_ASAP7_75t_SL g4614 ( 
.A(n_4271),
.B(n_3948),
.Y(n_4614)
);

INVx1_ASAP7_75t_SL g4615 ( 
.A(n_4259),
.Y(n_4615)
);

O2A1O1Ixp33_ASAP7_75t_L g4616 ( 
.A1(n_4558),
.A2(n_4236),
.B(n_857),
.C(n_863),
.Y(n_4616)
);

NOR2xp33_ASAP7_75t_L g4617 ( 
.A(n_4289),
.B(n_4079),
.Y(n_4617)
);

AND2x4_ASAP7_75t_L g4618 ( 
.A(n_4271),
.B(n_4008),
.Y(n_4618)
);

NOR2xp33_ASAP7_75t_L g4619 ( 
.A(n_4335),
.B(n_36),
.Y(n_4619)
);

CKINVDCx5p33_ASAP7_75t_R g4620 ( 
.A(n_4324),
.Y(n_4620)
);

OAI21xp33_ASAP7_75t_SL g4621 ( 
.A1(n_4259),
.A2(n_3940),
.B(n_4106),
.Y(n_4621)
);

AOI22xp5_ASAP7_75t_L g4622 ( 
.A1(n_4292),
.A2(n_4112),
.B1(n_4068),
.B2(n_3994),
.Y(n_4622)
);

AOI21xp5_ASAP7_75t_L g4623 ( 
.A1(n_4601),
.A2(n_4045),
.B(n_3924),
.Y(n_4623)
);

BUFx3_ASAP7_75t_L g4624 ( 
.A(n_4391),
.Y(n_4624)
);

AOI21xp5_ASAP7_75t_L g4625 ( 
.A1(n_4341),
.A2(n_4042),
.B(n_4026),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4433),
.B(n_4213),
.Y(n_4626)
);

OAI22xp5_ASAP7_75t_L g4627 ( 
.A1(n_4281),
.A2(n_4114),
.B1(n_4118),
.B2(n_4081),
.Y(n_4627)
);

INVx2_ASAP7_75t_SL g4628 ( 
.A(n_4545),
.Y(n_4628)
);

AND2x2_ASAP7_75t_L g4629 ( 
.A(n_4384),
.B(n_4189),
.Y(n_4629)
);

OAI22xp5_ASAP7_75t_L g4630 ( 
.A1(n_4281),
.A2(n_4019),
.B1(n_4076),
.B2(n_3925),
.Y(n_4630)
);

A2O1A1Ixp33_ASAP7_75t_L g4631 ( 
.A1(n_4586),
.A2(n_3965),
.B(n_3960),
.C(n_4163),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4453),
.B(n_4194),
.Y(n_4632)
);

NOR2xp67_ASAP7_75t_L g4633 ( 
.A(n_4334),
.B(n_3948),
.Y(n_4633)
);

O2A1O1Ixp33_ASAP7_75t_L g4634 ( 
.A1(n_4366),
.A2(n_872),
.B(n_874),
.C(n_856),
.Y(n_4634)
);

A2O1A1Ixp33_ASAP7_75t_L g4635 ( 
.A1(n_4408),
.A2(n_3965),
.B(n_3960),
.C(n_4163),
.Y(n_4635)
);

INVx3_ASAP7_75t_L g4636 ( 
.A(n_4271),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4457),
.B(n_4218),
.Y(n_4637)
);

INVx3_ASAP7_75t_L g4638 ( 
.A(n_4282),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4562),
.B(n_4231),
.Y(n_4639)
);

INVx4_ASAP7_75t_L g4640 ( 
.A(n_4565),
.Y(n_4640)
);

A2O1A1Ixp33_ASAP7_75t_L g4641 ( 
.A1(n_4451),
.A2(n_4199),
.B(n_4192),
.C(n_4188),
.Y(n_4641)
);

OAI22xp5_ASAP7_75t_L g4642 ( 
.A1(n_4329),
.A2(n_3962),
.B1(n_4147),
.B2(n_4144),
.Y(n_4642)
);

NOR2xp33_ASAP7_75t_L g4643 ( 
.A(n_4415),
.B(n_38),
.Y(n_4643)
);

NOR2xp33_ASAP7_75t_L g4644 ( 
.A(n_4311),
.B(n_42),
.Y(n_4644)
);

NOR2xp33_ASAP7_75t_L g4645 ( 
.A(n_4385),
.B(n_42),
.Y(n_4645)
);

NAND2x1p5_ASAP7_75t_L g4646 ( 
.A(n_4282),
.B(n_3998),
.Y(n_4646)
);

AOI21xp5_ASAP7_75t_L g4647 ( 
.A1(n_4341),
.A2(n_4253),
.B(n_4205),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4578),
.A2(n_4253),
.B(n_4205),
.Y(n_4648)
);

BUFx2_ASAP7_75t_L g4649 ( 
.A(n_4270),
.Y(n_4649)
);

OAI21xp5_ASAP7_75t_L g4650 ( 
.A1(n_4328),
.A2(n_4063),
.B(n_3934),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4499),
.B(n_4237),
.Y(n_4651)
);

AOI21xp5_ASAP7_75t_L g4652 ( 
.A1(n_4380),
.A2(n_4206),
.B(n_4201),
.Y(n_4652)
);

AND2x2_ASAP7_75t_L g4653 ( 
.A(n_4256),
.B(n_4296),
.Y(n_4653)
);

AOI22xp33_ASAP7_75t_L g4654 ( 
.A1(n_4292),
.A2(n_4436),
.B1(n_4501),
.B2(n_4599),
.Y(n_4654)
);

O2A1O1Ixp5_ASAP7_75t_L g4655 ( 
.A1(n_4302),
.A2(n_4107),
.B(n_4220),
.C(n_4183),
.Y(n_4655)
);

AND2x2_ASAP7_75t_L g4656 ( 
.A(n_4293),
.B(n_4185),
.Y(n_4656)
);

A2O1A1Ixp33_ASAP7_75t_SL g4657 ( 
.A1(n_4584),
.A2(n_872),
.B(n_877),
.C(n_856),
.Y(n_4657)
);

OAI22xp5_ASAP7_75t_L g4658 ( 
.A1(n_4261),
.A2(n_4169),
.B1(n_4185),
.B2(n_4097),
.Y(n_4658)
);

BUFx6f_ASAP7_75t_L g4659 ( 
.A(n_4446),
.Y(n_4659)
);

INVx4_ASAP7_75t_L g4660 ( 
.A(n_4565),
.Y(n_4660)
);

O2A1O1Ixp33_ASAP7_75t_L g4661 ( 
.A1(n_4429),
.A2(n_878),
.B(n_881),
.C(n_877),
.Y(n_4661)
);

NOR2xp33_ASAP7_75t_SL g4662 ( 
.A(n_4282),
.B(n_3998),
.Y(n_4662)
);

INVx1_ASAP7_75t_L g4663 ( 
.A(n_4572),
.Y(n_4663)
);

NAND2xp5_ASAP7_75t_SL g4664 ( 
.A(n_4390),
.B(n_4028),
.Y(n_4664)
);

BUFx8_ASAP7_75t_SL g4665 ( 
.A(n_4272),
.Y(n_4665)
);

NAND2x1p5_ASAP7_75t_L g4666 ( 
.A(n_4282),
.B(n_3998),
.Y(n_4666)
);

CKINVDCx6p67_ASAP7_75t_R g4667 ( 
.A(n_4262),
.Y(n_4667)
);

AND2x2_ASAP7_75t_L g4668 ( 
.A(n_4274),
.B(n_4185),
.Y(n_4668)
);

INVx2_ASAP7_75t_L g4669 ( 
.A(n_4418),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_SL g4670 ( 
.A(n_4347),
.B(n_4072),
.Y(n_4670)
);

NOR2xp33_ASAP7_75t_L g4671 ( 
.A(n_4331),
.B(n_43),
.Y(n_4671)
);

NOR2xp33_ASAP7_75t_L g4672 ( 
.A(n_4397),
.B(n_44),
.Y(n_4672)
);

AOI21xp5_ASAP7_75t_L g4673 ( 
.A1(n_4260),
.A2(n_4211),
.B(n_4119),
.Y(n_4673)
);

AOI21xp5_ASAP7_75t_L g4674 ( 
.A1(n_4583),
.A2(n_4212),
.B(n_3950),
.Y(n_4674)
);

A2O1A1Ixp33_ASAP7_75t_L g4675 ( 
.A1(n_4470),
.A2(n_878),
.B(n_883),
.C(n_881),
.Y(n_4675)
);

OAI22xp5_ASAP7_75t_L g4676 ( 
.A1(n_4350),
.A2(n_4094),
.B1(n_4180),
.B2(n_4097),
.Y(n_4676)
);

CKINVDCx20_ASAP7_75t_R g4677 ( 
.A(n_4417),
.Y(n_4677)
);

NAND2xp5_ASAP7_75t_SL g4678 ( 
.A(n_4347),
.B(n_4072),
.Y(n_4678)
);

OAI22xp5_ASAP7_75t_L g4679 ( 
.A1(n_4357),
.A2(n_4094),
.B1(n_4208),
.B2(n_4180),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4431),
.Y(n_4680)
);

AOI21xp5_ASAP7_75t_L g4681 ( 
.A1(n_4599),
.A2(n_3950),
.B(n_4208),
.Y(n_4681)
);

NAND2xp5_ASAP7_75t_SL g4682 ( 
.A(n_4347),
.B(n_4217),
.Y(n_4682)
);

AO21x1_ASAP7_75t_L g4683 ( 
.A1(n_4269),
.A2(n_895),
.B(n_883),
.Y(n_4683)
);

INVx3_ASAP7_75t_L g4684 ( 
.A(n_4347),
.Y(n_4684)
);

AO22x1_ASAP7_75t_L g4685 ( 
.A1(n_4360),
.A2(n_4103),
.B1(n_4105),
.B2(n_4095),
.Y(n_4685)
);

OAI22xp5_ASAP7_75t_L g4686 ( 
.A1(n_4356),
.A2(n_4529),
.B1(n_4439),
.B2(n_4550),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4525),
.B(n_4138),
.Y(n_4687)
);

AOI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_4490),
.A2(n_3056),
.B(n_3054),
.Y(n_4688)
);

A2O1A1Ixp33_ASAP7_75t_L g4689 ( 
.A1(n_4473),
.A2(n_895),
.B(n_911),
.C(n_901),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4525),
.B(n_4151),
.Y(n_4690)
);

O2A1O1Ixp33_ASAP7_75t_L g4691 ( 
.A1(n_4478),
.A2(n_4529),
.B(n_4334),
.C(n_4439),
.Y(n_4691)
);

NOR2xp33_ASAP7_75t_L g4692 ( 
.A(n_4475),
.B(n_44),
.Y(n_4692)
);

INVx1_ASAP7_75t_L g4693 ( 
.A(n_4469),
.Y(n_4693)
);

O2A1O1Ixp33_ASAP7_75t_L g4694 ( 
.A1(n_4472),
.A2(n_911),
.B(n_918),
.C(n_901),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_SL g4695 ( 
.A(n_4360),
.B(n_4151),
.Y(n_4695)
);

OAI21xp5_ASAP7_75t_L g4696 ( 
.A1(n_4382),
.A2(n_921),
.B(n_918),
.Y(n_4696)
);

OAI22xp5_ASAP7_75t_L g4697 ( 
.A1(n_4508),
.A2(n_4518),
.B1(n_4506),
.B2(n_4294),
.Y(n_4697)
);

OR2x6_ASAP7_75t_L g4698 ( 
.A(n_4435),
.B(n_4095),
.Y(n_4698)
);

NOR2xp33_ASAP7_75t_L g4699 ( 
.A(n_4488),
.B(n_46),
.Y(n_4699)
);

BUFx6f_ASAP7_75t_L g4700 ( 
.A(n_4446),
.Y(n_4700)
);

OAI21xp33_ASAP7_75t_L g4701 ( 
.A1(n_4267),
.A2(n_925),
.B(n_923),
.Y(n_4701)
);

OAI22xp5_ASAP7_75t_L g4702 ( 
.A1(n_4370),
.A2(n_925),
.B1(n_926),
.B2(n_923),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_SL g4703 ( 
.A(n_4360),
.B(n_4151),
.Y(n_4703)
);

NAND2xp5_ASAP7_75t_L g4704 ( 
.A(n_4560),
.B(n_4161),
.Y(n_4704)
);

O2A1O1Ixp33_ASAP7_75t_L g4705 ( 
.A1(n_4472),
.A2(n_926),
.B(n_930),
.C(n_928),
.Y(n_4705)
);

NAND2xp5_ASAP7_75t_L g4706 ( 
.A(n_4361),
.B(n_4161),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_SL g4707 ( 
.A(n_4360),
.B(n_4161),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_L g4708 ( 
.A(n_4361),
.B(n_928),
.Y(n_4708)
);

HB1xp67_ASAP7_75t_L g4709 ( 
.A(n_4268),
.Y(n_4709)
);

NOR2xp33_ASAP7_75t_L g4710 ( 
.A(n_4484),
.B(n_47),
.Y(n_4710)
);

AOI21xp5_ASAP7_75t_L g4711 ( 
.A1(n_4267),
.A2(n_3216),
.B(n_3215),
.Y(n_4711)
);

AOI21xp5_ASAP7_75t_L g4712 ( 
.A1(n_4489),
.A2(n_3216),
.B(n_3215),
.Y(n_4712)
);

INVx8_ASAP7_75t_L g4713 ( 
.A(n_4546),
.Y(n_4713)
);

BUFx6f_ASAP7_75t_L g4714 ( 
.A(n_4517),
.Y(n_4714)
);

AND2x2_ASAP7_75t_SL g4715 ( 
.A(n_4495),
.B(n_4095),
.Y(n_4715)
);

INVx2_ASAP7_75t_L g4716 ( 
.A(n_4442),
.Y(n_4716)
);

INVx2_ASAP7_75t_L g4717 ( 
.A(n_4445),
.Y(n_4717)
);

O2A1O1Ixp33_ASAP7_75t_L g4718 ( 
.A1(n_4482),
.A2(n_930),
.B(n_936),
.C(n_932),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4367),
.B(n_932),
.Y(n_4719)
);

AOI21xp5_ASAP7_75t_L g4720 ( 
.A1(n_4265),
.A2(n_3224),
.B(n_3217),
.Y(n_4720)
);

NAND2xp5_ASAP7_75t_SL g4721 ( 
.A(n_4509),
.B(n_4103),
.Y(n_4721)
);

NAND2xp33_ASAP7_75t_L g4722 ( 
.A(n_4287),
.B(n_859),
.Y(n_4722)
);

NAND2xp5_ASAP7_75t_L g4723 ( 
.A(n_4376),
.B(n_936),
.Y(n_4723)
);

AOI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_4354),
.A2(n_3240),
.B(n_3236),
.Y(n_4724)
);

INVx4_ASAP7_75t_L g4725 ( 
.A(n_4566),
.Y(n_4725)
);

INVx2_ASAP7_75t_L g4726 ( 
.A(n_4455),
.Y(n_4726)
);

CKINVDCx5p33_ASAP7_75t_R g4727 ( 
.A(n_4300),
.Y(n_4727)
);

INVx1_ASAP7_75t_L g4728 ( 
.A(n_4286),
.Y(n_4728)
);

AOI21xp5_ASAP7_75t_L g4729 ( 
.A1(n_4369),
.A2(n_4375),
.B(n_4419),
.Y(n_4729)
);

INVxp67_ASAP7_75t_SL g4730 ( 
.A(n_4568),
.Y(n_4730)
);

NAND2xp5_ASAP7_75t_L g4731 ( 
.A(n_4377),
.B(n_946),
.Y(n_4731)
);

A2O1A1Ixp33_ASAP7_75t_L g4732 ( 
.A1(n_4405),
.A2(n_950),
.B(n_952),
.C(n_948),
.Y(n_4732)
);

INVx2_ASAP7_75t_L g4733 ( 
.A(n_4468),
.Y(n_4733)
);

NAND2xp5_ASAP7_75t_SL g4734 ( 
.A(n_4404),
.B(n_4568),
.Y(n_4734)
);

OAI21xp33_ASAP7_75t_L g4735 ( 
.A1(n_4269),
.A2(n_950),
.B(n_948),
.Y(n_4735)
);

HB1xp67_ASAP7_75t_L g4736 ( 
.A(n_4479),
.Y(n_4736)
);

NOR2xp33_ASAP7_75t_L g4737 ( 
.A(n_4537),
.B(n_47),
.Y(n_4737)
);

OR2x2_ASAP7_75t_L g4738 ( 
.A(n_4532),
.B(n_4103),
.Y(n_4738)
);

AND2x4_ASAP7_75t_L g4739 ( 
.A(n_4278),
.B(n_4105),
.Y(n_4739)
);

O2A1O1Ixp33_ASAP7_75t_L g4740 ( 
.A1(n_4482),
.A2(n_953),
.B(n_956),
.C(n_952),
.Y(n_4740)
);

NAND2xp5_ASAP7_75t_L g4741 ( 
.A(n_4266),
.B(n_953),
.Y(n_4741)
);

OAI22xp5_ASAP7_75t_SL g4742 ( 
.A1(n_4312),
.A2(n_962),
.B1(n_963),
.B2(n_958),
.Y(n_4742)
);

OAI22xp5_ASAP7_75t_L g4743 ( 
.A1(n_4474),
.A2(n_962),
.B1(n_968),
.B2(n_963),
.Y(n_4743)
);

O2A1O1Ixp33_ASAP7_75t_L g4744 ( 
.A1(n_4464),
.A2(n_968),
.B(n_969),
.C(n_958),
.Y(n_4744)
);

BUFx6f_ASAP7_75t_L g4745 ( 
.A(n_4517),
.Y(n_4745)
);

NAND2xp5_ASAP7_75t_L g4746 ( 
.A(n_4532),
.B(n_4480),
.Y(n_4746)
);

NAND3xp33_ASAP7_75t_SL g4747 ( 
.A(n_4409),
.B(n_970),
.C(n_969),
.Y(n_4747)
);

INVxp67_ASAP7_75t_SL g4748 ( 
.A(n_4476),
.Y(n_4748)
);

HB1xp67_ASAP7_75t_L g4749 ( 
.A(n_4512),
.Y(n_4749)
);

CKINVDCx5p33_ASAP7_75t_R g4750 ( 
.A(n_4322),
.Y(n_4750)
);

O2A1O1Ixp33_ASAP7_75t_L g4751 ( 
.A1(n_4464),
.A2(n_971),
.B(n_972),
.C(n_970),
.Y(n_4751)
);

INVx1_ASAP7_75t_L g4752 ( 
.A(n_4295),
.Y(n_4752)
);

NAND2x1p5_ASAP7_75t_L g4753 ( 
.A(n_4485),
.B(n_3162),
.Y(n_4753)
);

AOI21xp5_ASAP7_75t_L g4754 ( 
.A1(n_4375),
.A2(n_4383),
.B(n_4416),
.Y(n_4754)
);

NOR2xp67_ASAP7_75t_SL g4755 ( 
.A(n_4546),
.B(n_3167),
.Y(n_4755)
);

INVx4_ASAP7_75t_SL g4756 ( 
.A(n_4494),
.Y(n_4756)
);

NAND2xp5_ASAP7_75t_L g4757 ( 
.A(n_4519),
.B(n_972),
.Y(n_4757)
);

NAND2xp5_ASAP7_75t_SL g4758 ( 
.A(n_4587),
.B(n_4228),
.Y(n_4758)
);

AOI22xp5_ASAP7_75t_L g4759 ( 
.A1(n_4312),
.A2(n_990),
.B1(n_991),
.B2(n_980),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_SL g4760 ( 
.A(n_4587),
.B(n_4228),
.Y(n_4760)
);

NAND2xp5_ASAP7_75t_L g4761 ( 
.A(n_4526),
.B(n_980),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4298),
.Y(n_4762)
);

AOI22xp5_ASAP7_75t_L g4763 ( 
.A1(n_4386),
.A2(n_991),
.B1(n_994),
.B2(n_990),
.Y(n_4763)
);

NAND2xp5_ASAP7_75t_SL g4764 ( 
.A(n_4587),
.B(n_3167),
.Y(n_4764)
);

BUFx6f_ASAP7_75t_L g4765 ( 
.A(n_4517),
.Y(n_4765)
);

NAND2xp5_ASAP7_75t_SL g4766 ( 
.A(n_4587),
.B(n_3167),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_SL g4767 ( 
.A(n_4587),
.B(n_3167),
.Y(n_4767)
);

INVx1_ASAP7_75t_SL g4768 ( 
.A(n_4392),
.Y(n_4768)
);

HB1xp67_ASAP7_75t_L g4769 ( 
.A(n_4465),
.Y(n_4769)
);

AND2x4_ASAP7_75t_L g4770 ( 
.A(n_4278),
.B(n_1418),
.Y(n_4770)
);

AND2x2_ASAP7_75t_L g4771 ( 
.A(n_4539),
.B(n_994),
.Y(n_4771)
);

AOI21x1_ASAP7_75t_L g4772 ( 
.A1(n_4454),
.A2(n_1424),
.B(n_1423),
.Y(n_4772)
);

AND2x4_ASAP7_75t_L g4773 ( 
.A(n_4291),
.B(n_4307),
.Y(n_4773)
);

NOR2xp33_ASAP7_75t_L g4774 ( 
.A(n_4516),
.B(n_49),
.Y(n_4774)
);

AOI22xp5_ASAP7_75t_L g4775 ( 
.A1(n_4389),
.A2(n_996),
.B1(n_1000),
.B2(n_995),
.Y(n_4775)
);

INVx3_ASAP7_75t_L g4776 ( 
.A(n_4291),
.Y(n_4776)
);

BUFx2_ASAP7_75t_L g4777 ( 
.A(n_4342),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4538),
.B(n_995),
.Y(n_4778)
);

AOI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4383),
.A2(n_3256),
.B(n_3242),
.Y(n_4779)
);

OAI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_4389),
.A2(n_1023),
.B(n_1011),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_SL g4781 ( 
.A(n_4263),
.B(n_3176),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_SL g4782 ( 
.A(n_4263),
.B(n_3176),
.Y(n_4782)
);

NOR2xp33_ASAP7_75t_L g4783 ( 
.A(n_4596),
.B(n_49),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_SL g4784 ( 
.A(n_4544),
.B(n_3176),
.Y(n_4784)
);

CKINVDCx20_ASAP7_75t_R g4785 ( 
.A(n_4447),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4542),
.B(n_1023),
.Y(n_4786)
);

CKINVDCx5p33_ASAP7_75t_R g4787 ( 
.A(n_4310),
.Y(n_4787)
);

BUFx2_ASAP7_75t_L g4788 ( 
.A(n_4342),
.Y(n_4788)
);

HB1xp67_ASAP7_75t_L g4789 ( 
.A(n_4465),
.Y(n_4789)
);

A2O1A1Ixp33_ASAP7_75t_L g4790 ( 
.A1(n_4602),
.A2(n_1034),
.B(n_1038),
.C(n_1029),
.Y(n_4790)
);

NOR2xp33_ASAP7_75t_L g4791 ( 
.A(n_4600),
.B(n_50),
.Y(n_4791)
);

INVx2_ASAP7_75t_L g4792 ( 
.A(n_4477),
.Y(n_4792)
);

OAI22xp5_ASAP7_75t_L g4793 ( 
.A1(n_4427),
.A2(n_1040),
.B1(n_1043),
.B2(n_1038),
.Y(n_4793)
);

INVx1_ASAP7_75t_L g4794 ( 
.A(n_4315),
.Y(n_4794)
);

NAND2xp33_ASAP7_75t_SL g4795 ( 
.A(n_4493),
.B(n_1040),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4551),
.B(n_1043),
.Y(n_4796)
);

A2O1A1Ixp33_ASAP7_75t_L g4797 ( 
.A1(n_4422),
.A2(n_1056),
.B(n_1059),
.C(n_1046),
.Y(n_4797)
);

AND2x4_ASAP7_75t_L g4798 ( 
.A(n_4307),
.B(n_1426),
.Y(n_4798)
);

BUFx12f_ASAP7_75t_L g4799 ( 
.A(n_4450),
.Y(n_4799)
);

A2O1A1Ixp33_ASAP7_75t_L g4800 ( 
.A1(n_4594),
.A2(n_1056),
.B(n_1059),
.C(n_1046),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4554),
.B(n_1061),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4557),
.B(n_1061),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4588),
.B(n_1064),
.Y(n_4803)
);

INVx1_ASAP7_75t_L g4804 ( 
.A(n_4321),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4593),
.B(n_1064),
.Y(n_4805)
);

NOR2xp33_ASAP7_75t_SL g4806 ( 
.A(n_4430),
.B(n_3091),
.Y(n_4806)
);

AOI21xp5_ASAP7_75t_L g4807 ( 
.A1(n_4388),
.A2(n_3220),
.B(n_2463),
.Y(n_4807)
);

AOI21xp5_ASAP7_75t_L g4808 ( 
.A1(n_4323),
.A2(n_3220),
.B(n_2463),
.Y(n_4808)
);

AOI21xp5_ASAP7_75t_L g4809 ( 
.A1(n_4330),
.A2(n_3220),
.B(n_3110),
.Y(n_4809)
);

NOR2xp33_ASAP7_75t_L g4810 ( 
.A(n_4503),
.B(n_50),
.Y(n_4810)
);

INVxp67_ASAP7_75t_SL g4811 ( 
.A(n_4513),
.Y(n_4811)
);

BUFx6f_ASAP7_75t_L g4812 ( 
.A(n_4355),
.Y(n_4812)
);

INVx2_ASAP7_75t_L g4813 ( 
.A(n_4498),
.Y(n_4813)
);

AND2x2_ASAP7_75t_L g4814 ( 
.A(n_4317),
.B(n_1065),
.Y(n_4814)
);

INVx2_ASAP7_75t_SL g4815 ( 
.A(n_4456),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4511),
.B(n_1065),
.Y(n_4816)
);

OAI21xp33_ASAP7_75t_L g4817 ( 
.A1(n_4598),
.A2(n_1068),
.B(n_1066),
.Y(n_4817)
);

AOI21xp5_ASAP7_75t_L g4818 ( 
.A1(n_4571),
.A2(n_3110),
.B(n_3107),
.Y(n_4818)
);

BUFx3_ASAP7_75t_L g4819 ( 
.A(n_4351),
.Y(n_4819)
);

BUFx6f_ASAP7_75t_L g4820 ( 
.A(n_4355),
.Y(n_4820)
);

OAI22xp5_ASAP7_75t_L g4821 ( 
.A1(n_4467),
.A2(n_1068),
.B1(n_1072),
.B2(n_1066),
.Y(n_4821)
);

OAI22xp5_ASAP7_75t_SL g4822 ( 
.A1(n_4530),
.A2(n_4603),
.B1(n_4299),
.B2(n_4497),
.Y(n_4822)
);

AOI21xp5_ASAP7_75t_L g4823 ( 
.A1(n_4575),
.A2(n_3117),
.B(n_3107),
.Y(n_4823)
);

OR2x2_ASAP7_75t_L g4824 ( 
.A(n_4520),
.B(n_1427),
.Y(n_4824)
);

INVx2_ASAP7_75t_L g4825 ( 
.A(n_4276),
.Y(n_4825)
);

AOI22x1_ASAP7_75t_L g4826 ( 
.A1(n_4255),
.A2(n_1072),
.B1(n_1073),
.B2(n_1071),
.Y(n_4826)
);

BUFx6f_ASAP7_75t_L g4827 ( 
.A(n_4355),
.Y(n_4827)
);

OR2x6_ASAP7_75t_L g4828 ( 
.A(n_4435),
.B(n_3117),
.Y(n_4828)
);

BUFx3_ASAP7_75t_L g4829 ( 
.A(n_4351),
.Y(n_4829)
);

OAI22xp5_ASAP7_75t_L g4830 ( 
.A1(n_4467),
.A2(n_1073),
.B1(n_1075),
.B2(n_1071),
.Y(n_4830)
);

NAND2xp5_ASAP7_75t_L g4831 ( 
.A(n_4531),
.B(n_1075),
.Y(n_4831)
);

INVxp67_ASAP7_75t_L g4832 ( 
.A(n_4400),
.Y(n_4832)
);

NAND2xp5_ASAP7_75t_L g4833 ( 
.A(n_4556),
.B(n_1079),
.Y(n_4833)
);

NOR3xp33_ASAP7_75t_L g4834 ( 
.A(n_4437),
.B(n_1080),
.C(n_1079),
.Y(n_4834)
);

INVx2_ASAP7_75t_L g4835 ( 
.A(n_4277),
.Y(n_4835)
);

NOR2xp33_ASAP7_75t_L g4836 ( 
.A(n_4258),
.B(n_51),
.Y(n_4836)
);

NOR2xp33_ASAP7_75t_L g4837 ( 
.A(n_4258),
.B(n_52),
.Y(n_4837)
);

AND2x4_ASAP7_75t_L g4838 ( 
.A(n_4491),
.B(n_1428),
.Y(n_4838)
);

INVx2_ASAP7_75t_L g4839 ( 
.A(n_4304),
.Y(n_4839)
);

NOR3xp33_ASAP7_75t_L g4840 ( 
.A(n_4437),
.B(n_1083),
.C(n_1080),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_SL g4841 ( 
.A(n_4580),
.B(n_3117),
.Y(n_4841)
);

A2O1A1Ixp33_ASAP7_75t_L g4842 ( 
.A1(n_4326),
.A2(n_1087),
.B(n_1089),
.C(n_1083),
.Y(n_4842)
);

AOI21xp5_ASAP7_75t_L g4843 ( 
.A1(n_4575),
.A2(n_3126),
.B(n_2835),
.Y(n_4843)
);

NAND2xp5_ASAP7_75t_L g4844 ( 
.A(n_4559),
.B(n_1087),
.Y(n_4844)
);

INVx2_ASAP7_75t_L g4845 ( 
.A(n_4305),
.Y(n_4845)
);

BUFx12f_ASAP7_75t_L g4846 ( 
.A(n_4421),
.Y(n_4846)
);

INVx3_ASAP7_75t_L g4847 ( 
.A(n_4591),
.Y(n_4847)
);

INVx1_ASAP7_75t_L g4848 ( 
.A(n_4343),
.Y(n_4848)
);

NOR2xp33_ASAP7_75t_L g4849 ( 
.A(n_4441),
.B(n_54),
.Y(n_4849)
);

O2A1O1Ixp33_ASAP7_75t_L g4850 ( 
.A1(n_4487),
.A2(n_1094),
.B(n_1097),
.C(n_1089),
.Y(n_4850)
);

AOI21xp5_ASAP7_75t_L g4851 ( 
.A1(n_4402),
.A2(n_3126),
.B(n_2875),
.Y(n_4851)
);

INVx3_ASAP7_75t_L g4852 ( 
.A(n_4591),
.Y(n_4852)
);

AOI21xp5_ASAP7_75t_L g4853 ( 
.A1(n_4402),
.A2(n_2875),
.B(n_2856),
.Y(n_4853)
);

OAI22xp5_ASAP7_75t_L g4854 ( 
.A1(n_4500),
.A2(n_1097),
.B1(n_1099),
.B2(n_1094),
.Y(n_4854)
);

OAI21x1_ASAP7_75t_L g4855 ( 
.A1(n_4403),
.A2(n_2511),
.B(n_2592),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4514),
.B(n_1099),
.Y(n_4856)
);

INVx2_ASAP7_75t_L g4857 ( 
.A(n_4318),
.Y(n_4857)
);

NOR2xp33_ASAP7_75t_L g4858 ( 
.A(n_4510),
.B(n_4521),
.Y(n_4858)
);

O2A1O1Ixp33_ASAP7_75t_L g4859 ( 
.A1(n_4487),
.A2(n_1104),
.B(n_1106),
.C(n_1103),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4573),
.B(n_1104),
.Y(n_4860)
);

O2A1O1Ixp33_ASAP7_75t_L g4861 ( 
.A1(n_4492),
.A2(n_4496),
.B(n_4500),
.C(n_4449),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_4353),
.Y(n_4862)
);

INVx1_ASAP7_75t_L g4863 ( 
.A(n_4362),
.Y(n_4863)
);

OAI22xp5_ASAP7_75t_L g4864 ( 
.A1(n_4492),
.A2(n_1111),
.B1(n_1112),
.B2(n_1106),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4373),
.B(n_1111),
.Y(n_4865)
);

NOR2xp33_ASAP7_75t_L g4866 ( 
.A(n_4521),
.B(n_4340),
.Y(n_4866)
);

CKINVDCx5p33_ASAP7_75t_R g4867 ( 
.A(n_4421),
.Y(n_4867)
);

INVx1_ASAP7_75t_L g4868 ( 
.A(n_4379),
.Y(n_4868)
);

AOI21xp5_ASAP7_75t_L g4869 ( 
.A1(n_4358),
.A2(n_2875),
.B(n_2856),
.Y(n_4869)
);

INVx1_ASAP7_75t_L g4870 ( 
.A(n_4387),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4398),
.B(n_1113),
.Y(n_4871)
);

INVx4_ASAP7_75t_L g4872 ( 
.A(n_4566),
.Y(n_4872)
);

AOI22xp33_ASAP7_75t_L g4873 ( 
.A1(n_4505),
.A2(n_2913),
.B1(n_2917),
.B2(n_2916),
.Y(n_4873)
);

A2O1A1Ixp33_ASAP7_75t_L g4874 ( 
.A1(n_4326),
.A2(n_1116),
.B(n_1118),
.C(n_1115),
.Y(n_4874)
);

AND2x2_ASAP7_75t_L g4875 ( 
.A(n_4325),
.B(n_1115),
.Y(n_4875)
);

AOI21xp5_ASAP7_75t_L g4876 ( 
.A1(n_4358),
.A2(n_2877),
.B(n_2856),
.Y(n_4876)
);

INVx2_ASAP7_75t_L g4877 ( 
.A(n_4332),
.Y(n_4877)
);

NAND2xp5_ASAP7_75t_SL g4878 ( 
.A(n_4485),
.B(n_2877),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4399),
.B(n_1116),
.Y(n_4879)
);

INVx3_ASAP7_75t_L g4880 ( 
.A(n_4491),
.Y(n_4880)
);

BUFx6f_ASAP7_75t_L g4881 ( 
.A(n_4363),
.Y(n_4881)
);

NAND3xp33_ASAP7_75t_L g4882 ( 
.A(n_4448),
.B(n_864),
.C(n_859),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_L g4883 ( 
.A(n_4423),
.B(n_859),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_SL g4884 ( 
.A(n_4502),
.B(n_2877),
.Y(n_4884)
);

INVx2_ASAP7_75t_L g4885 ( 
.A(n_4333),
.Y(n_4885)
);

BUFx6f_ASAP7_75t_L g4886 ( 
.A(n_4363),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4428),
.B(n_859),
.Y(n_4887)
);

OAI22xp5_ASAP7_75t_L g4888 ( 
.A1(n_4496),
.A2(n_2894),
.B1(n_2919),
.B2(n_2891),
.Y(n_4888)
);

OAI22xp5_ASAP7_75t_L g4889 ( 
.A1(n_4448),
.A2(n_2894),
.B1(n_2919),
.B2(n_2891),
.Y(n_4889)
);

O2A1O1Ixp5_ASAP7_75t_L g4890 ( 
.A1(n_4440),
.A2(n_1499),
.B(n_1514),
.C(n_1484),
.Y(n_4890)
);

NAND2xp5_ASAP7_75t_L g4891 ( 
.A(n_4444),
.B(n_859),
.Y(n_4891)
);

AND2x4_ASAP7_75t_L g4892 ( 
.A(n_4533),
.B(n_1484),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_SL g4893 ( 
.A(n_4502),
.B(n_2891),
.Y(n_4893)
);

AOI22xp33_ASAP7_75t_L g4894 ( 
.A1(n_4424),
.A2(n_2916),
.B1(n_2918),
.B2(n_2917),
.Y(n_4894)
);

AND2x2_ASAP7_75t_L g4895 ( 
.A(n_4547),
.B(n_864),
.Y(n_4895)
);

OR2x6_ASAP7_75t_L g4896 ( 
.A(n_4471),
.B(n_2843),
.Y(n_4896)
);

NAND2xp5_ASAP7_75t_SL g4897 ( 
.A(n_4502),
.B(n_2894),
.Y(n_4897)
);

INVx2_ASAP7_75t_L g4898 ( 
.A(n_4344),
.Y(n_4898)
);

OAI22xp5_ASAP7_75t_SL g4899 ( 
.A1(n_4299),
.A2(n_929),
.B1(n_938),
.B2(n_935),
.Y(n_4899)
);

INVx1_ASAP7_75t_L g4900 ( 
.A(n_4458),
.Y(n_4900)
);

INVx5_ASAP7_75t_L g4901 ( 
.A(n_4494),
.Y(n_4901)
);

OAI22xp5_ASAP7_75t_L g4902 ( 
.A1(n_4452),
.A2(n_2925),
.B1(n_2959),
.B2(n_2922),
.Y(n_4902)
);

A2O1A1Ixp33_ASAP7_75t_L g4903 ( 
.A1(n_4316),
.A2(n_939),
.B(n_941),
.C(n_940),
.Y(n_4903)
);

BUFx6f_ASAP7_75t_L g4904 ( 
.A(n_4363),
.Y(n_4904)
);

CKINVDCx5p33_ASAP7_75t_R g4905 ( 
.A(n_4421),
.Y(n_4905)
);

NAND2x1p5_ASAP7_75t_L g4906 ( 
.A(n_4502),
.B(n_2922),
.Y(n_4906)
);

INVx1_ASAP7_75t_L g4907 ( 
.A(n_4460),
.Y(n_4907)
);

INVx1_ASAP7_75t_L g4908 ( 
.A(n_4462),
.Y(n_4908)
);

AND2x2_ASAP7_75t_L g4909 ( 
.A(n_4547),
.B(n_4346),
.Y(n_4909)
);

BUFx4f_ASAP7_75t_L g4910 ( 
.A(n_4364),
.Y(n_4910)
);

AND2x2_ASAP7_75t_L g4911 ( 
.A(n_4346),
.B(n_864),
.Y(n_4911)
);

CKINVDCx5p33_ASAP7_75t_R g4912 ( 
.A(n_4257),
.Y(n_4912)
);

NOR2xp33_ASAP7_75t_L g4913 ( 
.A(n_4340),
.B(n_54),
.Y(n_4913)
);

BUFx2_ASAP7_75t_L g4914 ( 
.A(n_4394),
.Y(n_4914)
);

INVx2_ASAP7_75t_L g4915 ( 
.A(n_4349),
.Y(n_4915)
);

CKINVDCx5p33_ASAP7_75t_R g4916 ( 
.A(n_4285),
.Y(n_4916)
);

NAND2xp5_ASAP7_75t_L g4917 ( 
.A(n_4273),
.B(n_864),
.Y(n_4917)
);

BUFx6f_ASAP7_75t_L g4918 ( 
.A(n_4364),
.Y(n_4918)
);

NAND3xp33_ASAP7_75t_L g4919 ( 
.A(n_4459),
.B(n_927),
.C(n_864),
.Y(n_4919)
);

INVx3_ASAP7_75t_L g4920 ( 
.A(n_4533),
.Y(n_4920)
);

NAND2xp5_ASAP7_75t_SL g4921 ( 
.A(n_4364),
.B(n_2925),
.Y(n_4921)
);

AOI21xp5_ASAP7_75t_L g4922 ( 
.A1(n_4275),
.A2(n_2959),
.B(n_2925),
.Y(n_4922)
);

NAND2xp5_ASAP7_75t_SL g4923 ( 
.A(n_4365),
.B(n_2959),
.Y(n_4923)
);

AOI22xp33_ASAP7_75t_L g4924 ( 
.A1(n_4434),
.A2(n_2918),
.B1(n_2927),
.B2(n_2920),
.Y(n_4924)
);

BUFx6f_ASAP7_75t_L g4925 ( 
.A(n_4365),
.Y(n_4925)
);

O2A1O1Ixp33_ASAP7_75t_L g4926 ( 
.A1(n_4504),
.A2(n_2152),
.B(n_2161),
.C(n_2160),
.Y(n_4926)
);

INVx1_ASAP7_75t_L g4927 ( 
.A(n_4590),
.Y(n_4927)
);

AND2x4_ASAP7_75t_L g4928 ( 
.A(n_4430),
.B(n_1499),
.Y(n_4928)
);

AND2x2_ASAP7_75t_L g4929 ( 
.A(n_4394),
.B(n_864),
.Y(n_4929)
);

AOI21x1_ASAP7_75t_L g4930 ( 
.A1(n_4507),
.A2(n_1529),
.B(n_1514),
.Y(n_4930)
);

OR2x2_ASAP7_75t_L g4931 ( 
.A(n_4693),
.B(n_4339),
.Y(n_4931)
);

OAI22xp5_ASAP7_75t_L g4932 ( 
.A1(n_4635),
.A2(n_4264),
.B1(n_4299),
.B2(n_4471),
.Y(n_4932)
);

INVx1_ASAP7_75t_L g4933 ( 
.A(n_4663),
.Y(n_4933)
);

NAND2xp5_ASAP7_75t_L g4934 ( 
.A(n_4769),
.B(n_4789),
.Y(n_4934)
);

AOI22xp5_ASAP7_75t_L g4935 ( 
.A1(n_4722),
.A2(n_4308),
.B1(n_4345),
.B2(n_4348),
.Y(n_4935)
);

NAND2xp5_ASAP7_75t_L g4936 ( 
.A(n_4748),
.B(n_4279),
.Y(n_4936)
);

BUFx2_ASAP7_75t_L g4937 ( 
.A(n_4749),
.Y(n_4937)
);

NAND2xp5_ASAP7_75t_L g4938 ( 
.A(n_4811),
.B(n_4279),
.Y(n_4938)
);

AO31x2_ASAP7_75t_L g4939 ( 
.A1(n_4631),
.A2(n_4338),
.A3(n_4407),
.B(n_4425),
.Y(n_4939)
);

OAI22xp5_ASAP7_75t_L g4940 ( 
.A1(n_4691),
.A2(n_4483),
.B1(n_4471),
.B2(n_4507),
.Y(n_4940)
);

AOI21xp5_ASAP7_75t_SL g4941 ( 
.A1(n_4664),
.A2(n_4288),
.B(n_4280),
.Y(n_4941)
);

O2A1O1Ixp5_ASAP7_75t_SL g4942 ( 
.A1(n_4856),
.A2(n_4406),
.B(n_4410),
.C(n_4401),
.Y(n_4942)
);

CKINVDCx20_ASAP7_75t_R g4943 ( 
.A(n_4665),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_4615),
.B(n_4280),
.Y(n_4944)
);

A2O1A1Ixp33_ASAP7_75t_L g4945 ( 
.A1(n_4710),
.A2(n_4374),
.B(n_4438),
.C(n_4319),
.Y(n_4945)
);

INVx2_ASAP7_75t_L g4946 ( 
.A(n_4669),
.Y(n_4946)
);

NAND2xp5_ASAP7_75t_L g4947 ( 
.A(n_4615),
.B(n_4288),
.Y(n_4947)
);

INVx8_ASAP7_75t_L g4948 ( 
.A(n_4677),
.Y(n_4948)
);

AOI21x1_ASAP7_75t_L g4949 ( 
.A1(n_4917),
.A2(n_4466),
.B(n_4461),
.Y(n_4949)
);

NAND2xp5_ASAP7_75t_L g4950 ( 
.A(n_4709),
.B(n_4301),
.Y(n_4950)
);

OAI21xp5_ASAP7_75t_L g4951 ( 
.A1(n_4634),
.A2(n_4486),
.B(n_4543),
.Y(n_4951)
);

NAND2xp5_ASAP7_75t_L g4952 ( 
.A(n_4729),
.B(n_4303),
.Y(n_4952)
);

NOR2xp67_ASAP7_75t_SL g4953 ( 
.A(n_4605),
.B(n_4494),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4736),
.B(n_4515),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_4730),
.B(n_4515),
.Y(n_4955)
);

OAI21x1_ASAP7_75t_L g4956 ( 
.A1(n_4930),
.A2(n_4425),
.B(n_4407),
.Y(n_4956)
);

AOI21xp5_ASAP7_75t_L g4957 ( 
.A1(n_4623),
.A2(n_4420),
.B(n_4549),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4728),
.Y(n_4958)
);

AOI21xp5_ASAP7_75t_L g4959 ( 
.A1(n_4625),
.A2(n_4541),
.B(n_4283),
.Y(n_4959)
);

INVx2_ASAP7_75t_SL g4960 ( 
.A(n_4624),
.Y(n_4960)
);

O2A1O1Ixp5_ASAP7_75t_L g4961 ( 
.A1(n_4737),
.A2(n_4406),
.B(n_4410),
.C(n_4401),
.Y(n_4961)
);

OAI21x1_ASAP7_75t_L g4962 ( 
.A1(n_4652),
.A2(n_4563),
.B(n_4561),
.Y(n_4962)
);

AND2x6_ASAP7_75t_L g4963 ( 
.A(n_4618),
.B(n_4345),
.Y(n_4963)
);

AOI21xp5_ASAP7_75t_L g4964 ( 
.A1(n_4701),
.A2(n_4283),
.B(n_4561),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_4654),
.A2(n_4483),
.B1(n_4574),
.B2(n_4548),
.Y(n_4965)
);

OAI21x1_ASAP7_75t_SL g4966 ( 
.A1(n_4861),
.A2(n_4723),
.B(n_4719),
.Y(n_4966)
);

AO31x2_ASAP7_75t_L g4967 ( 
.A1(n_4683),
.A2(n_4563),
.A3(n_4604),
.B(n_4595),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4752),
.Y(n_4968)
);

OAI21x1_ASAP7_75t_L g4969 ( 
.A1(n_4647),
.A2(n_4604),
.B(n_4595),
.Y(n_4969)
);

HB1xp67_ASAP7_75t_L g4970 ( 
.A(n_4649),
.Y(n_4970)
);

INVx2_ASAP7_75t_L g4971 ( 
.A(n_4680),
.Y(n_4971)
);

AOI221xp5_ASAP7_75t_L g4972 ( 
.A1(n_4702),
.A2(n_4742),
.B1(n_4735),
.B2(n_4689),
.C(n_4675),
.Y(n_4972)
);

AOI22xp5_ASAP7_75t_L g4973 ( 
.A1(n_4701),
.A2(n_4348),
.B1(n_4314),
.B2(n_4412),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4754),
.B(n_4522),
.Y(n_4974)
);

NAND2xp5_ASAP7_75t_L g4975 ( 
.A(n_4611),
.B(n_4522),
.Y(n_4975)
);

BUFx10_ASAP7_75t_L g4976 ( 
.A(n_4750),
.Y(n_4976)
);

INVx2_ASAP7_75t_L g4977 ( 
.A(n_4716),
.Y(n_4977)
);

INVx5_ASAP7_75t_L g4978 ( 
.A(n_4608),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4626),
.B(n_4632),
.Y(n_4979)
);

CKINVDCx20_ASAP7_75t_R g4980 ( 
.A(n_4667),
.Y(n_4980)
);

A2O1A1Ixp33_ASAP7_75t_L g4981 ( 
.A1(n_4616),
.A2(n_4523),
.B(n_4314),
.C(n_4576),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4637),
.B(n_4527),
.Y(n_4982)
);

A2O1A1Ixp33_ASAP7_75t_L g4983 ( 
.A1(n_4849),
.A2(n_4430),
.B(n_4555),
.C(n_4426),
.Y(n_4983)
);

OA21x2_ASAP7_75t_L g4984 ( 
.A1(n_4648),
.A2(n_4555),
.B(n_4540),
.Y(n_4984)
);

NAND3x1_ASAP7_75t_L g4985 ( 
.A(n_4653),
.B(n_4574),
.C(n_4548),
.Y(n_4985)
);

OR2x2_ASAP7_75t_L g4986 ( 
.A(n_4927),
.B(n_4313),
.Y(n_4986)
);

CKINVDCx5p33_ASAP7_75t_R g4987 ( 
.A(n_4620),
.Y(n_4987)
);

OAI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_4834),
.A2(n_4536),
.B(n_4540),
.Y(n_4988)
);

INVx2_ASAP7_75t_SL g4989 ( 
.A(n_4628),
.Y(n_4989)
);

AO31x2_ASAP7_75t_L g4990 ( 
.A1(n_4673),
.A2(n_4552),
.A3(n_4536),
.B(n_4368),
.Y(n_4990)
);

INVx2_ASAP7_75t_L g4991 ( 
.A(n_4717),
.Y(n_4991)
);

BUFx6f_ASAP7_75t_L g4992 ( 
.A(n_4846),
.Y(n_4992)
);

A2O1A1Ixp33_ASAP7_75t_L g4993 ( 
.A1(n_4735),
.A2(n_4430),
.B(n_4337),
.C(n_4570),
.Y(n_4993)
);

NAND3xp33_ASAP7_75t_L g4994 ( 
.A(n_4621),
.B(n_4395),
.C(n_4359),
.Y(n_4994)
);

INVx3_ASAP7_75t_L g4995 ( 
.A(n_4847),
.Y(n_4995)
);

AOI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4606),
.A2(n_4432),
.B(n_4396),
.Y(n_4996)
);

OAI22x1_ASAP7_75t_L g4997 ( 
.A1(n_4787),
.A2(n_4564),
.B1(n_4412),
.B2(n_4535),
.Y(n_4997)
);

INVxp67_ASAP7_75t_SL g4998 ( 
.A(n_4633),
.Y(n_4998)
);

O2A1O1Ixp5_ASAP7_75t_L g4999 ( 
.A1(n_4734),
.A2(n_4359),
.B(n_4463),
.C(n_4443),
.Y(n_4999)
);

INVx1_ASAP7_75t_L g5000 ( 
.A(n_4762),
.Y(n_5000)
);

OAI21xp5_ASAP7_75t_L g5001 ( 
.A1(n_4840),
.A2(n_4585),
.B(n_4581),
.Y(n_5001)
);

NAND2xp5_ASAP7_75t_SL g5002 ( 
.A(n_4867),
.B(n_4285),
.Y(n_5002)
);

AND2x4_ASAP7_75t_L g5003 ( 
.A(n_4819),
.B(n_4290),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4686),
.A2(n_4463),
.B(n_4443),
.Y(n_5004)
);

AO31x2_ASAP7_75t_L g5005 ( 
.A1(n_4697),
.A2(n_4371),
.A3(n_4372),
.B(n_4352),
.Y(n_5005)
);

OAI21xp5_ASAP7_75t_L g5006 ( 
.A1(n_4790),
.A2(n_4585),
.B(n_943),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4639),
.B(n_4378),
.Y(n_5007)
);

OAI21xp5_ASAP7_75t_L g5008 ( 
.A1(n_4800),
.A2(n_945),
.B(n_942),
.Y(n_5008)
);

NOR2xp33_ASAP7_75t_L g5009 ( 
.A(n_4727),
.B(n_4534),
.Y(n_5009)
);

AND2x4_ASAP7_75t_L g5010 ( 
.A(n_4829),
.B(n_4290),
.Y(n_5010)
);

BUFx8_ASAP7_75t_L g5011 ( 
.A(n_4771),
.Y(n_5011)
);

O2A1O1Ixp5_ASAP7_75t_SL g5012 ( 
.A1(n_4731),
.A2(n_4865),
.B(n_4879),
.C(n_4871),
.Y(n_5012)
);

BUFx4f_ASAP7_75t_SL g5013 ( 
.A(n_4799),
.Y(n_5013)
);

NAND2xp5_ASAP7_75t_SL g5014 ( 
.A(n_4905),
.B(n_4640),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4768),
.B(n_4381),
.Y(n_5015)
);

NOR2xp33_ASAP7_75t_L g5016 ( 
.A(n_4643),
.B(n_4534),
.Y(n_5016)
);

NAND2xp5_ASAP7_75t_SL g5017 ( 
.A(n_4640),
.B(n_4290),
.Y(n_5017)
);

OAI21x1_ASAP7_75t_L g5018 ( 
.A1(n_4674),
.A2(n_4414),
.B(n_4413),
.Y(n_5018)
);

NAND2xp5_ASAP7_75t_L g5019 ( 
.A(n_4746),
.B(n_4481),
.Y(n_5019)
);

OR2x6_ASAP7_75t_L g5020 ( 
.A(n_4608),
.B(n_4306),
.Y(n_5020)
);

AOI21x1_ASAP7_75t_L g5021 ( 
.A1(n_4860),
.A2(n_4524),
.B(n_4589),
.Y(n_5021)
);

NAND2xp5_ASAP7_75t_SL g5022 ( 
.A(n_4660),
.B(n_4306),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_4609),
.B(n_4535),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_4794),
.B(n_4306),
.Y(n_5024)
);

OAI21x1_ASAP7_75t_L g5025 ( 
.A1(n_4807),
.A2(n_4320),
.B(n_2511),
.Y(n_5025)
);

INVx2_ASAP7_75t_SL g5026 ( 
.A(n_4815),
.Y(n_5026)
);

INVx4_ASAP7_75t_L g5027 ( 
.A(n_4660),
.Y(n_5027)
);

NOR2xp33_ASAP7_75t_R g5028 ( 
.A(n_4785),
.B(n_4365),
.Y(n_5028)
);

AO31x2_ASAP7_75t_L g5029 ( 
.A1(n_4883),
.A2(n_1572),
.A3(n_1529),
.B(n_3003),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4804),
.B(n_4327),
.Y(n_5030)
);

AND2x4_ASAP7_75t_L g5031 ( 
.A(n_4773),
.B(n_4327),
.Y(n_5031)
);

OAI21xp5_ASAP7_75t_L g5032 ( 
.A1(n_4797),
.A2(n_955),
.B(n_954),
.Y(n_5032)
);

OA21x2_ASAP7_75t_L g5033 ( 
.A1(n_4887),
.A2(n_4597),
.B(n_4589),
.Y(n_5033)
);

AND3x2_ASAP7_75t_L g5034 ( 
.A(n_4645),
.B(n_4662),
.C(n_4614),
.Y(n_5034)
);

AOI21x1_ASAP7_75t_L g5035 ( 
.A1(n_4741),
.A2(n_4597),
.B(n_4567),
.Y(n_5035)
);

NAND2xp5_ASAP7_75t_SL g5036 ( 
.A(n_4725),
.B(n_4336),
.Y(n_5036)
);

NAND2xp5_ASAP7_75t_SL g5037 ( 
.A(n_4725),
.B(n_4336),
.Y(n_5037)
);

AOI21xp5_ASAP7_75t_L g5038 ( 
.A1(n_4642),
.A2(n_4567),
.B(n_4553),
.Y(n_5038)
);

AOI21xp5_ASAP7_75t_L g5039 ( 
.A1(n_4614),
.A2(n_4569),
.B(n_4553),
.Y(n_5039)
);

OAI21x1_ASAP7_75t_L g5040 ( 
.A1(n_4646),
.A2(n_4666),
.B(n_4855),
.Y(n_5040)
);

AOI21xp5_ASAP7_75t_L g5041 ( 
.A1(n_4662),
.A2(n_4681),
.B(n_4764),
.Y(n_5041)
);

OAI21x1_ASAP7_75t_SL g5042 ( 
.A1(n_4872),
.A2(n_2171),
.B(n_2167),
.Y(n_5042)
);

NOR2xp33_ASAP7_75t_L g5043 ( 
.A(n_4692),
.B(n_4336),
.Y(n_5043)
);

AND2x2_ASAP7_75t_L g5044 ( 
.A(n_4656),
.B(n_4579),
.Y(n_5044)
);

AOI211x1_ASAP7_75t_L g5045 ( 
.A1(n_4708),
.A2(n_11),
.B(n_9),
.C(n_10),
.Y(n_5045)
);

AOI22xp33_ASAP7_75t_L g5046 ( 
.A1(n_4627),
.A2(n_4630),
.B1(n_4742),
.B2(n_4696),
.Y(n_5046)
);

AO22x2_ASAP7_75t_L g5047 ( 
.A1(n_4726),
.A2(n_4569),
.B1(n_4577),
.B2(n_4528),
.Y(n_5047)
);

OAI21xp5_ASAP7_75t_L g5048 ( 
.A1(n_4641),
.A2(n_960),
.B(n_959),
.Y(n_5048)
);

BUFx6f_ASAP7_75t_L g5049 ( 
.A(n_4812),
.Y(n_5049)
);

CKINVDCx5p33_ASAP7_75t_R g5050 ( 
.A(n_4912),
.Y(n_5050)
);

NOR2xp33_ASAP7_75t_L g5051 ( 
.A(n_4699),
.B(n_55),
.Y(n_5051)
);

INVx2_ASAP7_75t_SL g5052 ( 
.A(n_4629),
.Y(n_5052)
);

AOI21xp5_ASAP7_75t_L g5053 ( 
.A1(n_4766),
.A2(n_4577),
.B(n_2965),
.Y(n_5053)
);

NOR2xp33_ASAP7_75t_L g5054 ( 
.A(n_4672),
.B(n_55),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_4916),
.Y(n_5055)
);

AOI21xp5_ASAP7_75t_L g5056 ( 
.A1(n_4767),
.A2(n_4682),
.B(n_4851),
.Y(n_5056)
);

AO31x2_ASAP7_75t_L g5057 ( 
.A1(n_4891),
.A2(n_1572),
.A3(n_3006),
.B(n_3005),
.Y(n_5057)
);

AOI21xp5_ASAP7_75t_L g5058 ( 
.A1(n_4926),
.A2(n_2965),
.B(n_2963),
.Y(n_5058)
);

AND3x4_ASAP7_75t_L g5059 ( 
.A(n_4618),
.B(n_2171),
.C(n_2167),
.Y(n_5059)
);

HB1xp67_ASAP7_75t_L g5060 ( 
.A(n_4848),
.Y(n_5060)
);

BUFx3_ASAP7_75t_L g5061 ( 
.A(n_4617),
.Y(n_5061)
);

NAND2xp5_ASAP7_75t_L g5062 ( 
.A(n_4862),
.B(n_4579),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4863),
.B(n_4579),
.Y(n_5063)
);

BUFx6f_ASAP7_75t_L g5064 ( 
.A(n_4812),
.Y(n_5064)
);

O2A1O1Ixp5_ASAP7_75t_L g5065 ( 
.A1(n_4836),
.A2(n_2963),
.B(n_3026),
.C(n_2971),
.Y(n_5065)
);

AOI21xp5_ASAP7_75t_L g5066 ( 
.A1(n_4688),
.A2(n_3026),
.B(n_2971),
.Y(n_5066)
);

AOI221x1_ASAP7_75t_L g5067 ( 
.A1(n_4837),
.A2(n_4592),
.B1(n_1120),
.B2(n_1018),
.C(n_927),
.Y(n_5067)
);

BUFx10_ASAP7_75t_L g5068 ( 
.A(n_4913),
.Y(n_5068)
);

INVx3_ASAP7_75t_L g5069 ( 
.A(n_4847),
.Y(n_5069)
);

NAND2xp5_ASAP7_75t_L g5070 ( 
.A(n_4868),
.B(n_4870),
.Y(n_5070)
);

OAI21x1_ASAP7_75t_L g5071 ( 
.A1(n_4646),
.A2(n_3026),
.B(n_2971),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4900),
.B(n_4284),
.Y(n_5072)
);

INVx1_ASAP7_75t_SL g5073 ( 
.A(n_4706),
.Y(n_5073)
);

OR2x6_ASAP7_75t_L g5074 ( 
.A(n_4608),
.B(n_4284),
.Y(n_5074)
);

OAI21x1_ASAP7_75t_L g5075 ( 
.A1(n_4666),
.A2(n_3047),
.B(n_3041),
.Y(n_5075)
);

O2A1O1Ixp33_ASAP7_75t_L g5076 ( 
.A1(n_4657),
.A2(n_2131),
.B(n_2065),
.C(n_2068),
.Y(n_5076)
);

AOI21xp5_ASAP7_75t_L g5077 ( 
.A1(n_4853),
.A2(n_3047),
.B(n_3041),
.Y(n_5077)
);

NOR2xp33_ASAP7_75t_L g5078 ( 
.A(n_4858),
.B(n_4619),
.Y(n_5078)
);

BUFx10_ASAP7_75t_L g5079 ( 
.A(n_4810),
.Y(n_5079)
);

OR2x6_ASAP7_75t_L g5080 ( 
.A(n_4721),
.B(n_4284),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4907),
.Y(n_5081)
);

OAI21xp33_ASAP7_75t_SL g5082 ( 
.A1(n_4715),
.A2(n_12),
.B(n_14),
.Y(n_5082)
);

NAND3xp33_ASAP7_75t_L g5083 ( 
.A(n_4694),
.B(n_1018),
.C(n_927),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4908),
.Y(n_5084)
);

INVx4_ASAP7_75t_L g5085 ( 
.A(n_4812),
.Y(n_5085)
);

AOI21xp33_ASAP7_75t_L g5086 ( 
.A1(n_4705),
.A2(n_1018),
.B(n_927),
.Y(n_5086)
);

A2O1A1Ixp33_ASAP7_75t_L g5087 ( 
.A1(n_4718),
.A2(n_984),
.B(n_1017),
.C(n_974),
.Y(n_5087)
);

NAND2xp5_ASAP7_75t_SL g5088 ( 
.A(n_4622),
.B(n_927),
.Y(n_5088)
);

OAI21xp5_ASAP7_75t_L g5089 ( 
.A1(n_4882),
.A2(n_965),
.B(n_964),
.Y(n_5089)
);

O2A1O1Ixp33_ASAP7_75t_SL g5090 ( 
.A1(n_4774),
.A2(n_15),
.B(n_12),
.C(n_14),
.Y(n_5090)
);

NAND2xp5_ASAP7_75t_L g5091 ( 
.A(n_4832),
.B(n_4284),
.Y(n_5091)
);

NAND2xp5_ASAP7_75t_L g5092 ( 
.A(n_4651),
.B(n_1018),
.Y(n_5092)
);

AOI21x1_ASAP7_75t_L g5093 ( 
.A1(n_4757),
.A2(n_2068),
.B(n_2049),
.Y(n_5093)
);

AOI221xp5_ASAP7_75t_SL g5094 ( 
.A1(n_4732),
.A2(n_1120),
.B1(n_1018),
.B2(n_17),
.C(n_12),
.Y(n_5094)
);

HB1xp67_ASAP7_75t_L g5095 ( 
.A(n_4777),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4919),
.A2(n_3047),
.B(n_3041),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_L g5097 ( 
.A(n_4687),
.B(n_4690),
.Y(n_5097)
);

OAI21x1_ASAP7_75t_L g5098 ( 
.A1(n_4655),
.A2(n_3094),
.B(n_3069),
.Y(n_5098)
);

OAI21xp5_ASAP7_75t_SL g5099 ( 
.A1(n_4783),
.A2(n_1120),
.B(n_16),
.Y(n_5099)
);

HB1xp67_ASAP7_75t_L g5100 ( 
.A(n_4788),
.Y(n_5100)
);

INVx2_ASAP7_75t_SL g5101 ( 
.A(n_4909),
.Y(n_5101)
);

OAI21x1_ASAP7_75t_L g5102 ( 
.A1(n_4636),
.A2(n_3094),
.B(n_3069),
.Y(n_5102)
);

OAI21x1_ASAP7_75t_L g5103 ( 
.A1(n_4636),
.A2(n_3094),
.B(n_3069),
.Y(n_5103)
);

INVxp67_ASAP7_75t_L g5104 ( 
.A(n_4914),
.Y(n_5104)
);

AO31x2_ASAP7_75t_L g5105 ( 
.A1(n_4733),
.A2(n_3012),
.A3(n_3016),
.B(n_3006),
.Y(n_5105)
);

OAI21xp5_ASAP7_75t_SL g5106 ( 
.A1(n_4791),
.A2(n_1120),
.B(n_18),
.Y(n_5106)
);

INVx3_ASAP7_75t_L g5107 ( 
.A(n_4852),
.Y(n_5107)
);

HB1xp67_ASAP7_75t_L g5108 ( 
.A(n_4852),
.Y(n_5108)
);

AOI21xp5_ASAP7_75t_L g5109 ( 
.A1(n_4919),
.A2(n_3154),
.B(n_3112),
.Y(n_5109)
);

NAND2xp5_ASAP7_75t_L g5110 ( 
.A(n_4814),
.B(n_973),
.Y(n_5110)
);

NOR3xp33_ASAP7_75t_L g5111 ( 
.A(n_4740),
.B(n_4751),
.C(n_4744),
.Y(n_5111)
);

AOI22xp5_ASAP7_75t_L g5112 ( 
.A1(n_4899),
.A2(n_1001),
.B1(n_976),
.B2(n_2015),
.Y(n_5112)
);

OR2x2_ASAP7_75t_L g5113 ( 
.A(n_4668),
.B(n_1210),
.Y(n_5113)
);

AO31x2_ASAP7_75t_L g5114 ( 
.A1(n_4792),
.A2(n_4813),
.A3(n_4676),
.B(n_4658),
.Y(n_5114)
);

NAND2xp33_ASAP7_75t_L g5115 ( 
.A(n_4899),
.B(n_975),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_4704),
.Y(n_5116)
);

AOI21xp5_ASAP7_75t_L g5117 ( 
.A1(n_4758),
.A2(n_3154),
.B(n_3112),
.Y(n_5117)
);

BUFx2_ASAP7_75t_L g5118 ( 
.A(n_4776),
.Y(n_5118)
);

AOI21xp5_ASAP7_75t_L g5119 ( 
.A1(n_4760),
.A2(n_3154),
.B(n_3112),
.Y(n_5119)
);

OAI21x1_ASAP7_75t_L g5120 ( 
.A1(n_4638),
.A2(n_3214),
.B(n_3173),
.Y(n_5120)
);

NAND2xp5_ASAP7_75t_L g5121 ( 
.A(n_4875),
.B(n_977),
.Y(n_5121)
);

NOR2xp33_ASAP7_75t_L g5122 ( 
.A(n_4671),
.B(n_57),
.Y(n_5122)
);

INVx5_ASAP7_75t_L g5123 ( 
.A(n_4896),
.Y(n_5123)
);

AOI21xp5_ASAP7_75t_L g5124 ( 
.A1(n_4670),
.A2(n_3214),
.B(n_3173),
.Y(n_5124)
);

AND2x2_ASAP7_75t_L g5125 ( 
.A(n_4776),
.B(n_18),
.Y(n_5125)
);

AOI21xp5_ASAP7_75t_L g5126 ( 
.A1(n_4678),
.A2(n_3173),
.B(n_2867),
.Y(n_5126)
);

BUFx2_ASAP7_75t_L g5127 ( 
.A(n_4880),
.Y(n_5127)
);

NAND3xp33_ASAP7_75t_L g5128 ( 
.A(n_4850),
.B(n_4859),
.C(n_4759),
.Y(n_5128)
);

AOI21xp5_ASAP7_75t_L g5129 ( 
.A1(n_4784),
.A2(n_2867),
.B(n_2843),
.Y(n_5129)
);

OAI21x1_ASAP7_75t_L g5130 ( 
.A1(n_4684),
.A2(n_3016),
.B(n_3012),
.Y(n_5130)
);

OAI21xp5_ASAP7_75t_L g5131 ( 
.A1(n_4661),
.A2(n_4903),
.B(n_4874),
.Y(n_5131)
);

INVx3_ASAP7_75t_SL g5132 ( 
.A(n_4713),
.Y(n_5132)
);

INVx4_ASAP7_75t_L g5133 ( 
.A(n_4820),
.Y(n_5133)
);

OAI21x1_ASAP7_75t_L g5134 ( 
.A1(n_4684),
.A2(n_3025),
.B(n_3020),
.Y(n_5134)
);

NAND2xp5_ASAP7_75t_L g5135 ( 
.A(n_4761),
.B(n_981),
.Y(n_5135)
);

INVx3_ASAP7_75t_L g5136 ( 
.A(n_4880),
.Y(n_5136)
);

OAI21xp5_ASAP7_75t_L g5137 ( 
.A1(n_4842),
.A2(n_4793),
.B(n_4747),
.Y(n_5137)
);

OAI22xp5_ASAP7_75t_L g5138 ( 
.A1(n_4607),
.A2(n_985),
.B1(n_987),
.B2(n_986),
.Y(n_5138)
);

OA21x2_ASAP7_75t_L g5139 ( 
.A1(n_4778),
.A2(n_992),
.B(n_989),
.Y(n_5139)
);

OAI21x1_ASAP7_75t_L g5140 ( 
.A1(n_4650),
.A2(n_3025),
.B(n_3020),
.Y(n_5140)
);

INVx2_ASAP7_75t_L g5141 ( 
.A(n_4825),
.Y(n_5141)
);

AOI21xp5_ASAP7_75t_L g5142 ( 
.A1(n_4650),
.A2(n_2914),
.B(n_2890),
.Y(n_5142)
);

INVx1_ASAP7_75t_SL g5143 ( 
.A(n_4738),
.Y(n_5143)
);

NAND2xp5_ASAP7_75t_L g5144 ( 
.A(n_4786),
.B(n_993),
.Y(n_5144)
);

OAI21x1_ASAP7_75t_L g5145 ( 
.A1(n_4922),
.A2(n_4876),
.B(n_4869),
.Y(n_5145)
);

NAND3x1_ASAP7_75t_L g5146 ( 
.A(n_4644),
.B(n_18),
.C(n_19),
.Y(n_5146)
);

OAI22xp5_ASAP7_75t_L g5147 ( 
.A1(n_4612),
.A2(n_4826),
.B1(n_4763),
.B2(n_4627),
.Y(n_5147)
);

BUFx2_ASAP7_75t_L g5148 ( 
.A(n_4920),
.Y(n_5148)
);

OAI21xp5_ASAP7_75t_L g5149 ( 
.A1(n_4817),
.A2(n_1002),
.B(n_997),
.Y(n_5149)
);

AOI21xp5_ASAP7_75t_L g5150 ( 
.A1(n_4878),
.A2(n_2914),
.B(n_2890),
.Y(n_5150)
);

OAI21x1_ASAP7_75t_L g5151 ( 
.A1(n_4818),
.A2(n_3042),
.B(n_3040),
.Y(n_5151)
);

OAI22xp5_ASAP7_75t_L g5152 ( 
.A1(n_4775),
.A2(n_1004),
.B1(n_1009),
.B2(n_1003),
.Y(n_5152)
);

BUFx3_ASAP7_75t_L g5153 ( 
.A(n_4613),
.Y(n_5153)
);

NOR3xp33_ASAP7_75t_L g5154 ( 
.A(n_4821),
.B(n_1013),
.C(n_1010),
.Y(n_5154)
);

OAI21x1_ASAP7_75t_L g5155 ( 
.A1(n_4823),
.A2(n_3045),
.B(n_3043),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_L g5156 ( 
.A(n_4796),
.B(n_1015),
.Y(n_5156)
);

NOR2xp33_ASAP7_75t_R g5157 ( 
.A(n_4795),
.B(n_57),
.Y(n_5157)
);

AO31x2_ASAP7_75t_L g5158 ( 
.A1(n_4835),
.A2(n_3045),
.A3(n_3046),
.B(n_3043),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4801),
.B(n_1019),
.Y(n_5159)
);

INVx3_ASAP7_75t_L g5160 ( 
.A(n_4773),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_4802),
.B(n_4803),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_4805),
.B(n_1022),
.Y(n_5162)
);

NOR2xp33_ASAP7_75t_L g5163 ( 
.A(n_4866),
.B(n_59),
.Y(n_5163)
);

AOI21xp33_ASAP7_75t_L g5164 ( 
.A1(n_4830),
.A2(n_4864),
.B(n_4854),
.Y(n_5164)
);

OAI21x1_ASAP7_75t_L g5165 ( 
.A1(n_4753),
.A2(n_4703),
.B(n_4695),
.Y(n_5165)
);

AOI31xp67_ASAP7_75t_L g5166 ( 
.A1(n_4770),
.A2(n_1474),
.A3(n_1482),
.B(n_1471),
.Y(n_5166)
);

AOI22xp5_ASAP7_75t_L g5167 ( 
.A1(n_4822),
.A2(n_1001),
.B1(n_976),
.B2(n_2015),
.Y(n_5167)
);

AOI21xp5_ASAP7_75t_L g5168 ( 
.A1(n_4884),
.A2(n_2932),
.B(n_2924),
.Y(n_5168)
);

BUFx5_ASAP7_75t_L g5169 ( 
.A(n_4928),
.Y(n_5169)
);

OAI21x1_ASAP7_75t_L g5170 ( 
.A1(n_4707),
.A2(n_3052),
.B(n_3048),
.Y(n_5170)
);

A2O1A1Ixp33_ASAP7_75t_L g5171 ( 
.A1(n_4780),
.A2(n_1039),
.B(n_1054),
.C(n_1028),
.Y(n_5171)
);

OAI21xp33_ASAP7_75t_L g5172 ( 
.A1(n_4780),
.A2(n_4895),
.B(n_4911),
.Y(n_5172)
);

AO31x2_ASAP7_75t_L g5173 ( 
.A1(n_4839),
.A2(n_3060),
.A3(n_3061),
.B(n_3052),
.Y(n_5173)
);

OAI22xp5_ASAP7_75t_L g5174 ( 
.A1(n_4679),
.A2(n_1027),
.B1(n_1030),
.B2(n_1026),
.Y(n_5174)
);

AO31x2_ASAP7_75t_L g5175 ( 
.A1(n_4845),
.A2(n_3061),
.A3(n_3064),
.B(n_3060),
.Y(n_5175)
);

INVx2_ASAP7_75t_L g5176 ( 
.A(n_4857),
.Y(n_5176)
);

OAI21x1_ASAP7_75t_L g5177 ( 
.A1(n_4843),
.A2(n_3070),
.B(n_3064),
.Y(n_5177)
);

AO32x2_ASAP7_75t_L g5178 ( 
.A1(n_4822),
.A2(n_2839),
.A3(n_2836),
.B1(n_2828),
.B2(n_2924),
.Y(n_5178)
);

OAI21x1_ASAP7_75t_L g5179 ( 
.A1(n_4720),
.A2(n_3088),
.B(n_3073),
.Y(n_5179)
);

OAI21x1_ASAP7_75t_L g5180 ( 
.A1(n_4711),
.A2(n_3105),
.B(n_3088),
.Y(n_5180)
);

A2O1A1Ixp33_ASAP7_75t_L g5181 ( 
.A1(n_4610),
.A2(n_1063),
.B(n_1088),
.C(n_1042),
.Y(n_5181)
);

A2O1A1Ixp33_ASAP7_75t_L g5182 ( 
.A1(n_4743),
.A2(n_1069),
.B(n_1093),
.C(n_1044),
.Y(n_5182)
);

INVx2_ASAP7_75t_L g5183 ( 
.A(n_4877),
.Y(n_5183)
);

OA21x2_ASAP7_75t_L g5184 ( 
.A1(n_4816),
.A2(n_1035),
.B(n_1032),
.Y(n_5184)
);

INVx1_ASAP7_75t_L g5185 ( 
.A(n_4885),
.Y(n_5185)
);

NOR2xp67_ASAP7_75t_SL g5186 ( 
.A(n_4605),
.B(n_2391),
.Y(n_5186)
);

INVx3_ASAP7_75t_L g5187 ( 
.A(n_4605),
.Y(n_5187)
);

AOI21xp5_ASAP7_75t_L g5188 ( 
.A1(n_4893),
.A2(n_2939),
.B(n_2932),
.Y(n_5188)
);

BUFx12f_ASAP7_75t_L g5189 ( 
.A(n_4659),
.Y(n_5189)
);

AOI221xp5_ASAP7_75t_SL g5190 ( 
.A1(n_4888),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.C(n_22),
.Y(n_5190)
);

O2A1O1Ixp5_ASAP7_75t_SL g5191 ( 
.A1(n_4831),
.A2(n_2070),
.B(n_2072),
.C(n_2069),
.Y(n_5191)
);

NOR4xp25_ASAP7_75t_L g5192 ( 
.A(n_4833),
.B(n_1001),
.C(n_976),
.D(n_21),
.Y(n_5192)
);

A2O1A1Ixp33_ASAP7_75t_L g5193 ( 
.A1(n_4844),
.A2(n_1091),
.B(n_1107),
.C(n_1058),
.Y(n_5193)
);

AOI21xp5_ASAP7_75t_L g5194 ( 
.A1(n_4897),
.A2(n_2978),
.B(n_2939),
.Y(n_5194)
);

AOI22xp5_ASAP7_75t_L g5195 ( 
.A1(n_4838),
.A2(n_1001),
.B1(n_2052),
.B2(n_2015),
.Y(n_5195)
);

OAI21x1_ASAP7_75t_L g5196 ( 
.A1(n_4841),
.A2(n_3111),
.B(n_3108),
.Y(n_5196)
);

BUFx6f_ASAP7_75t_L g5197 ( 
.A(n_4820),
.Y(n_5197)
);

A2O1A1Ixp33_ASAP7_75t_L g5198 ( 
.A1(n_5099),
.A2(n_4910),
.B(n_4798),
.C(n_4700),
.Y(n_5198)
);

NAND2xp5_ASAP7_75t_L g5199 ( 
.A(n_4974),
.B(n_4929),
.Y(n_5199)
);

NAND2xp5_ASAP7_75t_L g5200 ( 
.A(n_4952),
.B(n_4892),
.Y(n_5200)
);

AOI22xp33_ASAP7_75t_L g5201 ( 
.A1(n_5046),
.A2(n_4894),
.B1(n_4924),
.B2(n_4928),
.Y(n_5201)
);

AND2x2_ASAP7_75t_L g5202 ( 
.A(n_5160),
.B(n_5101),
.Y(n_5202)
);

BUFx4f_ASAP7_75t_SL g5203 ( 
.A(n_4943),
.Y(n_5203)
);

AND2x2_ASAP7_75t_L g5204 ( 
.A(n_4937),
.B(n_4756),
.Y(n_5204)
);

CKINVDCx5p33_ASAP7_75t_R g5205 ( 
.A(n_4987),
.Y(n_5205)
);

BUFx2_ASAP7_75t_L g5206 ( 
.A(n_5028),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5113),
.Y(n_5207)
);

AND2x2_ASAP7_75t_L g5208 ( 
.A(n_4970),
.B(n_4756),
.Y(n_5208)
);

INVx2_ASAP7_75t_L g5209 ( 
.A(n_5018),
.Y(n_5209)
);

INVx3_ASAP7_75t_L g5210 ( 
.A(n_4995),
.Y(n_5210)
);

AOI21xp5_ASAP7_75t_L g5211 ( 
.A1(n_4964),
.A2(n_4910),
.B(n_4782),
.Y(n_5211)
);

INVx1_ASAP7_75t_L g5212 ( 
.A(n_5060),
.Y(n_5212)
);

CKINVDCx11_ASAP7_75t_R g5213 ( 
.A(n_4980),
.Y(n_5213)
);

AOI21xp5_ASAP7_75t_L g5214 ( 
.A1(n_5041),
.A2(n_4781),
.B(n_4685),
.Y(n_5214)
);

O2A1O1Ixp33_ASAP7_75t_L g5215 ( 
.A1(n_5106),
.A2(n_4889),
.B(n_4902),
.C(n_4824),
.Y(n_5215)
);

AOI21xp5_ASAP7_75t_L g5216 ( 
.A1(n_5147),
.A2(n_4809),
.B(n_4921),
.Y(n_5216)
);

AOI22xp33_ASAP7_75t_L g5217 ( 
.A1(n_5111),
.A2(n_4739),
.B1(n_4873),
.B2(n_4898),
.Y(n_5217)
);

AND2x4_ASAP7_75t_L g5218 ( 
.A(n_5123),
.B(n_4901),
.Y(n_5218)
);

OAI22xp33_ASAP7_75t_L g5219 ( 
.A1(n_5167),
.A2(n_4896),
.B1(n_4828),
.B2(n_4698),
.Y(n_5219)
);

NAND2x1p5_ASAP7_75t_L g5220 ( 
.A(n_4978),
.B(n_4901),
.Y(n_5220)
);

O2A1O1Ixp5_ASAP7_75t_L g5221 ( 
.A1(n_4961),
.A2(n_4923),
.B(n_4739),
.C(n_4808),
.Y(n_5221)
);

AOI22xp33_ASAP7_75t_L g5222 ( 
.A1(n_5139),
.A2(n_4915),
.B1(n_4698),
.B2(n_4714),
.Y(n_5222)
);

HB1xp67_ASAP7_75t_L g5223 ( 
.A(n_4934),
.Y(n_5223)
);

OR2x6_ASAP7_75t_L g5224 ( 
.A(n_5038),
.B(n_5080),
.Y(n_5224)
);

AOI21xp5_ASAP7_75t_L g5225 ( 
.A1(n_4941),
.A2(n_4896),
.B(n_4828),
.Y(n_5225)
);

BUFx10_ASAP7_75t_L g5226 ( 
.A(n_5163),
.Y(n_5226)
);

BUFx3_ASAP7_75t_L g5227 ( 
.A(n_4948),
.Y(n_5227)
);

CKINVDCx5p33_ASAP7_75t_R g5228 ( 
.A(n_5050),
.Y(n_5228)
);

INVx2_ASAP7_75t_L g5229 ( 
.A(n_5185),
.Y(n_5229)
);

AND2x2_ASAP7_75t_L g5230 ( 
.A(n_5095),
.B(n_4820),
.Y(n_5230)
);

NAND2xp5_ASAP7_75t_L g5231 ( 
.A(n_4936),
.B(n_4827),
.Y(n_5231)
);

INVx4_ASAP7_75t_L g5232 ( 
.A(n_5013),
.Y(n_5232)
);

AND2x2_ASAP7_75t_L g5233 ( 
.A(n_5100),
.B(n_4827),
.Y(n_5233)
);

AND2x2_ASAP7_75t_L g5234 ( 
.A(n_5052),
.B(n_4827),
.Y(n_5234)
);

INVx6_ASAP7_75t_L g5235 ( 
.A(n_4976),
.Y(n_5235)
);

INVx1_ASAP7_75t_L g5236 ( 
.A(n_5000),
.Y(n_5236)
);

BUFx2_ASAP7_75t_R g5237 ( 
.A(n_5055),
.Y(n_5237)
);

INVx1_ASAP7_75t_L g5238 ( 
.A(n_5084),
.Y(n_5238)
);

OR2x2_ASAP7_75t_L g5239 ( 
.A(n_4955),
.B(n_4828),
.Y(n_5239)
);

AOI21xp5_ASAP7_75t_L g5240 ( 
.A1(n_5056),
.A2(n_4806),
.B(n_4779),
.Y(n_5240)
);

BUFx2_ASAP7_75t_L g5241 ( 
.A(n_5108),
.Y(n_5241)
);

INVx3_ASAP7_75t_L g5242 ( 
.A(n_5069),
.Y(n_5242)
);

INVxp67_ASAP7_75t_SL g5243 ( 
.A(n_4984),
.Y(n_5243)
);

NAND2xp5_ASAP7_75t_SL g5244 ( 
.A(n_5068),
.B(n_4881),
.Y(n_5244)
);

AOI22xp33_ASAP7_75t_L g5245 ( 
.A1(n_5139),
.A2(n_4745),
.B1(n_4765),
.B2(n_4714),
.Y(n_5245)
);

INVx1_ASAP7_75t_L g5246 ( 
.A(n_4933),
.Y(n_5246)
);

AOI21xp5_ASAP7_75t_L g5247 ( 
.A1(n_4959),
.A2(n_4806),
.B(n_4713),
.Y(n_5247)
);

NAND2xp5_ASAP7_75t_L g5248 ( 
.A(n_4938),
.B(n_4881),
.Y(n_5248)
);

INVx2_ASAP7_75t_L g5249 ( 
.A(n_4946),
.Y(n_5249)
);

NAND2x1p5_ASAP7_75t_L g5250 ( 
.A(n_4978),
.B(n_4745),
.Y(n_5250)
);

INVx3_ASAP7_75t_L g5251 ( 
.A(n_5069),
.Y(n_5251)
);

INVx3_ASAP7_75t_SL g5252 ( 
.A(n_4976),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_4950),
.B(n_4979),
.Y(n_5253)
);

INVx1_ASAP7_75t_L g5254 ( 
.A(n_4933),
.Y(n_5254)
);

AOI22xp33_ASAP7_75t_L g5255 ( 
.A1(n_5184),
.A2(n_4765),
.B1(n_4745),
.B2(n_2356),
.Y(n_5255)
);

INVx2_ASAP7_75t_L g5256 ( 
.A(n_4971),
.Y(n_5256)
);

INVx1_ASAP7_75t_L g5257 ( 
.A(n_5070),
.Y(n_5257)
);

A2O1A1Ixp33_ASAP7_75t_L g5258 ( 
.A1(n_5082),
.A2(n_5051),
.B(n_5054),
.C(n_5122),
.Y(n_5258)
);

BUFx6f_ASAP7_75t_L g5259 ( 
.A(n_4992),
.Y(n_5259)
);

INVx3_ASAP7_75t_L g5260 ( 
.A(n_5107),
.Y(n_5260)
);

AOI22xp5_ASAP7_75t_L g5261 ( 
.A1(n_5138),
.A2(n_4765),
.B1(n_4904),
.B2(n_4886),
.Y(n_5261)
);

INVx1_ASAP7_75t_SL g5262 ( 
.A(n_5061),
.Y(n_5262)
);

INVx5_ASAP7_75t_SL g5263 ( 
.A(n_4992),
.Y(n_5263)
);

AOI21xp5_ASAP7_75t_L g5264 ( 
.A1(n_5088),
.A2(n_4906),
.B(n_4724),
.Y(n_5264)
);

INVx1_ASAP7_75t_L g5265 ( 
.A(n_4958),
.Y(n_5265)
);

NOR2xp33_ASAP7_75t_L g5266 ( 
.A(n_5078),
.B(n_5068),
.Y(n_5266)
);

OAI21xp5_ASAP7_75t_L g5267 ( 
.A1(n_5146),
.A2(n_4772),
.B(n_4890),
.Y(n_5267)
);

NAND2xp5_ASAP7_75t_L g5268 ( 
.A(n_4944),
.B(n_4886),
.Y(n_5268)
);

INVx2_ASAP7_75t_SL g5269 ( 
.A(n_4960),
.Y(n_5269)
);

OA21x2_ASAP7_75t_L g5270 ( 
.A1(n_5165),
.A2(n_4712),
.B(n_1041),
.Y(n_5270)
);

NAND2xp5_ASAP7_75t_L g5271 ( 
.A(n_4947),
.B(n_4904),
.Y(n_5271)
);

AND2x4_ASAP7_75t_L g5272 ( 
.A(n_5123),
.B(n_4904),
.Y(n_5272)
);

AOI222xp33_ASAP7_75t_L g5273 ( 
.A1(n_5048),
.A2(n_1050),
.B1(n_1047),
.B2(n_1052),
.C1(n_1048),
.C2(n_1037),
.Y(n_5273)
);

AOI21xp5_ASAP7_75t_L g5274 ( 
.A1(n_5065),
.A2(n_4925),
.B(n_4918),
.Y(n_5274)
);

BUFx12f_ASAP7_75t_L g5275 ( 
.A(n_5079),
.Y(n_5275)
);

OAI22xp5_ASAP7_75t_L g5276 ( 
.A1(n_5059),
.A2(n_4925),
.B1(n_4918),
.B2(n_1067),
.Y(n_5276)
);

A2O1A1Ixp33_ASAP7_75t_L g5277 ( 
.A1(n_4972),
.A2(n_1074),
.B(n_1081),
.C(n_1062),
.Y(n_5277)
);

BUFx6f_ASAP7_75t_L g5278 ( 
.A(n_5049),
.Y(n_5278)
);

AND2x4_ASAP7_75t_L g5279 ( 
.A(n_5123),
.B(n_4918),
.Y(n_5279)
);

BUFx2_ASAP7_75t_L g5280 ( 
.A(n_5118),
.Y(n_5280)
);

AND2x4_ASAP7_75t_L g5281 ( 
.A(n_5031),
.B(n_4998),
.Y(n_5281)
);

AO32x1_ASAP7_75t_L g5282 ( 
.A1(n_5027),
.A2(n_4965),
.A3(n_4940),
.B1(n_4932),
.B2(n_4989),
.Y(n_5282)
);

HB1xp67_ASAP7_75t_L g5283 ( 
.A(n_4954),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4968),
.Y(n_5284)
);

OR2x6_ASAP7_75t_L g5285 ( 
.A(n_5080),
.B(n_4925),
.Y(n_5285)
);

INVx1_ASAP7_75t_SL g5286 ( 
.A(n_5143),
.Y(n_5286)
);

AOI22xp33_ASAP7_75t_SL g5287 ( 
.A1(n_5184),
.A2(n_1101),
.B1(n_1082),
.B2(n_1085),
.Y(n_5287)
);

NAND2x1_ASAP7_75t_L g5288 ( 
.A(n_5127),
.B(n_4755),
.Y(n_5288)
);

INVx2_ASAP7_75t_SL g5289 ( 
.A(n_5026),
.Y(n_5289)
);

A2O1A1Ixp33_ASAP7_75t_L g5290 ( 
.A1(n_5094),
.A2(n_1092),
.B(n_1095),
.C(n_1084),
.Y(n_5290)
);

INVx1_ASAP7_75t_SL g5291 ( 
.A(n_5073),
.Y(n_5291)
);

AND2x2_ASAP7_75t_L g5292 ( 
.A(n_5104),
.B(n_19),
.Y(n_5292)
);

CKINVDCx20_ASAP7_75t_R g5293 ( 
.A(n_5011),
.Y(n_5293)
);

HB1xp67_ASAP7_75t_L g5294 ( 
.A(n_4931),
.Y(n_5294)
);

INVx3_ASAP7_75t_SL g5295 ( 
.A(n_5132),
.Y(n_5295)
);

OAI21xp5_ASAP7_75t_L g5296 ( 
.A1(n_5012),
.A2(n_1098),
.B(n_1096),
.Y(n_5296)
);

NOR2xp33_ASAP7_75t_L g5297 ( 
.A(n_5009),
.B(n_60),
.Y(n_5297)
);

OR2x6_ASAP7_75t_L g5298 ( 
.A(n_5004),
.B(n_5074),
.Y(n_5298)
);

NAND2xp5_ASAP7_75t_SL g5299 ( 
.A(n_4999),
.B(n_1225),
.Y(n_5299)
);

INVx2_ASAP7_75t_SL g5300 ( 
.A(n_5011),
.Y(n_5300)
);

INVx3_ASAP7_75t_L g5301 ( 
.A(n_5136),
.Y(n_5301)
);

AOI21xp5_ASAP7_75t_L g5302 ( 
.A1(n_4957),
.A2(n_4983),
.B(n_4993),
.Y(n_5302)
);

BUFx2_ASAP7_75t_L g5303 ( 
.A(n_5148),
.Y(n_5303)
);

OAI22xp5_ASAP7_75t_L g5304 ( 
.A1(n_5045),
.A2(n_1105),
.B1(n_1108),
.B2(n_1100),
.Y(n_5304)
);

BUFx3_ASAP7_75t_L g5305 ( 
.A(n_5043),
.Y(n_5305)
);

INVx6_ASAP7_75t_L g5306 ( 
.A(n_5189),
.Y(n_5306)
);

OR2x6_ASAP7_75t_L g5307 ( 
.A(n_5074),
.B(n_2978),
.Y(n_5307)
);

AND2x2_ASAP7_75t_L g5308 ( 
.A(n_5044),
.B(n_20),
.Y(n_5308)
);

A2O1A1Ixp33_ASAP7_75t_L g5309 ( 
.A1(n_5190),
.A2(n_1110),
.B(n_2070),
.C(n_2069),
.Y(n_5309)
);

BUFx6f_ASAP7_75t_L g5310 ( 
.A(n_5049),
.Y(n_5310)
);

AOI21xp5_ASAP7_75t_L g5311 ( 
.A1(n_5039),
.A2(n_2836),
.B(n_2828),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_4939),
.B(n_22),
.Y(n_5312)
);

NAND2x1_ASAP7_75t_L g5313 ( 
.A(n_5136),
.B(n_3446),
.Y(n_5313)
);

AND2x4_ASAP7_75t_L g5314 ( 
.A(n_5003),
.B(n_5010),
.Y(n_5314)
);

NAND2x1p5_ASAP7_75t_L g5315 ( 
.A(n_4978),
.B(n_2821),
.Y(n_5315)
);

INVx4_ASAP7_75t_L g5316 ( 
.A(n_5027),
.Y(n_5316)
);

O2A1O1Ixp33_ASAP7_75t_L g5317 ( 
.A1(n_5090),
.A2(n_2079),
.B(n_2083),
.C(n_2072),
.Y(n_5317)
);

NOR2xp67_ASAP7_75t_SL g5318 ( 
.A(n_4994),
.B(n_2391),
.Y(n_5318)
);

AND2x2_ASAP7_75t_L g5319 ( 
.A(n_5023),
.B(n_23),
.Y(n_5319)
);

OR2x2_ASAP7_75t_L g5320 ( 
.A(n_4975),
.B(n_4982),
.Y(n_5320)
);

BUFx6f_ASAP7_75t_L g5321 ( 
.A(n_5049),
.Y(n_5321)
);

NOR2xp33_ASAP7_75t_L g5322 ( 
.A(n_5016),
.B(n_61),
.Y(n_5322)
);

INVx3_ASAP7_75t_L g5323 ( 
.A(n_4985),
.Y(n_5323)
);

AND2x4_ASAP7_75t_L g5324 ( 
.A(n_5003),
.B(n_24),
.Y(n_5324)
);

INVx3_ASAP7_75t_L g5325 ( 
.A(n_5187),
.Y(n_5325)
);

O2A1O1Ixp33_ASAP7_75t_L g5326 ( 
.A1(n_4966),
.A2(n_2085),
.B(n_2095),
.C(n_2079),
.Y(n_5326)
);

INVx2_ASAP7_75t_SL g5327 ( 
.A(n_5015),
.Y(n_5327)
);

OAI21xp5_ASAP7_75t_L g5328 ( 
.A1(n_5192),
.A2(n_4942),
.B(n_5067),
.Y(n_5328)
);

A2O1A1Ixp33_ASAP7_75t_L g5329 ( 
.A1(n_4945),
.A2(n_2105),
.B(n_2104),
.C(n_2140),
.Y(n_5329)
);

O2A1O1Ixp33_ASAP7_75t_L g5330 ( 
.A1(n_5115),
.A2(n_2105),
.B(n_2104),
.C(n_26),
.Y(n_5330)
);

BUFx6f_ASAP7_75t_L g5331 ( 
.A(n_5064),
.Y(n_5331)
);

AOI21xp5_ASAP7_75t_L g5332 ( 
.A1(n_5142),
.A2(n_2299),
.B(n_2391),
.Y(n_5332)
);

INVx1_ASAP7_75t_SL g5333 ( 
.A(n_5157),
.Y(n_5333)
);

AOI21xp5_ASAP7_75t_L g5334 ( 
.A1(n_5145),
.A2(n_2299),
.B(n_2391),
.Y(n_5334)
);

INVx5_ASAP7_75t_L g5335 ( 
.A(n_5020),
.Y(n_5335)
);

AND2x4_ASAP7_75t_L g5336 ( 
.A(n_5010),
.B(n_24),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_SL g5337 ( 
.A(n_5161),
.B(n_1225),
.Y(n_5337)
);

AND2x2_ASAP7_75t_L g5338 ( 
.A(n_5081),
.B(n_25),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_L g5339 ( 
.A(n_4984),
.B(n_25),
.Y(n_5339)
);

OAI21xp5_ASAP7_75t_L g5340 ( 
.A1(n_5128),
.A2(n_2052),
.B(n_2015),
.Y(n_5340)
);

INVx2_ASAP7_75t_L g5341 ( 
.A(n_4977),
.Y(n_5341)
);

AND2x6_ASAP7_75t_L g5342 ( 
.A(n_4935),
.B(n_2821),
.Y(n_5342)
);

NOR2xp33_ASAP7_75t_L g5343 ( 
.A(n_5014),
.B(n_61),
.Y(n_5343)
);

OAI22xp5_ASAP7_75t_L g5344 ( 
.A1(n_5174),
.A2(n_2795),
.B1(n_2810),
.B2(n_2173),
.Y(n_5344)
);

A2O1A1Ixp33_ASAP7_75t_L g5345 ( 
.A1(n_5137),
.A2(n_30),
.B(n_26),
.C(n_29),
.Y(n_5345)
);

NAND2xp33_ASAP7_75t_L g5346 ( 
.A(n_5064),
.B(n_1240),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_5007),
.Y(n_5347)
);

AOI21xp5_ASAP7_75t_L g5348 ( 
.A1(n_5017),
.A2(n_2408),
.B(n_2402),
.Y(n_5348)
);

AOI22xp33_ASAP7_75t_L g5349 ( 
.A1(n_5131),
.A2(n_2356),
.B1(n_2341),
.B2(n_2149),
.Y(n_5349)
);

INVx1_ASAP7_75t_SL g5350 ( 
.A(n_5097),
.Y(n_5350)
);

AND2x4_ASAP7_75t_L g5351 ( 
.A(n_4963),
.B(n_29),
.Y(n_5351)
);

NAND2x1p5_ASAP7_75t_L g5352 ( 
.A(n_5186),
.B(n_2821),
.Y(n_5352)
);

AOI21xp5_ASAP7_75t_L g5353 ( 
.A1(n_5022),
.A2(n_2408),
.B(n_2402),
.Y(n_5353)
);

OR2x6_ASAP7_75t_SL g5354 ( 
.A(n_5091),
.B(n_29),
.Y(n_5354)
);

NOR2xp33_ASAP7_75t_L g5355 ( 
.A(n_5135),
.B(n_62),
.Y(n_5355)
);

INVx5_ASAP7_75t_L g5356 ( 
.A(n_5020),
.Y(n_5356)
);

OAI22xp5_ASAP7_75t_L g5357 ( 
.A1(n_4973),
.A2(n_4996),
.B1(n_5072),
.B2(n_5112),
.Y(n_5357)
);

BUFx6f_ASAP7_75t_L g5358 ( 
.A(n_5064),
.Y(n_5358)
);

NOR2xp33_ASAP7_75t_L g5359 ( 
.A(n_5144),
.B(n_62),
.Y(n_5359)
);

BUFx3_ASAP7_75t_L g5360 ( 
.A(n_5125),
.Y(n_5360)
);

INVx1_ASAP7_75t_L g5361 ( 
.A(n_4986),
.Y(n_5361)
);

OAI22xp5_ASAP7_75t_L g5362 ( 
.A1(n_4981),
.A2(n_2810),
.B1(n_2795),
.B2(n_2113),
.Y(n_5362)
);

AOI22xp33_ASAP7_75t_L g5363 ( 
.A1(n_5083),
.A2(n_5164),
.B1(n_5086),
.B2(n_5116),
.Y(n_5363)
);

AOI21xp5_ASAP7_75t_L g5364 ( 
.A1(n_5036),
.A2(n_2408),
.B(n_2402),
.Y(n_5364)
);

AND2x2_ASAP7_75t_L g5365 ( 
.A(n_5019),
.B(n_30),
.Y(n_5365)
);

INVx2_ASAP7_75t_L g5366 ( 
.A(n_4991),
.Y(n_5366)
);

AOI21x1_ASAP7_75t_L g5367 ( 
.A1(n_5092),
.A2(n_2488),
.B(n_2592),
.Y(n_5367)
);

BUFx2_ASAP7_75t_L g5368 ( 
.A(n_5153),
.Y(n_5368)
);

AND2x4_ASAP7_75t_L g5369 ( 
.A(n_4963),
.B(n_30),
.Y(n_5369)
);

AND2x4_ASAP7_75t_L g5370 ( 
.A(n_4963),
.B(n_31),
.Y(n_5370)
);

NAND2xp5_ASAP7_75t_L g5371 ( 
.A(n_4962),
.B(n_31),
.Y(n_5371)
);

BUFx6f_ASAP7_75t_L g5372 ( 
.A(n_5197),
.Y(n_5372)
);

AND2x4_ASAP7_75t_L g5373 ( 
.A(n_4963),
.B(n_32),
.Y(n_5373)
);

OAI22xp5_ASAP7_75t_L g5374 ( 
.A1(n_4951),
.A2(n_2810),
.B1(n_2795),
.B2(n_2113),
.Y(n_5374)
);

BUFx8_ASAP7_75t_L g5375 ( 
.A(n_5197),
.Y(n_5375)
);

NAND2xp5_ASAP7_75t_L g5376 ( 
.A(n_4969),
.B(n_32),
.Y(n_5376)
);

NAND2x1_ASAP7_75t_L g5377 ( 
.A(n_5187),
.B(n_1296),
.Y(n_5377)
);

OAI21x1_ASAP7_75t_L g5378 ( 
.A1(n_5021),
.A2(n_3121),
.B(n_2535),
.Y(n_5378)
);

OAI21xp33_ASAP7_75t_L g5379 ( 
.A1(n_5062),
.A2(n_1299),
.B(n_1296),
.Y(n_5379)
);

NAND2xp5_ASAP7_75t_L g5380 ( 
.A(n_5063),
.B(n_33),
.Y(n_5380)
);

INVx3_ASAP7_75t_L g5381 ( 
.A(n_5085),
.Y(n_5381)
);

INVx4_ASAP7_75t_L g5382 ( 
.A(n_5197),
.Y(n_5382)
);

A2O1A1Ixp33_ASAP7_75t_L g5383 ( 
.A1(n_5006),
.A2(n_33),
.B(n_34),
.C(n_1544),
.Y(n_5383)
);

AOI21xp5_ASAP7_75t_L g5384 ( 
.A1(n_5037),
.A2(n_2408),
.B(n_2402),
.Y(n_5384)
);

INVx3_ASAP7_75t_SL g5385 ( 
.A(n_5002),
.Y(n_5385)
);

AND2x2_ASAP7_75t_L g5386 ( 
.A(n_5024),
.B(n_33),
.Y(n_5386)
);

AND2x2_ASAP7_75t_L g5387 ( 
.A(n_5030),
.B(n_34),
.Y(n_5387)
);

OAI22xp5_ASAP7_75t_L g5388 ( 
.A1(n_5093),
.A2(n_2112),
.B1(n_2129),
.B2(n_2113),
.Y(n_5388)
);

O2A1O1Ixp5_ASAP7_75t_SL g5389 ( 
.A1(n_5110),
.A2(n_2129),
.B(n_2112),
.C(n_1992),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_4988),
.B(n_4990),
.Y(n_5390)
);

OR2x6_ASAP7_75t_L g5391 ( 
.A(n_5035),
.B(n_1299),
.Y(n_5391)
);

INVx1_ASAP7_75t_L g5392 ( 
.A(n_4990),
.Y(n_5392)
);

AND2x2_ASAP7_75t_L g5393 ( 
.A(n_5133),
.B(n_63),
.Y(n_5393)
);

HB1xp67_ASAP7_75t_L g5394 ( 
.A(n_5005),
.Y(n_5394)
);

INVx2_ASAP7_75t_SL g5395 ( 
.A(n_5133),
.Y(n_5395)
);

NOR2xp33_ASAP7_75t_L g5396 ( 
.A(n_5156),
.B(n_63),
.Y(n_5396)
);

INVx3_ASAP7_75t_L g5397 ( 
.A(n_5040),
.Y(n_5397)
);

CKINVDCx5p33_ASAP7_75t_R g5398 ( 
.A(n_4997),
.Y(n_5398)
);

HB1xp67_ASAP7_75t_L g5399 ( 
.A(n_5005),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_5141),
.Y(n_5400)
);

BUFx6f_ASAP7_75t_L g5401 ( 
.A(n_5034),
.Y(n_5401)
);

INVx2_ASAP7_75t_L g5402 ( 
.A(n_5176),
.Y(n_5402)
);

NOR2xp33_ASAP7_75t_L g5403 ( 
.A(n_5159),
.B(n_64),
.Y(n_5403)
);

HB1xp67_ASAP7_75t_L g5404 ( 
.A(n_5114),
.Y(n_5404)
);

BUFx6f_ASAP7_75t_L g5405 ( 
.A(n_4949),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5183),
.Y(n_5406)
);

NOR2xp33_ASAP7_75t_SL g5407 ( 
.A(n_5172),
.B(n_2927),
.Y(n_5407)
);

AOI21xp5_ASAP7_75t_L g5408 ( 
.A1(n_5089),
.A2(n_2447),
.B(n_2433),
.Y(n_5408)
);

AOI22xp5_ASAP7_75t_L g5409 ( 
.A1(n_5357),
.A2(n_5033),
.B1(n_5121),
.B2(n_5001),
.Y(n_5409)
);

AOI22xp33_ASAP7_75t_L g5410 ( 
.A1(n_5312),
.A2(n_5154),
.B1(n_5033),
.B2(n_5162),
.Y(n_5410)
);

CKINVDCx20_ASAP7_75t_R g5411 ( 
.A(n_5213),
.Y(n_5411)
);

INVx3_ASAP7_75t_L g5412 ( 
.A(n_5288),
.Y(n_5412)
);

INVx2_ASAP7_75t_L g5413 ( 
.A(n_5239),
.Y(n_5413)
);

INVx6_ASAP7_75t_L g5414 ( 
.A(n_5375),
.Y(n_5414)
);

OAI22xp33_ASAP7_75t_L g5415 ( 
.A1(n_5398),
.A2(n_5224),
.B1(n_5339),
.B2(n_5298),
.Y(n_5415)
);

INVx6_ASAP7_75t_L g5416 ( 
.A(n_5232),
.Y(n_5416)
);

OAI21xp33_ASAP7_75t_L g5417 ( 
.A1(n_5243),
.A2(n_5171),
.B(n_5087),
.Y(n_5417)
);

OAI22xp33_ASAP7_75t_L g5418 ( 
.A1(n_5224),
.A2(n_5298),
.B1(n_5240),
.B2(n_5407),
.Y(n_5418)
);

INVx4_ASAP7_75t_L g5419 ( 
.A(n_5232),
.Y(n_5419)
);

AOI22xp33_ASAP7_75t_L g5420 ( 
.A1(n_5328),
.A2(n_5047),
.B1(n_5149),
.B2(n_4956),
.Y(n_5420)
);

AOI22xp5_ASAP7_75t_L g5421 ( 
.A1(n_5362),
.A2(n_5342),
.B1(n_5359),
.B2(n_5355),
.Y(n_5421)
);

INVx2_ASAP7_75t_L g5422 ( 
.A(n_5209),
.Y(n_5422)
);

AOI22xp33_ASAP7_75t_L g5423 ( 
.A1(n_5207),
.A2(n_5008),
.B1(n_5152),
.B2(n_5032),
.Y(n_5423)
);

CKINVDCx6p67_ASAP7_75t_R g5424 ( 
.A(n_5293),
.Y(n_5424)
);

BUFx4f_ASAP7_75t_L g5425 ( 
.A(n_5259),
.Y(n_5425)
);

BUFx8_ASAP7_75t_L g5426 ( 
.A(n_5259),
.Y(n_5426)
);

INVx6_ASAP7_75t_L g5427 ( 
.A(n_5259),
.Y(n_5427)
);

AOI22xp33_ASAP7_75t_L g5428 ( 
.A1(n_5270),
.A2(n_5222),
.B1(n_5255),
.B2(n_5287),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_5236),
.Y(n_5429)
);

INVx4_ASAP7_75t_L g5430 ( 
.A(n_5203),
.Y(n_5430)
);

INVx8_ASAP7_75t_L g5431 ( 
.A(n_5275),
.Y(n_5431)
);

CKINVDCx5p33_ASAP7_75t_R g5432 ( 
.A(n_5205),
.Y(n_5432)
);

NAND2x1p5_ASAP7_75t_L g5433 ( 
.A(n_5351),
.B(n_4953),
.Y(n_5433)
);

CKINVDCx5p33_ASAP7_75t_R g5434 ( 
.A(n_5228),
.Y(n_5434)
);

CKINVDCx11_ASAP7_75t_R g5435 ( 
.A(n_5252),
.Y(n_5435)
);

AOI22xp33_ASAP7_75t_L g5436 ( 
.A1(n_5396),
.A2(n_5169),
.B1(n_5042),
.B2(n_5195),
.Y(n_5436)
);

INVx2_ASAP7_75t_L g5437 ( 
.A(n_5405),
.Y(n_5437)
);

NAND2xp5_ASAP7_75t_L g5438 ( 
.A(n_5283),
.B(n_4967),
.Y(n_5438)
);

INVx1_ASAP7_75t_L g5439 ( 
.A(n_5238),
.Y(n_5439)
);

INVx6_ASAP7_75t_L g5440 ( 
.A(n_5324),
.Y(n_5440)
);

AOI22xp5_ASAP7_75t_L g5441 ( 
.A1(n_5342),
.A2(n_5403),
.B1(n_5299),
.B2(n_5217),
.Y(n_5441)
);

BUFx10_ASAP7_75t_L g5442 ( 
.A(n_5343),
.Y(n_5442)
);

BUFx10_ASAP7_75t_L g5443 ( 
.A(n_5235),
.Y(n_5443)
);

INVx1_ASAP7_75t_SL g5444 ( 
.A(n_5237),
.Y(n_5444)
);

INVx3_ASAP7_75t_L g5445 ( 
.A(n_5281),
.Y(n_5445)
);

INVx1_ASAP7_75t_SL g5446 ( 
.A(n_5206),
.Y(n_5446)
);

NAND2xp5_ASAP7_75t_L g5447 ( 
.A(n_5199),
.B(n_4967),
.Y(n_5447)
);

AND2x2_ASAP7_75t_L g5448 ( 
.A(n_5281),
.B(n_5178),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_5257),
.B(n_4967),
.Y(n_5449)
);

INVx1_ASAP7_75t_SL g5450 ( 
.A(n_5262),
.Y(n_5450)
);

AOI22xp33_ASAP7_75t_L g5451 ( 
.A1(n_5390),
.A2(n_5169),
.B1(n_5140),
.B2(n_5025),
.Y(n_5451)
);

OAI22xp5_ASAP7_75t_L g5452 ( 
.A1(n_5302),
.A2(n_5053),
.B1(n_5193),
.B2(n_5077),
.Y(n_5452)
);

BUFx3_ASAP7_75t_L g5453 ( 
.A(n_5227),
.Y(n_5453)
);

BUFx2_ASAP7_75t_SL g5454 ( 
.A(n_5300),
.Y(n_5454)
);

AOI22xp33_ASAP7_75t_L g5455 ( 
.A1(n_5401),
.A2(n_5196),
.B1(n_5129),
.B2(n_5119),
.Y(n_5455)
);

CKINVDCx11_ASAP7_75t_R g5456 ( 
.A(n_5354),
.Y(n_5456)
);

NAND2x1p5_ASAP7_75t_L g5457 ( 
.A(n_5351),
.B(n_5071),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_5246),
.Y(n_5458)
);

INVx6_ASAP7_75t_L g5459 ( 
.A(n_5324),
.Y(n_5459)
);

INVx1_ASAP7_75t_SL g5460 ( 
.A(n_5333),
.Y(n_5460)
);

INVx2_ASAP7_75t_L g5461 ( 
.A(n_5229),
.Y(n_5461)
);

OAI22xp33_ASAP7_75t_L g5462 ( 
.A1(n_5391),
.A2(n_5058),
.B1(n_5109),
.B2(n_5096),
.Y(n_5462)
);

INVx6_ASAP7_75t_L g5463 ( 
.A(n_5336),
.Y(n_5463)
);

AND2x4_ASAP7_75t_L g5464 ( 
.A(n_5323),
.B(n_5102),
.Y(n_5464)
);

INVx1_ASAP7_75t_L g5465 ( 
.A(n_5254),
.Y(n_5465)
);

AOI22xp33_ASAP7_75t_SL g5466 ( 
.A1(n_5226),
.A2(n_5075),
.B1(n_5120),
.B2(n_5103),
.Y(n_5466)
);

OAI22xp5_ASAP7_75t_L g5467 ( 
.A1(n_5258),
.A2(n_5181),
.B1(n_5182),
.B2(n_5066),
.Y(n_5467)
);

INVx1_ASAP7_75t_SL g5468 ( 
.A(n_5295),
.Y(n_5468)
);

BUFx12f_ASAP7_75t_L g5469 ( 
.A(n_5306),
.Y(n_5469)
);

AOI22xp33_ASAP7_75t_L g5470 ( 
.A1(n_5342),
.A2(n_5117),
.B1(n_5098),
.B2(n_5126),
.Y(n_5470)
);

BUFx6f_ASAP7_75t_L g5471 ( 
.A(n_5377),
.Y(n_5471)
);

BUFx6f_ASAP7_75t_L g5472 ( 
.A(n_5278),
.Y(n_5472)
);

INVx1_ASAP7_75t_L g5473 ( 
.A(n_5212),
.Y(n_5473)
);

INVx6_ASAP7_75t_L g5474 ( 
.A(n_5336),
.Y(n_5474)
);

INVx1_ASAP7_75t_SL g5475 ( 
.A(n_5286),
.Y(n_5475)
);

INVx1_ASAP7_75t_L g5476 ( 
.A(n_5265),
.Y(n_5476)
);

AOI22xp33_ASAP7_75t_L g5477 ( 
.A1(n_5273),
.A2(n_5124),
.B1(n_5170),
.B2(n_5155),
.Y(n_5477)
);

BUFx8_ASAP7_75t_L g5478 ( 
.A(n_5292),
.Y(n_5478)
);

CKINVDCx20_ASAP7_75t_R g5479 ( 
.A(n_5263),
.Y(n_5479)
);

AOI22xp33_ASAP7_75t_SL g5480 ( 
.A1(n_5404),
.A2(n_5151),
.B1(n_5177),
.B2(n_5134),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_5284),
.Y(n_5481)
);

OAI22xp5_ASAP7_75t_L g5482 ( 
.A1(n_5198),
.A2(n_5168),
.B1(n_5188),
.B2(n_5150),
.Y(n_5482)
);

INVx6_ASAP7_75t_L g5483 ( 
.A(n_5306),
.Y(n_5483)
);

BUFx8_ASAP7_75t_L g5484 ( 
.A(n_5393),
.Y(n_5484)
);

AOI22xp5_ASAP7_75t_SL g5485 ( 
.A1(n_5266),
.A2(n_5194),
.B1(n_5191),
.B2(n_5166),
.Y(n_5485)
);

OAI21xp33_ASAP7_75t_L g5486 ( 
.A1(n_5345),
.A2(n_5076),
.B(n_5130),
.Y(n_5486)
);

INVx6_ASAP7_75t_L g5487 ( 
.A(n_5369),
.Y(n_5487)
);

INVx2_ASAP7_75t_L g5488 ( 
.A(n_5249),
.Y(n_5488)
);

BUFx2_ASAP7_75t_L g5489 ( 
.A(n_5314),
.Y(n_5489)
);

INVx5_ASAP7_75t_L g5490 ( 
.A(n_5285),
.Y(n_5490)
);

CKINVDCx6p67_ASAP7_75t_R g5491 ( 
.A(n_5385),
.Y(n_5491)
);

INVx2_ASAP7_75t_L g5492 ( 
.A(n_5256),
.Y(n_5492)
);

INVx2_ASAP7_75t_L g5493 ( 
.A(n_5341),
.Y(n_5493)
);

NAND2xp5_ASAP7_75t_L g5494 ( 
.A(n_5253),
.B(n_5294),
.Y(n_5494)
);

INVx2_ASAP7_75t_SL g5495 ( 
.A(n_5305),
.Y(n_5495)
);

INVx2_ASAP7_75t_SL g5496 ( 
.A(n_5230),
.Y(n_5496)
);

INVxp67_ASAP7_75t_L g5497 ( 
.A(n_5200),
.Y(n_5497)
);

BUFx10_ASAP7_75t_L g5498 ( 
.A(n_5297),
.Y(n_5498)
);

BUFx2_ASAP7_75t_SL g5499 ( 
.A(n_5269),
.Y(n_5499)
);

BUFx8_ASAP7_75t_L g5500 ( 
.A(n_5386),
.Y(n_5500)
);

INVx4_ASAP7_75t_L g5501 ( 
.A(n_5316),
.Y(n_5501)
);

BUFx10_ASAP7_75t_L g5502 ( 
.A(n_5322),
.Y(n_5502)
);

INVx3_ASAP7_75t_L g5503 ( 
.A(n_5316),
.Y(n_5503)
);

INVx2_ASAP7_75t_L g5504 ( 
.A(n_5366),
.Y(n_5504)
);

OAI22xp5_ASAP7_75t_L g5505 ( 
.A1(n_5369),
.A2(n_5029),
.B1(n_5057),
.B2(n_2129),
.Y(n_5505)
);

HB1xp67_ASAP7_75t_L g5506 ( 
.A(n_5223),
.Y(n_5506)
);

CKINVDCx20_ASAP7_75t_R g5507 ( 
.A(n_5360),
.Y(n_5507)
);

BUFx6f_ASAP7_75t_L g5508 ( 
.A(n_5278),
.Y(n_5508)
);

BUFx6f_ASAP7_75t_L g5509 ( 
.A(n_5278),
.Y(n_5509)
);

AOI22xp33_ASAP7_75t_SL g5510 ( 
.A1(n_5370),
.A2(n_5180),
.B1(n_5179),
.B2(n_2052),
.Y(n_5510)
);

OAI21xp5_ASAP7_75t_SL g5511 ( 
.A1(n_5309),
.A2(n_65),
.B(n_66),
.Y(n_5511)
);

INVx1_ASAP7_75t_SL g5512 ( 
.A(n_5291),
.Y(n_5512)
);

INVx3_ASAP7_75t_L g5513 ( 
.A(n_5325),
.Y(n_5513)
);

OAI21xp33_ASAP7_75t_L g5514 ( 
.A1(n_5277),
.A2(n_1553),
.B(n_1303),
.Y(n_5514)
);

AOI22xp33_ASAP7_75t_L g5515 ( 
.A1(n_5304),
.A2(n_2154),
.B1(n_2157),
.B2(n_2150),
.Y(n_5515)
);

BUFx12f_ASAP7_75t_L g5516 ( 
.A(n_5308),
.Y(n_5516)
);

AOI22xp33_ASAP7_75t_L g5517 ( 
.A1(n_5347),
.A2(n_2154),
.B1(n_2157),
.B2(n_2150),
.Y(n_5517)
);

OR2x2_ASAP7_75t_L g5518 ( 
.A(n_5320),
.B(n_5057),
.Y(n_5518)
);

BUFx6f_ASAP7_75t_L g5519 ( 
.A(n_5310),
.Y(n_5519)
);

AOI22xp33_ASAP7_75t_L g5520 ( 
.A1(n_5267),
.A2(n_2157),
.B1(n_2170),
.B2(n_2154),
.Y(n_5520)
);

CKINVDCx6p67_ASAP7_75t_R g5521 ( 
.A(n_5387),
.Y(n_5521)
);

BUFx10_ASAP7_75t_L g5522 ( 
.A(n_5370),
.Y(n_5522)
);

AND2x2_ASAP7_75t_L g5523 ( 
.A(n_5204),
.B(n_5029),
.Y(n_5523)
);

INVx2_ASAP7_75t_L g5524 ( 
.A(n_5400),
.Y(n_5524)
);

CKINVDCx11_ASAP7_75t_R g5525 ( 
.A(n_5368),
.Y(n_5525)
);

AOI22xp5_ASAP7_75t_L g5526 ( 
.A1(n_5219),
.A2(n_2052),
.B1(n_2058),
.B2(n_2015),
.Y(n_5526)
);

AOI22xp5_ASAP7_75t_L g5527 ( 
.A1(n_5373),
.A2(n_2058),
.B1(n_2075),
.B2(n_2052),
.Y(n_5527)
);

INVx6_ASAP7_75t_L g5528 ( 
.A(n_5335),
.Y(n_5528)
);

CKINVDCx6p67_ASAP7_75t_R g5529 ( 
.A(n_5380),
.Y(n_5529)
);

BUFx2_ASAP7_75t_L g5530 ( 
.A(n_5314),
.Y(n_5530)
);

BUFx2_ASAP7_75t_L g5531 ( 
.A(n_5280),
.Y(n_5531)
);

AND2x2_ASAP7_75t_L g5532 ( 
.A(n_5208),
.B(n_5105),
.Y(n_5532)
);

OAI22xp5_ASAP7_75t_L g5533 ( 
.A1(n_5214),
.A2(n_2736),
.B1(n_2775),
.B2(n_2732),
.Y(n_5533)
);

INVx2_ASAP7_75t_L g5534 ( 
.A(n_5402),
.Y(n_5534)
);

AOI22xp5_ASAP7_75t_L g5535 ( 
.A1(n_5245),
.A2(n_5350),
.B1(n_5371),
.B2(n_5376),
.Y(n_5535)
);

INVx6_ASAP7_75t_L g5536 ( 
.A(n_5335),
.Y(n_5536)
);

INVx6_ASAP7_75t_L g5537 ( 
.A(n_5335),
.Y(n_5537)
);

INVx2_ASAP7_75t_L g5538 ( 
.A(n_5394),
.Y(n_5538)
);

NAND2x1p5_ASAP7_75t_L g5539 ( 
.A(n_5356),
.B(n_2844),
.Y(n_5539)
);

AOI22xp33_ASAP7_75t_L g5540 ( 
.A1(n_5201),
.A2(n_2170),
.B1(n_2191),
.B2(n_2157),
.Y(n_5540)
);

OAI22xp33_ASAP7_75t_L g5541 ( 
.A1(n_5307),
.A2(n_2851),
.B1(n_2844),
.B2(n_2941),
.Y(n_5541)
);

INVx2_ASAP7_75t_L g5542 ( 
.A(n_5399),
.Y(n_5542)
);

AOI22xp33_ASAP7_75t_L g5543 ( 
.A1(n_5296),
.A2(n_5361),
.B1(n_5327),
.B2(n_5340),
.Y(n_5543)
);

INVx6_ASAP7_75t_L g5544 ( 
.A(n_5356),
.Y(n_5544)
);

INVx1_ASAP7_75t_L g5545 ( 
.A(n_5392),
.Y(n_5545)
);

OAI22xp5_ASAP7_75t_L g5546 ( 
.A1(n_5363),
.A2(n_5247),
.B1(n_5225),
.B2(n_5289),
.Y(n_5546)
);

HB1xp67_ASAP7_75t_L g5547 ( 
.A(n_5241),
.Y(n_5547)
);

AOI22xp33_ASAP7_75t_SL g5548 ( 
.A1(n_5282),
.A2(n_5365),
.B1(n_5338),
.B2(n_5319),
.Y(n_5548)
);

AOI22xp33_ASAP7_75t_L g5549 ( 
.A1(n_5406),
.A2(n_2191),
.B1(n_2193),
.B2(n_2170),
.Y(n_5549)
);

INVx2_ASAP7_75t_L g5550 ( 
.A(n_5397),
.Y(n_5550)
);

INVx6_ASAP7_75t_L g5551 ( 
.A(n_5356),
.Y(n_5551)
);

NAND2xp5_ASAP7_75t_SL g5552 ( 
.A(n_5303),
.B(n_1299),
.Y(n_5552)
);

AOI22xp33_ASAP7_75t_L g5553 ( 
.A1(n_5216),
.A2(n_2191),
.B1(n_2193),
.B2(n_2170),
.Y(n_5553)
);

BUFx3_ASAP7_75t_L g5554 ( 
.A(n_5233),
.Y(n_5554)
);

CKINVDCx20_ASAP7_75t_R g5555 ( 
.A(n_5244),
.Y(n_5555)
);

INVx1_ASAP7_75t_L g5556 ( 
.A(n_5231),
.Y(n_5556)
);

BUFx6f_ASAP7_75t_L g5557 ( 
.A(n_5310),
.Y(n_5557)
);

AOI22xp33_ASAP7_75t_L g5558 ( 
.A1(n_5211),
.A2(n_2224),
.B1(n_2229),
.B2(n_2193),
.Y(n_5558)
);

BUFx4f_ASAP7_75t_SL g5559 ( 
.A(n_5234),
.Y(n_5559)
);

AOI22xp33_ASAP7_75t_L g5560 ( 
.A1(n_5337),
.A2(n_2229),
.B1(n_2234),
.B2(n_2224),
.Y(n_5560)
);

BUFx4f_ASAP7_75t_SL g5561 ( 
.A(n_5310),
.Y(n_5561)
);

INVx1_ASAP7_75t_L g5562 ( 
.A(n_5248),
.Y(n_5562)
);

CKINVDCx6p67_ASAP7_75t_R g5563 ( 
.A(n_5321),
.Y(n_5563)
);

INVxp67_ASAP7_75t_L g5564 ( 
.A(n_5318),
.Y(n_5564)
);

INVx1_ASAP7_75t_SL g5565 ( 
.A(n_5268),
.Y(n_5565)
);

AOI22xp33_ASAP7_75t_L g5566 ( 
.A1(n_5349),
.A2(n_5388),
.B1(n_5374),
.B2(n_5379),
.Y(n_5566)
);

AND2x2_ASAP7_75t_L g5567 ( 
.A(n_5202),
.B(n_5105),
.Y(n_5567)
);

OAI22xp5_ASAP7_75t_L g5568 ( 
.A1(n_5261),
.A2(n_2736),
.B1(n_2775),
.B2(n_2732),
.Y(n_5568)
);

INVx2_ASAP7_75t_L g5569 ( 
.A(n_5221),
.Y(n_5569)
);

INVx1_ASAP7_75t_L g5570 ( 
.A(n_5271),
.Y(n_5570)
);

CKINVDCx6p67_ASAP7_75t_R g5571 ( 
.A(n_5321),
.Y(n_5571)
);

BUFx12f_ASAP7_75t_L g5572 ( 
.A(n_5321),
.Y(n_5572)
);

OAI22xp33_ASAP7_75t_L g5573 ( 
.A1(n_5220),
.A2(n_2851),
.B1(n_2844),
.B2(n_2941),
.Y(n_5573)
);

AOI22xp33_ASAP7_75t_SL g5574 ( 
.A1(n_5282),
.A2(n_2075),
.B1(n_2094),
.B2(n_2058),
.Y(n_5574)
);

CKINVDCx5p33_ASAP7_75t_R g5575 ( 
.A(n_5395),
.Y(n_5575)
);

INVx2_ASAP7_75t_L g5576 ( 
.A(n_5378),
.Y(n_5576)
);

CKINVDCx11_ASAP7_75t_R g5577 ( 
.A(n_5331),
.Y(n_5577)
);

AOI22xp33_ASAP7_75t_L g5578 ( 
.A1(n_5344),
.A2(n_2229),
.B1(n_2234),
.B2(n_2224),
.Y(n_5578)
);

OAI22xp33_ASAP7_75t_L g5579 ( 
.A1(n_5264),
.A2(n_2851),
.B1(n_2950),
.B2(n_2946),
.Y(n_5579)
);

INVx2_ASAP7_75t_SL g5580 ( 
.A(n_5210),
.Y(n_5580)
);

CKINVDCx11_ASAP7_75t_R g5581 ( 
.A(n_5331),
.Y(n_5581)
);

OAI22xp5_ASAP7_75t_L g5582 ( 
.A1(n_5421),
.A2(n_5290),
.B1(n_5215),
.B2(n_5383),
.Y(n_5582)
);

AO21x1_ASAP7_75t_L g5583 ( 
.A1(n_5569),
.A2(n_5330),
.B(n_5326),
.Y(n_5583)
);

OAI21xp5_ASAP7_75t_L g5584 ( 
.A1(n_5417),
.A2(n_5329),
.B(n_5276),
.Y(n_5584)
);

A2O1A1Ixp33_ASAP7_75t_L g5585 ( 
.A1(n_5548),
.A2(n_5332),
.B(n_5317),
.C(n_5274),
.Y(n_5585)
);

INVx1_ASAP7_75t_L g5586 ( 
.A(n_5476),
.Y(n_5586)
);

AOI22xp33_ASAP7_75t_L g5587 ( 
.A1(n_5574),
.A2(n_5408),
.B1(n_5218),
.B2(n_5334),
.Y(n_5587)
);

CKINVDCx20_ASAP7_75t_R g5588 ( 
.A(n_5411),
.Y(n_5588)
);

CKINVDCx20_ASAP7_75t_R g5589 ( 
.A(n_5424),
.Y(n_5589)
);

OAI221xp5_ASAP7_75t_L g5590 ( 
.A1(n_5420),
.A2(n_5250),
.B1(n_5313),
.B2(n_5311),
.C(n_5325),
.Y(n_5590)
);

OAI222xp33_ASAP7_75t_L g5591 ( 
.A1(n_5409),
.A2(n_5279),
.B1(n_5272),
.B2(n_5382),
.C1(n_5315),
.C2(n_5381),
.Y(n_5591)
);

INVx1_ASAP7_75t_SL g5592 ( 
.A(n_5456),
.Y(n_5592)
);

OA21x2_ASAP7_75t_L g5593 ( 
.A1(n_5449),
.A2(n_5438),
.B(n_5447),
.Y(n_5593)
);

INVx1_ASAP7_75t_L g5594 ( 
.A(n_5481),
.Y(n_5594)
);

NAND2xp5_ASAP7_75t_L g5595 ( 
.A(n_5506),
.B(n_5242),
.Y(n_5595)
);

OAI22xp5_ASAP7_75t_L g5596 ( 
.A1(n_5491),
.A2(n_5382),
.B1(n_5251),
.B2(n_5260),
.Y(n_5596)
);

AO221x1_ASAP7_75t_L g5597 ( 
.A1(n_5415),
.A2(n_5301),
.B1(n_5372),
.B2(n_5358),
.C(n_5279),
.Y(n_5597)
);

AND2x2_ASAP7_75t_SL g5598 ( 
.A(n_5425),
.B(n_5272),
.Y(n_5598)
);

NAND2x1p5_ASAP7_75t_L g5599 ( 
.A(n_5490),
.B(n_5358),
.Y(n_5599)
);

AOI22xp5_ASAP7_75t_L g5600 ( 
.A1(n_5511),
.A2(n_5346),
.B1(n_5372),
.B2(n_5352),
.Y(n_5600)
);

AOI22xp33_ASAP7_75t_L g5601 ( 
.A1(n_5428),
.A2(n_5353),
.B1(n_5364),
.B2(n_5348),
.Y(n_5601)
);

O2A1O1Ixp33_ASAP7_75t_L g5602 ( 
.A1(n_5467),
.A2(n_5384),
.B(n_67),
.C(n_65),
.Y(n_5602)
);

OAI22xp5_ASAP7_75t_L g5603 ( 
.A1(n_5441),
.A2(n_5367),
.B1(n_5389),
.B2(n_69),
.Y(n_5603)
);

AND2x2_ASAP7_75t_L g5604 ( 
.A(n_5489),
.B(n_66),
.Y(n_5604)
);

INVx1_ASAP7_75t_SL g5605 ( 
.A(n_5525),
.Y(n_5605)
);

OAI22xp33_ASAP7_75t_L g5606 ( 
.A1(n_5535),
.A2(n_2950),
.B1(n_2958),
.B2(n_2946),
.Y(n_5606)
);

CKINVDCx5p33_ASAP7_75t_R g5607 ( 
.A(n_5435),
.Y(n_5607)
);

AND2x2_ASAP7_75t_L g5608 ( 
.A(n_5530),
.B(n_68),
.Y(n_5608)
);

AOI22xp33_ASAP7_75t_L g5609 ( 
.A1(n_5437),
.A2(n_2229),
.B1(n_2234),
.B2(n_2224),
.Y(n_5609)
);

AOI221xp5_ASAP7_75t_L g5610 ( 
.A1(n_5410),
.A2(n_1406),
.B1(n_1465),
.B2(n_1303),
.C(n_1299),
.Y(n_5610)
);

CKINVDCx20_ASAP7_75t_R g5611 ( 
.A(n_5479),
.Y(n_5611)
);

NAND2xp5_ASAP7_75t_L g5612 ( 
.A(n_5497),
.B(n_5494),
.Y(n_5612)
);

AOI22xp33_ASAP7_75t_L g5613 ( 
.A1(n_5413),
.A2(n_2234),
.B1(n_2242),
.B2(n_2229),
.Y(n_5613)
);

AOI22xp33_ASAP7_75t_L g5614 ( 
.A1(n_5543),
.A2(n_2242),
.B1(n_2234),
.B2(n_2123),
.Y(n_5614)
);

AOI22xp33_ASAP7_75t_L g5615 ( 
.A1(n_5520),
.A2(n_2242),
.B1(n_2123),
.B2(n_2132),
.Y(n_5615)
);

OAI22xp33_ASAP7_75t_L g5616 ( 
.A1(n_5418),
.A2(n_2962),
.B1(n_2969),
.B2(n_2958),
.Y(n_5616)
);

AOI22xp33_ASAP7_75t_L g5617 ( 
.A1(n_5540),
.A2(n_2242),
.B1(n_2123),
.B2(n_2132),
.Y(n_5617)
);

AND2x2_ASAP7_75t_L g5618 ( 
.A(n_5445),
.B(n_68),
.Y(n_5618)
);

AND2x2_ASAP7_75t_L g5619 ( 
.A(n_5445),
.B(n_71),
.Y(n_5619)
);

OAI21xp5_ASAP7_75t_L g5620 ( 
.A1(n_5452),
.A2(n_2075),
.B(n_2058),
.Y(n_5620)
);

CKINVDCx8_ASAP7_75t_R g5621 ( 
.A(n_5454),
.Y(n_5621)
);

INVxp67_ASAP7_75t_L g5622 ( 
.A(n_5499),
.Y(n_5622)
);

OAI22xp5_ASAP7_75t_L g5623 ( 
.A1(n_5475),
.A2(n_75),
.B1(n_73),
.B2(n_74),
.Y(n_5623)
);

OAI22xp5_ASAP7_75t_L g5624 ( 
.A1(n_5512),
.A2(n_76),
.B1(n_73),
.B2(n_75),
.Y(n_5624)
);

OR2x2_ASAP7_75t_L g5625 ( 
.A(n_5473),
.B(n_5158),
.Y(n_5625)
);

INVx2_ASAP7_75t_L g5626 ( 
.A(n_5567),
.Y(n_5626)
);

AOI22xp33_ASAP7_75t_L g5627 ( 
.A1(n_5422),
.A2(n_5448),
.B1(n_5523),
.B2(n_5529),
.Y(n_5627)
);

AOI22xp33_ASAP7_75t_L g5628 ( 
.A1(n_5486),
.A2(n_2242),
.B1(n_2123),
.B2(n_2132),
.Y(n_5628)
);

OAI22xp5_ASAP7_75t_L g5629 ( 
.A1(n_5507),
.A2(n_81),
.B1(n_78),
.B2(n_80),
.Y(n_5629)
);

CKINVDCx5p33_ASAP7_75t_R g5630 ( 
.A(n_5432),
.Y(n_5630)
);

AND2x2_ASAP7_75t_L g5631 ( 
.A(n_5446),
.B(n_82),
.Y(n_5631)
);

AOI21xp5_ASAP7_75t_L g5632 ( 
.A1(n_5546),
.A2(n_1465),
.B(n_1406),
.Y(n_5632)
);

AOI22xp33_ASAP7_75t_L g5633 ( 
.A1(n_5514),
.A2(n_5442),
.B1(n_5502),
.B2(n_5532),
.Y(n_5633)
);

OAI22xp5_ASAP7_75t_L g5634 ( 
.A1(n_5521),
.A2(n_5459),
.B1(n_5463),
.B2(n_5440),
.Y(n_5634)
);

OAI22xp5_ASAP7_75t_L g5635 ( 
.A1(n_5440),
.A2(n_90),
.B1(n_86),
.B2(n_88),
.Y(n_5635)
);

INVx2_ASAP7_75t_L g5636 ( 
.A(n_5550),
.Y(n_5636)
);

BUFx4f_ASAP7_75t_SL g5637 ( 
.A(n_5469),
.Y(n_5637)
);

NOR2x1_ASAP7_75t_L g5638 ( 
.A(n_5419),
.B(n_86),
.Y(n_5638)
);

AOI22xp33_ASAP7_75t_L g5639 ( 
.A1(n_5442),
.A2(n_2123),
.B1(n_2132),
.B2(n_2109),
.Y(n_5639)
);

AND2x2_ASAP7_75t_L g5640 ( 
.A(n_5554),
.B(n_91),
.Y(n_5640)
);

NOR2x1_ASAP7_75t_R g5641 ( 
.A(n_5416),
.B(n_92),
.Y(n_5641)
);

BUFx6f_ASAP7_75t_L g5642 ( 
.A(n_5431),
.Y(n_5642)
);

AOI22xp33_ASAP7_75t_L g5643 ( 
.A1(n_5502),
.A2(n_2132),
.B1(n_2109),
.B2(n_2974),
.Y(n_5643)
);

OAI21x1_ASAP7_75t_L g5644 ( 
.A1(n_5412),
.A2(n_5173),
.B(n_5158),
.Y(n_5644)
);

HB1xp67_ASAP7_75t_L g5645 ( 
.A(n_5547),
.Y(n_5645)
);

OAI22xp5_ASAP7_75t_L g5646 ( 
.A1(n_5459),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_5646)
);

INVx4_ASAP7_75t_L g5647 ( 
.A(n_5431),
.Y(n_5647)
);

AOI22xp5_ASAP7_75t_L g5648 ( 
.A1(n_5423),
.A2(n_2075),
.B1(n_2094),
.B2(n_2058),
.Y(n_5648)
);

AND2x2_ASAP7_75t_L g5649 ( 
.A(n_5496),
.B(n_93),
.Y(n_5649)
);

OR2x2_ASAP7_75t_L g5650 ( 
.A(n_5531),
.B(n_5173),
.Y(n_5650)
);

NAND2xp33_ASAP7_75t_SL g5651 ( 
.A(n_5555),
.B(n_95),
.Y(n_5651)
);

AOI221xp5_ASAP7_75t_L g5652 ( 
.A1(n_5538),
.A2(n_1483),
.B1(n_1502),
.B2(n_1465),
.C(n_1406),
.Y(n_5652)
);

INVx2_ASAP7_75t_L g5653 ( 
.A(n_5542),
.Y(n_5653)
);

AOI22xp33_ASAP7_75t_L g5654 ( 
.A1(n_5498),
.A2(n_2109),
.B1(n_2981),
.B2(n_2977),
.Y(n_5654)
);

INVx2_ASAP7_75t_L g5655 ( 
.A(n_5488),
.Y(n_5655)
);

AOI22xp33_ASAP7_75t_SL g5656 ( 
.A1(n_5463),
.A2(n_2094),
.B1(n_2075),
.B2(n_2109),
.Y(n_5656)
);

NAND3xp33_ASAP7_75t_SL g5657 ( 
.A(n_5460),
.B(n_95),
.C(n_96),
.Y(n_5657)
);

NAND3xp33_ASAP7_75t_SL g5658 ( 
.A(n_5466),
.B(n_97),
.C(n_98),
.Y(n_5658)
);

AND2x2_ASAP7_75t_L g5659 ( 
.A(n_5563),
.B(n_97),
.Y(n_5659)
);

AOI22xp33_ASAP7_75t_L g5660 ( 
.A1(n_5498),
.A2(n_2992),
.B1(n_2999),
.B2(n_2982),
.Y(n_5660)
);

INVx2_ASAP7_75t_L g5661 ( 
.A(n_5492),
.Y(n_5661)
);

INVx2_ASAP7_75t_L g5662 ( 
.A(n_5493),
.Y(n_5662)
);

NAND3xp33_ASAP7_75t_L g5663 ( 
.A(n_5485),
.B(n_5552),
.C(n_5553),
.Y(n_5663)
);

AOI21xp5_ASAP7_75t_R g5664 ( 
.A1(n_5482),
.A2(n_98),
.B(n_99),
.Y(n_5664)
);

OAI221xp5_ASAP7_75t_L g5665 ( 
.A1(n_5477),
.A2(n_1483),
.B1(n_1502),
.B2(n_1465),
.C(n_1406),
.Y(n_5665)
);

INVx2_ASAP7_75t_L g5666 ( 
.A(n_5504),
.Y(n_5666)
);

BUFx6f_ASAP7_75t_L g5667 ( 
.A(n_5416),
.Y(n_5667)
);

OAI22xp5_ASAP7_75t_L g5668 ( 
.A1(n_5474),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_5668)
);

NAND2xp33_ASAP7_75t_R g5669 ( 
.A(n_5434),
.B(n_102),
.Y(n_5669)
);

NAND3xp33_ASAP7_75t_SL g5670 ( 
.A(n_5450),
.B(n_105),
.C(n_107),
.Y(n_5670)
);

INVx6_ASAP7_75t_L g5671 ( 
.A(n_5426),
.Y(n_5671)
);

CKINVDCx16_ASAP7_75t_R g5672 ( 
.A(n_5430),
.Y(n_5672)
);

AND2x2_ASAP7_75t_L g5673 ( 
.A(n_5571),
.B(n_105),
.Y(n_5673)
);

AO21x2_ASAP7_75t_L g5674 ( 
.A1(n_5545),
.A2(n_2032),
.B(n_2022),
.Y(n_5674)
);

NAND2x1p5_ASAP7_75t_L g5675 ( 
.A(n_5490),
.B(n_1483),
.Y(n_5675)
);

AOI21xp5_ASAP7_75t_L g5676 ( 
.A1(n_5444),
.A2(n_1502),
.B(n_1483),
.Y(n_5676)
);

INVx2_ASAP7_75t_L g5677 ( 
.A(n_5524),
.Y(n_5677)
);

CKINVDCx16_ASAP7_75t_R g5678 ( 
.A(n_5430),
.Y(n_5678)
);

CKINVDCx6p67_ASAP7_75t_R g5679 ( 
.A(n_5419),
.Y(n_5679)
);

INVx2_ASAP7_75t_L g5680 ( 
.A(n_5534),
.Y(n_5680)
);

OAI22xp5_ASAP7_75t_L g5681 ( 
.A1(n_5474),
.A2(n_110),
.B1(n_108),
.B2(n_109),
.Y(n_5681)
);

AOI21xp5_ASAP7_75t_L g5682 ( 
.A1(n_5425),
.A2(n_1516),
.B(n_1502),
.Y(n_5682)
);

OAI22xp5_ASAP7_75t_L g5683 ( 
.A1(n_5436),
.A2(n_5487),
.B1(n_5495),
.B2(n_5433),
.Y(n_5683)
);

INVx1_ASAP7_75t_L g5684 ( 
.A(n_5429),
.Y(n_5684)
);

OAI22xp33_ASAP7_75t_L g5685 ( 
.A1(n_5490),
.A2(n_1562),
.B1(n_1516),
.B2(n_2534),
.Y(n_5685)
);

AOI22xp33_ASAP7_75t_L g5686 ( 
.A1(n_5565),
.A2(n_2094),
.B1(n_2039),
.B2(n_2050),
.Y(n_5686)
);

OR2x2_ASAP7_75t_L g5687 ( 
.A(n_5556),
.B(n_5173),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5439),
.Y(n_5688)
);

OAI221xp5_ASAP7_75t_L g5689 ( 
.A1(n_5455),
.A2(n_1562),
.B1(n_1516),
.B2(n_2022),
.C(n_2062),
.Y(n_5689)
);

BUFx6f_ASAP7_75t_SL g5690 ( 
.A(n_5443),
.Y(n_5690)
);

NAND2xp5_ASAP7_75t_L g5691 ( 
.A(n_5562),
.B(n_110),
.Y(n_5691)
);

AND2x2_ASAP7_75t_L g5692 ( 
.A(n_5503),
.B(n_111),
.Y(n_5692)
);

AOI22xp33_ASAP7_75t_SL g5693 ( 
.A1(n_5516),
.A2(n_1562),
.B1(n_1516),
.B2(n_113),
.Y(n_5693)
);

A2O1A1Ixp33_ASAP7_75t_L g5694 ( 
.A1(n_5533),
.A2(n_114),
.B(n_111),
.C(n_112),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_5570),
.B(n_114),
.Y(n_5695)
);

OAI22xp5_ASAP7_75t_L g5696 ( 
.A1(n_5566),
.A2(n_117),
.B1(n_115),
.B2(n_116),
.Y(n_5696)
);

OAI221xp5_ASAP7_75t_L g5697 ( 
.A1(n_5518),
.A2(n_1562),
.B1(n_2064),
.B2(n_2062),
.C(n_1957),
.Y(n_5697)
);

INVx3_ASAP7_75t_L g5698 ( 
.A(n_5483),
.Y(n_5698)
);

INVx5_ASAP7_75t_L g5699 ( 
.A(n_5414),
.Y(n_5699)
);

BUFx3_ASAP7_75t_L g5700 ( 
.A(n_5484),
.Y(n_5700)
);

OAI22xp5_ASAP7_75t_L g5701 ( 
.A1(n_5564),
.A2(n_120),
.B1(n_118),
.B2(n_119),
.Y(n_5701)
);

CKINVDCx5p33_ASAP7_75t_R g5702 ( 
.A(n_5577),
.Y(n_5702)
);

CKINVDCx9p33_ASAP7_75t_R g5703 ( 
.A(n_5426),
.Y(n_5703)
);

AOI22xp33_ASAP7_75t_SL g5704 ( 
.A1(n_5500),
.A2(n_1562),
.B1(n_122),
.B2(n_118),
.Y(n_5704)
);

OAI22xp33_ASAP7_75t_L g5705 ( 
.A1(n_5457),
.A2(n_2535),
.B1(n_2542),
.B2(n_2534),
.Y(n_5705)
);

INVx1_ASAP7_75t_L g5706 ( 
.A(n_5458),
.Y(n_5706)
);

A2O1A1Ixp33_ASAP7_75t_L g5707 ( 
.A1(n_5526),
.A2(n_123),
.B(n_121),
.C(n_122),
.Y(n_5707)
);

OR2x2_ASAP7_75t_L g5708 ( 
.A(n_5465),
.B(n_5175),
.Y(n_5708)
);

AOI221xp5_ASAP7_75t_L g5709 ( 
.A1(n_5462),
.A2(n_128),
.B1(n_124),
.B2(n_127),
.C(n_129),
.Y(n_5709)
);

AND2x4_ASAP7_75t_L g5710 ( 
.A(n_5501),
.B(n_5464),
.Y(n_5710)
);

BUFx2_ASAP7_75t_L g5711 ( 
.A(n_5500),
.Y(n_5711)
);

AOI22xp5_ASAP7_75t_L g5712 ( 
.A1(n_5515),
.A2(n_2136),
.B1(n_2779),
.B2(n_2770),
.Y(n_5712)
);

OAI21x1_ASAP7_75t_L g5713 ( 
.A1(n_5513),
.A2(n_5175),
.B(n_2535),
.Y(n_5713)
);

AOI22xp33_ASAP7_75t_L g5714 ( 
.A1(n_5558),
.A2(n_2505),
.B1(n_2515),
.B2(n_2477),
.Y(n_5714)
);

AND2x2_ASAP7_75t_L g5715 ( 
.A(n_5427),
.B(n_128),
.Y(n_5715)
);

CKINVDCx11_ASAP7_75t_R g5716 ( 
.A(n_5468),
.Y(n_5716)
);

INVx2_ASAP7_75t_L g5717 ( 
.A(n_5461),
.Y(n_5717)
);

NAND2x1p5_ASAP7_75t_L g5718 ( 
.A(n_5471),
.B(n_2770),
.Y(n_5718)
);

INVx2_ASAP7_75t_L g5719 ( 
.A(n_5472),
.Y(n_5719)
);

AOI21xp5_ASAP7_75t_L g5720 ( 
.A1(n_5464),
.A2(n_129),
.B(n_130),
.Y(n_5720)
);

NAND2xp33_ASAP7_75t_R g5721 ( 
.A(n_5575),
.B(n_131),
.Y(n_5721)
);

OR2x2_ASAP7_75t_L g5722 ( 
.A(n_5580),
.B(n_5175),
.Y(n_5722)
);

AND2x4_ASAP7_75t_SL g5723 ( 
.A(n_5522),
.B(n_2505),
.Y(n_5723)
);

BUFx4f_ASAP7_75t_SL g5724 ( 
.A(n_5453),
.Y(n_5724)
);

AND2x2_ASAP7_75t_L g5725 ( 
.A(n_5427),
.B(n_132),
.Y(n_5725)
);

AOI22xp33_ASAP7_75t_L g5726 ( 
.A1(n_5505),
.A2(n_2522),
.B1(n_2515),
.B2(n_2770),
.Y(n_5726)
);

AND2x4_ASAP7_75t_L g5727 ( 
.A(n_5471),
.B(n_132),
.Y(n_5727)
);

INVx3_ASAP7_75t_L g5728 ( 
.A(n_5522),
.Y(n_5728)
);

INVx2_ASAP7_75t_L g5729 ( 
.A(n_5508),
.Y(n_5729)
);

INVx3_ASAP7_75t_L g5730 ( 
.A(n_5508),
.Y(n_5730)
);

AOI21xp5_ASAP7_75t_L g5731 ( 
.A1(n_5579),
.A2(n_135),
.B(n_136),
.Y(n_5731)
);

BUFx6f_ASAP7_75t_L g5732 ( 
.A(n_5581),
.Y(n_5732)
);

CKINVDCx16_ASAP7_75t_R g5733 ( 
.A(n_5572),
.Y(n_5733)
);

INVx4_ASAP7_75t_L g5734 ( 
.A(n_5561),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5576),
.Y(n_5735)
);

OR2x2_ASAP7_75t_L g5736 ( 
.A(n_5509),
.B(n_5519),
.Y(n_5736)
);

NAND2xp5_ASAP7_75t_L g5737 ( 
.A(n_5478),
.B(n_135),
.Y(n_5737)
);

OAI22xp5_ASAP7_75t_L g5738 ( 
.A1(n_5559),
.A2(n_141),
.B1(n_137),
.B2(n_139),
.Y(n_5738)
);

BUFx3_ASAP7_75t_L g5739 ( 
.A(n_5528),
.Y(n_5739)
);

BUFx3_ASAP7_75t_L g5740 ( 
.A(n_5528),
.Y(n_5740)
);

INVx2_ASAP7_75t_L g5741 ( 
.A(n_5519),
.Y(n_5741)
);

AOI22xp33_ASAP7_75t_L g5742 ( 
.A1(n_5583),
.A2(n_5537),
.B1(n_5544),
.B2(n_5536),
.Y(n_5742)
);

NAND2xp5_ASAP7_75t_L g5743 ( 
.A(n_5645),
.B(n_5451),
.Y(n_5743)
);

CKINVDCx16_ASAP7_75t_R g5744 ( 
.A(n_5721),
.Y(n_5744)
);

BUFx4f_ASAP7_75t_SL g5745 ( 
.A(n_5588),
.Y(n_5745)
);

OAI22xp5_ASAP7_75t_L g5746 ( 
.A1(n_5664),
.A2(n_5470),
.B1(n_5537),
.B2(n_5536),
.Y(n_5746)
);

OAI22xp33_ASAP7_75t_L g5747 ( 
.A1(n_5669),
.A2(n_5584),
.B1(n_5590),
.B2(n_5658),
.Y(n_5747)
);

NAND3xp33_ASAP7_75t_L g5748 ( 
.A(n_5696),
.B(n_5480),
.C(n_5578),
.Y(n_5748)
);

BUFx6f_ASAP7_75t_L g5749 ( 
.A(n_5642),
.Y(n_5749)
);

INVx3_ASAP7_75t_L g5750 ( 
.A(n_5732),
.Y(n_5750)
);

CKINVDCx11_ASAP7_75t_R g5751 ( 
.A(n_5611),
.Y(n_5751)
);

AOI22xp33_ASAP7_75t_L g5752 ( 
.A1(n_5651),
.A2(n_5551),
.B1(n_5517),
.B2(n_5549),
.Y(n_5752)
);

AOI22xp33_ASAP7_75t_SL g5753 ( 
.A1(n_5597),
.A2(n_5557),
.B1(n_5568),
.B2(n_5539),
.Y(n_5753)
);

CKINVDCx20_ASAP7_75t_R g5754 ( 
.A(n_5589),
.Y(n_5754)
);

OAI22xp5_ASAP7_75t_L g5755 ( 
.A1(n_5585),
.A2(n_5557),
.B1(n_5510),
.B2(n_5527),
.Y(n_5755)
);

NAND2xp5_ASAP7_75t_L g5756 ( 
.A(n_5691),
.B(n_5557),
.Y(n_5756)
);

OAI22xp5_ASAP7_75t_L g5757 ( 
.A1(n_5622),
.A2(n_5541),
.B1(n_5573),
.B2(n_5560),
.Y(n_5757)
);

INVx2_ASAP7_75t_L g5758 ( 
.A(n_5727),
.Y(n_5758)
);

AOI22xp33_ASAP7_75t_L g5759 ( 
.A1(n_5628),
.A2(n_2522),
.B1(n_2800),
.B2(n_2779),
.Y(n_5759)
);

CKINVDCx20_ASAP7_75t_R g5760 ( 
.A(n_5716),
.Y(n_5760)
);

AOI22xp33_ASAP7_75t_L g5761 ( 
.A1(n_5663),
.A2(n_2800),
.B1(n_2807),
.B2(n_2779),
.Y(n_5761)
);

OAI21xp5_ASAP7_75t_SL g5762 ( 
.A1(n_5592),
.A2(n_144),
.B(n_143),
.Y(n_5762)
);

AOI22xp33_ASAP7_75t_L g5763 ( 
.A1(n_5663),
.A2(n_2807),
.B1(n_2808),
.B2(n_2800),
.Y(n_5763)
);

INVx2_ASAP7_75t_L g5764 ( 
.A(n_5727),
.Y(n_5764)
);

BUFx6f_ASAP7_75t_SL g5765 ( 
.A(n_5642),
.Y(n_5765)
);

OAI22xp5_ASAP7_75t_L g5766 ( 
.A1(n_5627),
.A2(n_145),
.B1(n_142),
.B2(n_143),
.Y(n_5766)
);

NAND2xp33_ASAP7_75t_SL g5767 ( 
.A(n_5690),
.B(n_148),
.Y(n_5767)
);

AOI22xp33_ASAP7_75t_SL g5768 ( 
.A1(n_5683),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_5768)
);

INVx2_ASAP7_75t_L g5769 ( 
.A(n_5719),
.Y(n_5769)
);

CKINVDCx6p67_ASAP7_75t_R g5770 ( 
.A(n_5703),
.Y(n_5770)
);

AOI222xp33_ASAP7_75t_L g5771 ( 
.A1(n_5657),
.A2(n_175),
.B1(n_158),
.B2(n_185),
.C1(n_167),
.C2(n_149),
.Y(n_5771)
);

NAND2xp5_ASAP7_75t_L g5772 ( 
.A(n_5695),
.B(n_150),
.Y(n_5772)
);

AOI22xp5_ASAP7_75t_SL g5773 ( 
.A1(n_5582),
.A2(n_153),
.B1(n_151),
.B2(n_152),
.Y(n_5773)
);

OAI21xp5_ASAP7_75t_SL g5774 ( 
.A1(n_5582),
.A2(n_154),
.B(n_153),
.Y(n_5774)
);

AND2x2_ASAP7_75t_L g5775 ( 
.A(n_5598),
.B(n_152),
.Y(n_5775)
);

AOI22xp33_ASAP7_75t_L g5776 ( 
.A1(n_5665),
.A2(n_2808),
.B1(n_2807),
.B2(n_2064),
.Y(n_5776)
);

BUFx4f_ASAP7_75t_SL g5777 ( 
.A(n_5647),
.Y(n_5777)
);

AOI22xp33_ASAP7_75t_L g5778 ( 
.A1(n_5614),
.A2(n_2669),
.B1(n_2689),
.B2(n_2665),
.Y(n_5778)
);

NAND3xp33_ASAP7_75t_L g5779 ( 
.A(n_5696),
.B(n_155),
.C(n_158),
.Y(n_5779)
);

AOI22xp33_ASAP7_75t_L g5780 ( 
.A1(n_5717),
.A2(n_5655),
.B1(n_5662),
.B2(n_5661),
.Y(n_5780)
);

OAI21xp33_ASAP7_75t_L g5781 ( 
.A1(n_5612),
.A2(n_160),
.B(n_161),
.Y(n_5781)
);

OAI22xp5_ASAP7_75t_L g5782 ( 
.A1(n_5634),
.A2(n_163),
.B1(n_160),
.B2(n_162),
.Y(n_5782)
);

AOI22xp33_ASAP7_75t_L g5783 ( 
.A1(n_5666),
.A2(n_2694),
.B1(n_2698),
.B2(n_2689),
.Y(n_5783)
);

AND2x2_ASAP7_75t_L g5784 ( 
.A(n_5698),
.B(n_165),
.Y(n_5784)
);

BUFx12f_ASAP7_75t_L g5785 ( 
.A(n_5642),
.Y(n_5785)
);

INVx3_ASAP7_75t_L g5786 ( 
.A(n_5621),
.Y(n_5786)
);

INVx2_ASAP7_75t_SL g5787 ( 
.A(n_5607),
.Y(n_5787)
);

AOI22xp33_ASAP7_75t_SL g5788 ( 
.A1(n_5593),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_5788)
);

OAI22xp33_ASAP7_75t_L g5789 ( 
.A1(n_5600),
.A2(n_2657),
.B1(n_2577),
.B2(n_3155),
.Y(n_5789)
);

AOI22xp33_ASAP7_75t_SL g5790 ( 
.A1(n_5593),
.A2(n_5620),
.B1(n_5626),
.B2(n_5603),
.Y(n_5790)
);

AND2x2_ASAP7_75t_L g5791 ( 
.A(n_5698),
.B(n_172),
.Y(n_5791)
);

NOR2xp33_ASAP7_75t_L g5792 ( 
.A(n_5672),
.B(n_173),
.Y(n_5792)
);

OAI22xp5_ASAP7_75t_SL g5793 ( 
.A1(n_5733),
.A2(n_178),
.B1(n_174),
.B2(n_176),
.Y(n_5793)
);

BUFx6f_ASAP7_75t_L g5794 ( 
.A(n_5700),
.Y(n_5794)
);

INVx4_ASAP7_75t_L g5795 ( 
.A(n_5637),
.Y(n_5795)
);

AOI22xp33_ASAP7_75t_L g5796 ( 
.A1(n_5677),
.A2(n_5680),
.B1(n_5735),
.B2(n_5603),
.Y(n_5796)
);

OAI21xp33_ASAP7_75t_L g5797 ( 
.A1(n_5709),
.A2(n_181),
.B(n_182),
.Y(n_5797)
);

OAI21xp5_ASAP7_75t_SL g5798 ( 
.A1(n_5704),
.A2(n_182),
.B(n_183),
.Y(n_5798)
);

INVx5_ASAP7_75t_L g5799 ( 
.A(n_5647),
.Y(n_5799)
);

OAI22xp5_ASAP7_75t_L g5800 ( 
.A1(n_5633),
.A2(n_189),
.B1(n_187),
.B2(n_188),
.Y(n_5800)
);

AOI22xp33_ASAP7_75t_L g5801 ( 
.A1(n_5606),
.A2(n_5670),
.B1(n_5632),
.B2(n_5653),
.Y(n_5801)
);

INVx1_ASAP7_75t_L g5802 ( 
.A(n_5684),
.Y(n_5802)
);

INVx1_ASAP7_75t_L g5803 ( 
.A(n_5688),
.Y(n_5803)
);

OAI22xp33_ASAP7_75t_L g5804 ( 
.A1(n_5600),
.A2(n_2698),
.B1(n_2601),
.B2(n_190),
.Y(n_5804)
);

AOI22xp33_ASAP7_75t_SL g5805 ( 
.A1(n_5739),
.A2(n_190),
.B1(n_187),
.B2(n_188),
.Y(n_5805)
);

AOI22xp33_ASAP7_75t_L g5806 ( 
.A1(n_5697),
.A2(n_2010),
.B1(n_2029),
.B2(n_2000),
.Y(n_5806)
);

AOI22xp33_ASAP7_75t_SL g5807 ( 
.A1(n_5740),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_5807)
);

OAI21xp5_ASAP7_75t_SL g5808 ( 
.A1(n_5638),
.A2(n_191),
.B(n_192),
.Y(n_5808)
);

INVx3_ASAP7_75t_L g5809 ( 
.A(n_5671),
.Y(n_5809)
);

AOI22xp33_ASAP7_75t_SL g5810 ( 
.A1(n_5728),
.A2(n_203),
.B1(n_198),
.B2(n_199),
.Y(n_5810)
);

NAND2xp5_ASAP7_75t_L g5811 ( 
.A(n_5604),
.B(n_199),
.Y(n_5811)
);

AOI222xp33_ASAP7_75t_L g5812 ( 
.A1(n_5629),
.A2(n_208),
.B1(n_210),
.B2(n_206),
.C1(n_207),
.C2(n_209),
.Y(n_5812)
);

OAI21xp5_ASAP7_75t_L g5813 ( 
.A1(n_5720),
.A2(n_206),
.B(n_207),
.Y(n_5813)
);

AOI22xp33_ASAP7_75t_SL g5814 ( 
.A1(n_5629),
.A2(n_212),
.B1(n_209),
.B2(n_211),
.Y(n_5814)
);

AOI22xp33_ASAP7_75t_SL g5815 ( 
.A1(n_5608),
.A2(n_215),
.B1(n_212),
.B2(n_213),
.Y(n_5815)
);

AOI21xp33_ASAP7_75t_L g5816 ( 
.A1(n_5602),
.A2(n_216),
.B(n_217),
.Y(n_5816)
);

OAI22xp5_ASAP7_75t_SL g5817 ( 
.A1(n_5699),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_5817)
);

INVx1_ASAP7_75t_L g5818 ( 
.A(n_5706),
.Y(n_5818)
);

AOI22xp33_ASAP7_75t_L g5819 ( 
.A1(n_5610),
.A2(n_5616),
.B1(n_5601),
.B2(n_5689),
.Y(n_5819)
);

BUFx12f_ASAP7_75t_L g5820 ( 
.A(n_5702),
.Y(n_5820)
);

INVx4_ASAP7_75t_L g5821 ( 
.A(n_5699),
.Y(n_5821)
);

INVx1_ASAP7_75t_L g5822 ( 
.A(n_5586),
.Y(n_5822)
);

NOR2xp33_ASAP7_75t_L g5823 ( 
.A(n_5678),
.B(n_220),
.Y(n_5823)
);

BUFx6f_ASAP7_75t_L g5824 ( 
.A(n_5699),
.Y(n_5824)
);

AOI22xp33_ASAP7_75t_L g5825 ( 
.A1(n_5676),
.A2(n_2010),
.B1(n_2029),
.B2(n_2000),
.Y(n_5825)
);

NOR2xp33_ASAP7_75t_L g5826 ( 
.A(n_5605),
.B(n_225),
.Y(n_5826)
);

INVx1_ASAP7_75t_L g5827 ( 
.A(n_5594),
.Y(n_5827)
);

INVx2_ASAP7_75t_L g5828 ( 
.A(n_5729),
.Y(n_5828)
);

OAI21xp5_ASAP7_75t_SL g5829 ( 
.A1(n_5591),
.A2(n_227),
.B(n_228),
.Y(n_5829)
);

INVx2_ASAP7_75t_SL g5830 ( 
.A(n_5671),
.Y(n_5830)
);

AND2x2_ASAP7_75t_L g5831 ( 
.A(n_5741),
.B(n_230),
.Y(n_5831)
);

AOI22xp33_ASAP7_75t_L g5832 ( 
.A1(n_5636),
.A2(n_2044),
.B1(n_1474),
.B2(n_1482),
.Y(n_5832)
);

INVx2_ASAP7_75t_SL g5833 ( 
.A(n_5724),
.Y(n_5833)
);

OAI21xp5_ASAP7_75t_SL g5834 ( 
.A1(n_5711),
.A2(n_231),
.B(n_232),
.Y(n_5834)
);

NOR2x1_ASAP7_75t_L g5835 ( 
.A(n_5734),
.B(n_233),
.Y(n_5835)
);

INVx2_ASAP7_75t_L g5836 ( 
.A(n_5675),
.Y(n_5836)
);

INVx2_ASAP7_75t_L g5837 ( 
.A(n_5736),
.Y(n_5837)
);

NAND3xp33_ASAP7_75t_L g5838 ( 
.A(n_5623),
.B(n_235),
.C(n_236),
.Y(n_5838)
);

AOI222xp33_ASAP7_75t_L g5839 ( 
.A1(n_5624),
.A2(n_238),
.B1(n_240),
.B2(n_235),
.C1(n_237),
.C2(n_239),
.Y(n_5839)
);

OAI21xp33_ASAP7_75t_L g5840 ( 
.A1(n_5595),
.A2(n_237),
.B(n_238),
.Y(n_5840)
);

NAND2xp5_ASAP7_75t_L g5841 ( 
.A(n_5618),
.B(n_240),
.Y(n_5841)
);

OAI22xp5_ASAP7_75t_L g5842 ( 
.A1(n_5599),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_5842)
);

AOI22xp5_ASAP7_75t_L g5843 ( 
.A1(n_5648),
.A2(n_2488),
.B1(n_1956),
.B2(n_1973),
.Y(n_5843)
);

NAND2xp5_ASAP7_75t_L g5844 ( 
.A(n_5619),
.B(n_244),
.Y(n_5844)
);

AOI22xp33_ASAP7_75t_L g5845 ( 
.A1(n_5613),
.A2(n_2034),
.B1(n_2226),
.B2(n_2102),
.Y(n_5845)
);

BUFx3_ASAP7_75t_L g5846 ( 
.A(n_5630),
.Y(n_5846)
);

BUFx4f_ASAP7_75t_SL g5847 ( 
.A(n_5679),
.Y(n_5847)
);

AOI22xp33_ASAP7_75t_L g5848 ( 
.A1(n_5731),
.A2(n_2034),
.B1(n_2226),
.B2(n_2102),
.Y(n_5848)
);

OAI22xp5_ASAP7_75t_L g5849 ( 
.A1(n_5596),
.A2(n_250),
.B1(n_248),
.B2(n_249),
.Y(n_5849)
);

OAI22xp5_ASAP7_75t_L g5850 ( 
.A1(n_5587),
.A2(n_253),
.B1(n_248),
.B2(n_252),
.Y(n_5850)
);

AOI22xp33_ASAP7_75t_L g5851 ( 
.A1(n_5654),
.A2(n_2034),
.B1(n_2102),
.B2(n_2099),
.Y(n_5851)
);

AOI22xp33_ASAP7_75t_L g5852 ( 
.A1(n_5726),
.A2(n_2226),
.B1(n_2099),
.B2(n_2153),
.Y(n_5852)
);

AOI22xp33_ASAP7_75t_L g5853 ( 
.A1(n_5643),
.A2(n_2226),
.B1(n_2099),
.B2(n_2153),
.Y(n_5853)
);

AOI211xp5_ASAP7_75t_L g5854 ( 
.A1(n_5641),
.A2(n_256),
.B(n_254),
.C(n_255),
.Y(n_5854)
);

INVx3_ASAP7_75t_L g5855 ( 
.A(n_5667),
.Y(n_5855)
);

NAND2xp5_ASAP7_75t_L g5856 ( 
.A(n_5631),
.B(n_255),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5708),
.Y(n_5857)
);

INVx2_ASAP7_75t_L g5858 ( 
.A(n_5730),
.Y(n_5858)
);

BUFx4f_ASAP7_75t_SL g5859 ( 
.A(n_5667),
.Y(n_5859)
);

INVx1_ASAP7_75t_L g5860 ( 
.A(n_5692),
.Y(n_5860)
);

OAI222xp33_ASAP7_75t_L g5861 ( 
.A1(n_5701),
.A2(n_266),
.B1(n_268),
.B2(n_264),
.C1(n_265),
.C2(n_267),
.Y(n_5861)
);

INVx5_ASAP7_75t_L g5862 ( 
.A(n_5667),
.Y(n_5862)
);

AOI22xp5_ASAP7_75t_L g5863 ( 
.A1(n_5701),
.A2(n_5738),
.B1(n_5646),
.B2(n_5668),
.Y(n_5863)
);

OAI21xp5_ASAP7_75t_SL g5864 ( 
.A1(n_5737),
.A2(n_269),
.B(n_270),
.Y(n_5864)
);

AOI222xp33_ASAP7_75t_L g5865 ( 
.A1(n_5635),
.A2(n_5646),
.B1(n_5668),
.B2(n_5681),
.C1(n_5707),
.C2(n_5640),
.Y(n_5865)
);

AND2x2_ASAP7_75t_L g5866 ( 
.A(n_5710),
.B(n_270),
.Y(n_5866)
);

CKINVDCx5p33_ASAP7_75t_R g5867 ( 
.A(n_5690),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_5649),
.Y(n_5868)
);

INVx1_ASAP7_75t_L g5869 ( 
.A(n_5625),
.Y(n_5869)
);

AOI22xp33_ASAP7_75t_L g5870 ( 
.A1(n_5714),
.A2(n_5617),
.B1(n_5686),
.B2(n_5609),
.Y(n_5870)
);

OAI22xp5_ASAP7_75t_L g5871 ( 
.A1(n_5723),
.A2(n_273),
.B1(n_271),
.B2(n_272),
.Y(n_5871)
);

OAI22xp5_ASAP7_75t_L g5872 ( 
.A1(n_5693),
.A2(n_276),
.B1(n_272),
.B2(n_273),
.Y(n_5872)
);

OAI22xp5_ASAP7_75t_L g5873 ( 
.A1(n_5705),
.A2(n_279),
.B1(n_276),
.B2(n_277),
.Y(n_5873)
);

INVx1_ASAP7_75t_L g5874 ( 
.A(n_5715),
.Y(n_5874)
);

AOI22xp33_ASAP7_75t_L g5875 ( 
.A1(n_5639),
.A2(n_2100),
.B1(n_2098),
.B2(n_1995),
.Y(n_5875)
);

OAI22xp5_ASAP7_75t_L g5876 ( 
.A1(n_5681),
.A2(n_286),
.B1(n_281),
.B2(n_283),
.Y(n_5876)
);

BUFx3_ASAP7_75t_L g5877 ( 
.A(n_5760),
.Y(n_5877)
);

NAND2xp5_ASAP7_75t_L g5878 ( 
.A(n_5774),
.B(n_5725),
.Y(n_5878)
);

INVx4_ASAP7_75t_L g5879 ( 
.A(n_5795),
.Y(n_5879)
);

NAND2xp5_ASAP7_75t_L g5880 ( 
.A(n_5774),
.B(n_5659),
.Y(n_5880)
);

NAND2x1p5_ASAP7_75t_L g5881 ( 
.A(n_5835),
.B(n_5673),
.Y(n_5881)
);

BUFx2_ASAP7_75t_L g5882 ( 
.A(n_5754),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5802),
.Y(n_5883)
);

OAI221xp5_ASAP7_75t_SL g5884 ( 
.A1(n_5742),
.A2(n_5694),
.B1(n_5650),
.B2(n_5660),
.C(n_5712),
.Y(n_5884)
);

INVx1_ASAP7_75t_L g5885 ( 
.A(n_5803),
.Y(n_5885)
);

AND2x2_ASAP7_75t_L g5886 ( 
.A(n_5862),
.B(n_5718),
.Y(n_5886)
);

BUFx6f_ASAP7_75t_L g5887 ( 
.A(n_5751),
.Y(n_5887)
);

AND2x2_ASAP7_75t_L g5888 ( 
.A(n_5862),
.B(n_5722),
.Y(n_5888)
);

AOI22xp33_ASAP7_75t_SL g5889 ( 
.A1(n_5744),
.A2(n_5687),
.B1(n_5644),
.B2(n_5674),
.Y(n_5889)
);

INVx2_ASAP7_75t_L g5890 ( 
.A(n_5758),
.Y(n_5890)
);

INVx2_ASAP7_75t_L g5891 ( 
.A(n_5764),
.Y(n_5891)
);

OAI21xp5_ASAP7_75t_L g5892 ( 
.A1(n_5762),
.A2(n_5656),
.B(n_5682),
.Y(n_5892)
);

INVx1_ASAP7_75t_SL g5893 ( 
.A(n_5745),
.Y(n_5893)
);

AND2x2_ASAP7_75t_L g5894 ( 
.A(n_5750),
.B(n_5713),
.Y(n_5894)
);

INVx1_ASAP7_75t_L g5895 ( 
.A(n_5818),
.Y(n_5895)
);

AOI22xp33_ASAP7_75t_L g5896 ( 
.A1(n_5790),
.A2(n_5685),
.B1(n_5712),
.B2(n_5615),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5822),
.Y(n_5897)
);

OAI21xp5_ASAP7_75t_SL g5898 ( 
.A1(n_5834),
.A2(n_5762),
.B(n_5829),
.Y(n_5898)
);

INVxp67_ASAP7_75t_L g5899 ( 
.A(n_5773),
.Y(n_5899)
);

INVx1_ASAP7_75t_L g5900 ( 
.A(n_5827),
.Y(n_5900)
);

HB1xp67_ASAP7_75t_L g5901 ( 
.A(n_5837),
.Y(n_5901)
);

INVx2_ASAP7_75t_L g5902 ( 
.A(n_5855),
.Y(n_5902)
);

HB1xp67_ASAP7_75t_L g5903 ( 
.A(n_5769),
.Y(n_5903)
);

NOR2x1_ASAP7_75t_L g5904 ( 
.A(n_5834),
.B(n_287),
.Y(n_5904)
);

NAND2xp5_ASAP7_75t_L g5905 ( 
.A(n_5788),
.B(n_5652),
.Y(n_5905)
);

BUFx8_ASAP7_75t_L g5906 ( 
.A(n_5765),
.Y(n_5906)
);

INVx2_ASAP7_75t_L g5907 ( 
.A(n_5775),
.Y(n_5907)
);

BUFx2_ASAP7_75t_L g5908 ( 
.A(n_5859),
.Y(n_5908)
);

AND2x2_ASAP7_75t_L g5909 ( 
.A(n_5809),
.B(n_288),
.Y(n_5909)
);

HB1xp67_ASAP7_75t_L g5910 ( 
.A(n_5828),
.Y(n_5910)
);

AND2x2_ASAP7_75t_L g5911 ( 
.A(n_5786),
.B(n_289),
.Y(n_5911)
);

AND2x2_ASAP7_75t_L g5912 ( 
.A(n_5830),
.B(n_5770),
.Y(n_5912)
);

AND2x2_ASAP7_75t_L g5913 ( 
.A(n_5824),
.B(n_290),
.Y(n_5913)
);

INVx1_ASAP7_75t_L g5914 ( 
.A(n_5868),
.Y(n_5914)
);

NAND2xp5_ASAP7_75t_L g5915 ( 
.A(n_5796),
.B(n_291),
.Y(n_5915)
);

AND2x2_ASAP7_75t_L g5916 ( 
.A(n_5821),
.B(n_5866),
.Y(n_5916)
);

AND2x2_ASAP7_75t_L g5917 ( 
.A(n_5860),
.B(n_292),
.Y(n_5917)
);

INVx2_ASAP7_75t_L g5918 ( 
.A(n_5858),
.Y(n_5918)
);

NAND2xp5_ASAP7_75t_L g5919 ( 
.A(n_5864),
.B(n_5747),
.Y(n_5919)
);

INVx3_ASAP7_75t_L g5920 ( 
.A(n_5820),
.Y(n_5920)
);

BUFx2_ASAP7_75t_L g5921 ( 
.A(n_5867),
.Y(n_5921)
);

INVxp67_ASAP7_75t_L g5922 ( 
.A(n_5794),
.Y(n_5922)
);

OR2x2_ASAP7_75t_L g5923 ( 
.A(n_5743),
.B(n_294),
.Y(n_5923)
);

AOI22xp33_ASAP7_75t_L g5924 ( 
.A1(n_5748),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_5924)
);

INVx1_ASAP7_75t_SL g5925 ( 
.A(n_5767),
.Y(n_5925)
);

AND2x4_ASAP7_75t_L g5926 ( 
.A(n_5799),
.B(n_295),
.Y(n_5926)
);

INVx1_ASAP7_75t_L g5927 ( 
.A(n_5772),
.Y(n_5927)
);

AND2x2_ASAP7_75t_L g5928 ( 
.A(n_5749),
.B(n_296),
.Y(n_5928)
);

INVx2_ASAP7_75t_L g5929 ( 
.A(n_5836),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5874),
.Y(n_5930)
);

BUFx2_ASAP7_75t_L g5931 ( 
.A(n_5785),
.Y(n_5931)
);

OAI21xp5_ASAP7_75t_SL g5932 ( 
.A1(n_5829),
.A2(n_297),
.B(n_298),
.Y(n_5932)
);

AND2x4_ASAP7_75t_L g5933 ( 
.A(n_5799),
.B(n_297),
.Y(n_5933)
);

CKINVDCx14_ASAP7_75t_R g5934 ( 
.A(n_5795),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5857),
.Y(n_5935)
);

AND2x4_ASAP7_75t_L g5936 ( 
.A(n_5799),
.B(n_298),
.Y(n_5936)
);

AND2x4_ASAP7_75t_L g5937 ( 
.A(n_5833),
.B(n_299),
.Y(n_5937)
);

INVx1_ASAP7_75t_L g5938 ( 
.A(n_5869),
.Y(n_5938)
);

OAI21xp33_ASAP7_75t_L g5939 ( 
.A1(n_5863),
.A2(n_1999),
.B(n_300),
.Y(n_5939)
);

INVxp67_ASAP7_75t_SL g5940 ( 
.A(n_5854),
.Y(n_5940)
);

INVx4_ASAP7_75t_L g5941 ( 
.A(n_5794),
.Y(n_5941)
);

INVxp67_ASAP7_75t_L g5942 ( 
.A(n_5826),
.Y(n_5942)
);

AND2x4_ASAP7_75t_L g5943 ( 
.A(n_5787),
.B(n_301),
.Y(n_5943)
);

HB1xp67_ASAP7_75t_L g5944 ( 
.A(n_5748),
.Y(n_5944)
);

OR2x2_ASAP7_75t_L g5945 ( 
.A(n_5756),
.B(n_301),
.Y(n_5945)
);

INVx2_ASAP7_75t_SL g5946 ( 
.A(n_5846),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_5831),
.Y(n_5947)
);

AOI22xp33_ASAP7_75t_L g5948 ( 
.A1(n_5816),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.Y(n_5948)
);

INVx1_ASAP7_75t_L g5949 ( 
.A(n_5856),
.Y(n_5949)
);

NAND2xp5_ASAP7_75t_L g5950 ( 
.A(n_5808),
.B(n_306),
.Y(n_5950)
);

INVx1_ASAP7_75t_L g5951 ( 
.A(n_5784),
.Y(n_5951)
);

INVx4_ASAP7_75t_L g5952 ( 
.A(n_5777),
.Y(n_5952)
);

AND2x2_ASAP7_75t_L g5953 ( 
.A(n_5792),
.B(n_306),
.Y(n_5953)
);

INVx2_ASAP7_75t_SL g5954 ( 
.A(n_5847),
.Y(n_5954)
);

AND2x2_ASAP7_75t_L g5955 ( 
.A(n_5823),
.B(n_307),
.Y(n_5955)
);

HB1xp67_ASAP7_75t_L g5956 ( 
.A(n_5766),
.Y(n_5956)
);

BUFx2_ASAP7_75t_SL g5957 ( 
.A(n_5791),
.Y(n_5957)
);

INVxp67_ASAP7_75t_SL g5958 ( 
.A(n_5854),
.Y(n_5958)
);

AND2x4_ASAP7_75t_L g5959 ( 
.A(n_5841),
.B(n_311),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5844),
.Y(n_5960)
);

INVx2_ASAP7_75t_L g5961 ( 
.A(n_5811),
.Y(n_5961)
);

OR2x2_ASAP7_75t_L g5962 ( 
.A(n_5746),
.B(n_312),
.Y(n_5962)
);

INVx3_ASAP7_75t_L g5963 ( 
.A(n_5808),
.Y(n_5963)
);

BUFx2_ASAP7_75t_L g5964 ( 
.A(n_5813),
.Y(n_5964)
);

AND2x4_ASAP7_75t_L g5965 ( 
.A(n_5838),
.B(n_313),
.Y(n_5965)
);

AO31x2_ASAP7_75t_L g5966 ( 
.A1(n_5800),
.A2(n_316),
.A3(n_314),
.B(n_315),
.Y(n_5966)
);

INVx2_ASAP7_75t_L g5967 ( 
.A(n_5817),
.Y(n_5967)
);

AND2x2_ASAP7_75t_L g5968 ( 
.A(n_5753),
.B(n_314),
.Y(n_5968)
);

INVx2_ASAP7_75t_L g5969 ( 
.A(n_5757),
.Y(n_5969)
);

INVx4_ASAP7_75t_L g5970 ( 
.A(n_5793),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5779),
.Y(n_5971)
);

INVx2_ASAP7_75t_SL g5972 ( 
.A(n_5782),
.Y(n_5972)
);

NAND2xp5_ASAP7_75t_L g5973 ( 
.A(n_5865),
.B(n_316),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_5779),
.Y(n_5974)
);

NAND2xp5_ASAP7_75t_L g5975 ( 
.A(n_5768),
.B(n_317),
.Y(n_5975)
);

NAND2xp5_ASAP7_75t_L g5976 ( 
.A(n_5781),
.B(n_319),
.Y(n_5976)
);

AOI22xp33_ASAP7_75t_L g5977 ( 
.A1(n_5797),
.A2(n_323),
.B1(n_320),
.B2(n_322),
.Y(n_5977)
);

NOR2xp33_ASAP7_75t_L g5978 ( 
.A(n_5798),
.B(n_320),
.Y(n_5978)
);

NAND2xp5_ASAP7_75t_L g5979 ( 
.A(n_5840),
.B(n_323),
.Y(n_5979)
);

INVxp67_ASAP7_75t_SL g5980 ( 
.A(n_5850),
.Y(n_5980)
);

BUFx2_ASAP7_75t_L g5981 ( 
.A(n_5849),
.Y(n_5981)
);

OAI22xp5_ASAP7_75t_L g5982 ( 
.A1(n_5798),
.A2(n_327),
.B1(n_325),
.B2(n_326),
.Y(n_5982)
);

AND2x2_ASAP7_75t_L g5983 ( 
.A(n_5882),
.B(n_5755),
.Y(n_5983)
);

AND2x2_ASAP7_75t_L g5984 ( 
.A(n_5908),
.B(n_5810),
.Y(n_5984)
);

INVx2_ASAP7_75t_L g5985 ( 
.A(n_5877),
.Y(n_5985)
);

NAND2xp5_ASAP7_75t_L g5986 ( 
.A(n_5944),
.B(n_5940),
.Y(n_5986)
);

AND2x2_ASAP7_75t_L g5987 ( 
.A(n_5887),
.B(n_5815),
.Y(n_5987)
);

BUFx3_ASAP7_75t_L g5988 ( 
.A(n_5906),
.Y(n_5988)
);

INVx1_ASAP7_75t_L g5989 ( 
.A(n_5901),
.Y(n_5989)
);

OR2x6_ASAP7_75t_L g5990 ( 
.A(n_5973),
.B(n_5842),
.Y(n_5990)
);

HB1xp67_ASAP7_75t_L g5991 ( 
.A(n_5963),
.Y(n_5991)
);

AND2x2_ASAP7_75t_L g5992 ( 
.A(n_5912),
.B(n_5752),
.Y(n_5992)
);

HB1xp67_ASAP7_75t_L g5993 ( 
.A(n_5963),
.Y(n_5993)
);

AND2x2_ASAP7_75t_L g5994 ( 
.A(n_5921),
.B(n_5805),
.Y(n_5994)
);

AND2x4_ASAP7_75t_L g5995 ( 
.A(n_5922),
.B(n_5916),
.Y(n_5995)
);

BUFx3_ASAP7_75t_L g5996 ( 
.A(n_5906),
.Y(n_5996)
);

NAND2xp5_ASAP7_75t_L g5997 ( 
.A(n_5944),
.B(n_5771),
.Y(n_5997)
);

AND2x2_ASAP7_75t_L g5998 ( 
.A(n_5893),
.B(n_5807),
.Y(n_5998)
);

OR2x2_ASAP7_75t_L g5999 ( 
.A(n_5971),
.B(n_5974),
.Y(n_5999)
);

INVx2_ASAP7_75t_SL g6000 ( 
.A(n_5920),
.Y(n_6000)
);

INVx3_ASAP7_75t_L g6001 ( 
.A(n_5941),
.Y(n_6001)
);

AND2x2_ASAP7_75t_L g6002 ( 
.A(n_5922),
.B(n_5801),
.Y(n_6002)
);

AND2x2_ASAP7_75t_L g6003 ( 
.A(n_5931),
.B(n_5814),
.Y(n_6003)
);

NAND2xp5_ASAP7_75t_L g6004 ( 
.A(n_5940),
.B(n_5812),
.Y(n_6004)
);

HB1xp67_ASAP7_75t_L g6005 ( 
.A(n_5956),
.Y(n_6005)
);

NAND2xp5_ASAP7_75t_L g6006 ( 
.A(n_5958),
.B(n_5839),
.Y(n_6006)
);

INVx2_ASAP7_75t_L g6007 ( 
.A(n_5904),
.Y(n_6007)
);

INVx1_ASAP7_75t_L g6008 ( 
.A(n_5903),
.Y(n_6008)
);

INVx1_ASAP7_75t_L g6009 ( 
.A(n_5910),
.Y(n_6009)
);

NOR2x1_ASAP7_75t_L g6010 ( 
.A(n_5898),
.B(n_5861),
.Y(n_6010)
);

INVx2_ASAP7_75t_L g6011 ( 
.A(n_5965),
.Y(n_6011)
);

INVx2_ASAP7_75t_L g6012 ( 
.A(n_5970),
.Y(n_6012)
);

NAND2xp5_ASAP7_75t_L g6013 ( 
.A(n_5924),
.B(n_5780),
.Y(n_6013)
);

HB1xp67_ASAP7_75t_L g6014 ( 
.A(n_5956),
.Y(n_6014)
);

INVx3_ASAP7_75t_L g6015 ( 
.A(n_5952),
.Y(n_6015)
);

AO21x2_ASAP7_75t_L g6016 ( 
.A1(n_5919),
.A2(n_5876),
.B(n_5872),
.Y(n_6016)
);

NAND2xp5_ASAP7_75t_L g6017 ( 
.A(n_5924),
.B(n_5761),
.Y(n_6017)
);

INVx1_ASAP7_75t_L g6018 ( 
.A(n_5914),
.Y(n_6018)
);

INVx1_ASAP7_75t_L g6019 ( 
.A(n_5949),
.Y(n_6019)
);

OR2x2_ASAP7_75t_L g6020 ( 
.A(n_5880),
.B(n_5763),
.Y(n_6020)
);

BUFx3_ASAP7_75t_L g6021 ( 
.A(n_5920),
.Y(n_6021)
);

INVx1_ASAP7_75t_L g6022 ( 
.A(n_5883),
.Y(n_6022)
);

AOI221xp5_ASAP7_75t_L g6023 ( 
.A1(n_5919),
.A2(n_5873),
.B1(n_5819),
.B2(n_5789),
.C(n_5804),
.Y(n_6023)
);

OR2x2_ASAP7_75t_L g6024 ( 
.A(n_5880),
.B(n_5871),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5885),
.Y(n_6025)
);

HB1xp67_ASAP7_75t_L g6026 ( 
.A(n_5942),
.Y(n_6026)
);

INVx1_ASAP7_75t_L g6027 ( 
.A(n_5895),
.Y(n_6027)
);

INVx1_ASAP7_75t_L g6028 ( 
.A(n_5897),
.Y(n_6028)
);

INVx3_ASAP7_75t_L g6029 ( 
.A(n_5952),
.Y(n_6029)
);

HB1xp67_ASAP7_75t_L g6030 ( 
.A(n_5942),
.Y(n_6030)
);

BUFx3_ASAP7_75t_L g6031 ( 
.A(n_5937),
.Y(n_6031)
);

OR2x2_ASAP7_75t_L g6032 ( 
.A(n_5930),
.B(n_5981),
.Y(n_6032)
);

INVx1_ASAP7_75t_L g6033 ( 
.A(n_5900),
.Y(n_6033)
);

AND2x2_ASAP7_75t_L g6034 ( 
.A(n_5946),
.B(n_5870),
.Y(n_6034)
);

AND2x2_ASAP7_75t_L g6035 ( 
.A(n_5954),
.B(n_5848),
.Y(n_6035)
);

INVx2_ASAP7_75t_L g6036 ( 
.A(n_5964),
.Y(n_6036)
);

NOR3xp33_ASAP7_75t_L g6037 ( 
.A(n_5932),
.B(n_5843),
.C(n_5825),
.Y(n_6037)
);

INVx2_ASAP7_75t_L g6038 ( 
.A(n_5881),
.Y(n_6038)
);

INVx2_ASAP7_75t_L g6039 ( 
.A(n_5950),
.Y(n_6039)
);

AND2x4_ASAP7_75t_L g6040 ( 
.A(n_5951),
.B(n_5783),
.Y(n_6040)
);

OR2x2_ASAP7_75t_L g6041 ( 
.A(n_5927),
.B(n_5806),
.Y(n_6041)
);

AND2x2_ASAP7_75t_L g6042 ( 
.A(n_5911),
.B(n_5832),
.Y(n_6042)
);

INVx2_ASAP7_75t_L g6043 ( 
.A(n_5950),
.Y(n_6043)
);

INVx2_ASAP7_75t_L g6044 ( 
.A(n_5966),
.Y(n_6044)
);

HB1xp67_ASAP7_75t_L g6045 ( 
.A(n_5978),
.Y(n_6045)
);

AND2x2_ASAP7_75t_L g6046 ( 
.A(n_5934),
.B(n_5778),
.Y(n_6046)
);

OR2x2_ASAP7_75t_L g6047 ( 
.A(n_5980),
.B(n_5875),
.Y(n_6047)
);

AOI22xp33_ASAP7_75t_L g6048 ( 
.A1(n_5899),
.A2(n_5759),
.B1(n_5845),
.B2(n_5776),
.Y(n_6048)
);

INVx2_ASAP7_75t_L g6049 ( 
.A(n_5943),
.Y(n_6049)
);

AND2x2_ASAP7_75t_L g6050 ( 
.A(n_5943),
.B(n_5902),
.Y(n_6050)
);

BUFx6f_ASAP7_75t_L g6051 ( 
.A(n_5879),
.Y(n_6051)
);

AND2x2_ASAP7_75t_L g6052 ( 
.A(n_5957),
.B(n_5851),
.Y(n_6052)
);

AND2x2_ASAP7_75t_L g6053 ( 
.A(n_5886),
.B(n_5852),
.Y(n_6053)
);

AND2x2_ASAP7_75t_L g6054 ( 
.A(n_5925),
.B(n_5853),
.Y(n_6054)
);

BUFx3_ASAP7_75t_L g6055 ( 
.A(n_5988),
.Y(n_6055)
);

INVx2_ASAP7_75t_L g6056 ( 
.A(n_6031),
.Y(n_6056)
);

INVx2_ASAP7_75t_L g6057 ( 
.A(n_6021),
.Y(n_6057)
);

INVx3_ASAP7_75t_L g6058 ( 
.A(n_5996),
.Y(n_6058)
);

AO21x2_ASAP7_75t_L g6059 ( 
.A1(n_5986),
.A2(n_5915),
.B(n_5968),
.Y(n_6059)
);

AOI211xp5_ASAP7_75t_SL g6060 ( 
.A1(n_5986),
.A2(n_5991),
.B(n_5993),
.C(n_6005),
.Y(n_6060)
);

AND2x2_ASAP7_75t_L g6061 ( 
.A(n_5985),
.B(n_5918),
.Y(n_6061)
);

NAND2xp5_ASAP7_75t_L g6062 ( 
.A(n_6010),
.B(n_5978),
.Y(n_6062)
);

HB1xp67_ASAP7_75t_L g6063 ( 
.A(n_5993),
.Y(n_6063)
);

OAI22xp5_ASAP7_75t_L g6064 ( 
.A1(n_6005),
.A2(n_5878),
.B1(n_5972),
.B2(n_5962),
.Y(n_6064)
);

AND2x4_ASAP7_75t_L g6065 ( 
.A(n_5995),
.B(n_5947),
.Y(n_6065)
);

AND2x2_ASAP7_75t_L g6066 ( 
.A(n_5998),
.B(n_5926),
.Y(n_6066)
);

OAI21xp33_ASAP7_75t_L g6067 ( 
.A1(n_6014),
.A2(n_5939),
.B(n_5969),
.Y(n_6067)
);

INVx1_ASAP7_75t_L g6068 ( 
.A(n_6026),
.Y(n_6068)
);

INVx4_ASAP7_75t_L g6069 ( 
.A(n_6051),
.Y(n_6069)
);

INVx2_ASAP7_75t_L g6070 ( 
.A(n_5987),
.Y(n_6070)
);

INVx1_ASAP7_75t_L g6071 ( 
.A(n_6030),
.Y(n_6071)
);

INVx5_ASAP7_75t_L g6072 ( 
.A(n_6051),
.Y(n_6072)
);

NOR2xp33_ASAP7_75t_L g6073 ( 
.A(n_6045),
.B(n_5967),
.Y(n_6073)
);

AND2x4_ASAP7_75t_L g6074 ( 
.A(n_6049),
.B(n_5907),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_6030),
.Y(n_6075)
);

OR2x2_ASAP7_75t_L g6076 ( 
.A(n_6032),
.B(n_5935),
.Y(n_6076)
);

AND2x2_ASAP7_75t_L g6077 ( 
.A(n_6050),
.B(n_5926),
.Y(n_6077)
);

INVx2_ASAP7_75t_L g6078 ( 
.A(n_6007),
.Y(n_6078)
);

INVx2_ASAP7_75t_L g6079 ( 
.A(n_6000),
.Y(n_6079)
);

OR2x2_ASAP7_75t_L g6080 ( 
.A(n_6036),
.B(n_5938),
.Y(n_6080)
);

AND2x2_ASAP7_75t_L g6081 ( 
.A(n_5984),
.B(n_5933),
.Y(n_6081)
);

BUFx6f_ASAP7_75t_L g6082 ( 
.A(n_6051),
.Y(n_6082)
);

BUFx3_ASAP7_75t_L g6083 ( 
.A(n_6015),
.Y(n_6083)
);

AND2x2_ASAP7_75t_L g6084 ( 
.A(n_6029),
.B(n_5936),
.Y(n_6084)
);

OR2x2_ASAP7_75t_L g6085 ( 
.A(n_6036),
.B(n_5960),
.Y(n_6085)
);

AND2x2_ASAP7_75t_L g6086 ( 
.A(n_6029),
.B(n_5994),
.Y(n_6086)
);

NAND2xp5_ASAP7_75t_L g6087 ( 
.A(n_5997),
.B(n_5915),
.Y(n_6087)
);

INVxp67_ASAP7_75t_L g6088 ( 
.A(n_6012),
.Y(n_6088)
);

AOI22xp33_ASAP7_75t_L g6089 ( 
.A1(n_6006),
.A2(n_5961),
.B1(n_5923),
.B2(n_5878),
.Y(n_6089)
);

AND2x4_ASAP7_75t_L g6090 ( 
.A(n_6001),
.B(n_5909),
.Y(n_6090)
);

INVxp67_ASAP7_75t_L g6091 ( 
.A(n_6012),
.Y(n_6091)
);

INVx4_ASAP7_75t_L g6092 ( 
.A(n_6051),
.Y(n_6092)
);

INVx3_ASAP7_75t_L g6093 ( 
.A(n_6038),
.Y(n_6093)
);

INVx1_ASAP7_75t_L g6094 ( 
.A(n_5989),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_6008),
.Y(n_6095)
);

INVx1_ASAP7_75t_L g6096 ( 
.A(n_6009),
.Y(n_6096)
);

AND2x2_ASAP7_75t_L g6097 ( 
.A(n_6003),
.B(n_5992),
.Y(n_6097)
);

INVx2_ASAP7_75t_L g6098 ( 
.A(n_6044),
.Y(n_6098)
);

HB1xp67_ASAP7_75t_L g6099 ( 
.A(n_5999),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_6046),
.B(n_5928),
.Y(n_6100)
);

AND2x2_ASAP7_75t_L g6101 ( 
.A(n_6035),
.B(n_5983),
.Y(n_6101)
);

INVx1_ASAP7_75t_SL g6102 ( 
.A(n_6004),
.Y(n_6102)
);

AND2x4_ASAP7_75t_L g6103 ( 
.A(n_6011),
.B(n_5913),
.Y(n_6103)
);

AND2x2_ASAP7_75t_L g6104 ( 
.A(n_6034),
.B(n_5917),
.Y(n_6104)
);

NAND2x1_ASAP7_75t_L g6105 ( 
.A(n_6011),
.B(n_5888),
.Y(n_6105)
);

AO21x2_ASAP7_75t_L g6106 ( 
.A1(n_6006),
.A2(n_5975),
.B(n_5955),
.Y(n_6106)
);

NAND2xp5_ASAP7_75t_L g6107 ( 
.A(n_6016),
.B(n_5959),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_6039),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_6043),
.Y(n_6109)
);

BUFx2_ASAP7_75t_L g6110 ( 
.A(n_6024),
.Y(n_6110)
);

INVx2_ASAP7_75t_L g6111 ( 
.A(n_6055),
.Y(n_6111)
);

INVx2_ASAP7_75t_L g6112 ( 
.A(n_6055),
.Y(n_6112)
);

OAI221xp5_ASAP7_75t_L g6113 ( 
.A1(n_6062),
.A2(n_6013),
.B1(n_6037),
.B2(n_5990),
.C(n_5884),
.Y(n_6113)
);

OR2x2_ASAP7_75t_L g6114 ( 
.A(n_6110),
.B(n_6019),
.Y(n_6114)
);

INVx1_ASAP7_75t_L g6115 ( 
.A(n_6063),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_6063),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_6058),
.Y(n_6117)
);

INVxp67_ASAP7_75t_L g6118 ( 
.A(n_6101),
.Y(n_6118)
);

AOI31xp33_ASAP7_75t_L g6119 ( 
.A1(n_6060),
.A2(n_6002),
.A3(n_6018),
.B(n_6022),
.Y(n_6119)
);

OAI33xp33_ASAP7_75t_L g6120 ( 
.A1(n_6064),
.A2(n_6047),
.A3(n_6027),
.B1(n_6025),
.B2(n_6033),
.B3(n_6028),
.Y(n_6120)
);

NAND3xp33_ASAP7_75t_L g6121 ( 
.A(n_6099),
.B(n_5982),
.C(n_6023),
.Y(n_6121)
);

AOI22xp33_ASAP7_75t_L g6122 ( 
.A1(n_6102),
.A2(n_6017),
.B1(n_6020),
.B2(n_6054),
.Y(n_6122)
);

NAND2xp5_ASAP7_75t_L g6123 ( 
.A(n_6104),
.B(n_6040),
.Y(n_6123)
);

OAI33xp33_ASAP7_75t_L g6124 ( 
.A1(n_6064),
.A2(n_6041),
.A3(n_5975),
.B1(n_5976),
.B2(n_5979),
.B3(n_5891),
.Y(n_6124)
);

AOI22xp33_ASAP7_75t_L g6125 ( 
.A1(n_6087),
.A2(n_6106),
.B1(n_6059),
.B2(n_6089),
.Y(n_6125)
);

CKINVDCx5p33_ASAP7_75t_R g6126 ( 
.A(n_6083),
.Y(n_6126)
);

AOI222xp33_ASAP7_75t_L g6127 ( 
.A1(n_6087),
.A2(n_5892),
.B1(n_5979),
.B2(n_5977),
.C1(n_6048),
.C2(n_5948),
.Y(n_6127)
);

AO21x2_ASAP7_75t_L g6128 ( 
.A1(n_6107),
.A2(n_5953),
.B(n_6052),
.Y(n_6128)
);

AO21x2_ASAP7_75t_L g6129 ( 
.A1(n_6107),
.A2(n_5890),
.B(n_6053),
.Y(n_6129)
);

OAI221xp5_ASAP7_75t_L g6130 ( 
.A1(n_6089),
.A2(n_5889),
.B1(n_5896),
.B2(n_6048),
.C(n_5905),
.Y(n_6130)
);

AOI22xp33_ASAP7_75t_L g6131 ( 
.A1(n_6059),
.A2(n_5929),
.B1(n_6040),
.B2(n_6042),
.Y(n_6131)
);

AND2x4_ASAP7_75t_L g6132 ( 
.A(n_6077),
.B(n_5945),
.Y(n_6132)
);

CKINVDCx5p33_ASAP7_75t_R g6133 ( 
.A(n_6057),
.Y(n_6133)
);

BUFx10_ASAP7_75t_L g6134 ( 
.A(n_6082),
.Y(n_6134)
);

AND2x2_ASAP7_75t_L g6135 ( 
.A(n_6086),
.B(n_5894),
.Y(n_6135)
);

BUFx3_ASAP7_75t_L g6136 ( 
.A(n_6103),
.Y(n_6136)
);

BUFx3_ASAP7_75t_L g6137 ( 
.A(n_6103),
.Y(n_6137)
);

AND2x2_ASAP7_75t_L g6138 ( 
.A(n_6090),
.B(n_337),
.Y(n_6138)
);

OR2x2_ASAP7_75t_L g6139 ( 
.A(n_6085),
.B(n_338),
.Y(n_6139)
);

OAI21x1_ASAP7_75t_L g6140 ( 
.A1(n_6105),
.A2(n_339),
.B(n_341),
.Y(n_6140)
);

INVxp67_ASAP7_75t_L g6141 ( 
.A(n_6097),
.Y(n_6141)
);

OAI33xp33_ASAP7_75t_L g6142 ( 
.A1(n_6068),
.A2(n_339),
.A3(n_343),
.B1(n_348),
.B2(n_350),
.B3(n_351),
.Y(n_6142)
);

NAND2x1_ASAP7_75t_L g6143 ( 
.A(n_6090),
.B(n_343),
.Y(n_6143)
);

NAND3xp33_ASAP7_75t_L g6144 ( 
.A(n_6071),
.B(n_350),
.C(n_351),
.Y(n_6144)
);

OAI211xp5_ASAP7_75t_L g6145 ( 
.A1(n_6067),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_6145)
);

AOI21xp5_ASAP7_75t_L g6146 ( 
.A1(n_6067),
.A2(n_1966),
.B(n_353),
.Y(n_6146)
);

OAI21xp5_ASAP7_75t_SL g6147 ( 
.A1(n_6075),
.A2(n_6091),
.B(n_6088),
.Y(n_6147)
);

NOR2x1_ASAP7_75t_L g6148 ( 
.A(n_6069),
.B(n_358),
.Y(n_6148)
);

AND2x2_ASAP7_75t_L g6149 ( 
.A(n_6065),
.B(n_359),
.Y(n_6149)
);

OAI221xp5_ASAP7_75t_L g6150 ( 
.A1(n_6073),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.C(n_365),
.Y(n_6150)
);

OR2x2_ASAP7_75t_L g6151 ( 
.A(n_6076),
.B(n_367),
.Y(n_6151)
);

NAND3xp33_ASAP7_75t_L g6152 ( 
.A(n_6088),
.B(n_369),
.C(n_370),
.Y(n_6152)
);

AOI22xp33_ASAP7_75t_L g6153 ( 
.A1(n_6098),
.A2(n_1422),
.B1(n_1443),
.B2(n_1280),
.Y(n_6153)
);

INVx1_ASAP7_75t_SL g6154 ( 
.A(n_6066),
.Y(n_6154)
);

BUFx2_ASAP7_75t_L g6155 ( 
.A(n_6081),
.Y(n_6155)
);

AND2x2_ASAP7_75t_L g6156 ( 
.A(n_6155),
.B(n_6084),
.Y(n_6156)
);

AND2x2_ASAP7_75t_L g6157 ( 
.A(n_6141),
.B(n_6079),
.Y(n_6157)
);

AND2x4_ASAP7_75t_L g6158 ( 
.A(n_6136),
.B(n_6072),
.Y(n_6158)
);

INVx2_ASAP7_75t_L g6159 ( 
.A(n_6129),
.Y(n_6159)
);

OR2x2_ASAP7_75t_L g6160 ( 
.A(n_6118),
.B(n_6080),
.Y(n_6160)
);

OR2x2_ASAP7_75t_L g6161 ( 
.A(n_6114),
.B(n_6056),
.Y(n_6161)
);

AND2x2_ASAP7_75t_L g6162 ( 
.A(n_6154),
.B(n_6061),
.Y(n_6162)
);

NAND2xp5_ASAP7_75t_SL g6163 ( 
.A(n_6119),
.B(n_6072),
.Y(n_6163)
);

AND2x4_ASAP7_75t_L g6164 ( 
.A(n_6137),
.B(n_6069),
.Y(n_6164)
);

AND2x2_ASAP7_75t_L g6165 ( 
.A(n_6111),
.B(n_6092),
.Y(n_6165)
);

AND2x2_ASAP7_75t_L g6166 ( 
.A(n_6112),
.B(n_6092),
.Y(n_6166)
);

INVxp67_ASAP7_75t_L g6167 ( 
.A(n_6148),
.Y(n_6167)
);

AND2x4_ASAP7_75t_SL g6168 ( 
.A(n_6134),
.B(n_6074),
.Y(n_6168)
);

INVxp67_ASAP7_75t_SL g6169 ( 
.A(n_6125),
.Y(n_6169)
);

INVx2_ASAP7_75t_L g6170 ( 
.A(n_6128),
.Y(n_6170)
);

AND2x2_ASAP7_75t_L g6171 ( 
.A(n_6135),
.B(n_6100),
.Y(n_6171)
);

INVx1_ASAP7_75t_L g6172 ( 
.A(n_6139),
.Y(n_6172)
);

INVx1_ASAP7_75t_L g6173 ( 
.A(n_6123),
.Y(n_6173)
);

INVxp67_ASAP7_75t_L g6174 ( 
.A(n_6149),
.Y(n_6174)
);

INVx2_ASAP7_75t_L g6175 ( 
.A(n_6134),
.Y(n_6175)
);

INVx1_ASAP7_75t_L g6176 ( 
.A(n_6151),
.Y(n_6176)
);

AND2x2_ASAP7_75t_L g6177 ( 
.A(n_6117),
.B(n_6094),
.Y(n_6177)
);

NOR2xp33_ASAP7_75t_L g6178 ( 
.A(n_6121),
.B(n_6093),
.Y(n_6178)
);

AND2x2_ASAP7_75t_L g6179 ( 
.A(n_6126),
.B(n_6095),
.Y(n_6179)
);

INVx2_ASAP7_75t_L g6180 ( 
.A(n_6143),
.Y(n_6180)
);

INVx2_ASAP7_75t_L g6181 ( 
.A(n_6132),
.Y(n_6181)
);

INVx1_ASAP7_75t_L g6182 ( 
.A(n_6115),
.Y(n_6182)
);

INVx3_ASAP7_75t_L g6183 ( 
.A(n_6132),
.Y(n_6183)
);

AND2x2_ASAP7_75t_L g6184 ( 
.A(n_6133),
.B(n_6096),
.Y(n_6184)
);

NAND2xp5_ASAP7_75t_L g6185 ( 
.A(n_6138),
.B(n_6070),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_6116),
.Y(n_6186)
);

INVx3_ASAP7_75t_L g6187 ( 
.A(n_6140),
.Y(n_6187)
);

INVxp67_ASAP7_75t_SL g6188 ( 
.A(n_6152),
.Y(n_6188)
);

AND2x2_ASAP7_75t_L g6189 ( 
.A(n_6156),
.B(n_6171),
.Y(n_6189)
);

AND2x2_ASAP7_75t_L g6190 ( 
.A(n_6162),
.B(n_6147),
.Y(n_6190)
);

INVx1_ASAP7_75t_L g6191 ( 
.A(n_6183),
.Y(n_6191)
);

AND2x4_ASAP7_75t_L g6192 ( 
.A(n_6168),
.B(n_6078),
.Y(n_6192)
);

INVx1_ASAP7_75t_L g6193 ( 
.A(n_6159),
.Y(n_6193)
);

AOI22xp33_ASAP7_75t_SL g6194 ( 
.A1(n_6169),
.A2(n_6113),
.B1(n_6130),
.B2(n_6145),
.Y(n_6194)
);

AND2x2_ASAP7_75t_L g6195 ( 
.A(n_6157),
.B(n_6146),
.Y(n_6195)
);

NAND2xp5_ASAP7_75t_L g6196 ( 
.A(n_6178),
.B(n_6131),
.Y(n_6196)
);

NAND2xp5_ASAP7_75t_L g6197 ( 
.A(n_6178),
.B(n_6127),
.Y(n_6197)
);

INVx1_ASAP7_75t_L g6198 ( 
.A(n_6170),
.Y(n_6198)
);

INVx2_ASAP7_75t_L g6199 ( 
.A(n_6158),
.Y(n_6199)
);

AND2x2_ASAP7_75t_L g6200 ( 
.A(n_6184),
.B(n_6122),
.Y(n_6200)
);

AND2x4_ASAP7_75t_L g6201 ( 
.A(n_6181),
.B(n_6164),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_6170),
.Y(n_6202)
);

OR2x2_ASAP7_75t_L g6203 ( 
.A(n_6161),
.B(n_6144),
.Y(n_6203)
);

AND2x4_ASAP7_75t_L g6204 ( 
.A(n_6164),
.B(n_6180),
.Y(n_6204)
);

NOR2x1_ASAP7_75t_L g6205 ( 
.A(n_6163),
.B(n_6150),
.Y(n_6205)
);

NAND2xp5_ASAP7_75t_L g6206 ( 
.A(n_6188),
.B(n_6108),
.Y(n_6206)
);

NOR2xp33_ASAP7_75t_L g6207 ( 
.A(n_6167),
.B(n_6174),
.Y(n_6207)
);

INVx2_ASAP7_75t_L g6208 ( 
.A(n_6180),
.Y(n_6208)
);

INVx1_ASAP7_75t_L g6209 ( 
.A(n_6160),
.Y(n_6209)
);

AND2x4_ASAP7_75t_L g6210 ( 
.A(n_6165),
.B(n_6109),
.Y(n_6210)
);

INVx2_ASAP7_75t_L g6211 ( 
.A(n_6187),
.Y(n_6211)
);

NAND2xp5_ASAP7_75t_L g6212 ( 
.A(n_6189),
.B(n_6187),
.Y(n_6212)
);

AND2x4_ASAP7_75t_SL g6213 ( 
.A(n_6201),
.B(n_6166),
.Y(n_6213)
);

AND2x2_ASAP7_75t_L g6214 ( 
.A(n_6190),
.B(n_6173),
.Y(n_6214)
);

BUFx2_ASAP7_75t_L g6215 ( 
.A(n_6201),
.Y(n_6215)
);

AND2x2_ASAP7_75t_L g6216 ( 
.A(n_6200),
.B(n_6179),
.Y(n_6216)
);

INVx1_ASAP7_75t_L g6217 ( 
.A(n_6211),
.Y(n_6217)
);

NAND2xp5_ASAP7_75t_L g6218 ( 
.A(n_6204),
.B(n_6176),
.Y(n_6218)
);

AND2x4_ASAP7_75t_L g6219 ( 
.A(n_6192),
.B(n_6177),
.Y(n_6219)
);

INVx1_ASAP7_75t_L g6220 ( 
.A(n_6191),
.Y(n_6220)
);

OR2x2_ASAP7_75t_L g6221 ( 
.A(n_6203),
.B(n_6185),
.Y(n_6221)
);

XNOR2xp5_ASAP7_75t_L g6222 ( 
.A(n_6194),
.B(n_6172),
.Y(n_6222)
);

AOI22xp5_ASAP7_75t_L g6223 ( 
.A1(n_6196),
.A2(n_6124),
.B1(n_6120),
.B2(n_6142),
.Y(n_6223)
);

INVxp67_ASAP7_75t_L g6224 ( 
.A(n_6207),
.Y(n_6224)
);

NAND4xp75_ASAP7_75t_L g6225 ( 
.A(n_6205),
.B(n_6186),
.C(n_6182),
.D(n_6175),
.Y(n_6225)
);

INVx3_ASAP7_75t_L g6226 ( 
.A(n_6210),
.Y(n_6226)
);

INVx2_ASAP7_75t_L g6227 ( 
.A(n_6210),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_L g6228 ( 
.A(n_6215),
.B(n_6199),
.Y(n_6228)
);

OAI22xp33_ASAP7_75t_L g6229 ( 
.A1(n_6223),
.A2(n_6197),
.B1(n_6206),
.B2(n_6208),
.Y(n_6229)
);

CKINVDCx5p33_ASAP7_75t_R g6230 ( 
.A(n_6213),
.Y(n_6230)
);

NAND2xp5_ASAP7_75t_L g6231 ( 
.A(n_6219),
.B(n_6195),
.Y(n_6231)
);

NAND2xp5_ASAP7_75t_L g6232 ( 
.A(n_6226),
.B(n_6209),
.Y(n_6232)
);

AND2x2_ASAP7_75t_L g6233 ( 
.A(n_6216),
.B(n_6202),
.Y(n_6233)
);

NAND2xp33_ASAP7_75t_SL g6234 ( 
.A(n_6212),
.B(n_6198),
.Y(n_6234)
);

AND2x2_ASAP7_75t_L g6235 ( 
.A(n_6214),
.B(n_6193),
.Y(n_6235)
);

AND2x4_ASAP7_75t_L g6236 ( 
.A(n_6227),
.B(n_6153),
.Y(n_6236)
);

NAND2xp5_ASAP7_75t_L g6237 ( 
.A(n_6233),
.B(n_6222),
.Y(n_6237)
);

AND2x2_ASAP7_75t_L g6238 ( 
.A(n_6235),
.B(n_6230),
.Y(n_6238)
);

INVx1_ASAP7_75t_L g6239 ( 
.A(n_6228),
.Y(n_6239)
);

OR2x2_ASAP7_75t_L g6240 ( 
.A(n_6231),
.B(n_6218),
.Y(n_6240)
);

OAI33xp33_ASAP7_75t_L g6241 ( 
.A1(n_6229),
.A2(n_6217),
.A3(n_6220),
.B1(n_6224),
.B2(n_6221),
.B3(n_6225),
.Y(n_6241)
);

INVx1_ASAP7_75t_L g6242 ( 
.A(n_6232),
.Y(n_6242)
);

AND2x2_ASAP7_75t_L g6243 ( 
.A(n_6238),
.B(n_6236),
.Y(n_6243)
);

OR2x2_ASAP7_75t_L g6244 ( 
.A(n_6237),
.B(n_6234),
.Y(n_6244)
);

INVx1_ASAP7_75t_L g6245 ( 
.A(n_6240),
.Y(n_6245)
);

NAND2xp5_ASAP7_75t_L g6246 ( 
.A(n_6239),
.B(n_394),
.Y(n_6246)
);

BUFx3_ASAP7_75t_L g6247 ( 
.A(n_6242),
.Y(n_6247)
);

OR2x2_ASAP7_75t_L g6248 ( 
.A(n_6244),
.B(n_6241),
.Y(n_6248)
);

INVx1_ASAP7_75t_L g6249 ( 
.A(n_6245),
.Y(n_6249)
);

INVx2_ASAP7_75t_L g6250 ( 
.A(n_6247),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_6246),
.Y(n_6251)
);

INVx2_ASAP7_75t_L g6252 ( 
.A(n_6243),
.Y(n_6252)
);

AND2x4_ASAP7_75t_L g6253 ( 
.A(n_6243),
.B(n_405),
.Y(n_6253)
);

INVx1_ASAP7_75t_SL g6254 ( 
.A(n_6244),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_6252),
.Y(n_6255)
);

OAI21xp33_ASAP7_75t_SL g6256 ( 
.A1(n_6254),
.A2(n_406),
.B(n_407),
.Y(n_6256)
);

OR2x2_ASAP7_75t_L g6257 ( 
.A(n_6248),
.B(n_408),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_6250),
.B(n_409),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_6253),
.Y(n_6259)
);

INVx1_ASAP7_75t_L g6260 ( 
.A(n_6249),
.Y(n_6260)
);

NAND2xp5_ASAP7_75t_L g6261 ( 
.A(n_6251),
.B(n_416),
.Y(n_6261)
);

OR2x2_ASAP7_75t_L g6262 ( 
.A(n_6257),
.B(n_426),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_6259),
.Y(n_6263)
);

NOR2x1_ASAP7_75t_L g6264 ( 
.A(n_6260),
.B(n_427),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_6258),
.Y(n_6265)
);

HB1xp67_ASAP7_75t_L g6266 ( 
.A(n_6256),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_6261),
.Y(n_6267)
);

AND2x4_ASAP7_75t_L g6268 ( 
.A(n_6255),
.B(n_439),
.Y(n_6268)
);

OR2x2_ASAP7_75t_L g6269 ( 
.A(n_6266),
.B(n_440),
.Y(n_6269)
);

INVx1_ASAP7_75t_L g6270 ( 
.A(n_6264),
.Y(n_6270)
);

INVx2_ASAP7_75t_SL g6271 ( 
.A(n_6268),
.Y(n_6271)
);

INVx2_ASAP7_75t_SL g6272 ( 
.A(n_6268),
.Y(n_6272)
);

CKINVDCx16_ASAP7_75t_R g6273 ( 
.A(n_6265),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_6262),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_6263),
.Y(n_6275)
);

INVx1_ASAP7_75t_SL g6276 ( 
.A(n_6269),
.Y(n_6276)
);

INVx2_ASAP7_75t_L g6277 ( 
.A(n_6271),
.Y(n_6277)
);

NOR2x1_ASAP7_75t_L g6278 ( 
.A(n_6275),
.B(n_6267),
.Y(n_6278)
);

INVx8_ASAP7_75t_L g6279 ( 
.A(n_6273),
.Y(n_6279)
);

INVx2_ASAP7_75t_L g6280 ( 
.A(n_6272),
.Y(n_6280)
);

INVx1_ASAP7_75t_L g6281 ( 
.A(n_6270),
.Y(n_6281)
);

INVxp67_ASAP7_75t_L g6282 ( 
.A(n_6274),
.Y(n_6282)
);

INVx1_ASAP7_75t_L g6283 ( 
.A(n_6279),
.Y(n_6283)
);

O2A1O1Ixp33_ASAP7_75t_L g6284 ( 
.A1(n_6282),
.A2(n_450),
.B(n_454),
.C(n_455),
.Y(n_6284)
);

HB1xp67_ASAP7_75t_L g6285 ( 
.A(n_6278),
.Y(n_6285)
);

AOI22x1_ASAP7_75t_L g6286 ( 
.A1(n_6281),
.A2(n_455),
.B1(n_456),
.B2(n_457),
.Y(n_6286)
);

HB1xp67_ASAP7_75t_L g6287 ( 
.A(n_6277),
.Y(n_6287)
);

O2A1O1Ixp33_ASAP7_75t_L g6288 ( 
.A1(n_6280),
.A2(n_468),
.B(n_469),
.C(n_470),
.Y(n_6288)
);

OAI22x1_ASAP7_75t_L g6289 ( 
.A1(n_6276),
.A2(n_474),
.B1(n_475),
.B2(n_476),
.Y(n_6289)
);

OAI21xp33_ASAP7_75t_L g6290 ( 
.A1(n_6287),
.A2(n_482),
.B(n_483),
.Y(n_6290)
);

AOI221xp5_ASAP7_75t_L g6291 ( 
.A1(n_6283),
.A2(n_484),
.B1(n_485),
.B2(n_488),
.C(n_489),
.Y(n_6291)
);

A2O1A1Ixp33_ASAP7_75t_L g6292 ( 
.A1(n_6284),
.A2(n_498),
.B(n_499),
.C(n_502),
.Y(n_6292)
);

AOI221x1_ASAP7_75t_L g6293 ( 
.A1(n_6289),
.A2(n_503),
.B1(n_505),
.B2(n_506),
.C(n_507),
.Y(n_6293)
);

NAND3xp33_ASAP7_75t_L g6294 ( 
.A(n_6286),
.B(n_505),
.C(n_506),
.Y(n_6294)
);

AOI221xp5_ASAP7_75t_L g6295 ( 
.A1(n_6288),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.C(n_512),
.Y(n_6295)
);

AOI221xp5_ASAP7_75t_L g6296 ( 
.A1(n_6285),
.A2(n_515),
.B1(n_516),
.B2(n_517),
.C(n_518),
.Y(n_6296)
);

NAND4xp25_ASAP7_75t_L g6297 ( 
.A(n_6293),
.B(n_527),
.C(n_529),
.D(n_530),
.Y(n_6297)
);

AND2x4_ASAP7_75t_L g6298 ( 
.A(n_6294),
.B(n_6292),
.Y(n_6298)
);

AOI221xp5_ASAP7_75t_L g6299 ( 
.A1(n_6297),
.A2(n_6295),
.B1(n_6290),
.B2(n_6296),
.C(n_6291),
.Y(n_6299)
);

NAND2xp5_ASAP7_75t_L g6300 ( 
.A(n_6299),
.B(n_6298),
.Y(n_6300)
);

INVx1_ASAP7_75t_L g6301 ( 
.A(n_6300),
.Y(n_6301)
);

BUFx2_ASAP7_75t_L g6302 ( 
.A(n_6301),
.Y(n_6302)
);

HB1xp67_ASAP7_75t_L g6303 ( 
.A(n_6302),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_6303),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6304),
.Y(n_6305)
);

AOI22xp5_ASAP7_75t_L g6306 ( 
.A1(n_6304),
.A2(n_1463),
.B1(n_550),
.B2(n_552),
.Y(n_6306)
);

AO22x1_ASAP7_75t_L g6307 ( 
.A1(n_6304),
.A2(n_555),
.B1(n_556),
.B2(n_557),
.Y(n_6307)
);

OAI322xp33_ASAP7_75t_L g6308 ( 
.A1(n_6305),
.A2(n_556),
.A3(n_557),
.B1(n_558),
.B2(n_559),
.C1(n_560),
.C2(n_563),
.Y(n_6308)
);

AOI222xp33_ASAP7_75t_L g6309 ( 
.A1(n_6307),
.A2(n_566),
.B1(n_568),
.B2(n_569),
.C1(n_570),
.C2(n_571),
.Y(n_6309)
);

NAND3xp33_ASAP7_75t_SL g6310 ( 
.A(n_6306),
.B(n_573),
.C(n_576),
.Y(n_6310)
);

INVx1_ASAP7_75t_L g6311 ( 
.A(n_6310),
.Y(n_6311)
);

AOI22xp33_ASAP7_75t_L g6312 ( 
.A1(n_6309),
.A2(n_578),
.B1(n_579),
.B2(n_580),
.Y(n_6312)
);

AOI22xp33_ASAP7_75t_L g6313 ( 
.A1(n_6308),
.A2(n_581),
.B1(n_582),
.B2(n_583),
.Y(n_6313)
);

INVx1_ASAP7_75t_L g6314 ( 
.A(n_6311),
.Y(n_6314)
);

AND2x2_ASAP7_75t_L g6315 ( 
.A(n_6313),
.B(n_584),
.Y(n_6315)
);

BUFx2_ASAP7_75t_L g6316 ( 
.A(n_6314),
.Y(n_6316)
);

OAI22x1_ASAP7_75t_L g6317 ( 
.A1(n_6316),
.A2(n_6315),
.B1(n_6312),
.B2(n_585),
.Y(n_6317)
);

INVx1_ASAP7_75t_L g6318 ( 
.A(n_6317),
.Y(n_6318)
);

AOI22xp5_ASAP7_75t_L g6319 ( 
.A1(n_6318),
.A2(n_2002),
.B1(n_2055),
.B2(n_2053),
.Y(n_6319)
);

OAI21xp5_ASAP7_75t_L g6320 ( 
.A1(n_6319),
.A2(n_591),
.B(n_594),
.Y(n_6320)
);

AOI322xp5_ASAP7_75t_L g6321 ( 
.A1(n_6320),
.A2(n_595),
.A3(n_596),
.B1(n_598),
.B2(n_599),
.C1(n_600),
.C2(n_601),
.Y(n_6321)
);

INVx2_ASAP7_75t_L g6322 ( 
.A(n_6321),
.Y(n_6322)
);

AOI221xp5_ASAP7_75t_L g6323 ( 
.A1(n_6322),
.A2(n_2002),
.B1(n_1985),
.B2(n_1986),
.C(n_1989),
.Y(n_6323)
);

AOI21xp5_ASAP7_75t_L g6324 ( 
.A1(n_6323),
.A2(n_1981),
.B(n_1985),
.Y(n_6324)
);

AOI211xp5_ASAP7_75t_L g6325 ( 
.A1(n_6324),
.A2(n_1981),
.B(n_1986),
.C(n_1989),
.Y(n_6325)
);


endmodule