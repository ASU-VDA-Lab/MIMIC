module fake_ariane_1084_n_5396 (n_913, n_589, n_1174, n_691, n_423, n_603, n_373, n_1250, n_1169, n_789, n_850, n_610, n_245, n_96, n_319, n_49, n_690, n_416, n_1109, n_525, n_187, n_1238, n_817, n_924, n_781, n_189, n_717, n_72, n_952, n_864, n_1096, n_57, n_117, n_524, n_1214, n_634, n_1246, n_1138, n_214, n_764, n_462, n_1196, n_1181, n_32, n_410, n_1187, n_1131, n_1225, n_737, n_137, n_232, n_52, n_568, n_1088, n_77, n_766, n_377, n_520, n_870, n_279, n_945, n_958, n_813, n_419, n_146, n_270, n_338, n_995, n_285, n_1184, n_202, n_500, n_665, n_754, n_903, n_871, n_1073, n_239, n_402, n_54, n_829, n_1062, n_339, n_738, n_672, n_740, n_167, n_1018, n_69, n_259, n_953, n_143, n_1224, n_625, n_557, n_1107, n_989, n_242, n_645, n_331, n_559, n_267, n_495, n_350, n_381, n_795, n_721, n_1084, n_200, n_1241, n_821, n_561, n_770, n_507, n_486, n_901, n_569, n_1145, n_971, n_787, n_31, n_1195, n_518, n_1207, n_222, n_786, n_868, n_884, n_1034, n_1085, n_277, n_432, n_293, n_823, n_620, n_93, n_1074, n_859, n_108, n_587, n_693, n_863, n_303, n_1254, n_929, n_206, n_352, n_899, n_611, n_238, n_365, n_1013, n_136, n_334, n_192, n_661, n_300, n_533, n_104, n_438, n_16, n_440, n_273, n_1230, n_612, n_333, n_376, n_512, n_579, n_844, n_1012, n_1267, n_149, n_1213, n_237, n_780, n_1021, n_491, n_1142, n_1140, n_705, n_570, n_260, n_942, n_7, n_461, n_1121, n_209, n_490, n_17, n_225, n_1006, n_575, n_546, n_503, n_1112, n_700, n_1159, n_772, n_1216, n_1245, n_676, n_42, n_680, n_287, n_302, n_380, n_94, n_4, n_249, n_1108, n_355, n_212, n_65, n_123, n_444, n_851, n_257, n_652, n_475, n_135, n_947, n_930, n_1260, n_1179, n_468, n_102, n_182, n_696, n_482, n_798, n_577, n_407, n_27, n_916, n_912, n_460, n_366, n_762, n_1253, n_555, n_804, n_966, n_992, n_955, n_1182, n_794, n_78, n_514, n_418, n_513, n_288, n_179, n_1178, n_1026, n_306, n_92, n_203, n_436, n_150, n_324, n_669, n_931, n_619, n_337, n_437, n_111, n_21, n_274, n_967, n_1083, n_746, n_292, n_1079, n_615, n_1139, n_76, n_517, n_0, n_824, n_428, n_159, n_892, n_959, n_30, n_1101, n_563, n_144, n_990, n_867, n_1226, n_944, n_749, n_815, n_542, n_470, n_1240, n_1087, n_632, n_477, n_650, n_425, n_1155, n_1071, n_712, n_976, n_909, n_767, n_964, n_382, n_489, n_80, n_251, n_974, n_506, n_799, n_1147, n_397, n_471, n_351, n_965, n_155, n_934, n_1220, n_356, n_698, n_124, n_307, n_1209, n_1020, n_646, n_34, n_404, n_172, n_1058, n_347, n_1042, n_183, n_1234, n_479, n_299, n_836, n_564, n_133, n_66, n_205, n_1029, n_1247, n_760, n_522, n_20, n_367, n_1111, n_970, n_713, n_1255, n_598, n_345, n_1237, n_927, n_261, n_1095, n_370, n_706, n_286, n_776, n_424, n_85, n_130, n_466, n_1263, n_346, n_348, n_552, n_670, n_379, n_138, n_162, n_264, n_441, n_1032, n_1217, n_637, n_73, n_327, n_1259, n_1177, n_1231, n_980, n_905, n_207, n_720, n_926, n_41, n_194, n_1163, n_186, n_145, n_59, n_1173, n_1068, n_1198, n_487, n_90, n_855, n_158, n_808, n_553, n_814, n_578, n_405, n_120, n_320, n_1134, n_647, n_481, n_600, n_1053, n_529, n_502, n_218, n_247, n_1105, n_547, n_439, n_604, n_677, n_478, n_703, n_1061, n_326, n_681, n_227, n_874, n_707, n_11, n_129, n_126, n_983, n_590, n_699, n_727, n_301, n_545, n_1015, n_1162, n_536, n_325, n_688, n_636, n_427, n_1098, n_442, n_777, n_1080, n_920, n_1086, n_1092, n_986, n_1104, n_729, n_887, n_1122, n_1205, n_163, n_1132, n_390, n_1156, n_501, n_314, n_1120, n_1202, n_627, n_1188, n_233, n_957, n_388, n_1242, n_1218, n_221, n_321, n_86, n_861, n_877, n_1119, n_616, n_1055, n_1189, n_1089, n_281, n_262, n_735, n_297, n_1005, n_527, n_46, n_84, n_845, n_888, n_178, n_551, n_417, n_70, n_343, n_1222, n_582, n_755, n_1097, n_1219, n_710, n_534, n_1239, n_278, n_560, n_890, n_842, n_148, n_451, n_745, n_61, n_742, n_1081, n_1266, n_769, n_13, n_476, n_832, n_55, n_535, n_744, n_982, n_915, n_215, n_1075, n_454, n_298, n_1227, n_655, n_403, n_1007, n_657, n_837, n_812, n_606, n_951, n_862, n_659, n_509, n_666, n_430, n_1206, n_722, n_1171, n_1030, n_785, n_999, n_456, n_852, n_704, n_1060, n_1044, n_521, n_873, n_1243, n_342, n_358, n_608, n_1037, n_317, n_134, n_1257, n_1078, n_266, n_157, n_1161, n_811, n_624, n_791, n_876, n_618, n_1191, n_736, n_1025, n_1215, n_241, n_687, n_797, n_480, n_211, n_642, n_97, n_408, n_595, n_602, n_592, n_854, n_393, n_474, n_805, n_295, n_190, n_1072, n_695, n_64, n_180, n_730, n_386, n_516, n_1137, n_1258, n_197, n_640, n_463, n_943, n_1118, n_678, n_651, n_961, n_469, n_1046, n_726, n_1123, n_878, n_771, n_752, n_71, n_985, n_421, n_906, n_1180, n_283, n_806, n_649, n_374, n_643, n_226, n_682, n_36, n_819, n_586, n_686, n_605, n_1154, n_584, n_1130, n_349, n_756, n_1016, n_1149, n_979, n_2, n_897, n_949, n_515, n_807, n_891, n_885, n_198, n_1208, n_396, n_802, n_23, n_1151, n_554, n_960, n_1256, n_87, n_714, n_790, n_354, n_140, n_725, n_151, n_28, n_1009, n_230, n_1133, n_154, n_883, n_142, n_473, n_801, n_818, n_779, n_594, n_35, n_1052, n_272, n_833, n_879, n_1117, n_38, n_422, n_1269, n_597, n_75, n_1047, n_95, n_1050, n_566, n_152, n_169, n_106, n_1201, n_173, n_858, n_1185, n_335, n_1035, n_1143, n_344, n_426, n_433, n_398, n_62, n_210, n_1090, n_166, n_253, n_928, n_1153, n_271, n_465, n_825, n_1103, n_732, n_1192, n_128, n_224, n_82, n_894, n_420, n_562, n_748, n_510, n_1045, n_256, n_1160, n_1023, n_988, n_330, n_914, n_400, n_689, n_1116, n_282, n_328, n_368, n_467, n_644, n_1197, n_276, n_497, n_1165, n_168, n_81, n_538, n_576, n_843, n_511, n_455, n_429, n_588, n_638, n_1128, n_1048, n_775, n_667, n_1049, n_14, n_869, n_141, n_846, n_305, n_312, n_56, n_60, n_728, n_413, n_715, n_889, n_1066, n_935, n_685, n_911, n_361, n_89, n_623, n_1065, n_453, n_74, n_810, n_19, n_40, n_181, n_617, n_543, n_236, n_601, n_683, n_565, n_628, n_743, n_1194, n_907, n_660, n_464, n_962, n_941, n_1210, n_847, n_747, n_1135, n_918, n_107, n_639, n_452, n_673, n_1038, n_414, n_571, n_6, n_284, n_593, n_1164, n_37, n_58, n_609, n_1193, n_613, n_1022, n_1033, n_409, n_171, n_519, n_384, n_1166, n_1056, n_526, n_1040, n_674, n_1158, n_316, n_125, n_820, n_43, n_872, n_254, n_1157, n_234, n_848, n_280, n_629, n_161, n_532, n_763, n_99, n_540, n_216, n_692, n_5, n_984, n_223, n_750, n_834, n_800, n_395, n_621, n_213, n_67, n_1014, n_724, n_493, n_114, n_1100, n_585, n_875, n_827, n_697, n_622, n_296, n_880, n_793, n_1175, n_132, n_751, n_1027, n_1070, n_739, n_1028, n_1221, n_530, n_792, n_1262, n_580, n_494, n_434, n_975, n_229, n_394, n_923, n_1124, n_932, n_1183, n_981, n_1110, n_243, n_185, n_1204, n_994, n_973, n_268, n_972, n_164, n_184, n_856, n_1248, n_1176, n_1054, n_508, n_118, n_121, n_353, n_1057, n_191, n_978, n_1011, n_828, n_322, n_558, n_116, n_39, n_653, n_783, n_556, n_1127, n_170, n_160, n_119, n_1008, n_332, n_581, n_294, n_1024, n_830, n_176, n_987, n_936, n_541, n_499, n_788, n_12, n_908, n_1036, n_341, n_1270, n_109, n_1167, n_549, n_591, n_969, n_919, n_50, n_318, n_103, n_244, n_679, n_220, n_663, n_443, n_528, n_1200, n_387, n_406, n_826, n_139, n_391, n_940, n_1077, n_607, n_956, n_445, n_765, n_122, n_1268, n_385, n_917, n_1271, n_372, n_15, n_631, n_399, n_1170, n_1261, n_702, n_857, n_898, n_363, n_968, n_1067, n_1235, n_1064, n_633, n_900, n_1093, n_193, n_733, n_761, n_731, n_336, n_315, n_311, n_8, n_668, n_758, n_1106, n_47, n_153, n_18, n_648, n_784, n_269, n_816, n_835, n_446, n_1076, n_753, n_701, n_1003, n_1125, n_309, n_115, n_401, n_485, n_504, n_483, n_435, n_1141, n_291, n_822, n_1094, n_840, n_1099, n_839, n_79, n_3, n_759, n_567, n_91, n_240, n_369, n_44, n_1172, n_614, n_1212, n_831, n_778, n_48, n_188, n_323, n_550, n_997, n_635, n_694, n_1113, n_248, n_1152, n_921, n_1236, n_228, n_1265, n_671, n_1, n_1148, n_654, n_488, n_904, n_505, n_88, n_498, n_1059, n_684, n_1039, n_539, n_1150, n_977, n_449, n_392, n_459, n_1136, n_458, n_1190, n_1144, n_383, n_838, n_175, n_950, n_1017, n_711, n_734, n_723, n_658, n_630, n_53, n_362, n_310, n_709, n_24, n_809, n_235, n_881, n_1019, n_662, n_641, n_910, n_290, n_741, n_939, n_371, n_199, n_217, n_1114, n_708, n_308, n_1223, n_201, n_572, n_1199, n_865, n_10, n_1041, n_993, n_948, n_922, n_1004, n_448, n_860, n_1043, n_255, n_450, n_896, n_902, n_1031, n_853, n_716, n_196, n_774, n_933, n_596, n_954, n_1168, n_219, n_231, n_656, n_492, n_574, n_252, n_664, n_1229, n_68, n_415, n_63, n_544, n_1186, n_599, n_768, n_1091, n_537, n_1063, n_25, n_991, n_83, n_389, n_1126, n_195, n_938, n_895, n_110, n_304, n_583, n_1000, n_313, n_626, n_378, n_98, n_946, n_757, n_375, n_113, n_33, n_1146, n_1203, n_998, n_472, n_937, n_265, n_208, n_156, n_174, n_275, n_100, n_147, n_204, n_1232, n_996, n_1211, n_963, n_1264, n_51, n_1082, n_496, n_866, n_26, n_246, n_925, n_1001, n_1115, n_1002, n_105, n_1051, n_719, n_131, n_263, n_1102, n_360, n_1129, n_1252, n_250, n_773, n_165, n_1010, n_882, n_1249, n_101, n_803, n_329, n_718, n_340, n_289, n_9, n_112, n_45, n_548, n_523, n_457, n_177, n_782, n_364, n_258, n_431, n_1228, n_1244, n_411, n_484, n_849, n_22, n_29, n_357, n_412, n_1251, n_447, n_1233, n_893, n_841, n_886, n_1069, n_359, n_573, n_796, n_127, n_531, n_675, n_5396);

input n_913;
input n_589;
input n_1174;
input n_691;
input n_423;
input n_603;
input n_373;
input n_1250;
input n_1169;
input n_789;
input n_850;
input n_610;
input n_245;
input n_96;
input n_319;
input n_49;
input n_690;
input n_416;
input n_1109;
input n_525;
input n_187;
input n_1238;
input n_817;
input n_924;
input n_781;
input n_189;
input n_717;
input n_72;
input n_952;
input n_864;
input n_1096;
input n_57;
input n_117;
input n_524;
input n_1214;
input n_634;
input n_1246;
input n_1138;
input n_214;
input n_764;
input n_462;
input n_1196;
input n_1181;
input n_32;
input n_410;
input n_1187;
input n_1131;
input n_1225;
input n_737;
input n_137;
input n_232;
input n_52;
input n_568;
input n_1088;
input n_77;
input n_766;
input n_377;
input n_520;
input n_870;
input n_279;
input n_945;
input n_958;
input n_813;
input n_419;
input n_146;
input n_270;
input n_338;
input n_995;
input n_285;
input n_1184;
input n_202;
input n_500;
input n_665;
input n_754;
input n_903;
input n_871;
input n_1073;
input n_239;
input n_402;
input n_54;
input n_829;
input n_1062;
input n_339;
input n_738;
input n_672;
input n_740;
input n_167;
input n_1018;
input n_69;
input n_259;
input n_953;
input n_143;
input n_1224;
input n_625;
input n_557;
input n_1107;
input n_989;
input n_242;
input n_645;
input n_331;
input n_559;
input n_267;
input n_495;
input n_350;
input n_381;
input n_795;
input n_721;
input n_1084;
input n_200;
input n_1241;
input n_821;
input n_561;
input n_770;
input n_507;
input n_486;
input n_901;
input n_569;
input n_1145;
input n_971;
input n_787;
input n_31;
input n_1195;
input n_518;
input n_1207;
input n_222;
input n_786;
input n_868;
input n_884;
input n_1034;
input n_1085;
input n_277;
input n_432;
input n_293;
input n_823;
input n_620;
input n_93;
input n_1074;
input n_859;
input n_108;
input n_587;
input n_693;
input n_863;
input n_303;
input n_1254;
input n_929;
input n_206;
input n_352;
input n_899;
input n_611;
input n_238;
input n_365;
input n_1013;
input n_136;
input n_334;
input n_192;
input n_661;
input n_300;
input n_533;
input n_104;
input n_438;
input n_16;
input n_440;
input n_273;
input n_1230;
input n_612;
input n_333;
input n_376;
input n_512;
input n_579;
input n_844;
input n_1012;
input n_1267;
input n_149;
input n_1213;
input n_237;
input n_780;
input n_1021;
input n_491;
input n_1142;
input n_1140;
input n_705;
input n_570;
input n_260;
input n_942;
input n_7;
input n_461;
input n_1121;
input n_209;
input n_490;
input n_17;
input n_225;
input n_1006;
input n_575;
input n_546;
input n_503;
input n_1112;
input n_700;
input n_1159;
input n_772;
input n_1216;
input n_1245;
input n_676;
input n_42;
input n_680;
input n_287;
input n_302;
input n_380;
input n_94;
input n_4;
input n_249;
input n_1108;
input n_355;
input n_212;
input n_65;
input n_123;
input n_444;
input n_851;
input n_257;
input n_652;
input n_475;
input n_135;
input n_947;
input n_930;
input n_1260;
input n_1179;
input n_468;
input n_102;
input n_182;
input n_696;
input n_482;
input n_798;
input n_577;
input n_407;
input n_27;
input n_916;
input n_912;
input n_460;
input n_366;
input n_762;
input n_1253;
input n_555;
input n_804;
input n_966;
input n_992;
input n_955;
input n_1182;
input n_794;
input n_78;
input n_514;
input n_418;
input n_513;
input n_288;
input n_179;
input n_1178;
input n_1026;
input n_306;
input n_92;
input n_203;
input n_436;
input n_150;
input n_324;
input n_669;
input n_931;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_967;
input n_1083;
input n_746;
input n_292;
input n_1079;
input n_615;
input n_1139;
input n_76;
input n_517;
input n_0;
input n_824;
input n_428;
input n_159;
input n_892;
input n_959;
input n_30;
input n_1101;
input n_563;
input n_144;
input n_990;
input n_867;
input n_1226;
input n_944;
input n_749;
input n_815;
input n_542;
input n_470;
input n_1240;
input n_1087;
input n_632;
input n_477;
input n_650;
input n_425;
input n_1155;
input n_1071;
input n_712;
input n_976;
input n_909;
input n_767;
input n_964;
input n_382;
input n_489;
input n_80;
input n_251;
input n_974;
input n_506;
input n_799;
input n_1147;
input n_397;
input n_471;
input n_351;
input n_965;
input n_155;
input n_934;
input n_1220;
input n_356;
input n_698;
input n_124;
input n_307;
input n_1209;
input n_1020;
input n_646;
input n_34;
input n_404;
input n_172;
input n_1058;
input n_347;
input n_1042;
input n_183;
input n_1234;
input n_479;
input n_299;
input n_836;
input n_564;
input n_133;
input n_66;
input n_205;
input n_1029;
input n_1247;
input n_760;
input n_522;
input n_20;
input n_367;
input n_1111;
input n_970;
input n_713;
input n_1255;
input n_598;
input n_345;
input n_1237;
input n_927;
input n_261;
input n_1095;
input n_370;
input n_706;
input n_286;
input n_776;
input n_424;
input n_85;
input n_130;
input n_466;
input n_1263;
input n_346;
input n_348;
input n_552;
input n_670;
input n_379;
input n_138;
input n_162;
input n_264;
input n_441;
input n_1032;
input n_1217;
input n_637;
input n_73;
input n_327;
input n_1259;
input n_1177;
input n_1231;
input n_980;
input n_905;
input n_207;
input n_720;
input n_926;
input n_41;
input n_194;
input n_1163;
input n_186;
input n_145;
input n_59;
input n_1173;
input n_1068;
input n_1198;
input n_487;
input n_90;
input n_855;
input n_158;
input n_808;
input n_553;
input n_814;
input n_578;
input n_405;
input n_120;
input n_320;
input n_1134;
input n_647;
input n_481;
input n_600;
input n_1053;
input n_529;
input n_502;
input n_218;
input n_247;
input n_1105;
input n_547;
input n_439;
input n_604;
input n_677;
input n_478;
input n_703;
input n_1061;
input n_326;
input n_681;
input n_227;
input n_874;
input n_707;
input n_11;
input n_129;
input n_126;
input n_983;
input n_590;
input n_699;
input n_727;
input n_301;
input n_545;
input n_1015;
input n_1162;
input n_536;
input n_325;
input n_688;
input n_636;
input n_427;
input n_1098;
input n_442;
input n_777;
input n_1080;
input n_920;
input n_1086;
input n_1092;
input n_986;
input n_1104;
input n_729;
input n_887;
input n_1122;
input n_1205;
input n_163;
input n_1132;
input n_390;
input n_1156;
input n_501;
input n_314;
input n_1120;
input n_1202;
input n_627;
input n_1188;
input n_233;
input n_957;
input n_388;
input n_1242;
input n_1218;
input n_221;
input n_321;
input n_86;
input n_861;
input n_877;
input n_1119;
input n_616;
input n_1055;
input n_1189;
input n_1089;
input n_281;
input n_262;
input n_735;
input n_297;
input n_1005;
input n_527;
input n_46;
input n_84;
input n_845;
input n_888;
input n_178;
input n_551;
input n_417;
input n_70;
input n_343;
input n_1222;
input n_582;
input n_755;
input n_1097;
input n_1219;
input n_710;
input n_534;
input n_1239;
input n_278;
input n_560;
input n_890;
input n_842;
input n_148;
input n_451;
input n_745;
input n_61;
input n_742;
input n_1081;
input n_1266;
input n_769;
input n_13;
input n_476;
input n_832;
input n_55;
input n_535;
input n_744;
input n_982;
input n_915;
input n_215;
input n_1075;
input n_454;
input n_298;
input n_1227;
input n_655;
input n_403;
input n_1007;
input n_657;
input n_837;
input n_812;
input n_606;
input n_951;
input n_862;
input n_659;
input n_509;
input n_666;
input n_430;
input n_1206;
input n_722;
input n_1171;
input n_1030;
input n_785;
input n_999;
input n_456;
input n_852;
input n_704;
input n_1060;
input n_1044;
input n_521;
input n_873;
input n_1243;
input n_342;
input n_358;
input n_608;
input n_1037;
input n_317;
input n_134;
input n_1257;
input n_1078;
input n_266;
input n_157;
input n_1161;
input n_811;
input n_624;
input n_791;
input n_876;
input n_618;
input n_1191;
input n_736;
input n_1025;
input n_1215;
input n_241;
input n_687;
input n_797;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_602;
input n_592;
input n_854;
input n_393;
input n_474;
input n_805;
input n_295;
input n_190;
input n_1072;
input n_695;
input n_64;
input n_180;
input n_730;
input n_386;
input n_516;
input n_1137;
input n_1258;
input n_197;
input n_640;
input n_463;
input n_943;
input n_1118;
input n_678;
input n_651;
input n_961;
input n_469;
input n_1046;
input n_726;
input n_1123;
input n_878;
input n_771;
input n_752;
input n_71;
input n_985;
input n_421;
input n_906;
input n_1180;
input n_283;
input n_806;
input n_649;
input n_374;
input n_643;
input n_226;
input n_682;
input n_36;
input n_819;
input n_586;
input n_686;
input n_605;
input n_1154;
input n_584;
input n_1130;
input n_349;
input n_756;
input n_1016;
input n_1149;
input n_979;
input n_2;
input n_897;
input n_949;
input n_515;
input n_807;
input n_891;
input n_885;
input n_198;
input n_1208;
input n_396;
input n_802;
input n_23;
input n_1151;
input n_554;
input n_960;
input n_1256;
input n_87;
input n_714;
input n_790;
input n_354;
input n_140;
input n_725;
input n_151;
input n_28;
input n_1009;
input n_230;
input n_1133;
input n_154;
input n_883;
input n_142;
input n_473;
input n_801;
input n_818;
input n_779;
input n_594;
input n_35;
input n_1052;
input n_272;
input n_833;
input n_879;
input n_1117;
input n_38;
input n_422;
input n_1269;
input n_597;
input n_75;
input n_1047;
input n_95;
input n_1050;
input n_566;
input n_152;
input n_169;
input n_106;
input n_1201;
input n_173;
input n_858;
input n_1185;
input n_335;
input n_1035;
input n_1143;
input n_344;
input n_426;
input n_433;
input n_398;
input n_62;
input n_210;
input n_1090;
input n_166;
input n_253;
input n_928;
input n_1153;
input n_271;
input n_465;
input n_825;
input n_1103;
input n_732;
input n_1192;
input n_128;
input n_224;
input n_82;
input n_894;
input n_420;
input n_562;
input n_748;
input n_510;
input n_1045;
input n_256;
input n_1160;
input n_1023;
input n_988;
input n_330;
input n_914;
input n_400;
input n_689;
input n_1116;
input n_282;
input n_328;
input n_368;
input n_467;
input n_644;
input n_1197;
input n_276;
input n_497;
input n_1165;
input n_168;
input n_81;
input n_538;
input n_576;
input n_843;
input n_511;
input n_455;
input n_429;
input n_588;
input n_638;
input n_1128;
input n_1048;
input n_775;
input n_667;
input n_1049;
input n_14;
input n_869;
input n_141;
input n_846;
input n_305;
input n_312;
input n_56;
input n_60;
input n_728;
input n_413;
input n_715;
input n_889;
input n_1066;
input n_935;
input n_685;
input n_911;
input n_361;
input n_89;
input n_623;
input n_1065;
input n_453;
input n_74;
input n_810;
input n_19;
input n_40;
input n_181;
input n_617;
input n_543;
input n_236;
input n_601;
input n_683;
input n_565;
input n_628;
input n_743;
input n_1194;
input n_907;
input n_660;
input n_464;
input n_962;
input n_941;
input n_1210;
input n_847;
input n_747;
input n_1135;
input n_918;
input n_107;
input n_639;
input n_452;
input n_673;
input n_1038;
input n_414;
input n_571;
input n_6;
input n_284;
input n_593;
input n_1164;
input n_37;
input n_58;
input n_609;
input n_1193;
input n_613;
input n_1022;
input n_1033;
input n_409;
input n_171;
input n_519;
input n_384;
input n_1166;
input n_1056;
input n_526;
input n_1040;
input n_674;
input n_1158;
input n_316;
input n_125;
input n_820;
input n_43;
input n_872;
input n_254;
input n_1157;
input n_234;
input n_848;
input n_280;
input n_629;
input n_161;
input n_532;
input n_763;
input n_99;
input n_540;
input n_216;
input n_692;
input n_5;
input n_984;
input n_223;
input n_750;
input n_834;
input n_800;
input n_395;
input n_621;
input n_213;
input n_67;
input n_1014;
input n_724;
input n_493;
input n_114;
input n_1100;
input n_585;
input n_875;
input n_827;
input n_697;
input n_622;
input n_296;
input n_880;
input n_793;
input n_1175;
input n_132;
input n_751;
input n_1027;
input n_1070;
input n_739;
input n_1028;
input n_1221;
input n_530;
input n_792;
input n_1262;
input n_580;
input n_494;
input n_434;
input n_975;
input n_229;
input n_394;
input n_923;
input n_1124;
input n_932;
input n_1183;
input n_981;
input n_1110;
input n_243;
input n_185;
input n_1204;
input n_994;
input n_973;
input n_268;
input n_972;
input n_164;
input n_184;
input n_856;
input n_1248;
input n_1176;
input n_1054;
input n_508;
input n_118;
input n_121;
input n_353;
input n_1057;
input n_191;
input n_978;
input n_1011;
input n_828;
input n_322;
input n_558;
input n_116;
input n_39;
input n_653;
input n_783;
input n_556;
input n_1127;
input n_170;
input n_160;
input n_119;
input n_1008;
input n_332;
input n_581;
input n_294;
input n_1024;
input n_830;
input n_176;
input n_987;
input n_936;
input n_541;
input n_499;
input n_788;
input n_12;
input n_908;
input n_1036;
input n_341;
input n_1270;
input n_109;
input n_1167;
input n_549;
input n_591;
input n_969;
input n_919;
input n_50;
input n_318;
input n_103;
input n_244;
input n_679;
input n_220;
input n_663;
input n_443;
input n_528;
input n_1200;
input n_387;
input n_406;
input n_826;
input n_139;
input n_391;
input n_940;
input n_1077;
input n_607;
input n_956;
input n_445;
input n_765;
input n_122;
input n_1268;
input n_385;
input n_917;
input n_1271;
input n_372;
input n_15;
input n_631;
input n_399;
input n_1170;
input n_1261;
input n_702;
input n_857;
input n_898;
input n_363;
input n_968;
input n_1067;
input n_1235;
input n_1064;
input n_633;
input n_900;
input n_1093;
input n_193;
input n_733;
input n_761;
input n_731;
input n_336;
input n_315;
input n_311;
input n_8;
input n_668;
input n_758;
input n_1106;
input n_47;
input n_153;
input n_18;
input n_648;
input n_784;
input n_269;
input n_816;
input n_835;
input n_446;
input n_1076;
input n_753;
input n_701;
input n_1003;
input n_1125;
input n_309;
input n_115;
input n_401;
input n_485;
input n_504;
input n_483;
input n_435;
input n_1141;
input n_291;
input n_822;
input n_1094;
input n_840;
input n_1099;
input n_839;
input n_79;
input n_3;
input n_759;
input n_567;
input n_91;
input n_240;
input n_369;
input n_44;
input n_1172;
input n_614;
input n_1212;
input n_831;
input n_778;
input n_48;
input n_188;
input n_323;
input n_550;
input n_997;
input n_635;
input n_694;
input n_1113;
input n_248;
input n_1152;
input n_921;
input n_1236;
input n_228;
input n_1265;
input n_671;
input n_1;
input n_1148;
input n_654;
input n_488;
input n_904;
input n_505;
input n_88;
input n_498;
input n_1059;
input n_684;
input n_1039;
input n_539;
input n_1150;
input n_977;
input n_449;
input n_392;
input n_459;
input n_1136;
input n_458;
input n_1190;
input n_1144;
input n_383;
input n_838;
input n_175;
input n_950;
input n_1017;
input n_711;
input n_734;
input n_723;
input n_658;
input n_630;
input n_53;
input n_362;
input n_310;
input n_709;
input n_24;
input n_809;
input n_235;
input n_881;
input n_1019;
input n_662;
input n_641;
input n_910;
input n_290;
input n_741;
input n_939;
input n_371;
input n_199;
input n_217;
input n_1114;
input n_708;
input n_308;
input n_1223;
input n_201;
input n_572;
input n_1199;
input n_865;
input n_10;
input n_1041;
input n_993;
input n_948;
input n_922;
input n_1004;
input n_448;
input n_860;
input n_1043;
input n_255;
input n_450;
input n_896;
input n_902;
input n_1031;
input n_853;
input n_716;
input n_196;
input n_774;
input n_933;
input n_596;
input n_954;
input n_1168;
input n_219;
input n_231;
input n_656;
input n_492;
input n_574;
input n_252;
input n_664;
input n_1229;
input n_68;
input n_415;
input n_63;
input n_544;
input n_1186;
input n_599;
input n_768;
input n_1091;
input n_537;
input n_1063;
input n_25;
input n_991;
input n_83;
input n_389;
input n_1126;
input n_195;
input n_938;
input n_895;
input n_110;
input n_304;
input n_583;
input n_1000;
input n_313;
input n_626;
input n_378;
input n_98;
input n_946;
input n_757;
input n_375;
input n_113;
input n_33;
input n_1146;
input n_1203;
input n_998;
input n_472;
input n_937;
input n_265;
input n_208;
input n_156;
input n_174;
input n_275;
input n_100;
input n_147;
input n_204;
input n_1232;
input n_996;
input n_1211;
input n_963;
input n_1264;
input n_51;
input n_1082;
input n_496;
input n_866;
input n_26;
input n_246;
input n_925;
input n_1001;
input n_1115;
input n_1002;
input n_105;
input n_1051;
input n_719;
input n_131;
input n_263;
input n_1102;
input n_360;
input n_1129;
input n_1252;
input n_250;
input n_773;
input n_165;
input n_1010;
input n_882;
input n_1249;
input n_101;
input n_803;
input n_329;
input n_718;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_548;
input n_523;
input n_457;
input n_177;
input n_782;
input n_364;
input n_258;
input n_431;
input n_1228;
input n_1244;
input n_411;
input n_484;
input n_849;
input n_22;
input n_29;
input n_357;
input n_412;
input n_1251;
input n_447;
input n_1233;
input n_893;
input n_841;
input n_886;
input n_1069;
input n_359;
input n_573;
input n_796;
input n_127;
input n_531;
input n_675;

output n_5396;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_2182;
wire n_2680;
wire n_3264;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_5302;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_2646;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_2482;
wire n_1682;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_2663;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_4143;
wire n_4273;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_3482;
wire n_1900;
wire n_4268;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_4476;
wire n_2956;
wire n_5210;
wire n_2382;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5391;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_3549;
wire n_3914;
wire n_1692;
wire n_2611;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_2257;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_2019;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_2649;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_2697;
wire n_1817;
wire n_3704;
wire n_4296;
wire n_2677;
wire n_2483;
wire n_5088;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_5296;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_4292;
wire n_2118;
wire n_1490;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_2125;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_2707;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_3713;
wire n_1863;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_3944;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_2958;
wire n_1714;
wire n_4429;
wire n_3340;
wire n_5053;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_3864;
wire n_4694;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_2991;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_3740;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_4966;
wire n_2250;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_2610;
wire n_1593;
wire n_3715;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_3886;
wire n_2619;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_2613;
wire n_1517;
wire n_2647;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_3380;
wire n_2826;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_4355;
wire n_3818;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_3396;
wire n_4093;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_2561;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_3630;
wire n_1612;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2672;
wire n_2018;
wire n_2602;
wire n_2931;
wire n_3433;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_3786;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_4053;
wire n_3963;
wire n_3091;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_4083;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_5196;
wire n_2440;
wire n_2096;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_3633;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_2009;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1348;
wire n_2651;
wire n_2445;
wire n_2733;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_3457;
wire n_5384;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_5040;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_2148;
wire n_4663;
wire n_3296;
wire n_3762;
wire n_3794;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_3707;
wire n_3895;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_1581;
wire n_3058;
wire n_2047;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_5355;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_4120;
wire n_2880;
wire n_1313;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1339;
wire n_5116;
wire n_3771;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_2830;
wire n_4622;
wire n_4757;
wire n_1871;
wire n_4016;
wire n_3334;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_4591;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_2259;
wire n_5337;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_3181;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_1566;
wire n_2837;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_2248;
wire n_4660;
wire n_3081;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_2844;
wire n_1979;
wire n_4814;
wire n_2221;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_3150;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1652;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_1560;
wire n_2899;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_2685;
wire n_2061;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_4995;
wire n_4498;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_3234;
wire n_1351;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_3391;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_3240;
wire n_5066;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_5130;
wire n_4175;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5150;
wire n_5111;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_3257;
wire n_3730;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_4003;
wire n_1832;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5159;
wire n_4022;
wire n_2495;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_3031;
wire n_2335;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_3599;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_2218;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_3995;
wire n_3908;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_2266;
wire n_4324;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_3791;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1513;
wire n_1527;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_2486;
wire n_1897;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_5378;
wire n_4706;
wire n_3879;
wire n_2022;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_3317;
wire n_4835;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_4372;
wire n_4097;
wire n_4162;
wire n_5293;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_4960;
wire n_3738;
wire n_1380;
wire n_2020;
wire n_2310;
wire n_3600;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_3967;
wire n_4370;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_1968;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_4333;
wire n_5339;
wire n_2007;
wire n_3363;
wire n_1803;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_4217;
wire n_5277;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_3873;
wire n_4649;
wire n_2428;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_4999;
wire n_4592;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2817;
wire n_2773;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_5193;
wire n_4933;
wire n_4144;
wire n_2375;
wire n_3278;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5273;
wire n_2469;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1510;
wire n_3002;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_3681;
wire n_3970;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1941;
wire n_3637;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_2297;
wire n_1410;
wire n_4203;
wire n_1325;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_3674;
wire n_1638;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_3499;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5375;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_3075;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_4299;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_2731;
wire n_3703;
wire n_5265;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_3435;
wire n_2380;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_3856;
wire n_4038;
wire n_5316;
wire n_2735;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_4174;
wire n_5131;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1274;
wire n_4394;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_5333;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_3479;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_2755;
wire n_5109;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_3936;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_3078;
wire n_3971;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_2308;
wire n_1939;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_3983;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_2338;
wire n_5261;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_2660;
wire n_3426;
wire n_1859;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_5298;
wire n_3417;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1734;
wire n_1860;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_4545;
wire n_4758;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_4535;
wire n_4385;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1733;
wire n_4651;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_2353;
wire n_1429;
wire n_2528;
wire n_1778;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_3718;
wire n_3390;
wire n_2298;
wire n_4666;
wire n_4082;
wire n_2320;
wire n_3140;
wire n_3976;
wire n_2813;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_4377;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5270;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_4561;
wire n_3291;
wire n_1541;
wire n_1472;
wire n_2578;
wire n_2475;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_2845;
wire n_4151;
wire n_4412;
wire n_2036;
wire n_3358;
wire n_2533;
wire n_2003;
wire n_1307;
wire n_4682;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_3289;
wire n_1955;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_3620;
wire n_4601;
wire n_4518;
wire n_2767;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_2862;
wire n_4325;
wire n_2553;
wire n_2645;
wire n_1420;
wire n_4711;
wire n_2749;
wire n_4413;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_3131;
wire n_4138;
wire n_1973;
wire n_1444;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_4620;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_1645;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_2465;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_1834;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_4858;
wire n_1445;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_2409;
wire n_2966;
wire n_1720;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_2597;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_3032;
wire n_4886;
wire n_5172;
wire n_1477;
wire n_1982;
wire n_5311;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1273;
wire n_2982;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_4693;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_1891;
wire n_5348;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1725;
wire n_2318;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_3045;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_4047;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_2135;
wire n_4475;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_1503;
wire n_5295;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_2323;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_1988;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_2078;
wire n_4809;
wire n_4012;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_5368;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_2727;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_3698;
wire n_4513;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2549;
wire n_2499;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_2378;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_1483;
wire n_1363;
wire n_3467;
wire n_3179;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_3699;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_2801;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_3276;
wire n_3682;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2932;
wire n_2027;
wire n_3118;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_1467;
wire n_5209;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_3009;
wire n_5219;
wire n_3951;
wire n_3035;
wire n_4261;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_1388;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_1532;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_2916;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_5017;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_2091;
wire n_4312;
wire n_3789;
wire n_1658;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2725;
wire n_2667;
wire n_3746;
wire n_4537;
wire n_3694;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_2945;
wire n_1971;
wire n_3543;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_2698;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_4595;
wire n_2352;
wire n_5201;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_2174;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_1687;
wire n_4703;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1758;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_3677;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_4131;
wire n_4215;
wire n_2488;
wire n_1509;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_2169;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_4578;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_2724;
wire n_2258;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_2111;
wire n_3743;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_4749;
wire n_1845;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_4211;
wire n_3094;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_5034;
wire n_3312;
wire n_2451;
wire n_2913;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_4516;
wire n_5235;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1192),
.Y(n_1272)
);

CKINVDCx20_ASAP7_75t_R g1273 ( 
.A(n_1095),
.Y(n_1273)
);

BUFx10_ASAP7_75t_L g1274 ( 
.A(n_1014),
.Y(n_1274)
);

INVx2_ASAP7_75t_SL g1275 ( 
.A(n_979),
.Y(n_1275)
);

CKINVDCx5p33_ASAP7_75t_R g1276 ( 
.A(n_782),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1050),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_967),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_932),
.Y(n_1279)
);

BUFx5_ASAP7_75t_L g1280 ( 
.A(n_980),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1143),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_891),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_728),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1261),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1123),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_881),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_758),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_777),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1128),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1047),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1065),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_407),
.Y(n_1292)
);

BUFx2_ASAP7_75t_L g1293 ( 
.A(n_465),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_1152),
.Y(n_1294)
);

CKINVDCx20_ASAP7_75t_R g1295 ( 
.A(n_911),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_283),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1266),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1218),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_1042),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_268),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_1231),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_994),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1012),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_924),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_608),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_243),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_1212),
.Y(n_1307)
);

CKINVDCx5p33_ASAP7_75t_R g1308 ( 
.A(n_1183),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1072),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_1203),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_753),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_623),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1125),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_1082),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_150),
.Y(n_1315)
);

CKINVDCx5p33_ASAP7_75t_R g1316 ( 
.A(n_983),
.Y(n_1316)
);

BUFx6f_ASAP7_75t_L g1317 ( 
.A(n_1138),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_61),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_574),
.Y(n_1319)
);

BUFx6f_ASAP7_75t_L g1320 ( 
.A(n_250),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_926),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_784),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_703),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1106),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_367),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_900),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_729),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_821),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_366),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1137),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1111),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_188),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_509),
.Y(n_1333)
);

INVx1_ASAP7_75t_SL g1334 ( 
.A(n_403),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1209),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_525),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_459),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_1264),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1257),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_295),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_795),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1194),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1197),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_313),
.Y(n_1344)
);

CKINVDCx5p33_ASAP7_75t_R g1345 ( 
.A(n_930),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_986),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_189),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_889),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_662),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1130),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1085),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_359),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_888),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1071),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1247),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_398),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_57),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1190),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_612),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1131),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1066),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_958),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_943),
.Y(n_1363)
);

CKINVDCx16_ASAP7_75t_R g1364 ( 
.A(n_544),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_1243),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1078),
.Y(n_1366)
);

INVx1_ASAP7_75t_SL g1367 ( 
.A(n_1158),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_904),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_143),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_636),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_147),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_803),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_466),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_658),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1155),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1187),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_74),
.Y(n_1377)
);

INVx2_ASAP7_75t_SL g1378 ( 
.A(n_985),
.Y(n_1378)
);

CKINVDCx5p33_ASAP7_75t_R g1379 ( 
.A(n_700),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1080),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1079),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_331),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_236),
.Y(n_1383)
);

BUFx10_ASAP7_75t_L g1384 ( 
.A(n_1087),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1044),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_401),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_278),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_170),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_336),
.Y(n_1389)
);

CKINVDCx20_ASAP7_75t_R g1390 ( 
.A(n_1179),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_489),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_795),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_225),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_281),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_369),
.Y(n_1395)
);

BUFx6f_ASAP7_75t_L g1396 ( 
.A(n_180),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_663),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_954),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1221),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_376),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1016),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_19),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_415),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1160),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_756),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_300),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1170),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_860),
.Y(n_1408)
);

INVx1_ASAP7_75t_SL g1409 ( 
.A(n_1139),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_91),
.Y(n_1410)
);

CKINVDCx12_ASAP7_75t_R g1411 ( 
.A(n_942),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_325),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_166),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_973),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_607),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_1119),
.Y(n_1416)
);

CKINVDCx20_ASAP7_75t_R g1417 ( 
.A(n_1091),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_907),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1088),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_976),
.Y(n_1420)
);

BUFx2_ASAP7_75t_SL g1421 ( 
.A(n_928),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_519),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1093),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_900),
.Y(n_1424)
);

CKINVDCx14_ASAP7_75t_R g1425 ( 
.A(n_1052),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_440),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_818),
.Y(n_1427)
);

CKINVDCx5p33_ASAP7_75t_R g1428 ( 
.A(n_180),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_137),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1220),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_17),
.Y(n_1431)
);

CKINVDCx16_ASAP7_75t_R g1432 ( 
.A(n_93),
.Y(n_1432)
);

CKINVDCx16_ASAP7_75t_R g1433 ( 
.A(n_456),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_294),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_167),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_627),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_87),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_375),
.Y(n_1438)
);

CKINVDCx16_ASAP7_75t_R g1439 ( 
.A(n_441),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1248),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_280),
.Y(n_1441)
);

CKINVDCx20_ASAP7_75t_R g1442 ( 
.A(n_212),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_3),
.Y(n_1443)
);

INVx1_ASAP7_75t_SL g1444 ( 
.A(n_1237),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1148),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_518),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_993),
.Y(n_1447)
);

BUFx5_ASAP7_75t_L g1448 ( 
.A(n_1063),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_505),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_290),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1084),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_95),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_939),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_1263),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_226),
.Y(n_1455)
);

CKINVDCx5p33_ASAP7_75t_R g1456 ( 
.A(n_40),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_186),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_1240),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_698),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_995),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_372),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1108),
.Y(n_1462)
);

BUFx2_ASAP7_75t_L g1463 ( 
.A(n_711),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_120),
.Y(n_1464)
);

CKINVDCx16_ASAP7_75t_R g1465 ( 
.A(n_755),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_1176),
.Y(n_1466)
);

CKINVDCx20_ASAP7_75t_R g1467 ( 
.A(n_959),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1204),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_702),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_341),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1153),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_304),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_174),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_701),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_981),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_782),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_592),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_977),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_944),
.Y(n_1479)
);

BUFx10_ASAP7_75t_L g1480 ( 
.A(n_553),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_657),
.Y(n_1481)
);

CKINVDCx5p33_ASAP7_75t_R g1482 ( 
.A(n_869),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_150),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_675),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_1154),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1057),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1140),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1032),
.Y(n_1488)
);

INVx1_ASAP7_75t_SL g1489 ( 
.A(n_73),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_879),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1211),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_131),
.Y(n_1492)
);

BUFx2_ASAP7_75t_L g1493 ( 
.A(n_1055),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_716),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_1113),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1008),
.Y(n_1496)
);

CKINVDCx14_ASAP7_75t_R g1497 ( 
.A(n_1156),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_330),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_1124),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1224),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_274),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_462),
.Y(n_1502)
);

BUFx10_ASAP7_75t_L g1503 ( 
.A(n_917),
.Y(n_1503)
);

CKINVDCx14_ASAP7_75t_R g1504 ( 
.A(n_226),
.Y(n_1504)
);

CKINVDCx5p33_ASAP7_75t_R g1505 ( 
.A(n_559),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1232),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1162),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_184),
.Y(n_1508)
);

BUFx10_ASAP7_75t_L g1509 ( 
.A(n_1120),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_516),
.Y(n_1510)
);

BUFx6f_ASAP7_75t_L g1511 ( 
.A(n_592),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_739),
.Y(n_1512)
);

CKINVDCx16_ASAP7_75t_R g1513 ( 
.A(n_1129),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1046),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1070),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_138),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_582),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1033),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_105),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_69),
.Y(n_1520)
);

CKINVDCx5p33_ASAP7_75t_R g1521 ( 
.A(n_1115),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_238),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_11),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1244),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_662),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_628),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_950),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1000),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_781),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_931),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_873),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_203),
.Y(n_1532)
);

INVx1_ASAP7_75t_SL g1533 ( 
.A(n_1185),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_81),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_455),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1164),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_358),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_229),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_161),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_429),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_1242),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_222),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_619),
.Y(n_1543)
);

CKINVDCx20_ASAP7_75t_R g1544 ( 
.A(n_1073),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_354),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1105),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_694),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_864),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_756),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_81),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_832),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_489),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_609),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_605),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_239),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_946),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_925),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1172),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_20),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_633),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_185),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1245),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_963),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_851),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_63),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_991),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_745),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1056),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1167),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_240),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_946),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1045),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_564),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_797),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_154),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_953),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_955),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1122),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_951),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_205),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1141),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_386),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1250),
.Y(n_1583)
);

BUFx3_ASAP7_75t_L g1584 ( 
.A(n_1195),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_527),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_158),
.Y(n_1586)
);

CKINVDCx5p33_ASAP7_75t_R g1587 ( 
.A(n_783),
.Y(n_1587)
);

CKINVDCx5p33_ASAP7_75t_R g1588 ( 
.A(n_506),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_260),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_277),
.Y(n_1590)
);

CKINVDCx5p33_ASAP7_75t_R g1591 ( 
.A(n_153),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_1118),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_876),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_311),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_715),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_422),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_1168),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1181),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_737),
.Y(n_1599)
);

CKINVDCx5p33_ASAP7_75t_R g1600 ( 
.A(n_972),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_492),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1256),
.Y(n_1602)
);

CKINVDCx5p33_ASAP7_75t_R g1603 ( 
.A(n_483),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_814),
.Y(n_1604)
);

BUFx10_ASAP7_75t_L g1605 ( 
.A(n_308),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_625),
.Y(n_1606)
);

CKINVDCx20_ASAP7_75t_R g1607 ( 
.A(n_860),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_250),
.Y(n_1608)
);

CKINVDCx20_ASAP7_75t_R g1609 ( 
.A(n_205),
.Y(n_1609)
);

CKINVDCx5p33_ASAP7_75t_R g1610 ( 
.A(n_513),
.Y(n_1610)
);

BUFx8_ASAP7_75t_SL g1611 ( 
.A(n_689),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_704),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_945),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_956),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_492),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_367),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1249),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_141),
.Y(n_1618)
);

BUFx3_ASAP7_75t_L g1619 ( 
.A(n_326),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_893),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1159),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_32),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_962),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_791),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1007),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_974),
.Y(n_1626)
);

BUFx3_ASAP7_75t_L g1627 ( 
.A(n_1206),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1269),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1214),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_990),
.Y(n_1630)
);

CKINVDCx5p33_ASAP7_75t_R g1631 ( 
.A(n_455),
.Y(n_1631)
);

BUFx10_ASAP7_75t_L g1632 ( 
.A(n_366),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_49),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1114),
.Y(n_1634)
);

BUFx2_ASAP7_75t_L g1635 ( 
.A(n_300),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1104),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_960),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1135),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1142),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_817),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_464),
.Y(n_1641)
);

INVx2_ASAP7_75t_SL g1642 ( 
.A(n_1077),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_1134),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1234),
.Y(n_1644)
);

CKINVDCx5p33_ASAP7_75t_R g1645 ( 
.A(n_372),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_512),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1030),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_16),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_580),
.Y(n_1649)
);

CKINVDCx5p33_ASAP7_75t_R g1650 ( 
.A(n_786),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_365),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1133),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_907),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1201),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_538),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_225),
.Y(n_1656)
);

CKINVDCx5p33_ASAP7_75t_R g1657 ( 
.A(n_1217),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_802),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_992),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1198),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_332),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_1260),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_938),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_1210),
.Y(n_1664)
);

CKINVDCx20_ASAP7_75t_R g1665 ( 
.A(n_384),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_145),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1225),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_274),
.Y(n_1668)
);

BUFx3_ASAP7_75t_L g1669 ( 
.A(n_1233),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_696),
.Y(n_1670)
);

CKINVDCx5p33_ASAP7_75t_R g1671 ( 
.A(n_23),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_269),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_808),
.Y(n_1673)
);

CKINVDCx5p33_ASAP7_75t_R g1674 ( 
.A(n_1116),
.Y(n_1674)
);

INVx1_ASAP7_75t_SL g1675 ( 
.A(n_844),
.Y(n_1675)
);

CKINVDCx5p33_ASAP7_75t_R g1676 ( 
.A(n_314),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_133),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_471),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_190),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1161),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_59),
.Y(n_1681)
);

INVx1_ASAP7_75t_SL g1682 ( 
.A(n_1265),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_894),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_453),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_229),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_599),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_339),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_1048),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1098),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_963),
.Y(n_1690)
);

CKINVDCx5p33_ASAP7_75t_R g1691 ( 
.A(n_197),
.Y(n_1691)
);

CKINVDCx5p33_ASAP7_75t_R g1692 ( 
.A(n_821),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1230),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_313),
.Y(n_1694)
);

BUFx10_ASAP7_75t_L g1695 ( 
.A(n_1083),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_45),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_644),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1157),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_941),
.Y(n_1699)
);

BUFx3_ASAP7_75t_L g1700 ( 
.A(n_446),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_51),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1092),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_975),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_457),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_800),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_36),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1074),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1086),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1208),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1262),
.Y(n_1710)
);

CKINVDCx5p33_ASAP7_75t_R g1711 ( 
.A(n_691),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_660),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1268),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_220),
.Y(n_1714)
);

CKINVDCx20_ASAP7_75t_R g1715 ( 
.A(n_1017),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_359),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_771),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1270),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_458),
.Y(n_1719)
);

CKINVDCx5p33_ASAP7_75t_R g1720 ( 
.A(n_1097),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_96),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1019),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1241),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_748),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1202),
.Y(n_1725)
);

CKINVDCx5p33_ASAP7_75t_R g1726 ( 
.A(n_933),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_897),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1267),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_732),
.Y(n_1729)
);

INVx4_ASAP7_75t_R g1730 ( 
.A(n_1219),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_480),
.Y(n_1731)
);

CKINVDCx5p33_ASAP7_75t_R g1732 ( 
.A(n_1213),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1061),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_321),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1205),
.Y(n_1735)
);

CKINVDCx20_ASAP7_75t_R g1736 ( 
.A(n_303),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1174),
.Y(n_1737)
);

CKINVDCx14_ASAP7_75t_R g1738 ( 
.A(n_989),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_12),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_190),
.Y(n_1740)
);

BUFx10_ASAP7_75t_L g1741 ( 
.A(n_536),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1186),
.Y(n_1742)
);

CKINVDCx5p33_ASAP7_75t_R g1743 ( 
.A(n_1165),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_572),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_941),
.Y(n_1745)
);

CKINVDCx5p33_ASAP7_75t_R g1746 ( 
.A(n_985),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_822),
.Y(n_1747)
);

CKINVDCx5p33_ASAP7_75t_R g1748 ( 
.A(n_115),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_959),
.Y(n_1749)
);

CKINVDCx5p33_ASAP7_75t_R g1750 ( 
.A(n_1251),
.Y(n_1750)
);

CKINVDCx5p33_ASAP7_75t_R g1751 ( 
.A(n_837),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_482),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_377),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_461),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_320),
.Y(n_1755)
);

CKINVDCx5p33_ASAP7_75t_R g1756 ( 
.A(n_848),
.Y(n_1756)
);

CKINVDCx5p33_ASAP7_75t_R g1757 ( 
.A(n_934),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_91),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_547),
.Y(n_1759)
);

CKINVDCx16_ASAP7_75t_R g1760 ( 
.A(n_110),
.Y(n_1760)
);

INVx1_ASAP7_75t_SL g1761 ( 
.A(n_414),
.Y(n_1761)
);

CKINVDCx5p33_ASAP7_75t_R g1762 ( 
.A(n_1037),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1117),
.Y(n_1763)
);

CKINVDCx5p33_ASAP7_75t_R g1764 ( 
.A(n_289),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_645),
.Y(n_1765)
);

CKINVDCx20_ASAP7_75t_R g1766 ( 
.A(n_106),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1226),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_259),
.Y(n_1768)
);

CKINVDCx5p33_ASAP7_75t_R g1769 ( 
.A(n_399),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_948),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_493),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_656),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_130),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_965),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_854),
.Y(n_1775)
);

BUFx8_ASAP7_75t_SL g1776 ( 
.A(n_556),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1169),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_669),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_130),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_601),
.Y(n_1780)
);

CKINVDCx5p33_ASAP7_75t_R g1781 ( 
.A(n_927),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_710),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1110),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_774),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_107),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_388),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_855),
.Y(n_1787)
);

CKINVDCx5p33_ASAP7_75t_R g1788 ( 
.A(n_1010),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_435),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_459),
.Y(n_1790)
);

CKINVDCx5p33_ASAP7_75t_R g1791 ( 
.A(n_404),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_451),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_383),
.Y(n_1793)
);

CKINVDCx5p33_ASAP7_75t_R g1794 ( 
.A(n_731),
.Y(n_1794)
);

BUFx2_ASAP7_75t_L g1795 ( 
.A(n_1132),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_269),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1207),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1180),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1173),
.Y(n_1799)
);

CKINVDCx5p33_ASAP7_75t_R g1800 ( 
.A(n_1191),
.Y(n_1800)
);

BUFx5_ASAP7_75t_L g1801 ( 
.A(n_161),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_934),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1101),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_128),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1254),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_517),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_604),
.Y(n_1807)
);

CKINVDCx20_ASAP7_75t_R g1808 ( 
.A(n_177),
.Y(n_1808)
);

CKINVDCx5p33_ASAP7_75t_R g1809 ( 
.A(n_140),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1149),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_936),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_708),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1216),
.Y(n_1813)
);

BUFx6f_ASAP7_75t_L g1814 ( 
.A(n_970),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_319),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_971),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_913),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1076),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_987),
.Y(n_1819)
);

CKINVDCx5p33_ASAP7_75t_R g1820 ( 
.A(n_389),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1175),
.Y(n_1821)
);

CKINVDCx5p33_ASAP7_75t_R g1822 ( 
.A(n_610),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_140),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_630),
.Y(n_1824)
);

CKINVDCx20_ASAP7_75t_R g1825 ( 
.A(n_48),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_615),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1163),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_992),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_467),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_964),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_846),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_868),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_624),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_111),
.Y(n_1834)
);

CKINVDCx5p33_ASAP7_75t_R g1835 ( 
.A(n_1200),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_238),
.Y(n_1836)
);

BUFx10_ASAP7_75t_L g1837 ( 
.A(n_17),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_682),
.Y(n_1838)
);

CKINVDCx5p33_ASAP7_75t_R g1839 ( 
.A(n_1147),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1103),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_937),
.Y(n_1841)
);

CKINVDCx5p33_ASAP7_75t_R g1842 ( 
.A(n_354),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1051),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1094),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_563),
.Y(n_1845)
);

CKINVDCx5p33_ASAP7_75t_R g1846 ( 
.A(n_984),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1184),
.Y(n_1847)
);

CKINVDCx5p33_ASAP7_75t_R g1848 ( 
.A(n_1064),
.Y(n_1848)
);

CKINVDCx5p33_ASAP7_75t_R g1849 ( 
.A(n_1259),
.Y(n_1849)
);

CKINVDCx5p33_ASAP7_75t_R g1850 ( 
.A(n_383),
.Y(n_1850)
);

CKINVDCx5p33_ASAP7_75t_R g1851 ( 
.A(n_143),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1081),
.Y(n_1852)
);

CKINVDCx5p33_ASAP7_75t_R g1853 ( 
.A(n_421),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_145),
.Y(n_1854)
);

CKINVDCx5p33_ASAP7_75t_R g1855 ( 
.A(n_133),
.Y(n_1855)
);

INVx2_ASAP7_75t_SL g1856 ( 
.A(n_119),
.Y(n_1856)
);

CKINVDCx5p33_ASAP7_75t_R g1857 ( 
.A(n_978),
.Y(n_1857)
);

CKINVDCx5p33_ASAP7_75t_R g1858 ( 
.A(n_1005),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_355),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_802),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1150),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_673),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1228),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_99),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_168),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_935),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_759),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_965),
.Y(n_1868)
);

CKINVDCx5p33_ASAP7_75t_R g1869 ( 
.A(n_1053),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1166),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1253),
.Y(n_1871)
);

CKINVDCx5p33_ASAP7_75t_R g1872 ( 
.A(n_84),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1069),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1199),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_107),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_837),
.Y(n_1876)
);

CKINVDCx16_ASAP7_75t_R g1877 ( 
.A(n_899),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_187),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_607),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_955),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_236),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_766),
.Y(n_1882)
);

CKINVDCx5p33_ASAP7_75t_R g1883 ( 
.A(n_68),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_122),
.Y(n_1884)
);

INVx2_ASAP7_75t_SL g1885 ( 
.A(n_1235),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_979),
.Y(n_1886)
);

CKINVDCx5p33_ASAP7_75t_R g1887 ( 
.A(n_777),
.Y(n_1887)
);

BUFx6f_ASAP7_75t_L g1888 ( 
.A(n_256),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_488),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_484),
.Y(n_1890)
);

BUFx6f_ASAP7_75t_L g1891 ( 
.A(n_209),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_656),
.Y(n_1892)
);

CKINVDCx5p33_ASAP7_75t_R g1893 ( 
.A(n_957),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_155),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_578),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_449),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_116),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_888),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1127),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_457),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_605),
.Y(n_1901)
);

INVx3_ASAP7_75t_L g1902 ( 
.A(n_1151),
.Y(n_1902)
);

INVx1_ASAP7_75t_SL g1903 ( 
.A(n_103),
.Y(n_1903)
);

CKINVDCx5p33_ASAP7_75t_R g1904 ( 
.A(n_375),
.Y(n_1904)
);

CKINVDCx16_ASAP7_75t_R g1905 ( 
.A(n_961),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_856),
.Y(n_1906)
);

CKINVDCx5p33_ASAP7_75t_R g1907 ( 
.A(n_940),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_302),
.Y(n_1908)
);

CKINVDCx5p33_ASAP7_75t_R g1909 ( 
.A(n_921),
.Y(n_1909)
);

BUFx10_ASAP7_75t_L g1910 ( 
.A(n_1067),
.Y(n_1910)
);

BUFx10_ASAP7_75t_L g1911 ( 
.A(n_517),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1223),
.Y(n_1912)
);

CKINVDCx20_ASAP7_75t_R g1913 ( 
.A(n_0),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_604),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_969),
.Y(n_1915)
);

CKINVDCx5p33_ASAP7_75t_R g1916 ( 
.A(n_57),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_649),
.Y(n_1917)
);

CKINVDCx5p33_ASAP7_75t_R g1918 ( 
.A(n_546),
.Y(n_1918)
);

HB1xp67_ASAP7_75t_L g1919 ( 
.A(n_952),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_661),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1126),
.Y(n_1921)
);

CKINVDCx5p33_ASAP7_75t_R g1922 ( 
.A(n_264),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_20),
.Y(n_1923)
);

HB1xp67_ASAP7_75t_L g1924 ( 
.A(n_883),
.Y(n_1924)
);

BUFx10_ASAP7_75t_L g1925 ( 
.A(n_25),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_261),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_386),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_953),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_75),
.Y(n_1929)
);

CKINVDCx5p33_ASAP7_75t_R g1930 ( 
.A(n_540),
.Y(n_1930)
);

CKINVDCx5p33_ASAP7_75t_R g1931 ( 
.A(n_1058),
.Y(n_1931)
);

CKINVDCx5p33_ASAP7_75t_R g1932 ( 
.A(n_929),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1246),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1145),
.Y(n_1934)
);

BUFx3_ASAP7_75t_L g1935 ( 
.A(n_1107),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_973),
.Y(n_1936)
);

BUFx2_ASAP7_75t_L g1937 ( 
.A(n_1034),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_632),
.Y(n_1938)
);

CKINVDCx5p33_ASAP7_75t_R g1939 ( 
.A(n_1193),
.Y(n_1939)
);

CKINVDCx16_ASAP7_75t_R g1940 ( 
.A(n_1018),
.Y(n_1940)
);

CKINVDCx14_ASAP7_75t_R g1941 ( 
.A(n_968),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_151),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_933),
.Y(n_1943)
);

CKINVDCx5p33_ASAP7_75t_R g1944 ( 
.A(n_993),
.Y(n_1944)
);

CKINVDCx5p33_ASAP7_75t_R g1945 ( 
.A(n_135),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_982),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_732),
.Y(n_1947)
);

CKINVDCx5p33_ASAP7_75t_R g1948 ( 
.A(n_195),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_890),
.Y(n_1949)
);

BUFx2_ASAP7_75t_R g1950 ( 
.A(n_73),
.Y(n_1950)
);

CKINVDCx20_ASAP7_75t_R g1951 ( 
.A(n_302),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_644),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1049),
.Y(n_1953)
);

CKINVDCx5p33_ASAP7_75t_R g1954 ( 
.A(n_1178),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_547),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_289),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_664),
.Y(n_1957)
);

CKINVDCx5p33_ASAP7_75t_R g1958 ( 
.A(n_942),
.Y(n_1958)
);

CKINVDCx5p33_ASAP7_75t_R g1959 ( 
.A(n_828),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1112),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1146),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1236),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1060),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_293),
.Y(n_1964)
);

CKINVDCx5p33_ASAP7_75t_R g1965 ( 
.A(n_1100),
.Y(n_1965)
);

CKINVDCx20_ASAP7_75t_R g1966 ( 
.A(n_83),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_822),
.Y(n_1967)
);

CKINVDCx5p33_ASAP7_75t_R g1968 ( 
.A(n_654),
.Y(n_1968)
);

CKINVDCx5p33_ASAP7_75t_R g1969 ( 
.A(n_952),
.Y(n_1969)
);

BUFx2_ASAP7_75t_L g1970 ( 
.A(n_947),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_466),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1011),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_858),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_639),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_715),
.Y(n_1975)
);

BUFx6f_ASAP7_75t_L g1976 ( 
.A(n_1182),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1136),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_587),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_275),
.Y(n_1979)
);

CKINVDCx20_ASAP7_75t_R g1980 ( 
.A(n_132),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_981),
.Y(n_1981)
);

INVx1_ASAP7_75t_SL g1982 ( 
.A(n_544),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1038),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1171),
.Y(n_1984)
);

BUFx3_ASAP7_75t_L g1985 ( 
.A(n_346),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_139),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_772),
.Y(n_1987)
);

BUFx6f_ASAP7_75t_L g1988 ( 
.A(n_460),
.Y(n_1988)
);

BUFx2_ASAP7_75t_L g1989 ( 
.A(n_894),
.Y(n_1989)
);

CKINVDCx5p33_ASAP7_75t_R g1990 ( 
.A(n_755),
.Y(n_1990)
);

BUFx3_ASAP7_75t_L g1991 ( 
.A(n_534),
.Y(n_1991)
);

CKINVDCx5p33_ASAP7_75t_R g1992 ( 
.A(n_34),
.Y(n_1992)
);

CKINVDCx20_ASAP7_75t_R g1993 ( 
.A(n_1043),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_677),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_310),
.Y(n_1995)
);

CKINVDCx5p33_ASAP7_75t_R g1996 ( 
.A(n_1090),
.Y(n_1996)
);

CKINVDCx5p33_ASAP7_75t_R g1997 ( 
.A(n_1109),
.Y(n_1997)
);

INVx1_ASAP7_75t_SL g1998 ( 
.A(n_1054),
.Y(n_1998)
);

CKINVDCx5p33_ASAP7_75t_R g1999 ( 
.A(n_35),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1099),
.Y(n_2000)
);

CKINVDCx5p33_ASAP7_75t_R g2001 ( 
.A(n_188),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1189),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1062),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_778),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_524),
.Y(n_2005)
);

CKINVDCx5p33_ASAP7_75t_R g2006 ( 
.A(n_330),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_861),
.Y(n_2007)
);

CKINVDCx5p33_ASAP7_75t_R g2008 ( 
.A(n_714),
.Y(n_2008)
);

BUFx10_ASAP7_75t_L g2009 ( 
.A(n_1258),
.Y(n_2009)
);

CKINVDCx14_ASAP7_75t_R g2010 ( 
.A(n_422),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_643),
.Y(n_2011)
);

CKINVDCx5p33_ASAP7_75t_R g2012 ( 
.A(n_301),
.Y(n_2012)
);

INVx1_ASAP7_75t_SL g2013 ( 
.A(n_368),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_923),
.Y(n_2014)
);

BUFx2_ASAP7_75t_L g2015 ( 
.A(n_1255),
.Y(n_2015)
);

CKINVDCx5p33_ASAP7_75t_R g2016 ( 
.A(n_271),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_720),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_922),
.Y(n_2018)
);

CKINVDCx16_ASAP7_75t_R g2019 ( 
.A(n_971),
.Y(n_2019)
);

BUFx6f_ASAP7_75t_L g2020 ( 
.A(n_949),
.Y(n_2020)
);

CKINVDCx5p33_ASAP7_75t_R g2021 ( 
.A(n_488),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_761),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_974),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_111),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_412),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_815),
.Y(n_2026)
);

CKINVDCx5p33_ASAP7_75t_R g2027 ( 
.A(n_569),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_685),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_112),
.Y(n_2029)
);

INVx1_ASAP7_75t_SL g2030 ( 
.A(n_96),
.Y(n_2030)
);

CKINVDCx5p33_ASAP7_75t_R g2031 ( 
.A(n_1096),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1238),
.Y(n_2032)
);

CKINVDCx5p33_ASAP7_75t_R g2033 ( 
.A(n_543),
.Y(n_2033)
);

CKINVDCx5p33_ASAP7_75t_R g2034 ( 
.A(n_7),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1252),
.Y(n_2035)
);

CKINVDCx5p33_ASAP7_75t_R g2036 ( 
.A(n_932),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_867),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1239),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1144),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_323),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1089),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_0),
.Y(n_2042)
);

CKINVDCx5p33_ASAP7_75t_R g2043 ( 
.A(n_304),
.Y(n_2043)
);

CKINVDCx5p33_ASAP7_75t_R g2044 ( 
.A(n_1222),
.Y(n_2044)
);

BUFx6f_ASAP7_75t_L g2045 ( 
.A(n_804),
.Y(n_2045)
);

CKINVDCx5p33_ASAP7_75t_R g2046 ( 
.A(n_471),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_165),
.Y(n_2047)
);

BUFx10_ASAP7_75t_L g2048 ( 
.A(n_126),
.Y(n_2048)
);

BUFx6f_ASAP7_75t_L g2049 ( 
.A(n_1188),
.Y(n_2049)
);

CKINVDCx16_ASAP7_75t_R g2050 ( 
.A(n_1068),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_92),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_930),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_514),
.Y(n_2053)
);

CKINVDCx5p33_ASAP7_75t_R g2054 ( 
.A(n_1229),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_754),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_801),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_862),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_995),
.Y(n_2058)
);

CKINVDCx5p33_ASAP7_75t_R g2059 ( 
.A(n_975),
.Y(n_2059)
);

CKINVDCx5p33_ASAP7_75t_R g2060 ( 
.A(n_345),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_655),
.Y(n_2061)
);

CKINVDCx5p33_ASAP7_75t_R g2062 ( 
.A(n_1013),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_1196),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_37),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_668),
.Y(n_2065)
);

CKINVDCx5p33_ASAP7_75t_R g2066 ( 
.A(n_966),
.Y(n_2066)
);

INVx2_ASAP7_75t_L g2067 ( 
.A(n_231),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_649),
.Y(n_2068)
);

BUFx3_ASAP7_75t_L g2069 ( 
.A(n_882),
.Y(n_2069)
);

CKINVDCx20_ASAP7_75t_R g2070 ( 
.A(n_892),
.Y(n_2070)
);

CKINVDCx5p33_ASAP7_75t_R g2071 ( 
.A(n_224),
.Y(n_2071)
);

CKINVDCx20_ASAP7_75t_R g2072 ( 
.A(n_811),
.Y(n_2072)
);

INVxp67_ASAP7_75t_L g2073 ( 
.A(n_1002),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_442),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_502),
.Y(n_2075)
);

CKINVDCx5p33_ASAP7_75t_R g2076 ( 
.A(n_798),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_657),
.Y(n_2077)
);

CKINVDCx20_ASAP7_75t_R g2078 ( 
.A(n_1102),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1215),
.Y(n_2079)
);

INVx1_ASAP7_75t_SL g2080 ( 
.A(n_633),
.Y(n_2080)
);

CKINVDCx5p33_ASAP7_75t_R g2081 ( 
.A(n_799),
.Y(n_2081)
);

INVxp67_ASAP7_75t_L g2082 ( 
.A(n_305),
.Y(n_2082)
);

CKINVDCx5p33_ASAP7_75t_R g2083 ( 
.A(n_368),
.Y(n_2083)
);

CKINVDCx5p33_ASAP7_75t_R g2084 ( 
.A(n_520),
.Y(n_2084)
);

BUFx3_ASAP7_75t_L g2085 ( 
.A(n_1177),
.Y(n_2085)
);

CKINVDCx5p33_ASAP7_75t_R g2086 ( 
.A(n_247),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1271),
.Y(n_2087)
);

CKINVDCx5p33_ASAP7_75t_R g2088 ( 
.A(n_115),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_324),
.Y(n_2089)
);

INVx1_ASAP7_75t_L g2090 ( 
.A(n_199),
.Y(n_2090)
);

CKINVDCx5p33_ASAP7_75t_R g2091 ( 
.A(n_1059),
.Y(n_2091)
);

INVx2_ASAP7_75t_SL g2092 ( 
.A(n_494),
.Y(n_2092)
);

CKINVDCx5p33_ASAP7_75t_R g2093 ( 
.A(n_414),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1121),
.Y(n_2094)
);

INVx1_ASAP7_75t_SL g2095 ( 
.A(n_1075),
.Y(n_2095)
);

INVx2_ASAP7_75t_L g2096 ( 
.A(n_530),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_988),
.Y(n_2097)
);

BUFx6f_ASAP7_75t_L g2098 ( 
.A(n_137),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1227),
.Y(n_2099)
);

CKINVDCx20_ASAP7_75t_R g2100 ( 
.A(n_1504),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_1280),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1280),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1280),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1280),
.Y(n_2104)
);

INVx2_ASAP7_75t_L g2105 ( 
.A(n_1280),
.Y(n_2105)
);

INVxp33_ASAP7_75t_SL g2106 ( 
.A(n_1793),
.Y(n_2106)
);

INVxp33_ASAP7_75t_L g2107 ( 
.A(n_1919),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1801),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_1801),
.Y(n_2109)
);

INVxp67_ASAP7_75t_L g2110 ( 
.A(n_1293),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1801),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_1801),
.Y(n_2112)
);

INVxp67_ASAP7_75t_SL g2113 ( 
.A(n_1279),
.Y(n_2113)
);

INVxp67_ASAP7_75t_SL g2114 ( 
.A(n_1279),
.Y(n_2114)
);

CKINVDCx5p33_ASAP7_75t_R g2115 ( 
.A(n_1611),
.Y(n_2115)
);

INVx2_ASAP7_75t_L g2116 ( 
.A(n_1801),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1278),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1286),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1292),
.Y(n_2119)
);

CKINVDCx16_ASAP7_75t_R g2120 ( 
.A(n_1738),
.Y(n_2120)
);

HB1xp67_ASAP7_75t_L g2121 ( 
.A(n_1924),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1305),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1323),
.Y(n_2123)
);

INVxp67_ASAP7_75t_SL g2124 ( 
.A(n_1279),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1327),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1332),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_1340),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1346),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_1347),
.Y(n_2129)
);

CKINVDCx16_ASAP7_75t_R g2130 ( 
.A(n_1941),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1349),
.Y(n_2131)
);

INVxp33_ASAP7_75t_L g2132 ( 
.A(n_1776),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_1359),
.Y(n_2133)
);

INVxp33_ASAP7_75t_L g2134 ( 
.A(n_1329),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_1369),
.Y(n_2135)
);

CKINVDCx20_ASAP7_75t_R g2136 ( 
.A(n_2010),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1370),
.Y(n_2137)
);

CKINVDCx5p33_ASAP7_75t_R g2138 ( 
.A(n_1364),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1320),
.Y(n_2139)
);

INVxp33_ASAP7_75t_L g2140 ( 
.A(n_1463),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_1320),
.Y(n_2141)
);

INVxp33_ASAP7_75t_L g2142 ( 
.A(n_1516),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1382),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_1480),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_1320),
.Y(n_2145)
);

INVx2_ASAP7_75t_SL g2146 ( 
.A(n_1480),
.Y(n_2146)
);

NOR2xp67_ASAP7_75t_L g2147 ( 
.A(n_1449),
.B(n_1),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_1396),
.Y(n_2148)
);

CKINVDCx5p33_ASAP7_75t_R g2149 ( 
.A(n_1432),
.Y(n_2149)
);

INVx1_ASAP7_75t_L g2150 ( 
.A(n_1393),
.Y(n_2150)
);

INVxp33_ASAP7_75t_L g2151 ( 
.A(n_1590),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_1398),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1406),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1396),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_1413),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1415),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_1434),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_1447),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1457),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1459),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1461),
.Y(n_2161)
);

CKINVDCx5p33_ASAP7_75t_R g2162 ( 
.A(n_1433),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1472),
.Y(n_2163)
);

INVxp33_ASAP7_75t_L g2164 ( 
.A(n_1635),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_1439),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_1677),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1473),
.Y(n_2167)
);

HB1xp67_ASAP7_75t_L g2168 ( 
.A(n_1817),
.Y(n_2168)
);

INVx1_ASAP7_75t_L g2169 ( 
.A(n_1475),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_1396),
.Y(n_2170)
);

HB1xp67_ASAP7_75t_L g2171 ( 
.A(n_1970),
.Y(n_2171)
);

CKINVDCx16_ASAP7_75t_R g2172 ( 
.A(n_1465),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_1508),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1510),
.Y(n_2174)
);

CKINVDCx5p33_ASAP7_75t_R g2175 ( 
.A(n_1576),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1520),
.Y(n_2176)
);

BUFx3_ASAP7_75t_L g2177 ( 
.A(n_1493),
.Y(n_2177)
);

INVx1_ASAP7_75t_SL g2178 ( 
.A(n_1950),
.Y(n_2178)
);

INVxp67_ASAP7_75t_SL g2179 ( 
.A(n_1492),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_1531),
.Y(n_2180)
);

BUFx2_ASAP7_75t_L g2181 ( 
.A(n_1989),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1535),
.Y(n_2182)
);

INVxp67_ASAP7_75t_SL g2183 ( 
.A(n_1492),
.Y(n_2183)
);

BUFx6f_ASAP7_75t_L g2184 ( 
.A(n_1317),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1540),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1542),
.Y(n_2186)
);

CKINVDCx14_ASAP7_75t_R g2187 ( 
.A(n_1425),
.Y(n_2187)
);

INVx4_ASAP7_75t_R g2188 ( 
.A(n_1730),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1543),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1545),
.Y(n_2190)
);

INVx1_ASAP7_75t_SL g2191 ( 
.A(n_1295),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_1760),
.B(n_1),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1548),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1552),
.Y(n_2194)
);

CKINVDCx5p33_ASAP7_75t_R g2195 ( 
.A(n_1877),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1554),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1561),
.Y(n_2197)
);

CKINVDCx20_ASAP7_75t_R g2198 ( 
.A(n_1273),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_1563),
.Y(n_2199)
);

INVxp33_ASAP7_75t_SL g2200 ( 
.A(n_1421),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1566),
.Y(n_2201)
);

HB1xp67_ASAP7_75t_L g2202 ( 
.A(n_1905),
.Y(n_2202)
);

INVxp33_ASAP7_75t_SL g2203 ( 
.A(n_1276),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_1492),
.Y(n_2204)
);

BUFx3_ASAP7_75t_L g2205 ( 
.A(n_1795),
.Y(n_2205)
);

INVx1_ASAP7_75t_L g2206 ( 
.A(n_1571),
.Y(n_2206)
);

NOR2xp33_ASAP7_75t_L g2207 ( 
.A(n_1937),
.B(n_3),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_1577),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_1580),
.Y(n_2209)
);

INVxp33_ASAP7_75t_SL g2210 ( 
.A(n_1282),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_1582),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_1599),
.Y(n_2212)
);

BUFx3_ASAP7_75t_L g2213 ( 
.A(n_2015),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_1601),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_1612),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1615),
.Y(n_2216)
);

CKINVDCx14_ASAP7_75t_R g2217 ( 
.A(n_1497),
.Y(n_2217)
);

CKINVDCx5p33_ASAP7_75t_R g2218 ( 
.A(n_2019),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1616),
.Y(n_2219)
);

BUFx3_ASAP7_75t_L g2220 ( 
.A(n_1274),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1620),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1622),
.Y(n_2222)
);

INVxp67_ASAP7_75t_SL g2223 ( 
.A(n_1511),
.Y(n_2223)
);

CKINVDCx20_ASAP7_75t_R g2224 ( 
.A(n_1361),
.Y(n_2224)
);

INVxp67_ASAP7_75t_SL g2225 ( 
.A(n_1511),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1640),
.Y(n_2226)
);

CKINVDCx20_ASAP7_75t_R g2227 ( 
.A(n_1390),
.Y(n_2227)
);

HB1xp67_ASAP7_75t_L g2228 ( 
.A(n_1411),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_1648),
.Y(n_2229)
);

INVxp67_ASAP7_75t_SL g2230 ( 
.A(n_1511),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1655),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1656),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_1658),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1661),
.Y(n_2234)
);

BUFx3_ASAP7_75t_L g2235 ( 
.A(n_1274),
.Y(n_2235)
);

HB1xp67_ASAP7_75t_L g2236 ( 
.A(n_1287),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1668),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1672),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_1641),
.Y(n_2239)
);

CKINVDCx5p33_ASAP7_75t_R g2240 ( 
.A(n_1417),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1679),
.Y(n_2241)
);

BUFx6f_ASAP7_75t_L g2242 ( 
.A(n_1317),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_1681),
.Y(n_2243)
);

INVxp67_ASAP7_75t_SL g2244 ( 
.A(n_1641),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1684),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_1690),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_1466),
.Y(n_2247)
);

CKINVDCx5p33_ASAP7_75t_R g2248 ( 
.A(n_1491),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1696),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_1699),
.Y(n_2250)
);

INVxp33_ASAP7_75t_SL g2251 ( 
.A(n_1296),
.Y(n_2251)
);

BUFx2_ASAP7_75t_SL g2252 ( 
.A(n_1384),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1704),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_1705),
.Y(n_2254)
);

CKINVDCx20_ASAP7_75t_R g2255 ( 
.A(n_1544),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1706),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_1721),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_1734),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_1740),
.Y(n_2259)
);

INVxp33_ASAP7_75t_SL g2260 ( 
.A(n_1306),
.Y(n_2260)
);

INVxp33_ASAP7_75t_L g2261 ( 
.A(n_1283),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1772),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_1774),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1775),
.Y(n_2264)
);

INVxp67_ASAP7_75t_SL g2265 ( 
.A(n_1641),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1778),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_1779),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2184),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_2184),
.Y(n_2269)
);

BUFx6f_ASAP7_75t_L g2270 ( 
.A(n_2184),
.Y(n_2270)
);

INVx4_ASAP7_75t_L g2271 ( 
.A(n_2220),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2113),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2114),
.Y(n_2273)
);

BUFx3_ASAP7_75t_L g2274 ( 
.A(n_2235),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_2242),
.Y(n_2275)
);

INVx5_ASAP7_75t_L g2276 ( 
.A(n_2172),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_SL g2277 ( 
.A(n_2120),
.B(n_2130),
.Y(n_2277)
);

NAND2xp5_ASAP7_75t_L g2278 ( 
.A(n_2187),
.B(n_1289),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2217),
.B(n_1309),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2261),
.B(n_1294),
.Y(n_2280)
);

AND2x4_ASAP7_75t_L g2281 ( 
.A(n_2177),
.B(n_1352),
.Y(n_2281)
);

INVx2_ASAP7_75t_SL g2282 ( 
.A(n_2205),
.Y(n_2282)
);

INVxp67_ASAP7_75t_L g2283 ( 
.A(n_2252),
.Y(n_2283)
);

BUFx6f_ASAP7_75t_L g2284 ( 
.A(n_2242),
.Y(n_2284)
);

BUFx6f_ASAP7_75t_L g2285 ( 
.A(n_2242),
.Y(n_2285)
);

OAI22xp5_ASAP7_75t_L g2286 ( 
.A1(n_2110),
.A2(n_1302),
.B1(n_1403),
.B2(n_1315),
.Y(n_2286)
);

BUFx3_ASAP7_75t_L g2287 ( 
.A(n_2101),
.Y(n_2287)
);

AND2x4_ASAP7_75t_L g2288 ( 
.A(n_2213),
.B(n_2144),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2124),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_2179),
.B(n_1360),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_2139),
.Y(n_2291)
);

AOI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2106),
.A2(n_1467),
.B1(n_1519),
.B2(n_1442),
.Y(n_2292)
);

INVx4_ASAP7_75t_L g2293 ( 
.A(n_2138),
.Y(n_2293)
);

OAI21x1_ASAP7_75t_L g2294 ( 
.A1(n_2105),
.A2(n_1902),
.B(n_1598),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_2183),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2223),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2134),
.B(n_1513),
.Y(n_2297)
);

INVx4_ASAP7_75t_L g2298 ( 
.A(n_2149),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2225),
.B(n_1940),
.Y(n_2299)
);

INVx1_ASAP7_75t_L g2300 ( 
.A(n_2230),
.Y(n_2300)
);

INVx2_ASAP7_75t_L g2301 ( 
.A(n_2108),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2116),
.Y(n_2302)
);

BUFx3_ASAP7_75t_L g2303 ( 
.A(n_2102),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2244),
.Y(n_2304)
);

INVx3_ASAP7_75t_L g2305 ( 
.A(n_2141),
.Y(n_2305)
);

INVxp33_ASAP7_75t_SL g2306 ( 
.A(n_2240),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_2103),
.Y(n_2307)
);

INVx1_ASAP7_75t_L g2308 ( 
.A(n_2265),
.Y(n_2308)
);

INVx3_ASAP7_75t_L g2309 ( 
.A(n_2145),
.Y(n_2309)
);

INVx3_ASAP7_75t_L g2310 ( 
.A(n_2148),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2154),
.Y(n_2311)
);

BUFx6f_ASAP7_75t_L g2312 ( 
.A(n_2170),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2204),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2104),
.B(n_2050),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2109),
.Y(n_2315)
);

BUFx3_ASAP7_75t_L g2316 ( 
.A(n_2111),
.Y(n_2316)
);

INVx5_ASAP7_75t_L g2317 ( 
.A(n_2181),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2112),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_L g2319 ( 
.A(n_2239),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2140),
.B(n_1384),
.Y(n_2320)
);

BUFx6f_ASAP7_75t_L g2321 ( 
.A(n_2117),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_2118),
.Y(n_2322)
);

AND2x4_ASAP7_75t_L g2323 ( 
.A(n_2146),
.B(n_1372),
.Y(n_2323)
);

INVx1_ASAP7_75t_L g2324 ( 
.A(n_2119),
.Y(n_2324)
);

INVx5_ASAP7_75t_L g2325 ( 
.A(n_2192),
.Y(n_2325)
);

INVx5_ASAP7_75t_L g2326 ( 
.A(n_2142),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2122),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_L g2328 ( 
.A1(n_2151),
.A2(n_1570),
.B1(n_1606),
.B2(n_1530),
.Y(n_2328)
);

BUFx12f_ASAP7_75t_L g2329 ( 
.A(n_2115),
.Y(n_2329)
);

INVx4_ASAP7_75t_L g2330 ( 
.A(n_2162),
.Y(n_2330)
);

BUFx6f_ASAP7_75t_L g2331 ( 
.A(n_2123),
.Y(n_2331)
);

AND2x6_ASAP7_75t_L g2332 ( 
.A(n_2125),
.B(n_1431),
.Y(n_2332)
);

BUFx6f_ASAP7_75t_L g2333 ( 
.A(n_2126),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2127),
.Y(n_2334)
);

OA21x2_ASAP7_75t_L g2335 ( 
.A1(n_2128),
.A2(n_1290),
.B(n_1277),
.Y(n_2335)
);

AOI22xp5_ASAP7_75t_L g2336 ( 
.A1(n_2164),
.A2(n_1609),
.B1(n_1649),
.B2(n_1607),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2129),
.Y(n_2337)
);

BUFx2_ASAP7_75t_L g2338 ( 
.A(n_2165),
.Y(n_2338)
);

AND2x4_ASAP7_75t_L g2339 ( 
.A(n_2202),
.B(n_1437),
.Y(n_2339)
);

CKINVDCx6p67_ASAP7_75t_R g2340 ( 
.A(n_2100),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2131),
.Y(n_2341)
);

INVx5_ASAP7_75t_L g2342 ( 
.A(n_2132),
.Y(n_2342)
);

INVxp33_ASAP7_75t_SL g2343 ( 
.A(n_2247),
.Y(n_2343)
);

CKINVDCx5p33_ASAP7_75t_R g2344 ( 
.A(n_2248),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2133),
.Y(n_2345)
);

INVx5_ASAP7_75t_L g2346 ( 
.A(n_2107),
.Y(n_2346)
);

AND2x2_ASAP7_75t_SL g2347 ( 
.A(n_2207),
.B(n_1300),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_2135),
.Y(n_2348)
);

INVx2_ASAP7_75t_L g2349 ( 
.A(n_2137),
.Y(n_2349)
);

AOI22xp5_ASAP7_75t_L g2350 ( 
.A1(n_2175),
.A2(n_1683),
.B1(n_1716),
.B2(n_1665),
.Y(n_2350)
);

BUFx2_ASAP7_75t_L g2351 ( 
.A(n_2195),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2143),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2150),
.Y(n_2353)
);

BUFx6f_ASAP7_75t_L g2354 ( 
.A(n_2152),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_2218),
.Y(n_2355)
);

BUFx6f_ASAP7_75t_L g2356 ( 
.A(n_2153),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_2236),
.B(n_1446),
.Y(n_2357)
);

BUFx6f_ASAP7_75t_L g2358 ( 
.A(n_2155),
.Y(n_2358)
);

INVx2_ASAP7_75t_L g2359 ( 
.A(n_2156),
.Y(n_2359)
);

BUFx6f_ASAP7_75t_L g2360 ( 
.A(n_2157),
.Y(n_2360)
);

BUFx3_ASAP7_75t_L g2361 ( 
.A(n_2158),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2159),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2160),
.Y(n_2363)
);

BUFx3_ASAP7_75t_L g2364 ( 
.A(n_2161),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2163),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_2191),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2167),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2169),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2173),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2174),
.Y(n_2370)
);

INVx2_ASAP7_75t_L g2371 ( 
.A(n_2176),
.Y(n_2371)
);

AOI22xp5_ASAP7_75t_L g2372 ( 
.A1(n_2203),
.A2(n_1736),
.B1(n_1766),
.B2(n_1719),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2180),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_2182),
.Y(n_2374)
);

NOR2x1_ASAP7_75t_L g2375 ( 
.A(n_2185),
.B(n_1584),
.Y(n_2375)
);

AND2x4_ASAP7_75t_L g2376 ( 
.A(n_2166),
.B(n_2168),
.Y(n_2376)
);

INVx5_ASAP7_75t_L g2377 ( 
.A(n_2200),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_L g2378 ( 
.A(n_2186),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2189),
.Y(n_2379)
);

BUFx6f_ASAP7_75t_L g2380 ( 
.A(n_2190),
.Y(n_2380)
);

INVx5_ASAP7_75t_L g2381 ( 
.A(n_2136),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2193),
.Y(n_2382)
);

BUFx6f_ASAP7_75t_L g2383 ( 
.A(n_2194),
.Y(n_2383)
);

OR2x2_ASAP7_75t_L g2384 ( 
.A(n_2171),
.B(n_1780),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_L g2385 ( 
.A(n_2196),
.Y(n_2385)
);

INVxp67_ASAP7_75t_L g2386 ( 
.A(n_2228),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2197),
.B(n_1291),
.Y(n_2387)
);

INVx3_ASAP7_75t_L g2388 ( 
.A(n_2199),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2201),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_2206),
.Y(n_2390)
);

BUFx12f_ASAP7_75t_L g2391 ( 
.A(n_2188),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2210),
.B(n_1598),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2208),
.Y(n_2393)
);

BUFx8_ASAP7_75t_L g2394 ( 
.A(n_2209),
.Y(n_2394)
);

OAI22x1_ASAP7_75t_L g2395 ( 
.A1(n_2178),
.A2(n_1304),
.B1(n_1334),
.B2(n_1288),
.Y(n_2395)
);

BUFx2_ASAP7_75t_L g2396 ( 
.A(n_2198),
.Y(n_2396)
);

AND2x6_ASAP7_75t_L g2397 ( 
.A(n_2211),
.B(n_1575),
.Y(n_2397)
);

BUFx6f_ASAP7_75t_L g2398 ( 
.A(n_2212),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2214),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2215),
.B(n_1298),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2216),
.Y(n_2401)
);

INVx4_ASAP7_75t_L g2402 ( 
.A(n_2121),
.Y(n_2402)
);

HB1xp67_ASAP7_75t_L g2403 ( 
.A(n_2251),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2219),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2221),
.Y(n_2405)
);

INVx5_ASAP7_75t_L g2406 ( 
.A(n_2260),
.Y(n_2406)
);

BUFx8_ASAP7_75t_L g2407 ( 
.A(n_2222),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2226),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2229),
.B(n_1509),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_2231),
.Y(n_2410)
);

OA21x2_ASAP7_75t_L g2411 ( 
.A1(n_2232),
.A2(n_1313),
.B(n_1303),
.Y(n_2411)
);

AOI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_2147),
.A2(n_1825),
.B1(n_1880),
.B2(n_1808),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2233),
.Y(n_2413)
);

BUFx3_ASAP7_75t_L g2414 ( 
.A(n_2234),
.Y(n_2414)
);

INVx2_ASAP7_75t_L g2415 ( 
.A(n_2237),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2238),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2241),
.B(n_1331),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2243),
.B(n_1335),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2245),
.Y(n_2419)
);

CKINVDCx11_ASAP7_75t_R g2420 ( 
.A(n_2224),
.Y(n_2420)
);

AOI22xp5_ASAP7_75t_L g2421 ( 
.A1(n_2227),
.A2(n_1926),
.B1(n_1951),
.B2(n_1913),
.Y(n_2421)
);

BUFx2_ASAP7_75t_L g2422 ( 
.A(n_2255),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2246),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_2249),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2250),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2253),
.Y(n_2426)
);

CKINVDCx6p67_ASAP7_75t_R g2427 ( 
.A(n_2254),
.Y(n_2427)
);

AND2x4_ASAP7_75t_L g2428 ( 
.A(n_2256),
.B(n_1619),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_2257),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2258),
.Y(n_2430)
);

BUFx6f_ASAP7_75t_L g2431 ( 
.A(n_2259),
.Y(n_2431)
);

BUFx3_ASAP7_75t_L g2432 ( 
.A(n_2262),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2263),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2264),
.B(n_1339),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_2266),
.B(n_1902),
.Y(n_2435)
);

NAND2xp5_ASAP7_75t_L g2436 ( 
.A(n_2267),
.B(n_1342),
.Y(n_2436)
);

BUFx6f_ASAP7_75t_L g2437 ( 
.A(n_2184),
.Y(n_2437)
);

CKINVDCx5p33_ASAP7_75t_R g2438 ( 
.A(n_2240),
.Y(n_2438)
);

AND2x2_ASAP7_75t_L g2439 ( 
.A(n_2261),
.B(n_1509),
.Y(n_2439)
);

BUFx6f_ASAP7_75t_L g2440 ( 
.A(n_2184),
.Y(n_2440)
);

BUFx6f_ASAP7_75t_L g2441 ( 
.A(n_2184),
.Y(n_2441)
);

AND2x4_ASAP7_75t_L g2442 ( 
.A(n_2220),
.B(n_1700),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2184),
.Y(n_2443)
);

BUFx6f_ASAP7_75t_L g2444 ( 
.A(n_2184),
.Y(n_2444)
);

BUFx3_ASAP7_75t_L g2445 ( 
.A(n_2220),
.Y(n_2445)
);

AOI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_2106),
.A2(n_1974),
.B1(n_1980),
.B2(n_1966),
.Y(n_2446)
);

BUFx6f_ASAP7_75t_L g2447 ( 
.A(n_2184),
.Y(n_2447)
);

OAI21x1_ASAP7_75t_L g2448 ( 
.A1(n_2105),
.A2(n_1366),
.B(n_1350),
.Y(n_2448)
);

AND2x6_ASAP7_75t_L g2449 ( 
.A(n_2192),
.B(n_1985),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2113),
.Y(n_2450)
);

INVx2_ASAP7_75t_L g2451 ( 
.A(n_2184),
.Y(n_2451)
);

INVx3_ASAP7_75t_L g2452 ( 
.A(n_2220),
.Y(n_2452)
);

NAND2xp5_ASAP7_75t_L g2453 ( 
.A(n_2187),
.B(n_1375),
.Y(n_2453)
);

AOI22x1_ASAP7_75t_SL g2454 ( 
.A1(n_2198),
.A2(n_2070),
.B1(n_2072),
.B2(n_2056),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_2184),
.Y(n_2455)
);

OAI21x1_ASAP7_75t_L g2456 ( 
.A1(n_2105),
.A2(n_1404),
.B(n_1381),
.Y(n_2456)
);

BUFx6f_ASAP7_75t_L g2457 ( 
.A(n_2184),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2113),
.Y(n_2458)
);

BUFx3_ASAP7_75t_L g2459 ( 
.A(n_2220),
.Y(n_2459)
);

INVx2_ASAP7_75t_SL g2460 ( 
.A(n_2220),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2184),
.Y(n_2461)
);

INVx2_ASAP7_75t_L g2462 ( 
.A(n_2184),
.Y(n_2462)
);

BUFx6f_ASAP7_75t_L g2463 ( 
.A(n_2184),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2184),
.Y(n_2464)
);

CKINVDCx6p67_ASAP7_75t_R g2465 ( 
.A(n_2120),
.Y(n_2465)
);

BUFx3_ASAP7_75t_L g2466 ( 
.A(n_2220),
.Y(n_2466)
);

INVx5_ASAP7_75t_L g2467 ( 
.A(n_2172),
.Y(n_2467)
);

NAND2xp33_ASAP7_75t_SL g2468 ( 
.A(n_2192),
.B(n_1814),
.Y(n_2468)
);

AND2x6_ASAP7_75t_L g2469 ( 
.A(n_2192),
.B(n_1991),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2261),
.B(n_1695),
.Y(n_2470)
);

INVx2_ASAP7_75t_L g2471 ( 
.A(n_2184),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2184),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2113),
.Y(n_2473)
);

OAI22xp33_ASAP7_75t_R g2474 ( 
.A1(n_2178),
.A2(n_1785),
.B1(n_1787),
.B2(n_1782),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2184),
.Y(n_2475)
);

BUFx3_ASAP7_75t_L g2476 ( 
.A(n_2220),
.Y(n_2476)
);

OAI22xp5_ASAP7_75t_SL g2477 ( 
.A1(n_2198),
.A2(n_1422),
.B1(n_1441),
.B2(n_1377),
.Y(n_2477)
);

INVx3_ASAP7_75t_L g2478 ( 
.A(n_2220),
.Y(n_2478)
);

BUFx6f_ASAP7_75t_L g2479 ( 
.A(n_2184),
.Y(n_2479)
);

AND2x4_ASAP7_75t_L g2480 ( 
.A(n_2220),
.B(n_2069),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2261),
.B(n_1695),
.Y(n_2481)
);

AND2x4_ASAP7_75t_L g2482 ( 
.A(n_2220),
.B(n_1275),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2184),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2187),
.B(n_1430),
.Y(n_2484)
);

INVxp67_ASAP7_75t_L g2485 ( 
.A(n_2252),
.Y(n_2485)
);

AOI22x1_ASAP7_75t_SL g2486 ( 
.A1(n_2198),
.A2(n_1312),
.B1(n_1316),
.B2(n_1311),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2184),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2184),
.Y(n_2488)
);

INVx3_ASAP7_75t_L g2489 ( 
.A(n_2220),
.Y(n_2489)
);

BUFx6f_ASAP7_75t_L g2490 ( 
.A(n_2184),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2184),
.Y(n_2491)
);

BUFx8_ASAP7_75t_L g2492 ( 
.A(n_2181),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2261),
.B(n_1910),
.Y(n_2493)
);

INVx1_ASAP7_75t_L g2494 ( 
.A(n_2113),
.Y(n_2494)
);

CKINVDCx5p33_ASAP7_75t_R g2495 ( 
.A(n_2240),
.Y(n_2495)
);

BUFx3_ASAP7_75t_L g2496 ( 
.A(n_2220),
.Y(n_2496)
);

INVx3_ASAP7_75t_L g2497 ( 
.A(n_2220),
.Y(n_2497)
);

AND2x2_ASAP7_75t_L g2498 ( 
.A(n_2261),
.B(n_1910),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2187),
.B(n_1440),
.Y(n_2499)
);

OA21x2_ASAP7_75t_L g2500 ( 
.A1(n_2101),
.A2(n_1471),
.B(n_1468),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2184),
.Y(n_2501)
);

NAND2xp5_ASAP7_75t_L g2502 ( 
.A(n_2187),
.B(n_1487),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2184),
.Y(n_2503)
);

CKINVDCx5p33_ASAP7_75t_R g2504 ( 
.A(n_2240),
.Y(n_2504)
);

BUFx6f_ASAP7_75t_L g2505 ( 
.A(n_2184),
.Y(n_2505)
);

BUFx6f_ASAP7_75t_L g2506 ( 
.A(n_2184),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2184),
.Y(n_2507)
);

INVx3_ASAP7_75t_L g2508 ( 
.A(n_2220),
.Y(n_2508)
);

INVx5_ASAP7_75t_L g2509 ( 
.A(n_2172),
.Y(n_2509)
);

HB1xp67_ASAP7_75t_L g2510 ( 
.A(n_2202),
.Y(n_2510)
);

NOR2x1_ASAP7_75t_L g2511 ( 
.A(n_2220),
.B(n_1627),
.Y(n_2511)
);

OA21x2_ASAP7_75t_L g2512 ( 
.A1(n_2101),
.A2(n_1500),
.B(n_1496),
.Y(n_2512)
);

BUFx2_ASAP7_75t_L g2513 ( 
.A(n_2138),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2113),
.Y(n_2514)
);

BUFx3_ASAP7_75t_L g2515 ( 
.A(n_2220),
.Y(n_2515)
);

AND2x2_ASAP7_75t_L g2516 ( 
.A(n_2261),
.B(n_2009),
.Y(n_2516)
);

INVx4_ASAP7_75t_L g2517 ( 
.A(n_2220),
.Y(n_2517)
);

BUFx12f_ASAP7_75t_L g2518 ( 
.A(n_2115),
.Y(n_2518)
);

INVx5_ASAP7_75t_L g2519 ( 
.A(n_2172),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_L g2520 ( 
.A(n_2187),
.B(n_1506),
.Y(n_2520)
);

AND2x4_ASAP7_75t_L g2521 ( 
.A(n_2220),
.B(n_1378),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2113),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2187),
.B(n_1518),
.Y(n_2523)
);

OA21x2_ASAP7_75t_L g2524 ( 
.A1(n_2101),
.A2(n_1536),
.B(n_1528),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2220),
.Y(n_2525)
);

OA21x2_ASAP7_75t_L g2526 ( 
.A1(n_2101),
.A2(n_1562),
.B(n_1558),
.Y(n_2526)
);

NOR2xp33_ASAP7_75t_L g2527 ( 
.A(n_2220),
.B(n_2073),
.Y(n_2527)
);

BUFx6f_ASAP7_75t_L g2528 ( 
.A(n_2184),
.Y(n_2528)
);

BUFx6f_ASAP7_75t_L g2529 ( 
.A(n_2184),
.Y(n_2529)
);

BUFx3_ASAP7_75t_L g2530 ( 
.A(n_2220),
.Y(n_2530)
);

OAI22x1_ASAP7_75t_R g2531 ( 
.A1(n_2115),
.A2(n_1319),
.B1(n_1321),
.B2(n_1318),
.Y(n_2531)
);

BUFx6f_ASAP7_75t_L g2532 ( 
.A(n_2184),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_2220),
.B(n_1568),
.Y(n_2533)
);

INVx4_ASAP7_75t_L g2534 ( 
.A(n_2220),
.Y(n_2534)
);

HB1xp67_ASAP7_75t_L g2535 ( 
.A(n_2202),
.Y(n_2535)
);

AOI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_2106),
.A2(n_1583),
.B1(n_1643),
.B2(n_1578),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2202),
.Y(n_2537)
);

BUFx3_ASAP7_75t_L g2538 ( 
.A(n_2220),
.Y(n_2538)
);

OAI22xp5_ASAP7_75t_L g2539 ( 
.A1(n_2110),
.A2(n_2082),
.B1(n_1724),
.B2(n_1489),
.Y(n_2539)
);

INVxp67_ASAP7_75t_L g2540 ( 
.A(n_2252),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2113),
.Y(n_2541)
);

BUFx6f_ASAP7_75t_L g2542 ( 
.A(n_2184),
.Y(n_2542)
);

BUFx2_ASAP7_75t_L g2543 ( 
.A(n_2138),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_2240),
.Y(n_2544)
);

HB1xp67_ASAP7_75t_L g2545 ( 
.A(n_2202),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2113),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2113),
.Y(n_2547)
);

NAND2xp5_ASAP7_75t_L g2548 ( 
.A(n_2187),
.B(n_1569),
.Y(n_2548)
);

HB1xp67_ASAP7_75t_L g2549 ( 
.A(n_2202),
.Y(n_2549)
);

INVx3_ASAP7_75t_L g2550 ( 
.A(n_2220),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2220),
.B(n_1786),
.Y(n_2551)
);

AND2x2_ASAP7_75t_L g2552 ( 
.A(n_2261),
.B(n_2009),
.Y(n_2552)
);

BUFx6f_ASAP7_75t_L g2553 ( 
.A(n_2184),
.Y(n_2553)
);

BUFx3_ASAP7_75t_L g2554 ( 
.A(n_2220),
.Y(n_2554)
);

INVx1_ASAP7_75t_L g2555 ( 
.A(n_2113),
.Y(n_2555)
);

HB1xp67_ASAP7_75t_L g2556 ( 
.A(n_2202),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2184),
.Y(n_2557)
);

XNOR2x1_ASAP7_75t_L g2558 ( 
.A(n_2178),
.B(n_1481),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2113),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_L g2560 ( 
.A(n_2220),
.B(n_1572),
.Y(n_2560)
);

OAI21x1_ASAP7_75t_L g2561 ( 
.A1(n_2105),
.A2(n_1617),
.B(n_1581),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2113),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2184),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2113),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2187),
.B(n_1625),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2106),
.A2(n_1993),
.B1(n_2078),
.B2(n_1715),
.Y(n_2566)
);

INVx5_ASAP7_75t_L g2567 ( 
.A(n_2172),
.Y(n_2567)
);

BUFx8_ASAP7_75t_L g2568 ( 
.A(n_2181),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2184),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2113),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2184),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2113),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2113),
.Y(n_2573)
);

INVxp67_ASAP7_75t_L g2574 ( 
.A(n_2252),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_2220),
.B(n_1829),
.Y(n_2575)
);

BUFx6f_ASAP7_75t_L g2576 ( 
.A(n_2184),
.Y(n_2576)
);

BUFx6f_ASAP7_75t_L g2577 ( 
.A(n_2184),
.Y(n_2577)
);

BUFx6f_ASAP7_75t_L g2578 ( 
.A(n_2184),
.Y(n_2578)
);

CKINVDCx5p33_ASAP7_75t_R g2579 ( 
.A(n_2240),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_L g2580 ( 
.A(n_2184),
.Y(n_2580)
);

INVxp67_ASAP7_75t_L g2581 ( 
.A(n_2252),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2113),
.Y(n_2582)
);

INVx3_ASAP7_75t_L g2583 ( 
.A(n_2220),
.Y(n_2583)
);

AND2x4_ASAP7_75t_L g2584 ( 
.A(n_2220),
.B(n_1841),
.Y(n_2584)
);

INVx2_ASAP7_75t_L g2585 ( 
.A(n_2184),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2184),
.Y(n_2586)
);

INVx2_ASAP7_75t_L g2587 ( 
.A(n_2184),
.Y(n_2587)
);

OAI21x1_ASAP7_75t_L g2588 ( 
.A1(n_2105),
.A2(n_1634),
.B(n_1628),
.Y(n_2588)
);

BUFx6f_ASAP7_75t_L g2589 ( 
.A(n_2184),
.Y(n_2589)
);

OA21x2_ASAP7_75t_L g2590 ( 
.A1(n_2101),
.A2(n_1698),
.B(n_1644),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2220),
.Y(n_2591)
);

HB1xp67_ASAP7_75t_L g2592 ( 
.A(n_2202),
.Y(n_2592)
);

AND2x4_ASAP7_75t_L g2593 ( 
.A(n_2220),
.B(n_1856),
.Y(n_2593)
);

AOI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2106),
.A2(n_1534),
.B1(n_1560),
.B2(n_1512),
.Y(n_2594)
);

INVx2_ASAP7_75t_L g2595 ( 
.A(n_2184),
.Y(n_2595)
);

CKINVDCx5p33_ASAP7_75t_R g2596 ( 
.A(n_2344),
.Y(n_2596)
);

HB1xp67_ASAP7_75t_L g2597 ( 
.A(n_2326),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_2276),
.B(n_2040),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2322),
.Y(n_2599)
);

CKINVDCx5p33_ASAP7_75t_R g2600 ( 
.A(n_2438),
.Y(n_2600)
);

AND2x6_ASAP7_75t_L g2601 ( 
.A(n_2409),
.B(n_1707),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2346),
.Y(n_2602)
);

INVxp67_ASAP7_75t_L g2603 ( 
.A(n_2366),
.Y(n_2603)
);

CKINVDCx5p33_ASAP7_75t_R g2604 ( 
.A(n_2495),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2321),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2280),
.B(n_1503),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2341),
.Y(n_2607)
);

CKINVDCx5p33_ASAP7_75t_R g2608 ( 
.A(n_2504),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2301),
.Y(n_2609)
);

CKINVDCx5p33_ASAP7_75t_R g2610 ( 
.A(n_2544),
.Y(n_2610)
);

CKINVDCx20_ASAP7_75t_R g2611 ( 
.A(n_2420),
.Y(n_2611)
);

INVx2_ASAP7_75t_L g2612 ( 
.A(n_2302),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2297),
.B(n_1503),
.Y(n_2613)
);

INVxp67_ASAP7_75t_L g2614 ( 
.A(n_2439),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2291),
.Y(n_2615)
);

NAND2xp5_ASAP7_75t_SL g2616 ( 
.A(n_2392),
.B(n_1322),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2345),
.Y(n_2617)
);

NOR2x1_ASAP7_75t_L g2618 ( 
.A(n_2293),
.B(n_1669),
.Y(n_2618)
);

AND2x4_ASAP7_75t_L g2619 ( 
.A(n_2467),
.B(n_2092),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2349),
.Y(n_2620)
);

INVx3_ASAP7_75t_L g2621 ( 
.A(n_2331),
.Y(n_2621)
);

CKINVDCx5p33_ASAP7_75t_R g2622 ( 
.A(n_2579),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2359),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2338),
.Y(n_2624)
);

OR2x2_ASAP7_75t_L g2625 ( 
.A(n_2376),
.B(n_1675),
.Y(n_2625)
);

BUFx3_ASAP7_75t_L g2626 ( 
.A(n_2391),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2368),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2369),
.Y(n_2628)
);

HB1xp67_ASAP7_75t_L g2629 ( 
.A(n_2510),
.Y(n_2629)
);

CKINVDCx5p33_ASAP7_75t_R g2630 ( 
.A(n_2306),
.Y(n_2630)
);

INVxp67_ASAP7_75t_L g2631 ( 
.A(n_2470),
.Y(n_2631)
);

BUFx2_ASAP7_75t_L g2632 ( 
.A(n_2351),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2535),
.Y(n_2633)
);

CKINVDCx5p33_ASAP7_75t_R g2634 ( 
.A(n_2343),
.Y(n_2634)
);

INVx2_ASAP7_75t_L g2635 ( 
.A(n_2312),
.Y(n_2635)
);

XNOR2xp5_ASAP7_75t_L g2636 ( 
.A(n_2536),
.B(n_1697),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2319),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2311),
.Y(n_2638)
);

INVx2_ASAP7_75t_L g2639 ( 
.A(n_2313),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2305),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2309),
.Y(n_2641)
);

NOR2xp67_ASAP7_75t_L g2642 ( 
.A(n_2509),
.B(n_1524),
.Y(n_2642)
);

CKINVDCx5p33_ASAP7_75t_R g2643 ( 
.A(n_2329),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2371),
.Y(n_2644)
);

BUFx2_ASAP7_75t_L g2645 ( 
.A(n_2513),
.Y(n_2645)
);

HB1xp67_ASAP7_75t_L g2646 ( 
.A(n_2537),
.Y(n_2646)
);

BUFx2_ASAP7_75t_L g2647 ( 
.A(n_2543),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2481),
.B(n_1605),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2379),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2405),
.Y(n_2650)
);

CKINVDCx5p33_ASAP7_75t_R g2651 ( 
.A(n_2518),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2415),
.Y(n_2652)
);

CKINVDCx20_ASAP7_75t_R g2653 ( 
.A(n_2465),
.Y(n_2653)
);

INVx2_ASAP7_75t_L g2654 ( 
.A(n_2310),
.Y(n_2654)
);

INVx3_ASAP7_75t_L g2655 ( 
.A(n_2333),
.Y(n_2655)
);

HB1xp67_ASAP7_75t_L g2656 ( 
.A(n_2545),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2425),
.Y(n_2657)
);

BUFx3_ASAP7_75t_L g2658 ( 
.A(n_2274),
.Y(n_2658)
);

NOR2xp33_ASAP7_75t_R g2659 ( 
.A(n_2340),
.B(n_1272),
.Y(n_2659)
);

BUFx2_ASAP7_75t_L g2660 ( 
.A(n_2492),
.Y(n_2660)
);

AND2x4_ASAP7_75t_L g2661 ( 
.A(n_2519),
.B(n_2567),
.Y(n_2661)
);

CKINVDCx5p33_ASAP7_75t_R g2662 ( 
.A(n_2396),
.Y(n_2662)
);

BUFx6f_ASAP7_75t_L g2663 ( 
.A(n_2269),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2348),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2268),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2549),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2354),
.Y(n_2667)
);

INVx1_ASAP7_75t_L g2668 ( 
.A(n_2356),
.Y(n_2668)
);

CKINVDCx5p33_ASAP7_75t_R g2669 ( 
.A(n_2422),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2381),
.Y(n_2670)
);

CKINVDCx5p33_ASAP7_75t_R g2671 ( 
.A(n_2403),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2358),
.Y(n_2672)
);

INVx1_ASAP7_75t_L g2673 ( 
.A(n_2360),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2556),
.Y(n_2674)
);

XOR2xp5_ASAP7_75t_L g2675 ( 
.A(n_2558),
.B(n_1325),
.Y(n_2675)
);

CKINVDCx5p33_ASAP7_75t_R g2676 ( 
.A(n_2568),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2374),
.Y(n_2677)
);

AND2x6_ASAP7_75t_L g2678 ( 
.A(n_2493),
.B(n_1710),
.Y(n_2678)
);

CKINVDCx5p33_ASAP7_75t_R g2679 ( 
.A(n_2406),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2443),
.Y(n_2680)
);

OR2x2_ASAP7_75t_L g2681 ( 
.A(n_2592),
.B(n_1703),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2378),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2380),
.Y(n_2683)
);

BUFx2_ASAP7_75t_L g2684 ( 
.A(n_2317),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2383),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2385),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2398),
.Y(n_2687)
);

CKINVDCx5p33_ASAP7_75t_R g2688 ( 
.A(n_2355),
.Y(n_2688)
);

AND2x4_ASAP7_75t_L g2689 ( 
.A(n_2452),
.B(n_1761),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2451),
.Y(n_2690)
);

BUFx2_ASAP7_75t_L g2691 ( 
.A(n_2282),
.Y(n_2691)
);

INVx1_ASAP7_75t_L g2692 ( 
.A(n_2404),
.Y(n_2692)
);

BUFx6f_ASAP7_75t_L g2693 ( 
.A(n_2270),
.Y(n_2693)
);

OAI21x1_ASAP7_75t_L g2694 ( 
.A1(n_2294),
.A2(n_1718),
.B(n_1713),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2461),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2410),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2424),
.Y(n_2697)
);

OAI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2347),
.A2(n_1328),
.B1(n_1333),
.B2(n_1326),
.Y(n_2698)
);

CKINVDCx20_ASAP7_75t_R g2699 ( 
.A(n_2427),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2431),
.Y(n_2700)
);

CKINVDCx5p33_ASAP7_75t_R g2701 ( 
.A(n_2328),
.Y(n_2701)
);

INVx6_ASAP7_75t_L g2702 ( 
.A(n_2342),
.Y(n_2702)
);

NOR2xp33_ASAP7_75t_R g2703 ( 
.A(n_2478),
.B(n_1281),
.Y(n_2703)
);

INVx3_ASAP7_75t_L g2704 ( 
.A(n_2352),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2324),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2327),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2462),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2334),
.Y(n_2708)
);

INVx1_ASAP7_75t_L g2709 ( 
.A(n_2337),
.Y(n_2709)
);

HB1xp67_ASAP7_75t_L g2710 ( 
.A(n_2286),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2353),
.Y(n_2711)
);

AND2x2_ASAP7_75t_L g2712 ( 
.A(n_2498),
.B(n_1605),
.Y(n_2712)
);

INVx2_ASAP7_75t_L g2713 ( 
.A(n_2464),
.Y(n_2713)
);

CKINVDCx5p33_ASAP7_75t_R g2714 ( 
.A(n_2298),
.Y(n_2714)
);

NAND2xp33_ASAP7_75t_R g2715 ( 
.A(n_2288),
.B(n_1336),
.Y(n_2715)
);

INVx1_ASAP7_75t_L g2716 ( 
.A(n_2362),
.Y(n_2716)
);

CKINVDCx5p33_ASAP7_75t_R g2717 ( 
.A(n_2330),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_2445),
.Y(n_2718)
);

INVx2_ASAP7_75t_L g2719 ( 
.A(n_2471),
.Y(n_2719)
);

INVx1_ASAP7_75t_L g2720 ( 
.A(n_2363),
.Y(n_2720)
);

NAND2xp5_ASAP7_75t_L g2721 ( 
.A(n_2314),
.B(n_1367),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2472),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2365),
.Y(n_2723)
);

CKINVDCx5p33_ASAP7_75t_R g2724 ( 
.A(n_2459),
.Y(n_2724)
);

INVx3_ASAP7_75t_L g2725 ( 
.A(n_2361),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2475),
.Y(n_2726)
);

BUFx6f_ASAP7_75t_L g2727 ( 
.A(n_2275),
.Y(n_2727)
);

INVx3_ASAP7_75t_L g2728 ( 
.A(n_2364),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2466),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2367),
.Y(n_2730)
);

BUFx6f_ASAP7_75t_L g2731 ( 
.A(n_2284),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2370),
.Y(n_2732)
);

BUFx6f_ASAP7_75t_L g2733 ( 
.A(n_2285),
.Y(n_2733)
);

INVxp67_ASAP7_75t_L g2734 ( 
.A(n_2516),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2315),
.B(n_1409),
.Y(n_2735)
);

CKINVDCx5p33_ASAP7_75t_R g2736 ( 
.A(n_2476),
.Y(n_2736)
);

BUFx6f_ASAP7_75t_L g2737 ( 
.A(n_2437),
.Y(n_2737)
);

CKINVDCx5p33_ASAP7_75t_R g2738 ( 
.A(n_2496),
.Y(n_2738)
);

CKINVDCx5p33_ASAP7_75t_R g2739 ( 
.A(n_2515),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2373),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2382),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2389),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2483),
.Y(n_2743)
);

NAND2xp5_ASAP7_75t_SL g2744 ( 
.A(n_2283),
.B(n_1337),
.Y(n_2744)
);

INVx3_ASAP7_75t_L g2745 ( 
.A(n_2414),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2390),
.Y(n_2746)
);

INVx3_ASAP7_75t_L g2747 ( 
.A(n_2429),
.Y(n_2747)
);

NAND2xp33_ASAP7_75t_SL g2748 ( 
.A(n_2460),
.B(n_1341),
.Y(n_2748)
);

AND2x4_ASAP7_75t_L g2749 ( 
.A(n_2489),
.B(n_1771),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_2487),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2393),
.Y(n_2751)
);

BUFx6f_ASAP7_75t_L g2752 ( 
.A(n_2440),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2386),
.Y(n_2753)
);

BUFx6f_ASAP7_75t_L g2754 ( 
.A(n_2441),
.Y(n_2754)
);

CKINVDCx5p33_ASAP7_75t_R g2755 ( 
.A(n_2530),
.Y(n_2755)
);

INVx1_ASAP7_75t_L g2756 ( 
.A(n_2399),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_SL g2757 ( 
.A(n_2485),
.B(n_1344),
.Y(n_2757)
);

CKINVDCx5p33_ASAP7_75t_R g2758 ( 
.A(n_2538),
.Y(n_2758)
);

CKINVDCx20_ASAP7_75t_R g2759 ( 
.A(n_2566),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2401),
.Y(n_2760)
);

CKINVDCx20_ASAP7_75t_R g2761 ( 
.A(n_2554),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2488),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2491),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2408),
.Y(n_2764)
);

CKINVDCx20_ASAP7_75t_R g2765 ( 
.A(n_2421),
.Y(n_2765)
);

AND2x6_ASAP7_75t_L g2766 ( 
.A(n_2552),
.B(n_1725),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2413),
.Y(n_2767)
);

AND2x4_ASAP7_75t_L g2768 ( 
.A(n_2497),
.B(n_1823),
.Y(n_2768)
);

HB1xp67_ASAP7_75t_L g2769 ( 
.A(n_2320),
.Y(n_2769)
);

CKINVDCx5p33_ASAP7_75t_R g2770 ( 
.A(n_2377),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2318),
.B(n_1444),
.Y(n_2771)
);

NAND2xp5_ASAP7_75t_SL g2772 ( 
.A(n_2540),
.B(n_1345),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2501),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2508),
.B(n_1632),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2416),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2402),
.Y(n_2776)
);

INVx3_ASAP7_75t_L g2777 ( 
.A(n_2432),
.Y(n_2777)
);

CKINVDCx20_ASAP7_75t_R g2778 ( 
.A(n_2350),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2419),
.Y(n_2779)
);

OR2x6_ASAP7_75t_L g2780 ( 
.A(n_2277),
.B(n_1362),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2423),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_2525),
.Y(n_2782)
);

CKINVDCx5p33_ASAP7_75t_R g2783 ( 
.A(n_2550),
.Y(n_2783)
);

BUFx6f_ASAP7_75t_L g2784 ( 
.A(n_2444),
.Y(n_2784)
);

AND2x4_ASAP7_75t_L g2785 ( 
.A(n_2583),
.B(n_1903),
.Y(n_2785)
);

OA21x2_ASAP7_75t_L g2786 ( 
.A1(n_2448),
.A2(n_1735),
.B(n_1733),
.Y(n_2786)
);

CKINVDCx20_ASAP7_75t_R g2787 ( 
.A(n_2372),
.Y(n_2787)
);

NAND2xp33_ASAP7_75t_L g2788 ( 
.A(n_2449),
.B(n_1814),
.Y(n_2788)
);

INVx1_ASAP7_75t_L g2789 ( 
.A(n_2426),
.Y(n_2789)
);

NOR2xp33_ASAP7_75t_L g2790 ( 
.A(n_2453),
.B(n_2484),
.Y(n_2790)
);

NOR2xp33_ASAP7_75t_L g2791 ( 
.A(n_2499),
.B(n_1742),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2287),
.B(n_1533),
.Y(n_2792)
);

INVx2_ASAP7_75t_L g2793 ( 
.A(n_2503),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2433),
.Y(n_2794)
);

CKINVDCx5p33_ASAP7_75t_R g2795 ( 
.A(n_2591),
.Y(n_2795)
);

INVx1_ASAP7_75t_L g2796 ( 
.A(n_2272),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2430),
.B(n_1632),
.Y(n_2797)
);

NOR2xp33_ASAP7_75t_R g2798 ( 
.A(n_2468),
.B(n_1285),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2273),
.Y(n_2799)
);

CKINVDCx5p33_ASAP7_75t_R g2800 ( 
.A(n_2486),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2303),
.B(n_1682),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_R g2802 ( 
.A(n_2388),
.B(n_1297),
.Y(n_2802)
);

CKINVDCx5p33_ASAP7_75t_R g2803 ( 
.A(n_2574),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2339),
.B(n_1741),
.Y(n_2804)
);

INVx2_ASAP7_75t_L g2805 ( 
.A(n_2507),
.Y(n_2805)
);

CKINVDCx5p33_ASAP7_75t_R g2806 ( 
.A(n_2581),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_SL g2807 ( 
.A(n_2325),
.B(n_1348),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2289),
.Y(n_2808)
);

INVx1_ASAP7_75t_L g2809 ( 
.A(n_2295),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2296),
.Y(n_2810)
);

CKINVDCx5p33_ASAP7_75t_R g2811 ( 
.A(n_2271),
.Y(n_2811)
);

INVxp67_ASAP7_75t_SL g2812 ( 
.A(n_2307),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2300),
.Y(n_2813)
);

CKINVDCx5p33_ASAP7_75t_R g2814 ( 
.A(n_2517),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2304),
.Y(n_2815)
);

NAND2xp5_ASAP7_75t_L g2816 ( 
.A(n_2316),
.B(n_1798),
.Y(n_2816)
);

INVxp67_ASAP7_75t_L g2817 ( 
.A(n_2527),
.Y(n_2817)
);

AND2x6_ASAP7_75t_L g2818 ( 
.A(n_2375),
.B(n_1799),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2299),
.B(n_1899),
.Y(n_2819)
);

INVx1_ASAP7_75t_L g2820 ( 
.A(n_2308),
.Y(n_2820)
);

INVx2_ASAP7_75t_L g2821 ( 
.A(n_2563),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2450),
.B(n_1998),
.Y(n_2822)
);

OAI21x1_ASAP7_75t_L g2823 ( 
.A1(n_2456),
.A2(n_1810),
.B(n_1803),
.Y(n_2823)
);

CKINVDCx5p33_ASAP7_75t_R g2824 ( 
.A(n_2534),
.Y(n_2824)
);

OA21x2_ASAP7_75t_L g2825 ( 
.A1(n_2561),
.A2(n_1827),
.B(n_1818),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2447),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2458),
.Y(n_2827)
);

INVx3_ASAP7_75t_L g2828 ( 
.A(n_2455),
.Y(n_2828)
);

INVx1_ASAP7_75t_L g2829 ( 
.A(n_2473),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2494),
.Y(n_2830)
);

AND2x4_ASAP7_75t_L g2831 ( 
.A(n_2281),
.B(n_1982),
.Y(n_2831)
);

CKINVDCx20_ASAP7_75t_R g2832 ( 
.A(n_2292),
.Y(n_2832)
);

AOI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_2449),
.A2(n_2030),
.B1(n_2080),
.B2(n_2013),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2514),
.Y(n_2834)
);

INVx2_ASAP7_75t_L g2835 ( 
.A(n_2569),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2522),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2357),
.B(n_1741),
.Y(n_2837)
);

INVx1_ASAP7_75t_L g2838 ( 
.A(n_2541),
.Y(n_2838)
);

OA21x2_ASAP7_75t_L g2839 ( 
.A1(n_2588),
.A2(n_1844),
.B(n_1840),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2546),
.Y(n_2840)
);

NOR2xp33_ASAP7_75t_R g2841 ( 
.A(n_2547),
.B(n_1299),
.Y(n_2841)
);

INVxp67_ASAP7_75t_L g2842 ( 
.A(n_2533),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2555),
.Y(n_2843)
);

BUFx6f_ASAP7_75t_L g2844 ( 
.A(n_2457),
.Y(n_2844)
);

INVx1_ASAP7_75t_L g2845 ( 
.A(n_2559),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_2585),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2562),
.Y(n_2847)
);

CKINVDCx5p33_ASAP7_75t_R g2848 ( 
.A(n_2394),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2564),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2442),
.B(n_1837),
.Y(n_2850)
);

BUFx6f_ASAP7_75t_L g2851 ( 
.A(n_2463),
.Y(n_2851)
);

BUFx3_ASAP7_75t_L g2852 ( 
.A(n_2570),
.Y(n_2852)
);

AND2x4_ASAP7_75t_L g2853 ( 
.A(n_2480),
.B(n_1792),
.Y(n_2853)
);

CKINVDCx20_ASAP7_75t_R g2854 ( 
.A(n_2446),
.Y(n_2854)
);

CKINVDCx20_ASAP7_75t_R g2855 ( 
.A(n_2336),
.Y(n_2855)
);

INVx1_ASAP7_75t_L g2856 ( 
.A(n_2572),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2573),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2582),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2407),
.Y(n_2859)
);

INVx3_ASAP7_75t_L g2860 ( 
.A(n_2479),
.Y(n_2860)
);

INVx2_ASAP7_75t_L g2861 ( 
.A(n_2587),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2335),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2490),
.Y(n_2863)
);

INVx2_ASAP7_75t_L g2864 ( 
.A(n_2595),
.Y(n_2864)
);

AND2x2_ASAP7_75t_L g2865 ( 
.A(n_2594),
.B(n_1837),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2411),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2387),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2400),
.Y(n_2868)
);

AND2x4_ASAP7_75t_L g2869 ( 
.A(n_2323),
.B(n_1802),
.Y(n_2869)
);

AND2x4_ASAP7_75t_L g2870 ( 
.A(n_2482),
.B(n_1806),
.Y(n_2870)
);

NOR2xp33_ASAP7_75t_R g2871 ( 
.A(n_2502),
.B(n_2520),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2417),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2418),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2435),
.B(n_2095),
.Y(n_2874)
);

CKINVDCx5p33_ASAP7_75t_R g2875 ( 
.A(n_2454),
.Y(n_2875)
);

BUFx6f_ASAP7_75t_L g2876 ( 
.A(n_2505),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2434),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2523),
.B(n_1642),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2436),
.Y(n_2879)
);

INVx5_ASAP7_75t_L g2880 ( 
.A(n_2506),
.Y(n_2880)
);

INVx2_ASAP7_75t_L g2881 ( 
.A(n_2528),
.Y(n_2881)
);

INVx1_ASAP7_75t_L g2882 ( 
.A(n_2500),
.Y(n_2882)
);

CKINVDCx5p33_ASAP7_75t_R g2883 ( 
.A(n_2278),
.Y(n_2883)
);

CKINVDCx5p33_ASAP7_75t_R g2884 ( 
.A(n_2279),
.Y(n_2884)
);

CKINVDCx20_ASAP7_75t_R g2885 ( 
.A(n_2531),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2512),
.Y(n_2886)
);

BUFx2_ASAP7_75t_L g2887 ( 
.A(n_2469),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2524),
.Y(n_2888)
);

NAND3xp33_ASAP7_75t_L g2889 ( 
.A(n_2560),
.B(n_1356),
.C(n_1353),
.Y(n_2889)
);

INVx1_ASAP7_75t_L g2890 ( 
.A(n_2526),
.Y(n_2890)
);

NAND3xp33_ASAP7_75t_L g2891 ( 
.A(n_2539),
.B(n_1363),
.C(n_1357),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2590),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2529),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2548),
.B(n_1728),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2532),
.Y(n_2895)
);

HB1xp67_ASAP7_75t_L g2896 ( 
.A(n_2521),
.Y(n_2896)
);

NOR2xp33_ASAP7_75t_L g2897 ( 
.A(n_2565),
.B(n_1863),
.Y(n_2897)
);

CKINVDCx16_ASAP7_75t_R g2898 ( 
.A(n_2469),
.Y(n_2898)
);

INVx2_ASAP7_75t_L g2899 ( 
.A(n_2542),
.Y(n_2899)
);

NOR2xp33_ASAP7_75t_L g2900 ( 
.A(n_2290),
.B(n_2551),
.Y(n_2900)
);

CKINVDCx20_ASAP7_75t_R g2901 ( 
.A(n_2412),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2428),
.Y(n_2902)
);

HB1xp67_ASAP7_75t_L g2903 ( 
.A(n_2575),
.Y(n_2903)
);

INVx1_ASAP7_75t_L g2904 ( 
.A(n_2553),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2557),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2332),
.A2(n_1371),
.B1(n_1373),
.B2(n_1368),
.Y(n_2906)
);

CKINVDCx5p33_ASAP7_75t_R g2907 ( 
.A(n_2332),
.Y(n_2907)
);

CKINVDCx5p33_ASAP7_75t_R g2908 ( 
.A(n_2397),
.Y(n_2908)
);

INVx2_ASAP7_75t_SL g2909 ( 
.A(n_2584),
.Y(n_2909)
);

BUFx4f_ASAP7_75t_L g2910 ( 
.A(n_2661),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2796),
.Y(n_2911)
);

INVx2_ASAP7_75t_L g2912 ( 
.A(n_2609),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2612),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2799),
.Y(n_2914)
);

INVx6_ASAP7_75t_L g2915 ( 
.A(n_2702),
.Y(n_2915)
);

NAND3xp33_ASAP7_75t_L g2916 ( 
.A(n_2842),
.B(n_2384),
.C(n_2593),
.Y(n_2916)
);

NAND2xp5_ASAP7_75t_SL g2917 ( 
.A(n_2714),
.B(n_2511),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_L g2918 ( 
.A(n_2790),
.B(n_2477),
.Y(n_2918)
);

AOI22xp33_ASAP7_75t_L g2919 ( 
.A1(n_2710),
.A2(n_2397),
.B1(n_2474),
.B2(n_2395),
.Y(n_2919)
);

AND2x2_ASAP7_75t_L g2920 ( 
.A(n_2603),
.B(n_1911),
.Y(n_2920)
);

INVx1_ASAP7_75t_L g2921 ( 
.A(n_2808),
.Y(n_2921)
);

INVx1_ASAP7_75t_L g2922 ( 
.A(n_2809),
.Y(n_2922)
);

INVx3_ASAP7_75t_L g2923 ( 
.A(n_2658),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2810),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2813),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2638),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2624),
.B(n_1911),
.Y(n_2927)
);

INVx2_ASAP7_75t_SL g2928 ( 
.A(n_2774),
.Y(n_2928)
);

BUFx8_ASAP7_75t_SL g2929 ( 
.A(n_2611),
.Y(n_2929)
);

BUFx3_ASAP7_75t_L g2930 ( 
.A(n_2761),
.Y(n_2930)
);

INVx1_ASAP7_75t_L g2931 ( 
.A(n_2815),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_SL g2932 ( 
.A(n_2717),
.B(n_1374),
.Y(n_2932)
);

INVx3_ASAP7_75t_L g2933 ( 
.A(n_2663),
.Y(n_2933)
);

NAND3xp33_ASAP7_75t_L g2934 ( 
.A(n_2817),
.B(n_1383),
.C(n_1379),
.Y(n_2934)
);

NOR2xp33_ASAP7_75t_L g2935 ( 
.A(n_2883),
.B(n_1386),
.Y(n_2935)
);

INVx3_ASAP7_75t_L g2936 ( 
.A(n_2663),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2803),
.B(n_1387),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2639),
.Y(n_2938)
);

INVx4_ASAP7_75t_L g2939 ( 
.A(n_2718),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_SL g2940 ( 
.A(n_2806),
.B(n_1388),
.Y(n_2940)
);

INVx2_ASAP7_75t_L g2941 ( 
.A(n_2599),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_SL g2942 ( 
.A(n_2871),
.B(n_1389),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2867),
.B(n_1814),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2607),
.Y(n_2944)
);

AND2x2_ASAP7_75t_L g2945 ( 
.A(n_2632),
.B(n_1925),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2820),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2827),
.Y(n_2947)
);

INVx2_ASAP7_75t_L g2948 ( 
.A(n_2617),
.Y(n_2948)
);

NAND2xp5_ASAP7_75t_L g2949 ( 
.A(n_2868),
.B(n_1888),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2829),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2830),
.Y(n_2951)
);

INVx2_ASAP7_75t_L g2952 ( 
.A(n_2620),
.Y(n_2952)
);

INVx4_ASAP7_75t_L g2953 ( 
.A(n_2724),
.Y(n_2953)
);

INVx1_ASAP7_75t_L g2954 ( 
.A(n_2834),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2836),
.Y(n_2955)
);

AOI22xp33_ASAP7_75t_L g2956 ( 
.A1(n_2865),
.A2(n_2766),
.B1(n_2678),
.B2(n_2872),
.Y(n_2956)
);

NAND2xp5_ASAP7_75t_L g2957 ( 
.A(n_2873),
.B(n_1888),
.Y(n_2957)
);

INVx3_ASAP7_75t_L g2958 ( 
.A(n_2693),
.Y(n_2958)
);

AOI21x1_ASAP7_75t_L g2959 ( 
.A1(n_2882),
.A2(n_1873),
.B(n_1871),
.Y(n_2959)
);

INVx2_ASAP7_75t_L g2960 ( 
.A(n_2623),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2838),
.Y(n_2961)
);

AND2x6_ASAP7_75t_L g2962 ( 
.A(n_2877),
.B(n_1912),
.Y(n_2962)
);

INVx3_ASAP7_75t_L g2963 ( 
.A(n_2693),
.Y(n_2963)
);

AOI22xp5_ASAP7_75t_L g2964 ( 
.A1(n_2791),
.A2(n_1885),
.B1(n_1960),
.B2(n_1953),
.Y(n_2964)
);

AND2x2_ASAP7_75t_L g2965 ( 
.A(n_2645),
.B(n_1925),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2840),
.Y(n_2966)
);

AOI22xp5_ASAP7_75t_L g2967 ( 
.A1(n_2897),
.A2(n_1972),
.B1(n_1984),
.B2(n_1963),
.Y(n_2967)
);

BUFx6f_ASAP7_75t_SL g2968 ( 
.A(n_2626),
.Y(n_2968)
);

AOI22xp33_ASAP7_75t_SL g2969 ( 
.A1(n_2701),
.A2(n_2048),
.B1(n_1392),
.B2(n_1394),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_SL g2970 ( 
.A(n_2782),
.B(n_2783),
.Y(n_2970)
);

INVx1_ASAP7_75t_L g2971 ( 
.A(n_2843),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2879),
.B(n_1888),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_SL g2973 ( 
.A(n_2795),
.B(n_1391),
.Y(n_2973)
);

BUFx10_ASAP7_75t_L g2974 ( 
.A(n_2596),
.Y(n_2974)
);

BUFx2_ASAP7_75t_L g2975 ( 
.A(n_2647),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2691),
.B(n_2753),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2721),
.B(n_1891),
.Y(n_2977)
);

INVx2_ASAP7_75t_L g2978 ( 
.A(n_2627),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2727),
.Y(n_2979)
);

BUFx8_ASAP7_75t_SL g2980 ( 
.A(n_2643),
.Y(n_2980)
);

INVx1_ASAP7_75t_L g2981 ( 
.A(n_2845),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_L g2982 ( 
.A(n_2819),
.B(n_1891),
.Y(n_2982)
);

INVx3_ASAP7_75t_L g2983 ( 
.A(n_2727),
.Y(n_2983)
);

BUFx6f_ASAP7_75t_L g2984 ( 
.A(n_2731),
.Y(n_2984)
);

INVxp33_ASAP7_75t_SL g2985 ( 
.A(n_2600),
.Y(n_2985)
);

INVx1_ASAP7_75t_L g2986 ( 
.A(n_2847),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2874),
.B(n_1891),
.Y(n_2987)
);

NOR3xp33_ASAP7_75t_L g2988 ( 
.A(n_2671),
.B(n_1811),
.C(n_1807),
.Y(n_2988)
);

BUFx6f_ASAP7_75t_L g2989 ( 
.A(n_2731),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2849),
.Y(n_2990)
);

INVx4_ASAP7_75t_L g2991 ( 
.A(n_2729),
.Y(n_2991)
);

INVx2_ASAP7_75t_L g2992 ( 
.A(n_2628),
.Y(n_2992)
);

INVx8_ASAP7_75t_L g2993 ( 
.A(n_2670),
.Y(n_2993)
);

NAND2xp33_ASAP7_75t_SL g2994 ( 
.A(n_2604),
.B(n_1395),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2644),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2678),
.B(n_1988),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2856),
.Y(n_2997)
);

INVx5_ASAP7_75t_L g2998 ( 
.A(n_2660),
.Y(n_2998)
);

BUFx2_ASAP7_75t_L g2999 ( 
.A(n_2662),
.Y(n_2999)
);

AND2x6_ASAP7_75t_L g3000 ( 
.A(n_2648),
.B(n_2000),
.Y(n_3000)
);

BUFx6f_ASAP7_75t_L g3001 ( 
.A(n_2733),
.Y(n_3001)
);

INVx1_ASAP7_75t_L g3002 ( 
.A(n_2857),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2649),
.Y(n_3003)
);

BUFx10_ASAP7_75t_L g3004 ( 
.A(n_2608),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_L g3005 ( 
.A(n_2678),
.B(n_1988),
.Y(n_3005)
);

BUFx3_ASAP7_75t_L g3006 ( 
.A(n_2610),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2858),
.Y(n_3007)
);

INVx1_ASAP7_75t_L g3008 ( 
.A(n_2705),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2650),
.Y(n_3009)
);

OR2x6_ASAP7_75t_L g3010 ( 
.A(n_2887),
.B(n_1450),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_L g3011 ( 
.A(n_2766),
.B(n_1988),
.Y(n_3011)
);

NOR2xp33_ASAP7_75t_L g3012 ( 
.A(n_2884),
.B(n_2614),
.Y(n_3012)
);

AND2x2_ASAP7_75t_L g3013 ( 
.A(n_2797),
.B(n_2048),
.Y(n_3013)
);

INVx2_ASAP7_75t_L g3014 ( 
.A(n_2652),
.Y(n_3014)
);

INVx1_ASAP7_75t_L g3015 ( 
.A(n_2706),
.Y(n_3015)
);

INVx3_ASAP7_75t_L g3016 ( 
.A(n_2733),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2708),
.Y(n_3017)
);

BUFx6f_ASAP7_75t_L g3018 ( 
.A(n_2737),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2631),
.B(n_1397),
.Y(n_3019)
);

NAND2xp5_ASAP7_75t_L g3020 ( 
.A(n_2766),
.B(n_2900),
.Y(n_3020)
);

NOR2xp33_ASAP7_75t_L g3021 ( 
.A(n_2734),
.B(n_1400),
.Y(n_3021)
);

NAND2xp33_ASAP7_75t_L g3022 ( 
.A(n_2622),
.B(n_1402),
.Y(n_3022)
);

INVx1_ASAP7_75t_L g3023 ( 
.A(n_2709),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2769),
.B(n_1405),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_SL g3025 ( 
.A(n_2704),
.B(n_1408),
.Y(n_3025)
);

INVx4_ASAP7_75t_L g3026 ( 
.A(n_2736),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2657),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2640),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2725),
.B(n_1410),
.Y(n_3029)
);

INVx2_ASAP7_75t_SL g3030 ( 
.A(n_2689),
.Y(n_3030)
);

NOR2xp33_ASAP7_75t_L g3031 ( 
.A(n_2616),
.B(n_2629),
.Y(n_3031)
);

NAND2xp33_ASAP7_75t_SL g3032 ( 
.A(n_2630),
.B(n_1412),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2601),
.B(n_2020),
.Y(n_3033)
);

BUFx4f_ASAP7_75t_L g3034 ( 
.A(n_2684),
.Y(n_3034)
);

HB1xp67_ASAP7_75t_L g3035 ( 
.A(n_2633),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2641),
.Y(n_3036)
);

INVx1_ASAP7_75t_L g3037 ( 
.A(n_2711),
.Y(n_3037)
);

INVx1_ASAP7_75t_SL g3038 ( 
.A(n_2669),
.Y(n_3038)
);

OR2x6_ASAP7_75t_L g3039 ( 
.A(n_2780),
.B(n_1523),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2716),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2720),
.Y(n_3041)
);

AOI22x1_ASAP7_75t_L g3042 ( 
.A1(n_2723),
.A2(n_1418),
.B1(n_1420),
.B2(n_1414),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2730),
.Y(n_3043)
);

NOR2xp33_ASAP7_75t_L g3044 ( 
.A(n_2646),
.B(n_1424),
.Y(n_3044)
);

AND2x2_ASAP7_75t_L g3045 ( 
.A(n_2749),
.B(n_1816),
.Y(n_3045)
);

INVx3_ASAP7_75t_L g3046 ( 
.A(n_2737),
.Y(n_3046)
);

CKINVDCx5p33_ASAP7_75t_R g3047 ( 
.A(n_2634),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2732),
.Y(n_3048)
);

INVx2_ASAP7_75t_L g3049 ( 
.A(n_2654),
.Y(n_3049)
);

INVx2_ASAP7_75t_SL g3050 ( 
.A(n_2768),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2601),
.B(n_2020),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2601),
.B(n_2020),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2665),
.Y(n_3053)
);

INVx2_ASAP7_75t_SL g3054 ( 
.A(n_2785),
.Y(n_3054)
);

BUFx2_ASAP7_75t_L g3055 ( 
.A(n_2656),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2740),
.Y(n_3056)
);

INVx4_ASAP7_75t_L g3057 ( 
.A(n_2738),
.Y(n_3057)
);

OAI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2741),
.A2(n_1427),
.B1(n_1428),
.B2(n_1426),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2680),
.Y(n_3059)
);

AND2x2_ASAP7_75t_L g3060 ( 
.A(n_2613),
.B(n_1824),
.Y(n_3060)
);

INVx2_ASAP7_75t_L g3061 ( 
.A(n_2690),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2666),
.Y(n_3062)
);

INVx3_ASAP7_75t_L g3063 ( 
.A(n_2752),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2742),
.B(n_2045),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2695),
.Y(n_3065)
);

AND2x4_ASAP7_75t_L g3066 ( 
.A(n_2653),
.B(n_1831),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2746),
.Y(n_3067)
);

OR2x2_ASAP7_75t_L g3068 ( 
.A(n_2681),
.B(n_1832),
.Y(n_3068)
);

INVx6_ASAP7_75t_L g3069 ( 
.A(n_2880),
.Y(n_3069)
);

INVx2_ASAP7_75t_L g3070 ( 
.A(n_2707),
.Y(n_3070)
);

OR2x6_ASAP7_75t_L g3071 ( 
.A(n_2780),
.B(n_1537),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_2712),
.B(n_1838),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2713),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2674),
.B(n_1429),
.Y(n_3074)
);

INVx2_ASAP7_75t_L g3075 ( 
.A(n_2719),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2751),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2722),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2756),
.B(n_2045),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2760),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2764),
.B(n_2045),
.Y(n_3080)
);

BUFx3_ASAP7_75t_L g3081 ( 
.A(n_2739),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2767),
.Y(n_3082)
);

INVx4_ASAP7_75t_L g3083 ( 
.A(n_2755),
.Y(n_3083)
);

AOI22xp5_ASAP7_75t_L g3084 ( 
.A1(n_2788),
.A2(n_2032),
.B1(n_2035),
.B2(n_2002),
.Y(n_3084)
);

INVx2_ASAP7_75t_L g3085 ( 
.A(n_2726),
.Y(n_3085)
);

OAI21xp33_ASAP7_75t_SL g3086 ( 
.A1(n_2775),
.A2(n_1862),
.B(n_1845),
.Y(n_3086)
);

NAND2xp5_ASAP7_75t_L g3087 ( 
.A(n_2779),
.B(n_2098),
.Y(n_3087)
);

INVx2_ASAP7_75t_L g3088 ( 
.A(n_2743),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2781),
.Y(n_3089)
);

NAND2xp5_ASAP7_75t_L g3090 ( 
.A(n_2789),
.B(n_2098),
.Y(n_3090)
);

NOR2xp33_ASAP7_75t_L g3091 ( 
.A(n_2606),
.B(n_1435),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_SL g3092 ( 
.A(n_2728),
.B(n_1436),
.Y(n_3092)
);

BUFx2_ASAP7_75t_L g3093 ( 
.A(n_2688),
.Y(n_3093)
);

AND2x4_ASAP7_75t_L g3094 ( 
.A(n_2699),
.B(n_1866),
.Y(n_3094)
);

HB1xp67_ASAP7_75t_L g3095 ( 
.A(n_2758),
.Y(n_3095)
);

NAND2xp5_ASAP7_75t_L g3096 ( 
.A(n_2794),
.B(n_2098),
.Y(n_3096)
);

AOI22xp5_ASAP7_75t_L g3097 ( 
.A1(n_2812),
.A2(n_2094),
.B1(n_2041),
.B2(n_1301),
.Y(n_3097)
);

INVx2_ASAP7_75t_L g3098 ( 
.A(n_2750),
.Y(n_3098)
);

INVx2_ASAP7_75t_L g3099 ( 
.A(n_2762),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2852),
.Y(n_3100)
);

INVx2_ASAP7_75t_L g3101 ( 
.A(n_2763),
.Y(n_3101)
);

NAND2xp5_ASAP7_75t_L g3102 ( 
.A(n_2878),
.B(n_1438),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2773),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_SL g3104 ( 
.A(n_2745),
.B(n_1443),
.Y(n_3104)
);

INVx1_ASAP7_75t_L g3105 ( 
.A(n_2793),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2805),
.Y(n_3106)
);

NOR3xp33_ASAP7_75t_L g3107 ( 
.A(n_2698),
.B(n_1879),
.C(n_1875),
.Y(n_3107)
);

NOR3xp33_ASAP7_75t_L g3108 ( 
.A(n_2889),
.B(n_1884),
.C(n_1881),
.Y(n_3108)
);

INVxp67_ASAP7_75t_SL g3109 ( 
.A(n_2747),
.Y(n_3109)
);

BUFx6f_ASAP7_75t_L g3110 ( 
.A(n_2752),
.Y(n_3110)
);

AOI22xp33_ASAP7_75t_L g3111 ( 
.A1(n_2862),
.A2(n_1624),
.B1(n_1646),
.B2(n_1586),
.Y(n_3111)
);

INVx4_ASAP7_75t_L g3112 ( 
.A(n_2651),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_SL g3113 ( 
.A(n_2777),
.B(n_1452),
.Y(n_3113)
);

INVx3_ASAP7_75t_L g3114 ( 
.A(n_2754),
.Y(n_3114)
);

BUFx3_ASAP7_75t_L g3115 ( 
.A(n_2605),
.Y(n_3115)
);

INVxp67_ASAP7_75t_L g3116 ( 
.A(n_2625),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2821),
.Y(n_3117)
);

INVx2_ASAP7_75t_SL g3118 ( 
.A(n_2850),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_2703),
.B(n_1453),
.Y(n_3119)
);

INVx3_ASAP7_75t_L g3120 ( 
.A(n_2754),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2835),
.Y(n_3121)
);

INVx1_ASAP7_75t_L g3122 ( 
.A(n_2846),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2861),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2831),
.B(n_1889),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2784),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2864),
.Y(n_3126)
);

INVx3_ASAP7_75t_L g3127 ( 
.A(n_2784),
.Y(n_3127)
);

AOI21x1_ASAP7_75t_L g3128 ( 
.A1(n_2886),
.A2(n_1358),
.B(n_1284),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2776),
.B(n_1455),
.Y(n_3129)
);

NAND2xp5_ASAP7_75t_L g3130 ( 
.A(n_2894),
.B(n_1456),
.Y(n_3130)
);

NAND2xp5_ASAP7_75t_L g3131 ( 
.A(n_2792),
.B(n_1460),
.Y(n_3131)
);

AO22x2_ASAP7_75t_L g3132 ( 
.A1(n_2675),
.A2(n_1895),
.B1(n_1896),
.B2(n_1892),
.Y(n_3132)
);

INVx4_ASAP7_75t_L g3133 ( 
.A(n_2679),
.Y(n_3133)
);

AOI22xp33_ASAP7_75t_L g3134 ( 
.A1(n_2866),
.A2(n_1830),
.B1(n_1898),
.B2(n_1789),
.Y(n_3134)
);

BUFx6f_ASAP7_75t_L g3135 ( 
.A(n_2844),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_SL g3136 ( 
.A(n_2906),
.B(n_2802),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_SL g3137 ( 
.A(n_2833),
.B(n_1464),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2888),
.Y(n_3138)
);

INVx1_ASAP7_75t_L g3139 ( 
.A(n_2890),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2892),
.Y(n_3140)
);

AND2x2_ASAP7_75t_L g3141 ( 
.A(n_2804),
.B(n_1900),
.Y(n_3141)
);

INVx2_ASAP7_75t_L g3142 ( 
.A(n_2786),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_SL g3143 ( 
.A(n_2898),
.B(n_1469),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_SL g3144 ( 
.A(n_2811),
.B(n_1470),
.Y(n_3144)
);

INVx5_ASAP7_75t_L g3145 ( 
.A(n_2818),
.Y(n_3145)
);

INVx3_ASAP7_75t_L g3146 ( 
.A(n_2844),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2909),
.B(n_1474),
.Y(n_3147)
);

NOR2xp33_ASAP7_75t_L g3148 ( 
.A(n_2801),
.B(n_1476),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2822),
.Y(n_3149)
);

NAND2xp5_ASAP7_75t_L g3150 ( 
.A(n_2816),
.B(n_2735),
.Y(n_3150)
);

AND2x6_ASAP7_75t_L g3151 ( 
.A(n_3081),
.B(n_2837),
.Y(n_3151)
);

INVx5_ASAP7_75t_L g3152 ( 
.A(n_2929),
.Y(n_3152)
);

AND2x2_ASAP7_75t_SL g3153 ( 
.A(n_2918),
.B(n_2598),
.Y(n_3153)
);

BUFx3_ASAP7_75t_L g3154 ( 
.A(n_2930),
.Y(n_3154)
);

HB1xp67_ASAP7_75t_L g3155 ( 
.A(n_2975),
.Y(n_3155)
);

OR2x2_ASAP7_75t_SL g3156 ( 
.A(n_3095),
.B(n_2891),
.Y(n_3156)
);

CKINVDCx8_ASAP7_75t_R g3157 ( 
.A(n_3047),
.Y(n_3157)
);

INVx1_ASAP7_75t_L g3158 ( 
.A(n_2911),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_3149),
.B(n_2771),
.Y(n_3159)
);

AO22x2_ASAP7_75t_L g3160 ( 
.A1(n_3030),
.A2(n_2636),
.B1(n_2787),
.B2(n_2832),
.Y(n_3160)
);

CKINVDCx5p33_ASAP7_75t_R g3161 ( 
.A(n_2985),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2914),
.Y(n_3162)
);

NAND3xp33_ASAP7_75t_L g3163 ( 
.A(n_2935),
.B(n_2715),
.C(n_2770),
.Y(n_3163)
);

INVx1_ASAP7_75t_L g3164 ( 
.A(n_2921),
.Y(n_3164)
);

OAI22xp33_ASAP7_75t_L g3165 ( 
.A1(n_3038),
.A2(n_2967),
.B1(n_3093),
.B2(n_3006),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2922),
.Y(n_3166)
);

INVxp67_ASAP7_75t_L g3167 ( 
.A(n_3055),
.Y(n_3167)
);

BUFx2_ASAP7_75t_L g3168 ( 
.A(n_2999),
.Y(n_3168)
);

AND2x4_ASAP7_75t_L g3169 ( 
.A(n_2998),
.B(n_2902),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2924),
.Y(n_3170)
);

NAND3xp33_ASAP7_75t_L g3171 ( 
.A(n_3012),
.B(n_2824),
.C(n_2814),
.Y(n_3171)
);

BUFx3_ASAP7_75t_L g3172 ( 
.A(n_2915),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2925),
.Y(n_3173)
);

BUFx4f_ASAP7_75t_L g3174 ( 
.A(n_2993),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2931),
.Y(n_3175)
);

INVx3_ASAP7_75t_L g3176 ( 
.A(n_2980),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_3150),
.B(n_2907),
.Y(n_3177)
);

BUFx6f_ASAP7_75t_L g3178 ( 
.A(n_2979),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2946),
.Y(n_3179)
);

OR2x6_ASAP7_75t_L g3180 ( 
.A(n_2993),
.B(n_2597),
.Y(n_3180)
);

INVxp67_ASAP7_75t_L g3181 ( 
.A(n_2976),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2947),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_2950),
.Y(n_3183)
);

BUFx6f_ASAP7_75t_L g3184 ( 
.A(n_2979),
.Y(n_3184)
);

HB1xp67_ASAP7_75t_L g3185 ( 
.A(n_3035),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2962),
.B(n_2908),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2962),
.B(n_2841),
.Y(n_3187)
);

INVx2_ASAP7_75t_L g3188 ( 
.A(n_2912),
.Y(n_3188)
);

NAND2xp5_ASAP7_75t_L g3189 ( 
.A(n_2962),
.B(n_2869),
.Y(n_3189)
);

AND2x2_ASAP7_75t_L g3190 ( 
.A(n_3013),
.B(n_2896),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2951),
.Y(n_3191)
);

INVx2_ASAP7_75t_SL g3192 ( 
.A(n_2910),
.Y(n_3192)
);

BUFx6f_ASAP7_75t_L g3193 ( 
.A(n_2984),
.Y(n_3193)
);

INVx4_ASAP7_75t_SL g3194 ( 
.A(n_2968),
.Y(n_3194)
);

INVx2_ASAP7_75t_L g3195 ( 
.A(n_2913),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_3060),
.B(n_2903),
.Y(n_3196)
);

INVx2_ASAP7_75t_L g3197 ( 
.A(n_2926),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_SL g3198 ( 
.A(n_3020),
.B(n_2618),
.Y(n_3198)
);

BUFx6f_ASAP7_75t_L g3199 ( 
.A(n_2984),
.Y(n_3199)
);

INVx1_ASAP7_75t_L g3200 ( 
.A(n_2954),
.Y(n_3200)
);

OR2x2_ASAP7_75t_SL g3201 ( 
.A(n_2916),
.B(n_2885),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2955),
.Y(n_3202)
);

BUFx3_ASAP7_75t_L g3203 ( 
.A(n_3069),
.Y(n_3203)
);

INVx2_ASAP7_75t_L g3204 ( 
.A(n_2938),
.Y(n_3204)
);

BUFx2_ASAP7_75t_L g3205 ( 
.A(n_3062),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2961),
.Y(n_3206)
);

NOR2xp33_ASAP7_75t_L g3207 ( 
.A(n_3116),
.B(n_2759),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_2966),
.Y(n_3208)
);

AO21x2_ASAP7_75t_L g3209 ( 
.A1(n_3128),
.A2(n_2823),
.B(n_2694),
.Y(n_3209)
);

INVxp67_ASAP7_75t_SL g3210 ( 
.A(n_2923),
.Y(n_3210)
);

INVx1_ASAP7_75t_L g3211 ( 
.A(n_2971),
.Y(n_3211)
);

INVx2_ASAP7_75t_L g3212 ( 
.A(n_2941),
.Y(n_3212)
);

BUFx6f_ASAP7_75t_L g3213 ( 
.A(n_2989),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_L g3214 ( 
.A(n_3148),
.B(n_2818),
.Y(n_3214)
);

AND2x2_ASAP7_75t_L g3215 ( 
.A(n_3072),
.B(n_2920),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2974),
.Y(n_3216)
);

BUFx6f_ASAP7_75t_L g3217 ( 
.A(n_2989),
.Y(n_3217)
);

AND2x4_ASAP7_75t_L g3218 ( 
.A(n_2998),
.B(n_2621),
.Y(n_3218)
);

INVx3_ASAP7_75t_L g3219 ( 
.A(n_3004),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2981),
.Y(n_3220)
);

INVx1_ASAP7_75t_L g3221 ( 
.A(n_2986),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_SL g3222 ( 
.A(n_2939),
.B(n_2798),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2990),
.B(n_2818),
.Y(n_3223)
);

AO22x2_ASAP7_75t_L g3224 ( 
.A1(n_3050),
.A2(n_2854),
.B1(n_2778),
.B2(n_2855),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_2997),
.Y(n_3225)
);

INVx2_ASAP7_75t_L g3226 ( 
.A(n_2944),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_3001),
.Y(n_3227)
);

AND2x2_ASAP7_75t_L g3228 ( 
.A(n_2927),
.B(n_2870),
.Y(n_3228)
);

BUFx6f_ASAP7_75t_L g3229 ( 
.A(n_3001),
.Y(n_3229)
);

INVx1_ASAP7_75t_L g3230 ( 
.A(n_3002),
.Y(n_3230)
);

BUFx6f_ASAP7_75t_L g3231 ( 
.A(n_3018),
.Y(n_3231)
);

NOR2xp33_ASAP7_75t_L g3232 ( 
.A(n_2928),
.B(n_3031),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_2948),
.Y(n_3233)
);

INVx3_ASAP7_75t_L g3234 ( 
.A(n_2953),
.Y(n_3234)
);

AND2x2_ASAP7_75t_L g3235 ( 
.A(n_2945),
.B(n_2853),
.Y(n_3235)
);

BUFx2_ASAP7_75t_L g3236 ( 
.A(n_3010),
.Y(n_3236)
);

INVx2_ASAP7_75t_L g3237 ( 
.A(n_2952),
.Y(n_3237)
);

OR2x6_ASAP7_75t_L g3238 ( 
.A(n_2991),
.B(n_2602),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3007),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3008),
.Y(n_3240)
);

INVx2_ASAP7_75t_L g3241 ( 
.A(n_2960),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_3015),
.Y(n_3242)
);

INVxp67_ASAP7_75t_L g3243 ( 
.A(n_3044),
.Y(n_3243)
);

BUFx2_ASAP7_75t_L g3244 ( 
.A(n_3010),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_3026),
.B(n_2655),
.Y(n_3245)
);

NAND2xp5_ASAP7_75t_L g3246 ( 
.A(n_3091),
.B(n_2744),
.Y(n_3246)
);

AND2x4_ASAP7_75t_L g3247 ( 
.A(n_3057),
.B(n_3083),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_3017),
.B(n_2757),
.Y(n_3248)
);

NOR2xp33_ASAP7_75t_SL g3249 ( 
.A(n_3112),
.B(n_2676),
.Y(n_3249)
);

INVx1_ASAP7_75t_L g3250 ( 
.A(n_3023),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_2978),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_3037),
.B(n_2772),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_SL g3253 ( 
.A(n_2956),
.B(n_2619),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_L g3254 ( 
.A(n_3040),
.B(n_2642),
.Y(n_3254)
);

INVx3_ASAP7_75t_L g3255 ( 
.A(n_3018),
.Y(n_3255)
);

AO22x2_ASAP7_75t_L g3256 ( 
.A1(n_3054),
.A2(n_2765),
.B1(n_2901),
.B2(n_2667),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3041),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_3043),
.Y(n_3258)
);

NAND2xp5_ASAP7_75t_L g3259 ( 
.A(n_3048),
.B(n_2664),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_3056),
.Y(n_3260)
);

BUFx3_ASAP7_75t_L g3261 ( 
.A(n_3034),
.Y(n_3261)
);

OR2x2_ASAP7_75t_SL g3262 ( 
.A(n_3068),
.B(n_2848),
.Y(n_3262)
);

INVx2_ASAP7_75t_L g3263 ( 
.A(n_2992),
.Y(n_3263)
);

AOI22xp33_ASAP7_75t_L g3264 ( 
.A1(n_3107),
.A2(n_2668),
.B1(n_2673),
.B2(n_2672),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3067),
.Y(n_3265)
);

INVx1_ASAP7_75t_L g3266 ( 
.A(n_3076),
.Y(n_3266)
);

INVx2_ASAP7_75t_SL g3267 ( 
.A(n_3110),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3079),
.B(n_2677),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3082),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_3089),
.Y(n_3270)
);

AND2x4_ASAP7_75t_L g3271 ( 
.A(n_3118),
.B(n_3115),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2995),
.Y(n_3272)
);

INVx1_ASAP7_75t_L g3273 ( 
.A(n_3003),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3009),
.Y(n_3274)
);

INVx2_ASAP7_75t_L g3275 ( 
.A(n_3014),
.Y(n_3275)
);

INVx2_ASAP7_75t_L g3276 ( 
.A(n_3027),
.Y(n_3276)
);

INVx1_ASAP7_75t_L g3277 ( 
.A(n_3103),
.Y(n_3277)
);

OR2x2_ASAP7_75t_SL g3278 ( 
.A(n_2934),
.B(n_2859),
.Y(n_3278)
);

BUFx3_ASAP7_75t_L g3279 ( 
.A(n_3110),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_SL g3280 ( 
.A(n_3145),
.B(n_2659),
.Y(n_3280)
);

BUFx6f_ASAP7_75t_L g3281 ( 
.A(n_3125),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3105),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_3109),
.B(n_2682),
.Y(n_3283)
);

INVxp67_ASAP7_75t_L g3284 ( 
.A(n_3074),
.Y(n_3284)
);

OR2x2_ASAP7_75t_L g3285 ( 
.A(n_2965),
.B(n_2683),
.Y(n_3285)
);

NOR2xp33_ASAP7_75t_L g3286 ( 
.A(n_3129),
.B(n_2807),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_3000),
.B(n_2685),
.Y(n_3287)
);

NAND2xp5_ASAP7_75t_L g3288 ( 
.A(n_3000),
.B(n_2686),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3106),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3028),
.Y(n_3290)
);

AO22x2_ASAP7_75t_L g3291 ( 
.A1(n_2988),
.A2(n_2692),
.B1(n_2696),
.B2(n_2687),
.Y(n_3291)
);

INVx3_ASAP7_75t_L g3292 ( 
.A(n_3125),
.Y(n_3292)
);

INVx2_ASAP7_75t_L g3293 ( 
.A(n_3036),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3117),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3121),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3122),
.Y(n_3296)
);

AND2x4_ASAP7_75t_L g3297 ( 
.A(n_3133),
.B(n_2697),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3126),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3049),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3138),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3139),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_3000),
.B(n_2700),
.Y(n_3302)
);

CKINVDCx20_ASAP7_75t_R g3303 ( 
.A(n_2994),
.Y(n_3303)
);

INVx2_ASAP7_75t_L g3304 ( 
.A(n_3053),
.Y(n_3304)
);

AND2x6_ASAP7_75t_L g3305 ( 
.A(n_3141),
.B(n_2615),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_3059),
.Y(n_3306)
);

AND2x4_ASAP7_75t_L g3307 ( 
.A(n_3039),
.B(n_2635),
.Y(n_3307)
);

NAND2x1p5_ASAP7_75t_L g3308 ( 
.A(n_3135),
.B(n_2880),
.Y(n_3308)
);

AND2x2_ASAP7_75t_SL g3309 ( 
.A(n_2919),
.B(n_2851),
.Y(n_3309)
);

AND2x2_ASAP7_75t_L g3310 ( 
.A(n_3045),
.B(n_2826),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_SL g3311 ( 
.A(n_3165),
.B(n_2969),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_3212),
.Y(n_3312)
);

AOI22xp33_ASAP7_75t_L g3313 ( 
.A1(n_3309),
.A2(n_3132),
.B1(n_3071),
.B2(n_3039),
.Y(n_3313)
);

INVx2_ASAP7_75t_L g3314 ( 
.A(n_3226),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_SL g3315 ( 
.A1(n_3153),
.A2(n_3094),
.B1(n_3071),
.B2(n_3066),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_3243),
.B(n_3100),
.Y(n_3316)
);

INVx1_ASAP7_75t_L g3317 ( 
.A(n_3158),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3284),
.B(n_3021),
.Y(n_3318)
);

AND2x6_ASAP7_75t_SL g3319 ( 
.A(n_3180),
.B(n_3024),
.Y(n_3319)
);

OR2x6_ASAP7_75t_L g3320 ( 
.A(n_3172),
.B(n_3135),
.Y(n_3320)
);

AOI22xp33_ASAP7_75t_L g3321 ( 
.A1(n_3196),
.A2(n_3124),
.B1(n_3137),
.B2(n_3147),
.Y(n_3321)
);

AND2x4_ASAP7_75t_L g3322 ( 
.A(n_3261),
.B(n_2933),
.Y(n_3322)
);

NAND2xp5_ASAP7_75t_L g3323 ( 
.A(n_3232),
.B(n_3131),
.Y(n_3323)
);

BUFx12f_ASAP7_75t_L g3324 ( 
.A(n_3152),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_3162),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3164),
.Y(n_3326)
);

NOR2xp33_ASAP7_75t_L g3327 ( 
.A(n_3177),
.B(n_2970),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_3215),
.B(n_3136),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_3159),
.B(n_3102),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_L g3330 ( 
.A1(n_3207),
.A2(n_2964),
.B1(n_3108),
.B2(n_3065),
.Y(n_3330)
);

AOI22xp5_ASAP7_75t_L g3331 ( 
.A1(n_3286),
.A2(n_3022),
.B1(n_3032),
.B2(n_2942),
.Y(n_3331)
);

NOR2xp33_ASAP7_75t_L g3332 ( 
.A(n_3167),
.B(n_3130),
.Y(n_3332)
);

INVxp33_ASAP7_75t_L g3333 ( 
.A(n_3155),
.Y(n_3333)
);

INVx1_ASAP7_75t_L g3334 ( 
.A(n_3166),
.Y(n_3334)
);

OR2x6_ASAP7_75t_L g3335 ( 
.A(n_3192),
.B(n_3143),
.Y(n_3335)
);

INVx1_ASAP7_75t_SL g3336 ( 
.A(n_3205),
.Y(n_3336)
);

NAND2xp33_ASAP7_75t_SL g3337 ( 
.A(n_3161),
.B(n_2932),
.Y(n_3337)
);

NAND2xp5_ASAP7_75t_L g3338 ( 
.A(n_3181),
.B(n_3145),
.Y(n_3338)
);

NAND2xp5_ASAP7_75t_L g3339 ( 
.A(n_3246),
.B(n_3097),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3170),
.B(n_3173),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_3175),
.B(n_3111),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_3179),
.B(n_3134),
.Y(n_3342)
);

NAND3xp33_ASAP7_75t_L g3343 ( 
.A(n_3163),
.B(n_3042),
.C(n_3119),
.Y(n_3343)
);

INVx3_ASAP7_75t_L g3344 ( 
.A(n_3157),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_3233),
.Y(n_3345)
);

AOI21xp5_ASAP7_75t_L g3346 ( 
.A1(n_3214),
.A2(n_2949),
.B(n_2943),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_3182),
.B(n_3144),
.Y(n_3347)
);

INVx2_ASAP7_75t_SL g3348 ( 
.A(n_3174),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3183),
.B(n_2957),
.Y(n_3349)
);

INVx2_ASAP7_75t_SL g3350 ( 
.A(n_3203),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3191),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3200),
.Y(n_3352)
);

HB1xp67_ASAP7_75t_L g3353 ( 
.A(n_3185),
.Y(n_3353)
);

AND2x2_ASAP7_75t_L g3354 ( 
.A(n_3190),
.B(n_3058),
.Y(n_3354)
);

NAND2xp5_ASAP7_75t_L g3355 ( 
.A(n_3202),
.B(n_2972),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3206),
.B(n_2973),
.Y(n_3356)
);

CKINVDCx5p33_ASAP7_75t_R g3357 ( 
.A(n_3152),
.Y(n_3357)
);

NOR2x2_ASAP7_75t_L g3358 ( 
.A(n_3238),
.B(n_1917),
.Y(n_3358)
);

AND2x6_ASAP7_75t_SL g3359 ( 
.A(n_3218),
.B(n_2800),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_SL g3360 ( 
.A(n_3171),
.B(n_2937),
.Y(n_3360)
);

INVx2_ASAP7_75t_L g3361 ( 
.A(n_3237),
.Y(n_3361)
);

BUFx3_ASAP7_75t_L g3362 ( 
.A(n_3154),
.Y(n_3362)
);

AOI22xp33_ASAP7_75t_L g3363 ( 
.A1(n_3305),
.A2(n_3228),
.B1(n_3253),
.B2(n_3235),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3208),
.Y(n_3364)
);

INVx3_ASAP7_75t_L g3365 ( 
.A(n_3178),
.Y(n_3365)
);

OR2x2_ASAP7_75t_SL g3366 ( 
.A(n_3285),
.B(n_2851),
.Y(n_3366)
);

NAND2xp5_ASAP7_75t_L g3367 ( 
.A(n_3211),
.B(n_2940),
.Y(n_3367)
);

BUFx6f_ASAP7_75t_L g3368 ( 
.A(n_3178),
.Y(n_3368)
);

OR2x6_ASAP7_75t_L g3369 ( 
.A(n_3236),
.B(n_2936),
.Y(n_3369)
);

OAI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_3249),
.A2(n_3084),
.B1(n_2958),
.B2(n_2983),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_3220),
.B(n_3019),
.Y(n_3371)
);

NOR2xp33_ASAP7_75t_L g3372 ( 
.A(n_3168),
.B(n_2917),
.Y(n_3372)
);

NAND2xp5_ASAP7_75t_L g3373 ( 
.A(n_3221),
.B(n_2977),
.Y(n_3373)
);

INVx4_ASAP7_75t_L g3374 ( 
.A(n_3194),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_3305),
.A2(n_3070),
.B1(n_3073),
.B2(n_3061),
.Y(n_3375)
);

BUFx2_ASAP7_75t_L g3376 ( 
.A(n_3244),
.Y(n_3376)
);

AND2x4_ASAP7_75t_L g3377 ( 
.A(n_3279),
.B(n_2963),
.Y(n_3377)
);

CKINVDCx5p33_ASAP7_75t_R g3378 ( 
.A(n_3176),
.Y(n_3378)
);

NAND2xp5_ASAP7_75t_L g3379 ( 
.A(n_3225),
.B(n_3086),
.Y(n_3379)
);

INVx1_ASAP7_75t_L g3380 ( 
.A(n_3230),
.Y(n_3380)
);

NAND2xp5_ASAP7_75t_L g3381 ( 
.A(n_3239),
.B(n_3140),
.Y(n_3381)
);

BUFx3_ASAP7_75t_L g3382 ( 
.A(n_3184),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_3240),
.B(n_2982),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_3242),
.B(n_3250),
.Y(n_3384)
);

NAND2xp5_ASAP7_75t_L g3385 ( 
.A(n_3257),
.B(n_2996),
.Y(n_3385)
);

NAND2xp5_ASAP7_75t_L g3386 ( 
.A(n_3258),
.B(n_3005),
.Y(n_3386)
);

NAND2xp5_ASAP7_75t_L g3387 ( 
.A(n_3260),
.B(n_3011),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3265),
.Y(n_3388)
);

AND2x2_ASAP7_75t_L g3389 ( 
.A(n_3310),
.B(n_3016),
.Y(n_3389)
);

INVx5_ASAP7_75t_L g3390 ( 
.A(n_3151),
.Y(n_3390)
);

OR2x6_ASAP7_75t_L g3391 ( 
.A(n_3169),
.B(n_3046),
.Y(n_3391)
);

NAND3xp33_ASAP7_75t_L g3392 ( 
.A(n_3187),
.B(n_2987),
.C(n_3033),
.Y(n_3392)
);

NOR2xp33_ASAP7_75t_L g3393 ( 
.A(n_3189),
.B(n_3025),
.Y(n_3393)
);

AOI22xp33_ASAP7_75t_L g3394 ( 
.A1(n_3241),
.A2(n_3077),
.B1(n_3085),
.B2(n_3075),
.Y(n_3394)
);

NOR2xp33_ASAP7_75t_L g3395 ( 
.A(n_3186),
.B(n_3029),
.Y(n_3395)
);

BUFx3_ASAP7_75t_L g3396 ( 
.A(n_3184),
.Y(n_3396)
);

NOR2xp33_ASAP7_75t_L g3397 ( 
.A(n_3156),
.B(n_3092),
.Y(n_3397)
);

AOI22xp5_ASAP7_75t_L g3398 ( 
.A1(n_3303),
.A2(n_3151),
.B1(n_3271),
.B2(n_3210),
.Y(n_3398)
);

AOI22xp33_ASAP7_75t_L g3399 ( 
.A1(n_3251),
.A2(n_3098),
.B1(n_3099),
.B2(n_3088),
.Y(n_3399)
);

INVx2_ASAP7_75t_L g3400 ( 
.A(n_3263),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_L g3401 ( 
.A(n_3266),
.B(n_3051),
.Y(n_3401)
);

AOI22xp5_ASAP7_75t_L g3402 ( 
.A1(n_3267),
.A2(n_2748),
.B1(n_3052),
.B2(n_3104),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_SL g3403 ( 
.A(n_3193),
.B(n_3063),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3269),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3270),
.B(n_3101),
.Y(n_3405)
);

NAND2xp33_ASAP7_75t_L g3406 ( 
.A(n_3234),
.B(n_3113),
.Y(n_3406)
);

OAI22xp5_ASAP7_75t_SL g3407 ( 
.A1(n_3262),
.A2(n_3201),
.B1(n_3278),
.B2(n_2875),
.Y(n_3407)
);

NOR2xp33_ASAP7_75t_L g3408 ( 
.A(n_3248),
.B(n_3114),
.Y(n_3408)
);

INVxp67_ASAP7_75t_L g3409 ( 
.A(n_3193),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3300),
.B(n_3123),
.Y(n_3410)
);

NOR2xp33_ASAP7_75t_L g3411 ( 
.A(n_3252),
.B(n_3283),
.Y(n_3411)
);

INVx2_ASAP7_75t_L g3412 ( 
.A(n_3275),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_SL g3413 ( 
.A(n_3199),
.B(n_3120),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_3301),
.B(n_3127),
.Y(n_3414)
);

INVx2_ASAP7_75t_L g3415 ( 
.A(n_3276),
.Y(n_3415)
);

AOI22xp5_ASAP7_75t_L g3416 ( 
.A1(n_3247),
.A2(n_3146),
.B1(n_3078),
.B2(n_3080),
.Y(n_3416)
);

INVx3_ASAP7_75t_L g3417 ( 
.A(n_3199),
.Y(n_3417)
);

AND2x2_ASAP7_75t_L g3418 ( 
.A(n_3307),
.B(n_2876),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_L g3419 ( 
.A(n_3272),
.B(n_3064),
.Y(n_3419)
);

BUFx3_ASAP7_75t_L g3420 ( 
.A(n_3213),
.Y(n_3420)
);

INVx2_ASAP7_75t_L g3421 ( 
.A(n_3273),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_L g3422 ( 
.A(n_3274),
.B(n_3087),
.Y(n_3422)
);

INVx2_ASAP7_75t_L g3423 ( 
.A(n_3277),
.Y(n_3423)
);

NAND2x1_ASAP7_75t_L g3424 ( 
.A(n_3213),
.B(n_2825),
.Y(n_3424)
);

INVx1_ASAP7_75t_SL g3425 ( 
.A(n_3217),
.Y(n_3425)
);

INVx2_ASAP7_75t_SL g3426 ( 
.A(n_3217),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_SL g3427 ( 
.A(n_3227),
.B(n_3229),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3282),
.B(n_3090),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_3289),
.Y(n_3429)
);

AND2x2_ASAP7_75t_L g3430 ( 
.A(n_3224),
.B(n_2876),
.Y(n_3430)
);

CKINVDCx5p33_ASAP7_75t_R g3431 ( 
.A(n_3216),
.Y(n_3431)
);

NOR3xp33_ASAP7_75t_L g3432 ( 
.A(n_3222),
.B(n_3219),
.C(n_3254),
.Y(n_3432)
);

INVxp67_ASAP7_75t_SL g3433 ( 
.A(n_3227),
.Y(n_3433)
);

NOR2xp33_ASAP7_75t_L g3434 ( 
.A(n_3223),
.B(n_3096),
.Y(n_3434)
);

NOR2xp33_ASAP7_75t_L g3435 ( 
.A(n_3229),
.B(n_2637),
.Y(n_3435)
);

AND2x2_ASAP7_75t_L g3436 ( 
.A(n_3231),
.B(n_2828),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3294),
.B(n_1477),
.Y(n_3437)
);

BUFx2_ASAP7_75t_L g3438 ( 
.A(n_3231),
.Y(n_3438)
);

OR2x6_ASAP7_75t_L g3439 ( 
.A(n_3308),
.B(n_3281),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3295),
.B(n_1478),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_3296),
.Y(n_3441)
);

INVx5_ASAP7_75t_L g3442 ( 
.A(n_3281),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3298),
.B(n_1479),
.Y(n_3443)
);

INVx3_ASAP7_75t_L g3444 ( 
.A(n_3245),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_3290),
.B(n_1482),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3188),
.Y(n_3446)
);

NAND2xp33_ASAP7_75t_SL g3447 ( 
.A(n_3318),
.B(n_3280),
.Y(n_3447)
);

BUFx6f_ASAP7_75t_L g3448 ( 
.A(n_3362),
.Y(n_3448)
);

CKINVDCx16_ASAP7_75t_R g3449 ( 
.A(n_3324),
.Y(n_3449)
);

AND2x4_ASAP7_75t_L g3450 ( 
.A(n_3390),
.B(n_3255),
.Y(n_3450)
);

CKINVDCx5p33_ASAP7_75t_R g3451 ( 
.A(n_3357),
.Y(n_3451)
);

INVx5_ASAP7_75t_L g3452 ( 
.A(n_3320),
.Y(n_3452)
);

INVx1_ASAP7_75t_SL g3453 ( 
.A(n_3336),
.Y(n_3453)
);

INVx1_ASAP7_75t_L g3454 ( 
.A(n_3423),
.Y(n_3454)
);

AND2x6_ASAP7_75t_L g3455 ( 
.A(n_3398),
.B(n_3287),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3441),
.Y(n_3456)
);

INVx1_ASAP7_75t_L g3457 ( 
.A(n_3317),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3325),
.Y(n_3458)
);

BUFx6f_ASAP7_75t_L g3459 ( 
.A(n_3320),
.Y(n_3459)
);

NAND2x1p5_ASAP7_75t_L g3460 ( 
.A(n_3442),
.B(n_3292),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3326),
.Y(n_3461)
);

NOR2xp33_ASAP7_75t_L g3462 ( 
.A(n_3323),
.B(n_3288),
.Y(n_3462)
);

BUFx6f_ASAP7_75t_L g3463 ( 
.A(n_3442),
.Y(n_3463)
);

BUFx6f_ASAP7_75t_L g3464 ( 
.A(n_3368),
.Y(n_3464)
);

INVx2_ASAP7_75t_L g3465 ( 
.A(n_3421),
.Y(n_3465)
);

AOI22xp33_ASAP7_75t_L g3466 ( 
.A1(n_3311),
.A2(n_3160),
.B1(n_3256),
.B2(n_3197),
.Y(n_3466)
);

BUFx6f_ASAP7_75t_L g3467 ( 
.A(n_3368),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3334),
.Y(n_3468)
);

OR2x2_ASAP7_75t_SL g3469 ( 
.A(n_3339),
.B(n_3302),
.Y(n_3469)
);

INVx5_ASAP7_75t_L g3470 ( 
.A(n_3374),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3351),
.Y(n_3471)
);

AND2x2_ASAP7_75t_L g3472 ( 
.A(n_3354),
.B(n_3291),
.Y(n_3472)
);

CKINVDCx5p33_ASAP7_75t_R g3473 ( 
.A(n_3378),
.Y(n_3473)
);

BUFx3_ASAP7_75t_L g3474 ( 
.A(n_3382),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3352),
.Y(n_3475)
);

INVxp67_ASAP7_75t_L g3476 ( 
.A(n_3353),
.Y(n_3476)
);

AND2x4_ASAP7_75t_L g3477 ( 
.A(n_3390),
.B(n_3297),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_R g3478 ( 
.A(n_3344),
.B(n_2860),
.Y(n_3478)
);

INVx2_ASAP7_75t_L g3479 ( 
.A(n_3312),
.Y(n_3479)
);

INVx6_ASAP7_75t_L g3480 ( 
.A(n_3322),
.Y(n_3480)
);

BUFx2_ASAP7_75t_L g3481 ( 
.A(n_3391),
.Y(n_3481)
);

OR2x6_ASAP7_75t_L g3482 ( 
.A(n_3350),
.B(n_3259),
.Y(n_3482)
);

BUFx2_ASAP7_75t_L g3483 ( 
.A(n_3391),
.Y(n_3483)
);

INVxp67_ASAP7_75t_L g3484 ( 
.A(n_3389),
.Y(n_3484)
);

AND2x2_ASAP7_75t_L g3485 ( 
.A(n_3315),
.B(n_3299),
.Y(n_3485)
);

BUFx2_ASAP7_75t_L g3486 ( 
.A(n_3369),
.Y(n_3486)
);

INVx3_ASAP7_75t_L g3487 ( 
.A(n_3396),
.Y(n_3487)
);

INVx2_ASAP7_75t_SL g3488 ( 
.A(n_3439),
.Y(n_3488)
);

AOI22xp5_ASAP7_75t_L g3489 ( 
.A1(n_3332),
.A2(n_3264),
.B1(n_3268),
.B2(n_3198),
.Y(n_3489)
);

AND2x2_ASAP7_75t_L g3490 ( 
.A(n_3313),
.B(n_3293),
.Y(n_3490)
);

INVx2_ASAP7_75t_SL g3491 ( 
.A(n_3439),
.Y(n_3491)
);

AOI21xp33_ASAP7_75t_L g3492 ( 
.A1(n_3411),
.A2(n_3204),
.B(n_3195),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3329),
.B(n_3304),
.Y(n_3493)
);

AOI22xp5_ASAP7_75t_L g3494 ( 
.A1(n_3397),
.A2(n_1484),
.B1(n_1490),
.B2(n_1483),
.Y(n_3494)
);

NAND2x1p5_ASAP7_75t_L g3495 ( 
.A(n_3420),
.B(n_2863),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_L g3496 ( 
.A(n_3327),
.B(n_3306),
.Y(n_3496)
);

INVx2_ASAP7_75t_L g3497 ( 
.A(n_3314),
.Y(n_3497)
);

BUFx6f_ASAP7_75t_L g3498 ( 
.A(n_3377),
.Y(n_3498)
);

INVx1_ASAP7_75t_L g3499 ( 
.A(n_3364),
.Y(n_3499)
);

BUFx3_ASAP7_75t_L g3500 ( 
.A(n_3438),
.Y(n_3500)
);

HB1xp67_ASAP7_75t_L g3501 ( 
.A(n_3376),
.Y(n_3501)
);

AND2x4_ASAP7_75t_L g3502 ( 
.A(n_3348),
.B(n_2881),
.Y(n_3502)
);

OR2x6_ASAP7_75t_L g3503 ( 
.A(n_3369),
.B(n_2893),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3380),
.Y(n_3504)
);

NAND2xp33_ASAP7_75t_L g3505 ( 
.A(n_3331),
.B(n_1494),
.Y(n_3505)
);

NAND2x1p5_ASAP7_75t_L g3506 ( 
.A(n_3444),
.B(n_2904),
.Y(n_3506)
);

NOR3xp33_ASAP7_75t_SL g3507 ( 
.A(n_3431),
.B(n_1501),
.C(n_1498),
.Y(n_3507)
);

AOI22xp33_ASAP7_75t_L g3508 ( 
.A1(n_3430),
.A2(n_2905),
.B1(n_2899),
.B2(n_2895),
.Y(n_3508)
);

NAND2xp33_ASAP7_75t_SL g3509 ( 
.A(n_3360),
.B(n_1502),
.Y(n_3509)
);

NOR3xp33_ASAP7_75t_SL g3510 ( 
.A(n_3337),
.B(n_1517),
.C(n_1505),
.Y(n_3510)
);

INVxp67_ASAP7_75t_L g3511 ( 
.A(n_3418),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3388),
.Y(n_3512)
);

INVx3_ASAP7_75t_L g3513 ( 
.A(n_3365),
.Y(n_3513)
);

BUFx12f_ASAP7_75t_L g3514 ( 
.A(n_3359),
.Y(n_3514)
);

BUFx6f_ASAP7_75t_L g3515 ( 
.A(n_3426),
.Y(n_3515)
);

NAND2xp5_ASAP7_75t_SL g3516 ( 
.A(n_3328),
.B(n_3142),
.Y(n_3516)
);

NOR3xp33_ASAP7_75t_SL g3517 ( 
.A(n_3343),
.B(n_1525),
.C(n_1522),
.Y(n_3517)
);

INVx2_ASAP7_75t_L g3518 ( 
.A(n_3345),
.Y(n_3518)
);

INVx2_ASAP7_75t_L g3519 ( 
.A(n_3361),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3404),
.Y(n_3520)
);

INVx2_ASAP7_75t_L g3521 ( 
.A(n_3400),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_3408),
.B(n_1526),
.Y(n_3522)
);

NOR2x1_ASAP7_75t_L g3523 ( 
.A(n_3316),
.B(n_3417),
.Y(n_3523)
);

AOI22xp5_ASAP7_75t_L g3524 ( 
.A1(n_3363),
.A2(n_3321),
.B1(n_3372),
.B2(n_3393),
.Y(n_3524)
);

OAI221xp5_ASAP7_75t_L g3525 ( 
.A1(n_3330),
.A2(n_3367),
.B1(n_3356),
.B2(n_3347),
.C(n_3371),
.Y(n_3525)
);

AOI22xp5_ASAP7_75t_L g3526 ( 
.A1(n_3370),
.A2(n_1529),
.B1(n_1532),
.B2(n_1527),
.Y(n_3526)
);

HB1xp67_ASAP7_75t_L g3527 ( 
.A(n_3333),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_SL g3528 ( 
.A(n_3416),
.B(n_2959),
.Y(n_3528)
);

BUFx3_ASAP7_75t_L g3529 ( 
.A(n_3436),
.Y(n_3529)
);

CKINVDCx5p33_ASAP7_75t_R g3530 ( 
.A(n_3319),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3340),
.Y(n_3531)
);

AOI22xp5_ASAP7_75t_L g3532 ( 
.A1(n_3407),
.A2(n_1539),
.B1(n_1547),
.B2(n_1538),
.Y(n_3532)
);

NAND2xp5_ASAP7_75t_L g3533 ( 
.A(n_3384),
.B(n_1549),
.Y(n_3533)
);

NAND2xp5_ASAP7_75t_L g3534 ( 
.A(n_3381),
.B(n_1550),
.Y(n_3534)
);

NOR3xp33_ASAP7_75t_SL g3535 ( 
.A(n_3395),
.B(n_1553),
.C(n_1551),
.Y(n_3535)
);

AND2x4_ASAP7_75t_L g3536 ( 
.A(n_3433),
.B(n_2571),
.Y(n_3536)
);

NOR2xp33_ASAP7_75t_L g3537 ( 
.A(n_3425),
.B(n_1555),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_3335),
.A2(n_1557),
.B1(n_1559),
.B2(n_1556),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3429),
.Y(n_3539)
);

INVx1_ASAP7_75t_L g3540 ( 
.A(n_3405),
.Y(n_3540)
);

NAND2xp5_ASAP7_75t_L g3541 ( 
.A(n_3379),
.B(n_1564),
.Y(n_3541)
);

HB1xp67_ASAP7_75t_L g3542 ( 
.A(n_3409),
.Y(n_3542)
);

BUFx10_ASAP7_75t_L g3543 ( 
.A(n_3435),
.Y(n_3543)
);

AOI21xp5_ASAP7_75t_L g3544 ( 
.A1(n_3346),
.A2(n_3209),
.B(n_2839),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_3338),
.B(n_1565),
.Y(n_3545)
);

INVx2_ASAP7_75t_L g3546 ( 
.A(n_3412),
.Y(n_3546)
);

HB1xp67_ASAP7_75t_L g3547 ( 
.A(n_3414),
.Y(n_3547)
);

NAND2xp5_ASAP7_75t_L g3548 ( 
.A(n_3415),
.B(n_1567),
.Y(n_3548)
);

AOI22xp5_ASAP7_75t_L g3549 ( 
.A1(n_3335),
.A2(n_1574),
.B1(n_1579),
.B2(n_1573),
.Y(n_3549)
);

NAND2x1p5_ASAP7_75t_L g3550 ( 
.A(n_3427),
.B(n_2576),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3410),
.B(n_1585),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3446),
.Y(n_3552)
);

AO22x1_ASAP7_75t_L g3553 ( 
.A1(n_3432),
.A2(n_1588),
.B1(n_1589),
.B2(n_1587),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3341),
.Y(n_3554)
);

AOI22xp5_ASAP7_75t_L g3555 ( 
.A1(n_3406),
.A2(n_1593),
.B1(n_1594),
.B2(n_1591),
.Y(n_3555)
);

BUFx6f_ASAP7_75t_L g3556 ( 
.A(n_3403),
.Y(n_3556)
);

CKINVDCx16_ASAP7_75t_R g3557 ( 
.A(n_3366),
.Y(n_3557)
);

NAND2x1p5_ASAP7_75t_L g3558 ( 
.A(n_3452),
.B(n_3413),
.Y(n_3558)
);

BUFx6f_ASAP7_75t_L g3559 ( 
.A(n_3463),
.Y(n_3559)
);

BUFx2_ASAP7_75t_L g3560 ( 
.A(n_3501),
.Y(n_3560)
);

AOI21xp5_ASAP7_75t_L g3561 ( 
.A1(n_3505),
.A2(n_3434),
.B(n_3424),
.Y(n_3561)
);

A2O1A1Ixp33_ASAP7_75t_L g3562 ( 
.A1(n_3462),
.A2(n_3402),
.B(n_3349),
.C(n_3355),
.Y(n_3562)
);

INVx1_ASAP7_75t_L g3563 ( 
.A(n_3454),
.Y(n_3563)
);

OAI22xp33_ASAP7_75t_L g3564 ( 
.A1(n_3526),
.A2(n_3342),
.B1(n_3386),
.B2(n_3385),
.Y(n_3564)
);

BUFx3_ASAP7_75t_L g3565 ( 
.A(n_3448),
.Y(n_3565)
);

NAND2xp5_ASAP7_75t_SL g3566 ( 
.A(n_3524),
.B(n_3392),
.Y(n_3566)
);

AOI21xp5_ASAP7_75t_L g3567 ( 
.A1(n_3544),
.A2(n_3401),
.B(n_3387),
.Y(n_3567)
);

NOR2xp67_ASAP7_75t_SL g3568 ( 
.A(n_3470),
.B(n_3373),
.Y(n_3568)
);

INVxp67_ASAP7_75t_SL g3569 ( 
.A(n_3476),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3456),
.Y(n_3570)
);

OAI21xp5_ASAP7_75t_L g3571 ( 
.A1(n_3522),
.A2(n_3440),
.B(n_3437),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3457),
.Y(n_3572)
);

OR2x2_ASAP7_75t_L g3573 ( 
.A(n_3472),
.B(n_3443),
.Y(n_3573)
);

BUFx6f_ASAP7_75t_L g3574 ( 
.A(n_3463),
.Y(n_3574)
);

AOI22xp5_ASAP7_75t_L g3575 ( 
.A1(n_3509),
.A2(n_3375),
.B1(n_3383),
.B2(n_3445),
.Y(n_3575)
);

AOI22xp33_ASAP7_75t_L g3576 ( 
.A1(n_3490),
.A2(n_3466),
.B1(n_3485),
.B2(n_3455),
.Y(n_3576)
);

AOI21x1_ASAP7_75t_L g3577 ( 
.A1(n_3528),
.A2(n_3422),
.B(n_3419),
.Y(n_3577)
);

OAI222xp33_ASAP7_75t_L g3578 ( 
.A1(n_3557),
.A2(n_3428),
.B1(n_3399),
.B2(n_3394),
.C1(n_1928),
.C2(n_1923),
.Y(n_3578)
);

OAI21x1_ASAP7_75t_L g3579 ( 
.A1(n_3516),
.A2(n_1515),
.B(n_1507),
.Y(n_3579)
);

NOR2xp33_ASAP7_75t_L g3580 ( 
.A(n_3473),
.B(n_1595),
.Y(n_3580)
);

OAI21xp5_ASAP7_75t_L g3581 ( 
.A1(n_3494),
.A2(n_1927),
.B(n_1906),
.Y(n_3581)
);

OAI21x1_ASAP7_75t_L g3582 ( 
.A1(n_3458),
.A2(n_1709),
.B(n_1660),
.Y(n_3582)
);

NAND2xp5_ASAP7_75t_L g3583 ( 
.A(n_3531),
.B(n_1929),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3493),
.B(n_1936),
.Y(n_3584)
);

INVx1_ASAP7_75t_SL g3585 ( 
.A(n_3453),
.Y(n_3585)
);

OAI21x1_ASAP7_75t_L g3586 ( 
.A1(n_3461),
.A2(n_1797),
.B(n_1723),
.Y(n_3586)
);

OAI21xp5_ASAP7_75t_L g3587 ( 
.A1(n_3541),
.A2(n_1967),
.B(n_1964),
.Y(n_3587)
);

INVx2_ASAP7_75t_SL g3588 ( 
.A(n_3480),
.Y(n_3588)
);

AOI21xp5_ASAP7_75t_L g3589 ( 
.A1(n_3447),
.A2(n_1861),
.B(n_1813),
.Y(n_3589)
);

OAI21x1_ASAP7_75t_L g3590 ( 
.A1(n_3468),
.A2(n_1961),
.B(n_1870),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3465),
.Y(n_3591)
);

OAI21x1_ASAP7_75t_L g3592 ( 
.A1(n_3471),
.A2(n_2038),
.B(n_1977),
.Y(n_3592)
);

AND2x2_ASAP7_75t_L g3593 ( 
.A(n_3484),
.B(n_1971),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_3540),
.B(n_1973),
.Y(n_3594)
);

BUFx12f_ASAP7_75t_L g3595 ( 
.A(n_3451),
.Y(n_3595)
);

AND2x2_ASAP7_75t_L g3596 ( 
.A(n_3529),
.B(n_1978),
.Y(n_3596)
);

AO31x2_ASAP7_75t_L g3597 ( 
.A1(n_3554),
.A2(n_2079),
.A3(n_2087),
.B(n_2063),
.Y(n_3597)
);

AOI21xp5_ASAP7_75t_L g3598 ( 
.A1(n_3496),
.A2(n_1986),
.B(n_1979),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3525),
.A2(n_2004),
.B(n_1987),
.Y(n_3599)
);

AOI221xp5_ASAP7_75t_SL g3600 ( 
.A1(n_3545),
.A2(n_2011),
.B1(n_2026),
.B2(n_2024),
.C(n_2014),
.Y(n_3600)
);

NAND2x1p5_ASAP7_75t_L g3601 ( 
.A(n_3452),
.B(n_3358),
.Y(n_3601)
);

OAI21xp5_ASAP7_75t_L g3602 ( 
.A1(n_3489),
.A2(n_2042),
.B(n_2029),
.Y(n_3602)
);

INVx4_ASAP7_75t_L g3603 ( 
.A(n_3470),
.Y(n_3603)
);

OAI21x1_ASAP7_75t_L g3604 ( 
.A1(n_3475),
.A2(n_2051),
.B(n_2047),
.Y(n_3604)
);

O2A1O1Ixp5_ASAP7_75t_L g3605 ( 
.A1(n_3553),
.A2(n_2053),
.B(n_2057),
.C(n_2052),
.Y(n_3605)
);

OAI21xp5_ASAP7_75t_L g3606 ( 
.A1(n_3555),
.A2(n_2061),
.B(n_2058),
.Y(n_3606)
);

INVx4_ASAP7_75t_L g3607 ( 
.A(n_3448),
.Y(n_3607)
);

OAI21xp5_ASAP7_75t_L g3608 ( 
.A1(n_3534),
.A2(n_2068),
.B(n_2064),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3499),
.A2(n_2075),
.B(n_2074),
.Y(n_3609)
);

NAND2xp5_ASAP7_75t_L g3610 ( 
.A(n_3547),
.B(n_2090),
.Y(n_3610)
);

A2O1A1Ixp33_ASAP7_75t_L g3611 ( 
.A1(n_3517),
.A2(n_2097),
.B(n_1938),
.C(n_2037),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_L g3612 ( 
.A(n_3527),
.B(n_1596),
.Y(n_3612)
);

BUFx4f_ASAP7_75t_SL g3613 ( 
.A(n_3514),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3504),
.B(n_1600),
.Y(n_3614)
);

AOI21xp5_ASAP7_75t_L g3615 ( 
.A1(n_3492),
.A2(n_2067),
.B(n_1943),
.Y(n_3615)
);

INVx3_ASAP7_75t_L g3616 ( 
.A(n_3464),
.Y(n_3616)
);

INVx1_ASAP7_75t_L g3617 ( 
.A(n_3512),
.Y(n_3617)
);

AOI21x1_ASAP7_75t_L g3618 ( 
.A1(n_3520),
.A2(n_2096),
.B(n_2577),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3539),
.Y(n_3619)
);

INVx3_ASAP7_75t_L g3620 ( 
.A(n_3464),
.Y(n_3620)
);

NAND2xp5_ASAP7_75t_L g3621 ( 
.A(n_3511),
.B(n_3542),
.Y(n_3621)
);

INVx2_ASAP7_75t_L g3622 ( 
.A(n_3479),
.Y(n_3622)
);

OAI21xp5_ASAP7_75t_L g3623 ( 
.A1(n_3533),
.A2(n_1604),
.B(n_1603),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_3523),
.A2(n_1343),
.B(n_1317),
.Y(n_3624)
);

INVx3_ASAP7_75t_L g3625 ( 
.A(n_3467),
.Y(n_3625)
);

OAI21x1_ASAP7_75t_L g3626 ( 
.A1(n_3550),
.A2(n_1448),
.B(n_997),
.Y(n_3626)
);

AND2x4_ASAP7_75t_L g3627 ( 
.A(n_3474),
.B(n_2578),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_3500),
.B(n_1608),
.Y(n_3628)
);

OAI21x1_ASAP7_75t_L g3629 ( 
.A1(n_3497),
.A2(n_3519),
.B(n_3518),
.Y(n_3629)
);

AO21x1_ASAP7_75t_L g3630 ( 
.A1(n_3551),
.A2(n_1448),
.B(n_1935),
.Y(n_3630)
);

AOI21x1_ASAP7_75t_L g3631 ( 
.A1(n_3548),
.A2(n_3486),
.B(n_3482),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_L g3632 ( 
.A1(n_3521),
.A2(n_1448),
.B(n_998),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3481),
.B(n_1610),
.Y(n_3633)
);

OAI21xp5_ASAP7_75t_L g3634 ( 
.A1(n_3535),
.A2(n_1614),
.B(n_1613),
.Y(n_3634)
);

INVx6_ASAP7_75t_L g3635 ( 
.A(n_3459),
.Y(n_3635)
);

AOI21xp5_ASAP7_75t_L g3636 ( 
.A1(n_3546),
.A2(n_3552),
.B(n_3469),
.Y(n_3636)
);

AND2x4_ASAP7_75t_L g3637 ( 
.A(n_3477),
.B(n_2580),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_3556),
.A2(n_1693),
.B(n_1343),
.Y(n_3638)
);

AOI21xp5_ASAP7_75t_L g3639 ( 
.A1(n_3556),
.A2(n_1693),
.B(n_1343),
.Y(n_3639)
);

INVx2_ASAP7_75t_SL g3640 ( 
.A(n_3498),
.Y(n_3640)
);

AND2x2_ASAP7_75t_L g3641 ( 
.A(n_3483),
.B(n_1618),
.Y(n_3641)
);

OAI21xp33_ASAP7_75t_L g3642 ( 
.A1(n_3532),
.A2(n_1626),
.B(n_1623),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3488),
.B(n_1630),
.Y(n_3643)
);

NAND2xp5_ASAP7_75t_L g3644 ( 
.A(n_3491),
.B(n_1631),
.Y(n_3644)
);

A2O1A1Ixp33_ASAP7_75t_L g3645 ( 
.A1(n_3510),
.A2(n_2085),
.B(n_1637),
.C(n_1645),
.Y(n_3645)
);

OAI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_3537),
.A2(n_1650),
.B(n_1633),
.Y(n_3646)
);

NAND2xp5_ASAP7_75t_L g3647 ( 
.A(n_3455),
.B(n_1651),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3455),
.B(n_1653),
.Y(n_3648)
);

AO31x2_ASAP7_75t_L g3649 ( 
.A1(n_3508),
.A2(n_3543),
.A3(n_3507),
.B(n_3506),
.Y(n_3649)
);

INVx3_ASAP7_75t_L g3650 ( 
.A(n_3467),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3459),
.B(n_1659),
.Y(n_3651)
);

NAND3xp33_ASAP7_75t_L g3652 ( 
.A(n_3538),
.B(n_3549),
.C(n_3530),
.Y(n_3652)
);

OAI21x1_ASAP7_75t_L g3653 ( 
.A1(n_3460),
.A2(n_3513),
.B(n_3487),
.Y(n_3653)
);

AOI21x1_ASAP7_75t_L g3654 ( 
.A1(n_3450),
.A2(n_2589),
.B(n_2586),
.Y(n_3654)
);

INVx5_ASAP7_75t_L g3655 ( 
.A(n_3498),
.Y(n_3655)
);

OAI21x1_ASAP7_75t_L g3656 ( 
.A1(n_3495),
.A2(n_1448),
.B(n_999),
.Y(n_3656)
);

OAI21x1_ASAP7_75t_SL g3657 ( 
.A1(n_3449),
.A2(n_2),
.B(n_4),
.Y(n_3657)
);

BUFx2_ASAP7_75t_L g3658 ( 
.A(n_3515),
.Y(n_3658)
);

AOI21x1_ASAP7_75t_L g3659 ( 
.A1(n_3503),
.A2(n_1448),
.B(n_1693),
.Y(n_3659)
);

OAI21x1_ASAP7_75t_L g3660 ( 
.A1(n_3515),
.A2(n_1001),
.B(n_996),
.Y(n_3660)
);

OAI22x1_ASAP7_75t_L g3661 ( 
.A1(n_3536),
.A2(n_1666),
.B1(n_1670),
.B2(n_1663),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3502),
.A2(n_1852),
.B(n_1708),
.Y(n_3662)
);

OAI21x1_ASAP7_75t_L g3663 ( 
.A1(n_3478),
.A2(n_1004),
.B(n_1003),
.Y(n_3663)
);

OAI21x1_ASAP7_75t_L g3664 ( 
.A1(n_3544),
.A2(n_1009),
.B(n_1006),
.Y(n_3664)
);

INVx2_ASAP7_75t_L g3665 ( 
.A(n_3465),
.Y(n_3665)
);

A2O1A1Ixp33_ASAP7_75t_L g3666 ( 
.A1(n_3505),
.A2(n_1673),
.B(n_1676),
.C(n_1671),
.Y(n_3666)
);

INVx1_ASAP7_75t_L g3667 ( 
.A(n_3454),
.Y(n_3667)
);

OAI21x1_ASAP7_75t_L g3668 ( 
.A1(n_3544),
.A2(n_1020),
.B(n_1015),
.Y(n_3668)
);

AOI21xp5_ASAP7_75t_L g3669 ( 
.A1(n_3505),
.A2(n_1852),
.B(n_1708),
.Y(n_3669)
);

AOI21xp5_ASAP7_75t_L g3670 ( 
.A1(n_3561),
.A2(n_3567),
.B(n_3669),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3591),
.Y(n_3671)
);

BUFx2_ASAP7_75t_L g3672 ( 
.A(n_3560),
.Y(n_3672)
);

AOI21xp5_ASAP7_75t_L g3673 ( 
.A1(n_3566),
.A2(n_1685),
.B(n_1678),
.Y(n_3673)
);

AND2x4_ASAP7_75t_L g3674 ( 
.A(n_3585),
.B(n_1021),
.Y(n_3674)
);

AOI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3562),
.A2(n_1687),
.B(n_1686),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3569),
.B(n_1691),
.Y(n_3676)
);

BUFx2_ASAP7_75t_SL g3677 ( 
.A(n_3655),
.Y(n_3677)
);

INVx2_ASAP7_75t_L g3678 ( 
.A(n_3665),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_SL g3679 ( 
.A(n_3564),
.B(n_1307),
.Y(n_3679)
);

BUFx3_ASAP7_75t_L g3680 ( 
.A(n_3565),
.Y(n_3680)
);

NAND2xp5_ASAP7_75t_L g3681 ( 
.A(n_3572),
.B(n_1692),
.Y(n_3681)
);

INVx2_ASAP7_75t_SL g3682 ( 
.A(n_3635),
.Y(n_3682)
);

OR2x2_ASAP7_75t_L g3683 ( 
.A(n_3617),
.B(n_2),
.Y(n_3683)
);

AND2x2_ASAP7_75t_L g3684 ( 
.A(n_3573),
.B(n_4),
.Y(n_3684)
);

BUFx2_ASAP7_75t_L g3685 ( 
.A(n_3658),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_L g3686 ( 
.A1(n_3577),
.A2(n_1852),
.B(n_1708),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3622),
.Y(n_3687)
);

BUFx12f_ASAP7_75t_L g3688 ( 
.A(n_3595),
.Y(n_3688)
);

INVx1_ASAP7_75t_L g3689 ( 
.A(n_3619),
.Y(n_3689)
);

NAND2xp5_ASAP7_75t_SL g3690 ( 
.A(n_3647),
.B(n_1308),
.Y(n_3690)
);

INVx2_ASAP7_75t_SL g3691 ( 
.A(n_3635),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3621),
.B(n_1694),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3563),
.Y(n_3693)
);

AND2x2_ASAP7_75t_L g3694 ( 
.A(n_3596),
.B(n_5),
.Y(n_3694)
);

OR2x2_ASAP7_75t_L g3695 ( 
.A(n_3570),
.B(n_5),
.Y(n_3695)
);

CKINVDCx11_ASAP7_75t_R g3696 ( 
.A(n_3559),
.Y(n_3696)
);

AOI22xp33_ASAP7_75t_L g3697 ( 
.A1(n_3576),
.A2(n_1711),
.B1(n_1712),
.B2(n_1701),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3602),
.A2(n_1717),
.B1(n_1726),
.B2(n_1714),
.Y(n_3698)
);

NAND2xp33_ASAP7_75t_L g3699 ( 
.A(n_3666),
.B(n_1727),
.Y(n_3699)
);

BUFx6f_ASAP7_75t_L g3700 ( 
.A(n_3559),
.Y(n_3700)
);

AOI21xp5_ASAP7_75t_L g3701 ( 
.A1(n_3664),
.A2(n_1731),
.B(n_1729),
.Y(n_3701)
);

OA21x2_ASAP7_75t_L g3702 ( 
.A1(n_3630),
.A2(n_1744),
.B(n_1739),
.Y(n_3702)
);

INVx3_ASAP7_75t_L g3703 ( 
.A(n_3574),
.Y(n_3703)
);

OAI21x1_ASAP7_75t_SL g3704 ( 
.A1(n_3648),
.A2(n_6),
.B(n_7),
.Y(n_3704)
);

OR2x2_ASAP7_75t_L g3705 ( 
.A(n_3667),
.B(n_3610),
.Y(n_3705)
);

INVx2_ASAP7_75t_L g3706 ( 
.A(n_3629),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3593),
.B(n_1745),
.Y(n_3707)
);

BUFx3_ASAP7_75t_L g3708 ( 
.A(n_3574),
.Y(n_3708)
);

O2A1O1Ixp33_ASAP7_75t_SL g3709 ( 
.A1(n_3645),
.A2(n_9),
.B(n_6),
.C(n_8),
.Y(n_3709)
);

INVx6_ASAP7_75t_L g3710 ( 
.A(n_3655),
.Y(n_3710)
);

HB1xp67_ASAP7_75t_L g3711 ( 
.A(n_3631),
.Y(n_3711)
);

BUFx6f_ASAP7_75t_L g3712 ( 
.A(n_3588),
.Y(n_3712)
);

HAxp5_ASAP7_75t_L g3713 ( 
.A(n_3600),
.B(n_1746),
.CON(n_3713),
.SN(n_3713)
);

O2A1O1Ixp33_ASAP7_75t_SL g3714 ( 
.A1(n_3571),
.A2(n_3611),
.B(n_3608),
.C(n_3587),
.Y(n_3714)
);

HB1xp67_ASAP7_75t_L g3715 ( 
.A(n_3597),
.Y(n_3715)
);

AOI221xp5_ASAP7_75t_L g3716 ( 
.A1(n_3599),
.A2(n_1749),
.B1(n_1751),
.B2(n_1748),
.C(n_1747),
.Y(n_3716)
);

BUFx3_ASAP7_75t_L g3717 ( 
.A(n_3607),
.Y(n_3717)
);

AOI21xp5_ASAP7_75t_L g3718 ( 
.A1(n_3668),
.A2(n_1753),
.B(n_1752),
.Y(n_3718)
);

AND2x2_ASAP7_75t_L g3719 ( 
.A(n_3616),
.B(n_8),
.Y(n_3719)
);

INVx3_ASAP7_75t_L g3720 ( 
.A(n_3603),
.Y(n_3720)
);

INVx3_ASAP7_75t_L g3721 ( 
.A(n_3620),
.Y(n_3721)
);

NAND3xp33_ASAP7_75t_L g3722 ( 
.A(n_3589),
.B(n_1755),
.C(n_1754),
.Y(n_3722)
);

BUFx2_ASAP7_75t_L g3723 ( 
.A(n_3653),
.Y(n_3723)
);

AND2x2_ASAP7_75t_L g3724 ( 
.A(n_3625),
.B(n_9),
.Y(n_3724)
);

INVx2_ASAP7_75t_SL g3725 ( 
.A(n_3650),
.Y(n_3725)
);

NAND2xp5_ASAP7_75t_L g3726 ( 
.A(n_3584),
.B(n_1756),
.Y(n_3726)
);

AOI22xp33_ASAP7_75t_L g3727 ( 
.A1(n_3652),
.A2(n_1758),
.B1(n_1759),
.B2(n_1757),
.Y(n_3727)
);

OR2x2_ASAP7_75t_L g3728 ( 
.A(n_3583),
.B(n_10),
.Y(n_3728)
);

NAND2xp33_ASAP7_75t_L g3729 ( 
.A(n_3642),
.B(n_1764),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3636),
.Y(n_3730)
);

OR2x2_ASAP7_75t_L g3731 ( 
.A(n_3594),
.B(n_10),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_3568),
.B(n_1765),
.Y(n_3732)
);

INVxp67_ASAP7_75t_L g3733 ( 
.A(n_3641),
.Y(n_3733)
);

HB1xp67_ASAP7_75t_L g3734 ( 
.A(n_3597),
.Y(n_3734)
);

BUFx3_ASAP7_75t_L g3735 ( 
.A(n_3640),
.Y(n_3735)
);

INVx1_ASAP7_75t_L g3736 ( 
.A(n_3604),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3649),
.B(n_11),
.Y(n_3737)
);

OAI22xp33_ASAP7_75t_L g3738 ( 
.A1(n_3575),
.A2(n_1769),
.B1(n_1770),
.B2(n_1768),
.Y(n_3738)
);

CKINVDCx5p33_ASAP7_75t_R g3739 ( 
.A(n_3613),
.Y(n_3739)
);

INVx2_ASAP7_75t_SL g3740 ( 
.A(n_3627),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3609),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3618),
.Y(n_3742)
);

OAI21xp5_ASAP7_75t_L g3743 ( 
.A1(n_3605),
.A2(n_3623),
.B(n_3646),
.Y(n_3743)
);

NAND2xp5_ASAP7_75t_L g3744 ( 
.A(n_3598),
.B(n_1773),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3632),
.Y(n_3745)
);

NOR2xp33_ASAP7_75t_SL g3746 ( 
.A(n_3580),
.B(n_1781),
.Y(n_3746)
);

BUFx3_ASAP7_75t_L g3747 ( 
.A(n_3637),
.Y(n_3747)
);

NOR2xp33_ASAP7_75t_L g3748 ( 
.A(n_3628),
.B(n_1784),
.Y(n_3748)
);

CKINVDCx8_ASAP7_75t_R g3749 ( 
.A(n_3601),
.Y(n_3749)
);

AOI21xp5_ASAP7_75t_L g3750 ( 
.A1(n_3662),
.A2(n_1791),
.B(n_1790),
.Y(n_3750)
);

INVx3_ASAP7_75t_SL g3751 ( 
.A(n_3661),
.Y(n_3751)
);

NOR2x1_ASAP7_75t_SL g3752 ( 
.A(n_3659),
.B(n_1976),
.Y(n_3752)
);

CKINVDCx5p33_ASAP7_75t_R g3753 ( 
.A(n_3651),
.Y(n_3753)
);

INVx3_ASAP7_75t_L g3754 ( 
.A(n_3558),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3615),
.Y(n_3755)
);

INVx2_ASAP7_75t_SL g3756 ( 
.A(n_3649),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_L g3757 ( 
.A(n_3614),
.B(n_1794),
.Y(n_3757)
);

INVx3_ASAP7_75t_L g3758 ( 
.A(n_3654),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3582),
.Y(n_3759)
);

AOI22xp33_ASAP7_75t_L g3760 ( 
.A1(n_3581),
.A2(n_1804),
.B1(n_1809),
.B2(n_1796),
.Y(n_3760)
);

AOI21xp5_ASAP7_75t_L g3761 ( 
.A1(n_3624),
.A2(n_1815),
.B(n_1812),
.Y(n_3761)
);

BUFx6f_ASAP7_75t_L g3762 ( 
.A(n_3663),
.Y(n_3762)
);

AOI21xp5_ASAP7_75t_SL g3763 ( 
.A1(n_3638),
.A2(n_1314),
.B(n_1310),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3586),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3590),
.Y(n_3765)
);

AO21x2_ASAP7_75t_L g3766 ( 
.A1(n_3715),
.A2(n_3639),
.B(n_3592),
.Y(n_3766)
);

BUFx2_ASAP7_75t_L g3767 ( 
.A(n_3672),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3693),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3689),
.Y(n_3769)
);

INVxp67_ASAP7_75t_SL g3770 ( 
.A(n_3730),
.Y(n_3770)
);

OAI21x1_ASAP7_75t_L g3771 ( 
.A1(n_3670),
.A2(n_3686),
.B(n_3745),
.Y(n_3771)
);

AO21x2_ASAP7_75t_L g3772 ( 
.A1(n_3734),
.A2(n_3742),
.B(n_3711),
.Y(n_3772)
);

INVxp67_ASAP7_75t_SL g3773 ( 
.A(n_3723),
.Y(n_3773)
);

AND2x2_ASAP7_75t_L g3774 ( 
.A(n_3685),
.B(n_3633),
.Y(n_3774)
);

OAI21x1_ASAP7_75t_L g3775 ( 
.A1(n_3759),
.A2(n_3579),
.B(n_3626),
.Y(n_3775)
);

OAI21x1_ASAP7_75t_L g3776 ( 
.A1(n_3764),
.A2(n_3656),
.B(n_3660),
.Y(n_3776)
);

NOR2xp33_ASAP7_75t_L g3777 ( 
.A(n_3746),
.B(n_3612),
.Y(n_3777)
);

AOI21xp5_ASAP7_75t_L g3778 ( 
.A1(n_3679),
.A2(n_3714),
.B(n_3743),
.Y(n_3778)
);

OA21x2_ASAP7_75t_L g3779 ( 
.A1(n_3756),
.A2(n_3657),
.B(n_3606),
.Y(n_3779)
);

NAND2x1p5_ASAP7_75t_L g3780 ( 
.A(n_3700),
.B(n_3643),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3705),
.Y(n_3781)
);

NAND2x1p5_ASAP7_75t_L g3782 ( 
.A(n_3700),
.B(n_3644),
.Y(n_3782)
);

CKINVDCx16_ASAP7_75t_R g3783 ( 
.A(n_3688),
.Y(n_3783)
);

OAI21x1_ASAP7_75t_L g3784 ( 
.A1(n_3755),
.A2(n_3578),
.B(n_3634),
.Y(n_3784)
);

NOR2xp33_ASAP7_75t_L g3785 ( 
.A(n_3717),
.B(n_12),
.Y(n_3785)
);

BUFx6f_ASAP7_75t_L g3786 ( 
.A(n_3712),
.Y(n_3786)
);

INVxp67_ASAP7_75t_L g3787 ( 
.A(n_3725),
.Y(n_3787)
);

INVx1_ASAP7_75t_L g3788 ( 
.A(n_3671),
.Y(n_3788)
);

OAI21x1_ASAP7_75t_L g3789 ( 
.A1(n_3758),
.A2(n_2049),
.B(n_1976),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3678),
.Y(n_3790)
);

AO21x2_ASAP7_75t_L g3791 ( 
.A1(n_3765),
.A2(n_1330),
.B(n_1324),
.Y(n_3791)
);

CKINVDCx20_ASAP7_75t_R g3792 ( 
.A(n_3696),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3687),
.Y(n_3793)
);

NOR2xp33_ASAP7_75t_L g3794 ( 
.A(n_3712),
.B(n_13),
.Y(n_3794)
);

AOI22xp33_ASAP7_75t_L g3795 ( 
.A1(n_3697),
.A2(n_2049),
.B1(n_1976),
.B2(n_1820),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3736),
.Y(n_3796)
);

INVx3_ASAP7_75t_SL g3797 ( 
.A(n_3739),
.Y(n_3797)
);

INVx2_ASAP7_75t_L g3798 ( 
.A(n_3706),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3741),
.Y(n_3799)
);

OAI21x1_ASAP7_75t_L g3800 ( 
.A1(n_3701),
.A2(n_2049),
.B(n_1023),
.Y(n_3800)
);

O2A1O1Ixp33_ASAP7_75t_L g3801 ( 
.A1(n_3729),
.A2(n_1822),
.B(n_1826),
.C(n_1819),
.Y(n_3801)
);

AO21x2_ASAP7_75t_L g3802 ( 
.A1(n_3752),
.A2(n_3738),
.B(n_3704),
.Y(n_3802)
);

NAND2xp5_ASAP7_75t_L g3803 ( 
.A(n_3684),
.B(n_13),
.Y(n_3803)
);

BUFx3_ASAP7_75t_L g3804 ( 
.A(n_3680),
.Y(n_3804)
);

AOI22xp33_ASAP7_75t_L g3805 ( 
.A1(n_3737),
.A2(n_1833),
.B1(n_1834),
.B2(n_1828),
.Y(n_3805)
);

OAI21xp5_ASAP7_75t_L g3806 ( 
.A1(n_3675),
.A2(n_1842),
.B(n_1836),
.Y(n_3806)
);

OAI21x1_ASAP7_75t_L g3807 ( 
.A1(n_3718),
.A2(n_1024),
.B(n_1022),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3702),
.A2(n_1026),
.B(n_1025),
.Y(n_3808)
);

OAI22xp5_ASAP7_75t_L g3809 ( 
.A1(n_3727),
.A2(n_1850),
.B1(n_1851),
.B2(n_1846),
.Y(n_3809)
);

O2A1O1Ixp33_ASAP7_75t_L g3810 ( 
.A1(n_3699),
.A2(n_1854),
.B(n_1855),
.C(n_1853),
.Y(n_3810)
);

INVx2_ASAP7_75t_L g3811 ( 
.A(n_3695),
.Y(n_3811)
);

A2O1A1Ixp33_ASAP7_75t_L g3812 ( 
.A1(n_3748),
.A2(n_1859),
.B(n_1860),
.C(n_1857),
.Y(n_3812)
);

O2A1O1Ixp33_ASAP7_75t_L g3813 ( 
.A1(n_3709),
.A2(n_1865),
.B(n_1867),
.C(n_1864),
.Y(n_3813)
);

AO21x1_ASAP7_75t_L g3814 ( 
.A1(n_3683),
.A2(n_14),
.B(n_15),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_L g3815 ( 
.A(n_3708),
.B(n_14),
.Y(n_3815)
);

OAI21x1_ASAP7_75t_L g3816 ( 
.A1(n_3720),
.A2(n_3754),
.B(n_3750),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3762),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3762),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3728),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3694),
.B(n_15),
.Y(n_3820)
);

AND2x4_ASAP7_75t_L g3821 ( 
.A(n_3735),
.B(n_1027),
.Y(n_3821)
);

OAI21x1_ASAP7_75t_L g3822 ( 
.A1(n_3721),
.A2(n_1029),
.B(n_1028),
.Y(n_3822)
);

BUFx6f_ASAP7_75t_L g3823 ( 
.A(n_3710),
.Y(n_3823)
);

BUFx3_ASAP7_75t_L g3824 ( 
.A(n_3747),
.Y(n_3824)
);

NAND2xp5_ASAP7_75t_L g3825 ( 
.A(n_3731),
.B(n_16),
.Y(n_3825)
);

AND2x2_ASAP7_75t_L g3826 ( 
.A(n_3733),
.B(n_18),
.Y(n_3826)
);

OR2x2_ASAP7_75t_L g3827 ( 
.A(n_3676),
.B(n_18),
.Y(n_3827)
);

OAI21xp33_ASAP7_75t_L g3828 ( 
.A1(n_3744),
.A2(n_1872),
.B(n_1868),
.Y(n_3828)
);

INVx5_ASAP7_75t_L g3829 ( 
.A(n_3710),
.Y(n_3829)
);

AO21x2_ASAP7_75t_L g3830 ( 
.A1(n_3732),
.A2(n_1351),
.B(n_1338),
.Y(n_3830)
);

OAI21x1_ASAP7_75t_L g3831 ( 
.A1(n_3761),
.A2(n_1035),
.B(n_1031),
.Y(n_3831)
);

OAI21x1_ASAP7_75t_L g3832 ( 
.A1(n_3703),
.A2(n_1039),
.B(n_1036),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_3692),
.B(n_19),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3681),
.Y(n_3834)
);

AOI31xp33_ASAP7_75t_L g3835 ( 
.A1(n_3740),
.A2(n_1878),
.A3(n_1882),
.B(n_1876),
.Y(n_3835)
);

INVx2_ASAP7_75t_L g3836 ( 
.A(n_3674),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3719),
.Y(n_3837)
);

NAND2x1p5_ASAP7_75t_L g3838 ( 
.A(n_3682),
.B(n_1040),
.Y(n_3838)
);

BUFx12f_ASAP7_75t_L g3839 ( 
.A(n_3753),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3691),
.Y(n_3840)
);

AND2x4_ASAP7_75t_L g3841 ( 
.A(n_3724),
.B(n_1041),
.Y(n_3841)
);

INVx6_ASAP7_75t_L g3842 ( 
.A(n_3677),
.Y(n_3842)
);

OAI22xp5_ASAP7_75t_SL g3843 ( 
.A1(n_3792),
.A2(n_3751),
.B1(n_3749),
.B2(n_3698),
.Y(n_3843)
);

OAI22xp33_ASAP7_75t_L g3844 ( 
.A1(n_3778),
.A2(n_3722),
.B1(n_3726),
.B2(n_3707),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3767),
.B(n_3757),
.Y(n_3845)
);

INVxp67_ASAP7_75t_L g3846 ( 
.A(n_3840),
.Y(n_3846)
);

NOR2xp33_ASAP7_75t_L g3847 ( 
.A(n_3839),
.B(n_3690),
.Y(n_3847)
);

NOR2x1_ASAP7_75t_SL g3848 ( 
.A(n_3829),
.B(n_3763),
.Y(n_3848)
);

BUFx3_ASAP7_75t_L g3849 ( 
.A(n_3804),
.Y(n_3849)
);

NOR2x1_ASAP7_75t_L g3850 ( 
.A(n_3824),
.B(n_3673),
.Y(n_3850)
);

INVx3_ASAP7_75t_L g3851 ( 
.A(n_3823),
.Y(n_3851)
);

OAI21xp5_ASAP7_75t_SL g3852 ( 
.A1(n_3813),
.A2(n_3760),
.B(n_3716),
.Y(n_3852)
);

NAND3xp33_ASAP7_75t_L g3853 ( 
.A(n_3805),
.B(n_3834),
.C(n_3770),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_L g3854 ( 
.A(n_3768),
.B(n_1883),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3790),
.Y(n_3855)
);

INVx1_ASAP7_75t_L g3856 ( 
.A(n_3769),
.Y(n_3856)
);

AND2x4_ASAP7_75t_L g3857 ( 
.A(n_3829),
.B(n_21),
.Y(n_3857)
);

OAI22xp5_ASAP7_75t_L g3858 ( 
.A1(n_3825),
.A2(n_3713),
.B1(n_1887),
.B2(n_1890),
.Y(n_3858)
);

BUFx6f_ASAP7_75t_L g3859 ( 
.A(n_3786),
.Y(n_3859)
);

INVx4_ASAP7_75t_L g3860 ( 
.A(n_3786),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3811),
.B(n_1886),
.Y(n_3861)
);

CKINVDCx11_ASAP7_75t_R g3862 ( 
.A(n_3797),
.Y(n_3862)
);

OR2x6_ASAP7_75t_L g3863 ( 
.A(n_3842),
.B(n_21),
.Y(n_3863)
);

AND2x4_ASAP7_75t_L g3864 ( 
.A(n_3781),
.B(n_22),
.Y(n_3864)
);

AOI21xp5_ASAP7_75t_L g3865 ( 
.A1(n_3773),
.A2(n_1894),
.B(n_1893),
.Y(n_3865)
);

BUFx2_ASAP7_75t_L g3866 ( 
.A(n_3787),
.Y(n_3866)
);

CKINVDCx6p67_ASAP7_75t_R g3867 ( 
.A(n_3783),
.Y(n_3867)
);

INVx1_ASAP7_75t_L g3868 ( 
.A(n_3796),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3774),
.B(n_22),
.Y(n_3869)
);

OAI21x1_ASAP7_75t_L g3870 ( 
.A1(n_3771),
.A2(n_23),
.B(n_24),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_SL g3871 ( 
.A(n_3823),
.B(n_1897),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3799),
.Y(n_3872)
);

INVx4_ASAP7_75t_L g3873 ( 
.A(n_3821),
.Y(n_3873)
);

INVx3_ASAP7_75t_L g3874 ( 
.A(n_3780),
.Y(n_3874)
);

BUFx8_ASAP7_75t_SL g3875 ( 
.A(n_3820),
.Y(n_3875)
);

AOI22xp33_ASAP7_75t_L g3876 ( 
.A1(n_3814),
.A2(n_1904),
.B1(n_1907),
.B2(n_1901),
.Y(n_3876)
);

AND2x2_ASAP7_75t_L g3877 ( 
.A(n_3837),
.B(n_24),
.Y(n_3877)
);

INVx3_ASAP7_75t_L g3878 ( 
.A(n_3782),
.Y(n_3878)
);

AOI22xp33_ASAP7_75t_L g3879 ( 
.A1(n_3779),
.A2(n_3791),
.B1(n_3819),
.B2(n_3836),
.Y(n_3879)
);

INVx1_ASAP7_75t_L g3880 ( 
.A(n_3788),
.Y(n_3880)
);

NAND2xp5_ASAP7_75t_L g3881 ( 
.A(n_3826),
.B(n_1908),
.Y(n_3881)
);

AOI22xp33_ASAP7_75t_L g3882 ( 
.A1(n_3828),
.A2(n_3784),
.B1(n_3777),
.B2(n_3806),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_L g3883 ( 
.A(n_3793),
.B(n_3817),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_L g3884 ( 
.A(n_3818),
.B(n_1909),
.Y(n_3884)
);

AND2x2_ASAP7_75t_L g3885 ( 
.A(n_3794),
.B(n_25),
.Y(n_3885)
);

INVx3_ASAP7_75t_L g3886 ( 
.A(n_3816),
.Y(n_3886)
);

CKINVDCx16_ASAP7_75t_R g3887 ( 
.A(n_3785),
.Y(n_3887)
);

INVxp67_ASAP7_75t_SL g3888 ( 
.A(n_3798),
.Y(n_3888)
);

AND2x2_ASAP7_75t_L g3889 ( 
.A(n_3803),
.B(n_26),
.Y(n_3889)
);

OAI22xp5_ASAP7_75t_L g3890 ( 
.A1(n_3827),
.A2(n_1915),
.B1(n_1916),
.B2(n_1914),
.Y(n_3890)
);

NAND3xp33_ASAP7_75t_SL g3891 ( 
.A(n_3833),
.B(n_2093),
.C(n_2089),
.Y(n_3891)
);

OAI22xp5_ASAP7_75t_L g3892 ( 
.A1(n_3812),
.A2(n_1920),
.B1(n_1922),
.B2(n_1918),
.Y(n_3892)
);

AOI22xp33_ASAP7_75t_L g3893 ( 
.A1(n_3830),
.A2(n_3802),
.B1(n_3795),
.B2(n_3800),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3772),
.Y(n_3894)
);

INVx3_ASAP7_75t_L g3895 ( 
.A(n_3841),
.Y(n_3895)
);

OR2x6_ASAP7_75t_L g3896 ( 
.A(n_3838),
.B(n_26),
.Y(n_3896)
);

INVx1_ASAP7_75t_L g3897 ( 
.A(n_3766),
.Y(n_3897)
);

CKINVDCx6p67_ASAP7_75t_R g3898 ( 
.A(n_3835),
.Y(n_3898)
);

BUFx2_ASAP7_75t_L g3899 ( 
.A(n_3815),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_L g3900 ( 
.A(n_3810),
.B(n_27),
.Y(n_3900)
);

INVx2_ASAP7_75t_L g3901 ( 
.A(n_3776),
.Y(n_3901)
);

INVx2_ASAP7_75t_L g3902 ( 
.A(n_3775),
.Y(n_3902)
);

CKINVDCx16_ASAP7_75t_R g3903 ( 
.A(n_3809),
.Y(n_3903)
);

OR2x6_ASAP7_75t_L g3904 ( 
.A(n_3822),
.B(n_27),
.Y(n_3904)
);

CKINVDCx11_ASAP7_75t_R g3905 ( 
.A(n_3801),
.Y(n_3905)
);

O2A1O1Ixp5_ASAP7_75t_SL g3906 ( 
.A1(n_3808),
.A2(n_30),
.B(n_28),
.C(n_29),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_3807),
.B(n_1930),
.Y(n_3907)
);

AOI21xp33_ASAP7_75t_L g3908 ( 
.A1(n_3832),
.A2(n_1942),
.B(n_1932),
.Y(n_3908)
);

BUFx6f_ASAP7_75t_L g3909 ( 
.A(n_3831),
.Y(n_3909)
);

AOI22xp33_ASAP7_75t_L g3910 ( 
.A1(n_3789),
.A2(n_1945),
.B1(n_1946),
.B2(n_1944),
.Y(n_3910)
);

NAND2xp33_ASAP7_75t_R g3911 ( 
.A(n_3777),
.B(n_28),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_3767),
.B(n_1947),
.Y(n_3912)
);

BUFx6f_ASAP7_75t_L g3913 ( 
.A(n_3786),
.Y(n_3913)
);

AOI22xp5_ASAP7_75t_L g3914 ( 
.A1(n_3778),
.A2(n_1949),
.B1(n_1952),
.B2(n_1948),
.Y(n_3914)
);

AND2x2_ASAP7_75t_L g3915 ( 
.A(n_3767),
.B(n_29),
.Y(n_3915)
);

INVx1_ASAP7_75t_L g3916 ( 
.A(n_3769),
.Y(n_3916)
);

INVx1_ASAP7_75t_L g3917 ( 
.A(n_3769),
.Y(n_3917)
);

AOI21xp5_ASAP7_75t_L g3918 ( 
.A1(n_3778),
.A2(n_1956),
.B(n_1955),
.Y(n_3918)
);

NAND2x1_ASAP7_75t_L g3919 ( 
.A(n_3767),
.B(n_30),
.Y(n_3919)
);

NAND2x1p5_ASAP7_75t_L g3920 ( 
.A(n_3829),
.B(n_31),
.Y(n_3920)
);

AND2x4_ASAP7_75t_L g3921 ( 
.A(n_3767),
.B(n_31),
.Y(n_3921)
);

INVx1_ASAP7_75t_L g3922 ( 
.A(n_3868),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_L g3923 ( 
.A(n_3867),
.B(n_32),
.Y(n_3923)
);

INVx1_ASAP7_75t_L g3924 ( 
.A(n_3872),
.Y(n_3924)
);

BUFx6f_ASAP7_75t_L g3925 ( 
.A(n_3862),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3856),
.Y(n_3926)
);

INVx1_ASAP7_75t_L g3927 ( 
.A(n_3916),
.Y(n_3927)
);

AND2x2_ASAP7_75t_L g3928 ( 
.A(n_3866),
.B(n_33),
.Y(n_3928)
);

AO21x2_ASAP7_75t_L g3929 ( 
.A1(n_3897),
.A2(n_1958),
.B(n_1957),
.Y(n_3929)
);

INVx2_ASAP7_75t_L g3930 ( 
.A(n_3855),
.Y(n_3930)
);

BUFx6f_ASAP7_75t_L g3931 ( 
.A(n_3849),
.Y(n_3931)
);

INVx1_ASAP7_75t_L g3932 ( 
.A(n_3917),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3880),
.Y(n_3933)
);

INVx1_ASAP7_75t_L g3934 ( 
.A(n_3883),
.Y(n_3934)
);

HB1xp67_ASAP7_75t_L g3935 ( 
.A(n_3846),
.Y(n_3935)
);

INVx1_ASAP7_75t_L g3936 ( 
.A(n_3894),
.Y(n_3936)
);

AO21x2_ASAP7_75t_L g3937 ( 
.A1(n_3901),
.A2(n_1968),
.B(n_1959),
.Y(n_3937)
);

OR2x2_ASAP7_75t_L g3938 ( 
.A(n_3845),
.B(n_33),
.Y(n_3938)
);

INVx1_ASAP7_75t_L g3939 ( 
.A(n_3888),
.Y(n_3939)
);

INVx2_ASAP7_75t_L g3940 ( 
.A(n_3886),
.Y(n_3940)
);

BUFx2_ASAP7_75t_L g3941 ( 
.A(n_3860),
.Y(n_3941)
);

AND2x2_ASAP7_75t_L g3942 ( 
.A(n_3899),
.B(n_34),
.Y(n_3942)
);

INVx2_ASAP7_75t_L g3943 ( 
.A(n_3902),
.Y(n_3943)
);

INVx2_ASAP7_75t_L g3944 ( 
.A(n_3874),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3853),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_3854),
.Y(n_3946)
);

AOI21xp5_ASAP7_75t_L g3947 ( 
.A1(n_3893),
.A2(n_1975),
.B(n_1969),
.Y(n_3947)
);

BUFx5_ASAP7_75t_L g3948 ( 
.A(n_3857),
.Y(n_3948)
);

AO21x2_ASAP7_75t_L g3949 ( 
.A1(n_3912),
.A2(n_1990),
.B(n_1981),
.Y(n_3949)
);

INVx3_ASAP7_75t_L g3950 ( 
.A(n_3851),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3877),
.Y(n_3951)
);

AND2x4_ASAP7_75t_L g3952 ( 
.A(n_3895),
.B(n_35),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_3915),
.Y(n_3953)
);

OAI21xp5_ASAP7_75t_L g3954 ( 
.A1(n_3882),
.A2(n_1994),
.B(n_1992),
.Y(n_3954)
);

OAI21x1_ASAP7_75t_SL g3955 ( 
.A1(n_3873),
.A2(n_36),
.B(n_37),
.Y(n_3955)
);

INVx3_ASAP7_75t_L g3956 ( 
.A(n_3859),
.Y(n_3956)
);

INVx1_ASAP7_75t_L g3957 ( 
.A(n_3878),
.Y(n_3957)
);

AO21x2_ASAP7_75t_L g3958 ( 
.A1(n_3861),
.A2(n_1999),
.B(n_1995),
.Y(n_3958)
);

INVx1_ASAP7_75t_L g3959 ( 
.A(n_3864),
.Y(n_3959)
);

INVx2_ASAP7_75t_L g3960 ( 
.A(n_3909),
.Y(n_3960)
);

INVx1_ASAP7_75t_L g3961 ( 
.A(n_3870),
.Y(n_3961)
);

INVx1_ASAP7_75t_L g3962 ( 
.A(n_3884),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3909),
.Y(n_3963)
);

AND2x2_ASAP7_75t_L g3964 ( 
.A(n_3887),
.B(n_38),
.Y(n_3964)
);

AO31x2_ASAP7_75t_L g3965 ( 
.A1(n_3847),
.A2(n_3848),
.A3(n_3900),
.B(n_3890),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3879),
.Y(n_3966)
);

INVx2_ASAP7_75t_L g3967 ( 
.A(n_3859),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3869),
.B(n_38),
.Y(n_3968)
);

INVx1_ASAP7_75t_L g3969 ( 
.A(n_3921),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_3913),
.Y(n_3970)
);

INVx1_ASAP7_75t_L g3971 ( 
.A(n_3913),
.Y(n_3971)
);

OA21x2_ASAP7_75t_L g3972 ( 
.A1(n_3865),
.A2(n_2005),
.B(n_2001),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3919),
.Y(n_3973)
);

BUFx2_ASAP7_75t_L g3974 ( 
.A(n_3863),
.Y(n_3974)
);

INVx2_ASAP7_75t_L g3975 ( 
.A(n_3904),
.Y(n_3975)
);

INVx1_ASAP7_75t_L g3976 ( 
.A(n_3850),
.Y(n_3976)
);

INVx2_ASAP7_75t_L g3977 ( 
.A(n_3904),
.Y(n_3977)
);

OR2x6_ASAP7_75t_L g3978 ( 
.A(n_3863),
.B(n_3843),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_3889),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3885),
.Y(n_3980)
);

OAI21x1_ASAP7_75t_L g3981 ( 
.A1(n_3906),
.A2(n_39),
.B(n_40),
.Y(n_3981)
);

HB1xp67_ASAP7_75t_L g3982 ( 
.A(n_3881),
.Y(n_3982)
);

INVx3_ASAP7_75t_L g3983 ( 
.A(n_3875),
.Y(n_3983)
);

INVx3_ASAP7_75t_L g3984 ( 
.A(n_3920),
.Y(n_3984)
);

AO21x2_ASAP7_75t_L g3985 ( 
.A1(n_3907),
.A2(n_3844),
.B(n_3908),
.Y(n_3985)
);

OR2x6_ASAP7_75t_L g3986 ( 
.A(n_3896),
.B(n_39),
.Y(n_3986)
);

INVx3_ASAP7_75t_L g3987 ( 
.A(n_3896),
.Y(n_3987)
);

INVx1_ASAP7_75t_L g3988 ( 
.A(n_3903),
.Y(n_3988)
);

AND2x4_ASAP7_75t_L g3989 ( 
.A(n_3871),
.B(n_41),
.Y(n_3989)
);

OAI22xp33_ASAP7_75t_L g3990 ( 
.A1(n_3988),
.A2(n_3911),
.B1(n_3898),
.B2(n_3914),
.Y(n_3990)
);

OR2x2_ASAP7_75t_L g3991 ( 
.A(n_3945),
.B(n_3876),
.Y(n_3991)
);

BUFx2_ASAP7_75t_L g3992 ( 
.A(n_3925),
.Y(n_3992)
);

INVx1_ASAP7_75t_L g3993 ( 
.A(n_3934),
.Y(n_3993)
);

AOI22xp33_ASAP7_75t_L g3994 ( 
.A1(n_3966),
.A2(n_3905),
.B1(n_3858),
.B2(n_3918),
.Y(n_3994)
);

AOI22xp33_ASAP7_75t_L g3995 ( 
.A1(n_3985),
.A2(n_3891),
.B1(n_3892),
.B2(n_3910),
.Y(n_3995)
);

AND2x2_ASAP7_75t_L g3996 ( 
.A(n_3950),
.B(n_3941),
.Y(n_3996)
);

INVx1_ASAP7_75t_L g3997 ( 
.A(n_3922),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3976),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3946),
.B(n_3852),
.Y(n_3999)
);

AOI22xp33_ASAP7_75t_L g4000 ( 
.A1(n_3954),
.A2(n_2007),
.B1(n_2008),
.B2(n_2006),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3924),
.Y(n_4001)
);

AOI22xp33_ASAP7_75t_L g4002 ( 
.A1(n_3947),
.A2(n_2016),
.B1(n_2017),
.B2(n_2012),
.Y(n_4002)
);

OAI33xp33_ASAP7_75t_L g4003 ( 
.A1(n_3962),
.A2(n_2023),
.A3(n_2021),
.B1(n_2025),
.B2(n_2022),
.B3(n_2018),
.Y(n_4003)
);

AOI21xp33_ASAP7_75t_L g4004 ( 
.A1(n_3961),
.A2(n_2028),
.B(n_2027),
.Y(n_4004)
);

HB1xp67_ASAP7_75t_L g4005 ( 
.A(n_3926),
.Y(n_4005)
);

AO21x2_ASAP7_75t_L g4006 ( 
.A1(n_3940),
.A2(n_41),
.B(n_42),
.Y(n_4006)
);

OAI21xp5_ASAP7_75t_L g4007 ( 
.A1(n_3964),
.A2(n_2034),
.B(n_2033),
.Y(n_4007)
);

AOI221xp5_ASAP7_75t_L g4008 ( 
.A1(n_3982),
.A2(n_2046),
.B1(n_2055),
.B2(n_2043),
.C(n_2036),
.Y(n_4008)
);

OAI22xp33_ASAP7_75t_L g4009 ( 
.A1(n_3978),
.A2(n_2088),
.B1(n_2066),
.B2(n_2060),
.Y(n_4009)
);

AOI22xp33_ASAP7_75t_L g4010 ( 
.A1(n_3975),
.A2(n_2065),
.B1(n_2071),
.B2(n_2059),
.Y(n_4010)
);

BUFx2_ASAP7_75t_L g4011 ( 
.A(n_3948),
.Y(n_4011)
);

AOI22xp33_ASAP7_75t_L g4012 ( 
.A1(n_3977),
.A2(n_2077),
.B1(n_2081),
.B2(n_2076),
.Y(n_4012)
);

OAI22xp33_ASAP7_75t_L g4013 ( 
.A1(n_3986),
.A2(n_2084),
.B1(n_2086),
.B2(n_2083),
.Y(n_4013)
);

OAI22xp33_ASAP7_75t_L g4014 ( 
.A1(n_3974),
.A2(n_2039),
.B1(n_2044),
.B2(n_2031),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3967),
.B(n_42),
.Y(n_4015)
);

INVx2_ASAP7_75t_L g4016 ( 
.A(n_3943),
.Y(n_4016)
);

O2A1O1Ixp5_ASAP7_75t_L g4017 ( 
.A1(n_3973),
.A2(n_45),
.B(n_43),
.C(n_44),
.Y(n_4017)
);

OAI22xp5_ASAP7_75t_SL g4018 ( 
.A1(n_3923),
.A2(n_46),
.B1(n_43),
.B2(n_44),
.Y(n_4018)
);

OAI21xp33_ASAP7_75t_L g4019 ( 
.A1(n_3928),
.A2(n_3933),
.B(n_3932),
.Y(n_4019)
);

INVx1_ASAP7_75t_L g4020 ( 
.A(n_3927),
.Y(n_4020)
);

AO31x2_ASAP7_75t_L g4021 ( 
.A1(n_3936),
.A2(n_3963),
.A3(n_3960),
.B(n_3944),
.Y(n_4021)
);

AOI22xp33_ASAP7_75t_L g4022 ( 
.A1(n_3929),
.A2(n_1355),
.B1(n_1365),
.B2(n_1354),
.Y(n_4022)
);

OA21x2_ASAP7_75t_L g4023 ( 
.A1(n_3939),
.A2(n_3930),
.B(n_3969),
.Y(n_4023)
);

INVx2_ASAP7_75t_L g4024 ( 
.A(n_3935),
.Y(n_4024)
);

OAI221xp5_ASAP7_75t_SL g4025 ( 
.A1(n_3938),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.C(n_49),
.Y(n_4025)
);

AOI22xp5_ASAP7_75t_L g4026 ( 
.A1(n_3937),
.A2(n_1380),
.B1(n_1385),
.B2(n_1376),
.Y(n_4026)
);

AOI22xp33_ASAP7_75t_L g4027 ( 
.A1(n_3958),
.A2(n_1401),
.B1(n_1407),
.B2(n_1399),
.Y(n_4027)
);

BUFx6f_ASAP7_75t_L g4028 ( 
.A(n_3931),
.Y(n_4028)
);

AOI221xp5_ASAP7_75t_L g4029 ( 
.A1(n_3949),
.A2(n_3955),
.B1(n_3942),
.B2(n_3989),
.C(n_3951),
.Y(n_4029)
);

OR2x6_ASAP7_75t_L g4030 ( 
.A(n_3952),
.B(n_47),
.Y(n_4030)
);

AOI21xp5_ASAP7_75t_L g4031 ( 
.A1(n_3957),
.A2(n_1419),
.B(n_1416),
.Y(n_4031)
);

OAI221xp5_ASAP7_75t_L g4032 ( 
.A1(n_3972),
.A2(n_3987),
.B1(n_3979),
.B2(n_3953),
.C(n_3980),
.Y(n_4032)
);

OAI21x1_ASAP7_75t_L g4033 ( 
.A1(n_3970),
.A2(n_50),
.B(n_51),
.Y(n_4033)
);

NAND3xp33_ASAP7_75t_L g4034 ( 
.A(n_3971),
.B(n_1445),
.C(n_1423),
.Y(n_4034)
);

AOI22xp33_ASAP7_75t_L g4035 ( 
.A1(n_3959),
.A2(n_1454),
.B1(n_1458),
.B2(n_1451),
.Y(n_4035)
);

INVx3_ASAP7_75t_L g4036 ( 
.A(n_3948),
.Y(n_4036)
);

NOR2x1_ASAP7_75t_SL g4037 ( 
.A(n_3968),
.B(n_50),
.Y(n_4037)
);

OAI22xp33_ASAP7_75t_L g4038 ( 
.A1(n_3984),
.A2(n_3956),
.B1(n_3983),
.B2(n_3965),
.Y(n_4038)
);

OAI22xp5_ASAP7_75t_L g4039 ( 
.A1(n_3948),
.A2(n_1965),
.B1(n_1983),
.B2(n_1962),
.Y(n_4039)
);

AOI221xp5_ASAP7_75t_L g4040 ( 
.A1(n_3981),
.A2(n_1486),
.B1(n_1488),
.B2(n_1485),
.C(n_1462),
.Y(n_4040)
);

OAI221xp5_ASAP7_75t_L g4041 ( 
.A1(n_3954),
.A2(n_1514),
.B1(n_1521),
.B2(n_1499),
.C(n_1495),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3950),
.B(n_52),
.Y(n_4042)
);

OAI21xp5_ASAP7_75t_L g4043 ( 
.A1(n_3945),
.A2(n_1546),
.B(n_1541),
.Y(n_4043)
);

AOI221xp5_ASAP7_75t_L g4044 ( 
.A1(n_3945),
.A2(n_1602),
.B1(n_1621),
.B2(n_1597),
.C(n_1592),
.Y(n_4044)
);

AOI22xp33_ASAP7_75t_L g4045 ( 
.A1(n_3966),
.A2(n_1636),
.B1(n_1638),
.B2(n_1629),
.Y(n_4045)
);

INVx8_ASAP7_75t_L g4046 ( 
.A(n_3986),
.Y(n_4046)
);

AOI22xp33_ASAP7_75t_L g4047 ( 
.A1(n_3966),
.A2(n_1647),
.B1(n_1652),
.B2(n_1639),
.Y(n_4047)
);

AOI22xp33_ASAP7_75t_L g4048 ( 
.A1(n_3966),
.A2(n_1657),
.B1(n_1662),
.B2(n_1654),
.Y(n_4048)
);

AOI21xp5_ASAP7_75t_SL g4049 ( 
.A1(n_3976),
.A2(n_1667),
.B(n_1664),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_L g4050 ( 
.A(n_3945),
.B(n_52),
.Y(n_4050)
);

AO21x2_ASAP7_75t_L g4051 ( 
.A1(n_3976),
.A2(n_53),
.B(n_54),
.Y(n_4051)
);

INVx1_ASAP7_75t_L g4052 ( 
.A(n_3934),
.Y(n_4052)
);

AOI22xp33_ASAP7_75t_L g4053 ( 
.A1(n_3966),
.A2(n_1680),
.B1(n_1688),
.B2(n_1674),
.Y(n_4053)
);

BUFx6f_ASAP7_75t_L g4054 ( 
.A(n_3925),
.Y(n_4054)
);

OR2x2_ASAP7_75t_L g4055 ( 
.A(n_3945),
.B(n_53),
.Y(n_4055)
);

OAI22xp33_ASAP7_75t_L g4056 ( 
.A1(n_3988),
.A2(n_1954),
.B1(n_1996),
.B2(n_1939),
.Y(n_4056)
);

AOI22xp33_ASAP7_75t_SL g4057 ( 
.A1(n_3985),
.A2(n_1702),
.B1(n_1720),
.B2(n_1689),
.Y(n_4057)
);

AND2x2_ASAP7_75t_L g4058 ( 
.A(n_3950),
.B(n_54),
.Y(n_4058)
);

AOI22xp33_ASAP7_75t_L g4059 ( 
.A1(n_3966),
.A2(n_1732),
.B1(n_1737),
.B2(n_1722),
.Y(n_4059)
);

OAI31xp33_ASAP7_75t_L g4060 ( 
.A1(n_3945),
.A2(n_58),
.A3(n_59),
.B(n_56),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3934),
.Y(n_4061)
);

OR2x2_ASAP7_75t_L g4062 ( 
.A(n_3945),
.B(n_55),
.Y(n_4062)
);

INVx2_ASAP7_75t_L g4063 ( 
.A(n_3976),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_L g4064 ( 
.A(n_3945),
.B(n_55),
.Y(n_4064)
);

A2O1A1Ixp33_ASAP7_75t_L g4065 ( 
.A1(n_3954),
.A2(n_1750),
.B(n_1762),
.C(n_1743),
.Y(n_4065)
);

AOI22xp33_ASAP7_75t_L g4066 ( 
.A1(n_3966),
.A2(n_1767),
.B1(n_1777),
.B2(n_1763),
.Y(n_4066)
);

OAI21x1_ASAP7_75t_L g4067 ( 
.A1(n_3940),
.A2(n_56),
.B(n_58),
.Y(n_4067)
);

OAI211xp5_ASAP7_75t_SL g4068 ( 
.A1(n_3945),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_4068)
);

AOI22xp33_ASAP7_75t_L g4069 ( 
.A1(n_3966),
.A2(n_1788),
.B1(n_1800),
.B2(n_1783),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3934),
.Y(n_4070)
);

HB1xp67_ASAP7_75t_L g4071 ( 
.A(n_3976),
.Y(n_4071)
);

NAND4xp25_ASAP7_75t_L g4072 ( 
.A(n_3923),
.B(n_63),
.C(n_60),
.D(n_62),
.Y(n_4072)
);

OAI221xp5_ASAP7_75t_L g4073 ( 
.A1(n_3954),
.A2(n_1835),
.B1(n_1839),
.B2(n_1821),
.C(n_1805),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3976),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3976),
.Y(n_4075)
);

INVx2_ASAP7_75t_L g4076 ( 
.A(n_3976),
.Y(n_4076)
);

AOI22xp33_ASAP7_75t_L g4077 ( 
.A1(n_3966),
.A2(n_1847),
.B1(n_1848),
.B2(n_1843),
.Y(n_4077)
);

CKINVDCx14_ASAP7_75t_R g4078 ( 
.A(n_3925),
.Y(n_4078)
);

AO21x2_ASAP7_75t_L g4079 ( 
.A1(n_3976),
.A2(n_64),
.B(n_65),
.Y(n_4079)
);

NAND2x1_ASAP7_75t_L g4080 ( 
.A(n_3976),
.B(n_64),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3934),
.Y(n_4081)
);

HB1xp67_ASAP7_75t_L g4082 ( 
.A(n_3976),
.Y(n_4082)
);

OAI22xp5_ASAP7_75t_L g4083 ( 
.A1(n_3945),
.A2(n_2003),
.B1(n_2054),
.B2(n_1997),
.Y(n_4083)
);

OAI211xp5_ASAP7_75t_L g4084 ( 
.A1(n_3923),
.A2(n_67),
.B(n_65),
.C(n_66),
.Y(n_4084)
);

AOI22xp33_ASAP7_75t_SL g4085 ( 
.A1(n_3985),
.A2(n_1858),
.B1(n_1869),
.B2(n_1849),
.Y(n_4085)
);

OA21x2_ASAP7_75t_L g4086 ( 
.A1(n_3945),
.A2(n_1921),
.B(n_1874),
.Y(n_4086)
);

AOI22xp33_ASAP7_75t_L g4087 ( 
.A1(n_3966),
.A2(n_1933),
.B1(n_1934),
.B2(n_1931),
.Y(n_4087)
);

AOI221xp5_ASAP7_75t_L g4088 ( 
.A1(n_3945),
.A2(n_2099),
.B1(n_2091),
.B2(n_2062),
.C(n_68),
.Y(n_4088)
);

OR2x6_ASAP7_75t_L g4089 ( 
.A(n_3978),
.B(n_66),
.Y(n_4089)
);

AOI222xp33_ASAP7_75t_L g4090 ( 
.A1(n_3954),
.A2(n_70),
.B1(n_72),
.B2(n_67),
.C1(n_69),
.C2(n_71),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3976),
.Y(n_4091)
);

NAND3xp33_ASAP7_75t_L g4092 ( 
.A(n_3945),
.B(n_70),
.C(n_71),
.Y(n_4092)
);

INVxp67_ASAP7_75t_SL g4093 ( 
.A(n_3976),
.Y(n_4093)
);

AOI22xp5_ASAP7_75t_SL g4094 ( 
.A1(n_3988),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.Y(n_4094)
);

AOI21xp5_ASAP7_75t_L g4095 ( 
.A1(n_3985),
.A2(n_76),
.B(n_77),
.Y(n_4095)
);

INVx1_ASAP7_75t_SL g4096 ( 
.A(n_3983),
.Y(n_4096)
);

AOI22xp33_ASAP7_75t_SL g4097 ( 
.A1(n_3985),
.A2(n_85),
.B1(n_94),
.B2(n_76),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3945),
.B(n_77),
.Y(n_4098)
);

AOI22xp33_ASAP7_75t_L g4099 ( 
.A1(n_3966),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.Y(n_4099)
);

OAI211xp5_ASAP7_75t_L g4100 ( 
.A1(n_3923),
.A2(n_80),
.B(n_78),
.C(n_79),
.Y(n_4100)
);

NAND3xp33_ASAP7_75t_L g4101 ( 
.A(n_3945),
.B(n_82),
.C(n_83),
.Y(n_4101)
);

NAND3xp33_ASAP7_75t_L g4102 ( 
.A(n_3945),
.B(n_82),
.C(n_84),
.Y(n_4102)
);

AOI22xp33_ASAP7_75t_SL g4103 ( 
.A1(n_3985),
.A2(n_94),
.B1(n_103),
.B2(n_85),
.Y(n_4103)
);

AOI22xp33_ASAP7_75t_L g4104 ( 
.A1(n_3966),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_4104)
);

INVx1_ASAP7_75t_L g4105 ( 
.A(n_3934),
.Y(n_4105)
);

AOI21xp5_ASAP7_75t_L g4106 ( 
.A1(n_3985),
.A2(n_86),
.B(n_88),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_4005),
.Y(n_4107)
);

INVx1_ASAP7_75t_L g4108 ( 
.A(n_3997),
.Y(n_4108)
);

AND2x2_ASAP7_75t_L g4109 ( 
.A(n_3996),
.B(n_89),
.Y(n_4109)
);

INVx1_ASAP7_75t_L g4110 ( 
.A(n_4001),
.Y(n_4110)
);

HB1xp67_ASAP7_75t_L g4111 ( 
.A(n_4024),
.Y(n_4111)
);

CKINVDCx16_ASAP7_75t_R g4112 ( 
.A(n_4078),
.Y(n_4112)
);

INVx1_ASAP7_75t_L g4113 ( 
.A(n_4020),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_4011),
.B(n_89),
.Y(n_4114)
);

INVx1_ASAP7_75t_L g4115 ( 
.A(n_3993),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_L g4116 ( 
.A(n_3999),
.B(n_90),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_4052),
.Y(n_4117)
);

AOI22xp33_ASAP7_75t_L g4118 ( 
.A1(n_4095),
.A2(n_93),
.B1(n_90),
.B2(n_92),
.Y(n_4118)
);

INVx1_ASAP7_75t_L g4119 ( 
.A(n_4061),
.Y(n_4119)
);

AOI22xp33_ASAP7_75t_L g4120 ( 
.A1(n_4106),
.A2(n_98),
.B1(n_95),
.B2(n_97),
.Y(n_4120)
);

INVx1_ASAP7_75t_L g4121 ( 
.A(n_4070),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4081),
.Y(n_4122)
);

AND2x2_ASAP7_75t_L g4123 ( 
.A(n_4036),
.B(n_97),
.Y(n_4123)
);

AND2x2_ASAP7_75t_L g4124 ( 
.A(n_4071),
.B(n_98),
.Y(n_4124)
);

NOR2xp33_ASAP7_75t_L g4125 ( 
.A(n_4096),
.B(n_99),
.Y(n_4125)
);

INVx1_ASAP7_75t_L g4126 ( 
.A(n_4105),
.Y(n_4126)
);

AND2x2_ASAP7_75t_L g4127 ( 
.A(n_4082),
.B(n_100),
.Y(n_4127)
);

OR2x2_ASAP7_75t_L g4128 ( 
.A(n_4055),
.B(n_100),
.Y(n_4128)
);

OAI21xp5_ASAP7_75t_L g4129 ( 
.A1(n_4057),
.A2(n_101),
.B(n_102),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_4023),
.Y(n_4130)
);

HB1xp67_ASAP7_75t_L g4131 ( 
.A(n_3998),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_3992),
.B(n_101),
.Y(n_4132)
);

HB1xp67_ASAP7_75t_L g4133 ( 
.A(n_4063),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4074),
.Y(n_4134)
);

OR2x2_ASAP7_75t_L g4135 ( 
.A(n_4062),
.B(n_102),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_4075),
.Y(n_4136)
);

AOI22xp33_ASAP7_75t_L g4137 ( 
.A1(n_3991),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_4137)
);

INVx2_ASAP7_75t_L g4138 ( 
.A(n_4021),
.Y(n_4138)
);

OR2x2_ASAP7_75t_L g4139 ( 
.A(n_4076),
.B(n_4091),
.Y(n_4139)
);

OAI22xp5_ASAP7_75t_L g4140 ( 
.A1(n_4038),
.A2(n_109),
.B1(n_104),
.B2(n_108),
.Y(n_4140)
);

AND2x2_ASAP7_75t_L g4141 ( 
.A(n_4093),
.B(n_108),
.Y(n_4141)
);

OR2x2_ASAP7_75t_L g4142 ( 
.A(n_4050),
.B(n_109),
.Y(n_4142)
);

AND2x2_ASAP7_75t_L g4143 ( 
.A(n_4019),
.B(n_110),
.Y(n_4143)
);

OR2x2_ASAP7_75t_L g4144 ( 
.A(n_4064),
.B(n_112),
.Y(n_4144)
);

INVx3_ASAP7_75t_L g4145 ( 
.A(n_4054),
.Y(n_4145)
);

OR2x2_ASAP7_75t_L g4146 ( 
.A(n_4098),
.B(n_113),
.Y(n_4146)
);

HB1xp67_ASAP7_75t_L g4147 ( 
.A(n_4006),
.Y(n_4147)
);

INVx2_ASAP7_75t_SL g4148 ( 
.A(n_4046),
.Y(n_4148)
);

AND2x2_ASAP7_75t_L g4149 ( 
.A(n_4042),
.B(n_4058),
.Y(n_4149)
);

AND2x2_ASAP7_75t_L g4150 ( 
.A(n_4028),
.B(n_4037),
.Y(n_4150)
);

AND2x2_ASAP7_75t_L g4151 ( 
.A(n_4028),
.B(n_113),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4085),
.B(n_4086),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_4021),
.Y(n_4153)
);

OR2x2_ASAP7_75t_L g4154 ( 
.A(n_4032),
.B(n_114),
.Y(n_4154)
);

BUFx2_ASAP7_75t_L g4155 ( 
.A(n_4046),
.Y(n_4155)
);

INVxp67_ASAP7_75t_SL g4156 ( 
.A(n_3990),
.Y(n_4156)
);

AND2x4_ASAP7_75t_L g4157 ( 
.A(n_4054),
.B(n_114),
.Y(n_4157)
);

AND2x2_ASAP7_75t_L g4158 ( 
.A(n_4029),
.B(n_116),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_4067),
.Y(n_4159)
);

INVx2_ASAP7_75t_L g4160 ( 
.A(n_4016),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4051),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_SL g4162 ( 
.A(n_4009),
.B(n_117),
.Y(n_4162)
);

NAND2xp5_ASAP7_75t_L g4163 ( 
.A(n_4079),
.B(n_117),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4015),
.Y(n_4164)
);

BUFx2_ASAP7_75t_SL g4165 ( 
.A(n_4039),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_L g4166 ( 
.A(n_4097),
.B(n_118),
.Y(n_4166)
);

AND2x4_ASAP7_75t_L g4167 ( 
.A(n_4089),
.B(n_118),
.Y(n_4167)
);

INVx1_ASAP7_75t_SL g4168 ( 
.A(n_4089),
.Y(n_4168)
);

INVx1_ASAP7_75t_L g4169 ( 
.A(n_4092),
.Y(n_4169)
);

AND2x2_ASAP7_75t_L g4170 ( 
.A(n_4030),
.B(n_119),
.Y(n_4170)
);

HB1xp67_ASAP7_75t_L g4171 ( 
.A(n_4101),
.Y(n_4171)
);

INVx1_ASAP7_75t_L g4172 ( 
.A(n_4102),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4033),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4080),
.Y(n_4174)
);

INVx1_ASAP7_75t_L g4175 ( 
.A(n_4017),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4103),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_4094),
.B(n_120),
.Y(n_4177)
);

AND2x2_ASAP7_75t_L g4178 ( 
.A(n_4030),
.B(n_121),
.Y(n_4178)
);

OR2x2_ASAP7_75t_L g4179 ( 
.A(n_4072),
.B(n_121),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4045),
.B(n_122),
.Y(n_4180)
);

AND2x2_ASAP7_75t_L g4181 ( 
.A(n_4007),
.B(n_123),
.Y(n_4181)
);

AND2x2_ASAP7_75t_L g4182 ( 
.A(n_4010),
.B(n_123),
.Y(n_4182)
);

INVx2_ASAP7_75t_L g4183 ( 
.A(n_4018),
.Y(n_4183)
);

AND2x2_ASAP7_75t_L g4184 ( 
.A(n_4012),
.B(n_3994),
.Y(n_4184)
);

NOR2x1_ASAP7_75t_L g4185 ( 
.A(n_4014),
.B(n_124),
.Y(n_4185)
);

AND2x4_ASAP7_75t_SL g4186 ( 
.A(n_4035),
.B(n_124),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4043),
.B(n_125),
.Y(n_4187)
);

NAND2xp5_ASAP7_75t_L g4188 ( 
.A(n_4047),
.B(n_125),
.Y(n_4188)
);

INVx2_ASAP7_75t_L g4189 ( 
.A(n_4083),
.Y(n_4189)
);

AND2x4_ASAP7_75t_L g4190 ( 
.A(n_4034),
.B(n_3995),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_SL g4191 ( 
.A(n_4056),
.B(n_126),
.Y(n_4191)
);

INVx1_ASAP7_75t_L g4192 ( 
.A(n_4068),
.Y(n_4192)
);

INVx2_ASAP7_75t_L g4193 ( 
.A(n_4026),
.Y(n_4193)
);

INVx2_ASAP7_75t_L g4194 ( 
.A(n_4049),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4099),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4104),
.Y(n_4196)
);

OR2x2_ASAP7_75t_L g4197 ( 
.A(n_4025),
.B(n_127),
.Y(n_4197)
);

NOR2xp33_ASAP7_75t_L g4198 ( 
.A(n_4003),
.B(n_127),
.Y(n_4198)
);

INVx1_ASAP7_75t_L g4199 ( 
.A(n_4084),
.Y(n_4199)
);

OR2x2_ASAP7_75t_L g4200 ( 
.A(n_4060),
.B(n_4048),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_4100),
.B(n_128),
.Y(n_4201)
);

OR2x2_ASAP7_75t_L g4202 ( 
.A(n_4053),
.B(n_129),
.Y(n_4202)
);

INVxp67_ASAP7_75t_SL g4203 ( 
.A(n_4013),
.Y(n_4203)
);

BUFx3_ASAP7_75t_L g4204 ( 
.A(n_4041),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4004),
.Y(n_4205)
);

HB1xp67_ASAP7_75t_L g4206 ( 
.A(n_4088),
.Y(n_4206)
);

OR2x2_ASAP7_75t_L g4207 ( 
.A(n_4059),
.B(n_129),
.Y(n_4207)
);

AND2x2_ASAP7_75t_L g4208 ( 
.A(n_4031),
.B(n_131),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_4066),
.B(n_132),
.Y(n_4209)
);

INVx2_ASAP7_75t_L g4210 ( 
.A(n_4073),
.Y(n_4210)
);

OR2x2_ASAP7_75t_L g4211 ( 
.A(n_4069),
.B(n_134),
.Y(n_4211)
);

INVx1_ASAP7_75t_L g4212 ( 
.A(n_4077),
.Y(n_4212)
);

AOI22xp33_ASAP7_75t_SL g4213 ( 
.A1(n_4090),
.A2(n_136),
.B1(n_134),
.B2(n_135),
.Y(n_4213)
);

AND2x2_ASAP7_75t_L g4214 ( 
.A(n_4087),
.B(n_136),
.Y(n_4214)
);

BUFx12f_ASAP7_75t_L g4215 ( 
.A(n_4008),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_4040),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_4022),
.B(n_138),
.Y(n_4217)
);

AND2x2_ASAP7_75t_L g4218 ( 
.A(n_4027),
.B(n_4044),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_4000),
.B(n_139),
.Y(n_4219)
);

OR2x2_ASAP7_75t_L g4220 ( 
.A(n_4002),
.B(n_141),
.Y(n_4220)
);

AND2x4_ASAP7_75t_L g4221 ( 
.A(n_4065),
.B(n_142),
.Y(n_4221)
);

INVxp67_ASAP7_75t_SL g4222 ( 
.A(n_3999),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_3999),
.B(n_142),
.Y(n_4223)
);

NOR2x1_ASAP7_75t_L g4224 ( 
.A(n_4038),
.B(n_144),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_4005),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_3999),
.B(n_144),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4023),
.Y(n_4227)
);

OR2x2_ASAP7_75t_L g4228 ( 
.A(n_4024),
.B(n_146),
.Y(n_4228)
);

AND2x2_ASAP7_75t_L g4229 ( 
.A(n_3996),
.B(n_146),
.Y(n_4229)
);

INVx2_ASAP7_75t_L g4230 ( 
.A(n_4023),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_3999),
.B(n_147),
.Y(n_4231)
);

INVx2_ASAP7_75t_L g4232 ( 
.A(n_4023),
.Y(n_4232)
);

INVx1_ASAP7_75t_L g4233 ( 
.A(n_4005),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_4005),
.Y(n_4234)
);

AND2x2_ASAP7_75t_L g4235 ( 
.A(n_3996),
.B(n_148),
.Y(n_4235)
);

AND2x2_ASAP7_75t_L g4236 ( 
.A(n_3996),
.B(n_148),
.Y(n_4236)
);

AND2x2_ASAP7_75t_L g4237 ( 
.A(n_3996),
.B(n_149),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_4023),
.Y(n_4238)
);

INVx2_ASAP7_75t_L g4239 ( 
.A(n_4023),
.Y(n_4239)
);

NOR2xp33_ASAP7_75t_L g4240 ( 
.A(n_4078),
.B(n_149),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3999),
.B(n_151),
.Y(n_4241)
);

OR2x2_ASAP7_75t_L g4242 ( 
.A(n_4024),
.B(n_152),
.Y(n_4242)
);

NOR2xp67_ASAP7_75t_L g4243 ( 
.A(n_4036),
.B(n_152),
.Y(n_4243)
);

INVx2_ASAP7_75t_SL g4244 ( 
.A(n_4046),
.Y(n_4244)
);

HB1xp67_ASAP7_75t_L g4245 ( 
.A(n_4005),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_3999),
.B(n_153),
.Y(n_4246)
);

INVx1_ASAP7_75t_L g4247 ( 
.A(n_4005),
.Y(n_4247)
);

BUFx2_ASAP7_75t_L g4248 ( 
.A(n_4078),
.Y(n_4248)
);

INVx1_ASAP7_75t_L g4249 ( 
.A(n_4005),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4005),
.Y(n_4250)
);

OR2x6_ASAP7_75t_SL g4251 ( 
.A(n_3991),
.B(n_154),
.Y(n_4251)
);

AND2x4_ASAP7_75t_L g4252 ( 
.A(n_3996),
.B(n_155),
.Y(n_4252)
);

INVx2_ASAP7_75t_L g4253 ( 
.A(n_4023),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4005),
.Y(n_4254)
);

HB1xp67_ASAP7_75t_L g4255 ( 
.A(n_4005),
.Y(n_4255)
);

AOI22xp33_ASAP7_75t_L g4256 ( 
.A1(n_4095),
.A2(n_158),
.B1(n_156),
.B2(n_157),
.Y(n_4256)
);

AND2x4_ASAP7_75t_L g4257 ( 
.A(n_3996),
.B(n_156),
.Y(n_4257)
);

AND2x2_ASAP7_75t_L g4258 ( 
.A(n_3996),
.B(n_157),
.Y(n_4258)
);

NAND2xp5_ASAP7_75t_L g4259 ( 
.A(n_3999),
.B(n_159),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_4005),
.Y(n_4260)
);

HB1xp67_ASAP7_75t_L g4261 ( 
.A(n_4005),
.Y(n_4261)
);

AND2x4_ASAP7_75t_L g4262 ( 
.A(n_3996),
.B(n_159),
.Y(n_4262)
);

BUFx3_ASAP7_75t_L g4263 ( 
.A(n_4054),
.Y(n_4263)
);

INVx1_ASAP7_75t_L g4264 ( 
.A(n_4005),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_3996),
.B(n_160),
.Y(n_4265)
);

BUFx2_ASAP7_75t_L g4266 ( 
.A(n_4078),
.Y(n_4266)
);

INVx2_ASAP7_75t_L g4267 ( 
.A(n_4023),
.Y(n_4267)
);

OAI22xp5_ASAP7_75t_L g4268 ( 
.A1(n_3991),
.A2(n_163),
.B1(n_160),
.B2(n_162),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4108),
.Y(n_4269)
);

BUFx3_ASAP7_75t_L g4270 ( 
.A(n_4248),
.Y(n_4270)
);

OAI22xp5_ASAP7_75t_L g4271 ( 
.A1(n_4224),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4222),
.B(n_164),
.Y(n_4272)
);

AO21x2_ASAP7_75t_L g4273 ( 
.A1(n_4156),
.A2(n_165),
.B(n_166),
.Y(n_4273)
);

OR2x2_ASAP7_75t_L g4274 ( 
.A(n_4107),
.B(n_167),
.Y(n_4274)
);

NOR2xp33_ASAP7_75t_L g4275 ( 
.A(n_4112),
.B(n_168),
.Y(n_4275)
);

INVx2_ASAP7_75t_L g4276 ( 
.A(n_4155),
.Y(n_4276)
);

AND2x2_ASAP7_75t_L g4277 ( 
.A(n_4266),
.B(n_169),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4174),
.B(n_169),
.Y(n_4278)
);

AOI22xp33_ASAP7_75t_L g4279 ( 
.A1(n_4190),
.A2(n_4215),
.B1(n_4204),
.B2(n_4206),
.Y(n_4279)
);

AOI22xp33_ASAP7_75t_SL g4280 ( 
.A1(n_4161),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_4280)
);

BUFx3_ASAP7_75t_L g4281 ( 
.A(n_4263),
.Y(n_4281)
);

NOR2xp33_ASAP7_75t_R g4282 ( 
.A(n_4148),
.B(n_171),
.Y(n_4282)
);

AND2x4_ASAP7_75t_L g4283 ( 
.A(n_4244),
.B(n_172),
.Y(n_4283)
);

NAND2xp5_ASAP7_75t_L g4284 ( 
.A(n_4171),
.B(n_4175),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4110),
.Y(n_4285)
);

OAI22xp5_ASAP7_75t_L g4286 ( 
.A1(n_4140),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_4286)
);

AOI221xp5_ASAP7_75t_L g4287 ( 
.A1(n_4158),
.A2(n_176),
.B1(n_173),
.B2(n_175),
.C(n_177),
.Y(n_4287)
);

OAI221xp5_ASAP7_75t_L g4288 ( 
.A1(n_4152),
.A2(n_179),
.B1(n_176),
.B2(n_178),
.C(n_181),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_4141),
.B(n_178),
.Y(n_4289)
);

INVxp67_ASAP7_75t_L g4290 ( 
.A(n_4165),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_L g4291 ( 
.A(n_4245),
.B(n_179),
.Y(n_4291)
);

AND2x2_ASAP7_75t_L g4292 ( 
.A(n_4111),
.B(n_181),
.Y(n_4292)
);

NAND2xp5_ASAP7_75t_L g4293 ( 
.A(n_4255),
.B(n_182),
.Y(n_4293)
);

OAI31xp33_ASAP7_75t_L g4294 ( 
.A1(n_4147),
.A2(n_184),
.A3(n_182),
.B(n_183),
.Y(n_4294)
);

OAI22xp5_ASAP7_75t_L g4295 ( 
.A1(n_4251),
.A2(n_4169),
.B1(n_4172),
.B2(n_4199),
.Y(n_4295)
);

INVx1_ASAP7_75t_L g4296 ( 
.A(n_4113),
.Y(n_4296)
);

OAI221xp5_ASAP7_75t_L g4297 ( 
.A1(n_4154),
.A2(n_186),
.B1(n_183),
.B2(n_185),
.C(n_187),
.Y(n_4297)
);

AOI31xp67_ASAP7_75t_L g4298 ( 
.A1(n_4138),
.A2(n_192),
.A3(n_189),
.B(n_191),
.Y(n_4298)
);

HB1xp67_ASAP7_75t_L g4299 ( 
.A(n_4261),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4115),
.Y(n_4300)
);

INVx1_ASAP7_75t_L g4301 ( 
.A(n_4117),
.Y(n_4301)
);

NAND4xp25_ASAP7_75t_SL g4302 ( 
.A(n_4177),
.B(n_193),
.C(n_191),
.D(n_192),
.Y(n_4302)
);

OAI33xp33_ASAP7_75t_L g4303 ( 
.A1(n_4176),
.A2(n_195),
.A3(n_197),
.B1(n_193),
.B2(n_194),
.B3(n_196),
.Y(n_4303)
);

INVx3_ASAP7_75t_L g4304 ( 
.A(n_4145),
.Y(n_4304)
);

NAND2xp5_ASAP7_75t_SL g4305 ( 
.A(n_4243),
.B(n_194),
.Y(n_4305)
);

OAI222xp33_ASAP7_75t_L g4306 ( 
.A1(n_4130),
.A2(n_222),
.B1(n_206),
.B2(n_233),
.C1(n_214),
.C2(n_196),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4119),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4121),
.Y(n_4308)
);

NAND4xp25_ASAP7_75t_L g4309 ( 
.A(n_4125),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_4309)
);

NOR2xp33_ASAP7_75t_R g4310 ( 
.A(n_4240),
.B(n_198),
.Y(n_4310)
);

CKINVDCx6p67_ASAP7_75t_R g4311 ( 
.A(n_4170),
.Y(n_4311)
);

OAI221xp5_ASAP7_75t_L g4312 ( 
.A1(n_4163),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.C(n_203),
.Y(n_4312)
);

AOI221xp5_ASAP7_75t_L g4313 ( 
.A1(n_4268),
.A2(n_204),
.B1(n_201),
.B2(n_202),
.C(n_206),
.Y(n_4313)
);

INVxp67_ASAP7_75t_SL g4314 ( 
.A(n_4203),
.Y(n_4314)
);

AND2x2_ASAP7_75t_L g4315 ( 
.A(n_4149),
.B(n_204),
.Y(n_4315)
);

OAI222xp33_ASAP7_75t_L g4316 ( 
.A1(n_4227),
.A2(n_235),
.B1(n_215),
.B2(n_245),
.C1(n_224),
.C2(n_207),
.Y(n_4316)
);

INVx1_ASAP7_75t_L g4317 ( 
.A(n_4122),
.Y(n_4317)
);

INVx1_ASAP7_75t_L g4318 ( 
.A(n_4126),
.Y(n_4318)
);

OR2x2_ASAP7_75t_L g4319 ( 
.A(n_4225),
.B(n_4233),
.Y(n_4319)
);

BUFx10_ASAP7_75t_L g4320 ( 
.A(n_4167),
.Y(n_4320)
);

NAND3xp33_ASAP7_75t_SL g4321 ( 
.A(n_4168),
.B(n_207),
.C(n_208),
.Y(n_4321)
);

OAI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_4197),
.A2(n_210),
.B1(n_208),
.B2(n_209),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_4234),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_4153),
.Y(n_4324)
);

INVx1_ASAP7_75t_L g4325 ( 
.A(n_4247),
.Y(n_4325)
);

OAI321xp33_ASAP7_75t_L g4326 ( 
.A1(n_4230),
.A2(n_212),
.A3(n_214),
.B1(n_210),
.B2(n_211),
.C(n_213),
.Y(n_4326)
);

AND2x2_ASAP7_75t_L g4327 ( 
.A(n_4150),
.B(n_211),
.Y(n_4327)
);

OR2x6_ASAP7_75t_L g4328 ( 
.A(n_4132),
.B(n_213),
.Y(n_4328)
);

HB1xp67_ASAP7_75t_L g4329 ( 
.A(n_4173),
.Y(n_4329)
);

AND2x2_ASAP7_75t_L g4330 ( 
.A(n_4109),
.B(n_215),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_4229),
.B(n_216),
.Y(n_4331)
);

OAI211xp5_ASAP7_75t_SL g4332 ( 
.A1(n_4192),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_4332)
);

INVx2_ASAP7_75t_L g4333 ( 
.A(n_4139),
.Y(n_4333)
);

AOI22xp5_ASAP7_75t_L g4334 ( 
.A1(n_4195),
.A2(n_219),
.B1(n_217),
.B2(n_218),
.Y(n_4334)
);

INVx2_ASAP7_75t_L g4335 ( 
.A(n_4228),
.Y(n_4335)
);

AOI22xp33_ASAP7_75t_L g4336 ( 
.A1(n_4196),
.A2(n_221),
.B1(n_219),
.B2(n_220),
.Y(n_4336)
);

OR2x2_ASAP7_75t_L g4337 ( 
.A(n_4249),
.B(n_221),
.Y(n_4337)
);

INVx2_ASAP7_75t_L g4338 ( 
.A(n_4242),
.Y(n_4338)
);

OR2x2_ASAP7_75t_L g4339 ( 
.A(n_4250),
.B(n_223),
.Y(n_4339)
);

AOI222xp33_ASAP7_75t_L g4340 ( 
.A1(n_4201),
.A2(n_254),
.B1(n_235),
.B2(n_262),
.C1(n_245),
.C2(n_223),
.Y(n_4340)
);

BUFx3_ASAP7_75t_L g4341 ( 
.A(n_4252),
.Y(n_4341)
);

OAI211xp5_ASAP7_75t_L g4342 ( 
.A1(n_4213),
.A2(n_230),
.B(n_227),
.C(n_228),
.Y(n_4342)
);

AOI222xp33_ASAP7_75t_L g4343 ( 
.A1(n_4166),
.A2(n_257),
.B1(n_239),
.B2(n_265),
.C1(n_248),
.C2(n_227),
.Y(n_4343)
);

OA21x2_ASAP7_75t_L g4344 ( 
.A1(n_4232),
.A2(n_228),
.B(n_230),
.Y(n_4344)
);

AOI21xp5_ASAP7_75t_L g4345 ( 
.A1(n_4116),
.A2(n_231),
.B(n_232),
.Y(n_4345)
);

AND2x4_ASAP7_75t_L g4346 ( 
.A(n_4164),
.B(n_232),
.Y(n_4346)
);

OAI31xp33_ASAP7_75t_SL g4347 ( 
.A1(n_4143),
.A2(n_237),
.A3(n_233),
.B(n_234),
.Y(n_4347)
);

AND2x2_ASAP7_75t_L g4348 ( 
.A(n_4235),
.B(n_234),
.Y(n_4348)
);

OR2x2_ASAP7_75t_L g4349 ( 
.A(n_4254),
.B(n_237),
.Y(n_4349)
);

INVx1_ASAP7_75t_L g4350 ( 
.A(n_4260),
.Y(n_4350)
);

HB1xp67_ASAP7_75t_L g4351 ( 
.A(n_4264),
.Y(n_4351)
);

OAI22xp5_ASAP7_75t_L g4352 ( 
.A1(n_4223),
.A2(n_242),
.B1(n_240),
.B2(n_241),
.Y(n_4352)
);

AOI22xp5_ASAP7_75t_L g4353 ( 
.A1(n_4210),
.A2(n_243),
.B1(n_241),
.B2(n_242),
.Y(n_4353)
);

AND2x2_ASAP7_75t_L g4354 ( 
.A(n_4236),
.B(n_244),
.Y(n_4354)
);

AND2x4_ASAP7_75t_L g4355 ( 
.A(n_4257),
.B(n_244),
.Y(n_4355)
);

NAND3xp33_ASAP7_75t_L g4356 ( 
.A(n_4118),
.B(n_246),
.C(n_247),
.Y(n_4356)
);

CKINVDCx20_ASAP7_75t_R g4357 ( 
.A(n_4151),
.Y(n_4357)
);

INVx3_ASAP7_75t_L g4358 ( 
.A(n_4262),
.Y(n_4358)
);

INVx2_ASAP7_75t_L g4359 ( 
.A(n_4159),
.Y(n_4359)
);

AO21x2_ASAP7_75t_L g4360 ( 
.A1(n_4226),
.A2(n_4241),
.B(n_4231),
.Y(n_4360)
);

OAI211xp5_ASAP7_75t_L g4361 ( 
.A1(n_4179),
.A2(n_249),
.B(n_246),
.C(n_248),
.Y(n_4361)
);

INVx3_ASAP7_75t_L g4362 ( 
.A(n_4157),
.Y(n_4362)
);

AND2x4_ASAP7_75t_L g4363 ( 
.A(n_4237),
.B(n_249),
.Y(n_4363)
);

CKINVDCx5p33_ASAP7_75t_R g4364 ( 
.A(n_4194),
.Y(n_4364)
);

OAI221xp5_ASAP7_75t_L g4365 ( 
.A1(n_4185),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.C(n_254),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4131),
.Y(n_4366)
);

INVx2_ASAP7_75t_L g4367 ( 
.A(n_4160),
.Y(n_4367)
);

INVxp33_ASAP7_75t_L g4368 ( 
.A(n_4184),
.Y(n_4368)
);

OAI221xp5_ASAP7_75t_L g4369 ( 
.A1(n_4120),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.C(n_255),
.Y(n_4369)
);

NAND2xp33_ASAP7_75t_R g4370 ( 
.A(n_4183),
.B(n_255),
.Y(n_4370)
);

AND2x2_ASAP7_75t_L g4371 ( 
.A(n_4258),
.B(n_4265),
.Y(n_4371)
);

INVx3_ASAP7_75t_L g4372 ( 
.A(n_4114),
.Y(n_4372)
);

OAI222xp33_ASAP7_75t_L g4373 ( 
.A1(n_4238),
.A2(n_282),
.B1(n_264),
.B2(n_291),
.C1(n_273),
.C2(n_256),
.Y(n_4373)
);

OR2x2_ASAP7_75t_L g4374 ( 
.A(n_4134),
.B(n_257),
.Y(n_4374)
);

OAI221xp5_ASAP7_75t_L g4375 ( 
.A1(n_4256),
.A2(n_260),
.B1(n_258),
.B2(n_259),
.C(n_261),
.Y(n_4375)
);

INVxp67_ASAP7_75t_L g4376 ( 
.A(n_4200),
.Y(n_4376)
);

INVx2_ASAP7_75t_L g4377 ( 
.A(n_4239),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_4133),
.Y(n_4378)
);

OA21x2_ASAP7_75t_L g4379 ( 
.A1(n_4253),
.A2(n_258),
.B(n_262),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4124),
.B(n_4127),
.Y(n_4380)
);

CKINVDCx20_ASAP7_75t_R g4381 ( 
.A(n_4246),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_L g4382 ( 
.A(n_4259),
.B(n_263),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_4136),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_4267),
.Y(n_4384)
);

OAI22xp5_ASAP7_75t_L g4385 ( 
.A1(n_4189),
.A2(n_266),
.B1(n_263),
.B2(n_265),
.Y(n_4385)
);

OAI221xp5_ASAP7_75t_SL g4386 ( 
.A1(n_4137),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.C(n_270),
.Y(n_4386)
);

OAI22xp5_ASAP7_75t_SL g4387 ( 
.A1(n_4216),
.A2(n_271),
.B1(n_267),
.B2(n_270),
.Y(n_4387)
);

NAND2xp5_ASAP7_75t_SL g4388 ( 
.A(n_4123),
.B(n_272),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_4128),
.B(n_272),
.Y(n_4389)
);

NAND2xp33_ASAP7_75t_SL g4390 ( 
.A(n_4178),
.B(n_273),
.Y(n_4390)
);

AND2x4_ASAP7_75t_L g4391 ( 
.A(n_4135),
.B(n_275),
.Y(n_4391)
);

AND2x4_ASAP7_75t_L g4392 ( 
.A(n_4142),
.B(n_276),
.Y(n_4392)
);

AOI22xp33_ASAP7_75t_SL g4393 ( 
.A1(n_4221),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_4393)
);

INVx1_ASAP7_75t_L g4394 ( 
.A(n_4144),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_4205),
.Y(n_4395)
);

INVx1_ASAP7_75t_SL g4396 ( 
.A(n_4146),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4212),
.B(n_279),
.Y(n_4397)
);

NOR2x1_ASAP7_75t_L g4398 ( 
.A(n_4162),
.B(n_279),
.Y(n_4398)
);

AOI222xp33_ASAP7_75t_L g4399 ( 
.A1(n_4198),
.A2(n_308),
.B1(n_288),
.B2(n_317),
.C1(n_297),
.C2(n_280),
.Y(n_4399)
);

AOI22xp33_ASAP7_75t_L g4400 ( 
.A1(n_4193),
.A2(n_283),
.B1(n_281),
.B2(n_282),
.Y(n_4400)
);

AND2x2_ASAP7_75t_L g4401 ( 
.A(n_4181),
.B(n_284),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4180),
.Y(n_4402)
);

HB1xp67_ASAP7_75t_L g4403 ( 
.A(n_4188),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4209),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4187),
.B(n_284),
.Y(n_4405)
);

NOR2xp33_ASAP7_75t_L g4406 ( 
.A(n_4218),
.B(n_285),
.Y(n_4406)
);

OR2x2_ASAP7_75t_L g4407 ( 
.A(n_4217),
.B(n_285),
.Y(n_4407)
);

AND2x2_ASAP7_75t_L g4408 ( 
.A(n_4208),
.B(n_286),
.Y(n_4408)
);

NOR4xp25_ASAP7_75t_L g4409 ( 
.A(n_4191),
.B(n_288),
.C(n_286),
.D(n_287),
.Y(n_4409)
);

INVx1_ASAP7_75t_L g4410 ( 
.A(n_4202),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4207),
.Y(n_4411)
);

OAI22xp5_ASAP7_75t_L g4412 ( 
.A1(n_4211),
.A2(n_291),
.B1(n_287),
.B2(n_290),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_4220),
.Y(n_4413)
);

AOI22xp33_ASAP7_75t_L g4414 ( 
.A1(n_4129),
.A2(n_294),
.B1(n_292),
.B2(n_293),
.Y(n_4414)
);

AOI22xp33_ASAP7_75t_L g4415 ( 
.A1(n_4186),
.A2(n_296),
.B1(n_292),
.B2(n_295),
.Y(n_4415)
);

INVx2_ASAP7_75t_L g4416 ( 
.A(n_4214),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4219),
.Y(n_4417)
);

AND2x2_ASAP7_75t_L g4418 ( 
.A(n_4182),
.B(n_296),
.Y(n_4418)
);

OA21x2_ASAP7_75t_L g4419 ( 
.A1(n_4130),
.A2(n_297),
.B(n_298),
.Y(n_4419)
);

AOI22xp33_ASAP7_75t_L g4420 ( 
.A1(n_4190),
.A2(n_301),
.B1(n_298),
.B2(n_299),
.Y(n_4420)
);

INVx2_ASAP7_75t_L g4421 ( 
.A(n_4155),
.Y(n_4421)
);

OAI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4222),
.A2(n_312),
.B1(n_321),
.B2(n_299),
.Y(n_4422)
);

INVx1_ASAP7_75t_L g4423 ( 
.A(n_4108),
.Y(n_4423)
);

NAND3xp33_ASAP7_75t_L g4424 ( 
.A(n_4224),
.B(n_303),
.C(n_305),
.Y(n_4424)
);

NOR2xp33_ASAP7_75t_L g4425 ( 
.A(n_4112),
.B(n_306),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_4190),
.A2(n_309),
.B1(n_306),
.B2(n_307),
.Y(n_4426)
);

INVx3_ASAP7_75t_L g4427 ( 
.A(n_4112),
.Y(n_4427)
);

INVx2_ASAP7_75t_L g4428 ( 
.A(n_4155),
.Y(n_4428)
);

INVx2_ASAP7_75t_L g4429 ( 
.A(n_4155),
.Y(n_4429)
);

AND2x2_ASAP7_75t_L g4430 ( 
.A(n_4112),
.B(n_307),
.Y(n_4430)
);

INVxp67_ASAP7_75t_SL g4431 ( 
.A(n_4224),
.Y(n_4431)
);

OAI33xp33_ASAP7_75t_L g4432 ( 
.A1(n_4175),
.A2(n_311),
.A3(n_314),
.B1(n_309),
.B2(n_310),
.B3(n_312),
.Y(n_4432)
);

AOI221xp5_ASAP7_75t_L g4433 ( 
.A1(n_4222),
.A2(n_317),
.B1(n_315),
.B2(n_316),
.C(n_318),
.Y(n_4433)
);

NAND2xp5_ASAP7_75t_L g4434 ( 
.A(n_4222),
.B(n_315),
.Y(n_4434)
);

AND2x2_ASAP7_75t_L g4435 ( 
.A(n_4112),
.B(n_316),
.Y(n_4435)
);

AND2x6_ASAP7_75t_SL g4436 ( 
.A(n_4240),
.B(n_318),
.Y(n_4436)
);

AOI22xp33_ASAP7_75t_L g4437 ( 
.A1(n_4190),
.A2(n_322),
.B1(n_319),
.B2(n_320),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4108),
.Y(n_4438)
);

OAI211xp5_ASAP7_75t_L g4439 ( 
.A1(n_4224),
.A2(n_324),
.B(n_322),
.C(n_323),
.Y(n_4439)
);

NOR2x1_ASAP7_75t_SL g4440 ( 
.A(n_4174),
.B(n_325),
.Y(n_4440)
);

OAI31xp33_ASAP7_75t_L g4441 ( 
.A1(n_4140),
.A2(n_328),
.A3(n_326),
.B(n_327),
.Y(n_4441)
);

A2O1A1Ixp33_ASAP7_75t_L g4442 ( 
.A1(n_4224),
.A2(n_329),
.B(n_327),
.C(n_328),
.Y(n_4442)
);

AND2x2_ASAP7_75t_L g4443 ( 
.A(n_4112),
.B(n_329),
.Y(n_4443)
);

INVx2_ASAP7_75t_SL g4444 ( 
.A(n_4112),
.Y(n_4444)
);

INVx4_ASAP7_75t_L g4445 ( 
.A(n_4112),
.Y(n_4445)
);

NOR2x2_ASAP7_75t_L g4446 ( 
.A(n_4183),
.B(n_331),
.Y(n_4446)
);

AOI22xp33_ASAP7_75t_L g4447 ( 
.A1(n_4190),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_4447)
);

NAND2xp33_ASAP7_75t_SL g4448 ( 
.A(n_4248),
.B(n_333),
.Y(n_4448)
);

AO21x2_ASAP7_75t_L g4449 ( 
.A1(n_4156),
.A2(n_334),
.B(n_335),
.Y(n_4449)
);

AO21x2_ASAP7_75t_L g4450 ( 
.A1(n_4156),
.A2(n_335),
.B(n_336),
.Y(n_4450)
);

OA21x2_ASAP7_75t_L g4451 ( 
.A1(n_4130),
.A2(n_337),
.B(n_338),
.Y(n_4451)
);

AOI22xp33_ASAP7_75t_SL g4452 ( 
.A1(n_4156),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.Y(n_4452)
);

OAI221xp5_ASAP7_75t_L g4453 ( 
.A1(n_4224),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.C(n_343),
.Y(n_4453)
);

AOI33xp33_ASAP7_75t_L g4454 ( 
.A1(n_4192),
.A2(n_343),
.A3(n_345),
.B1(n_340),
.B2(n_342),
.B3(n_344),
.Y(n_4454)
);

AND2x4_ASAP7_75t_SL g4455 ( 
.A(n_4150),
.B(n_344),
.Y(n_4455)
);

INVx2_ASAP7_75t_L g4456 ( 
.A(n_4155),
.Y(n_4456)
);

BUFx3_ASAP7_75t_L g4457 ( 
.A(n_4248),
.Y(n_4457)
);

INVx1_ASAP7_75t_L g4458 ( 
.A(n_4108),
.Y(n_4458)
);

INVx1_ASAP7_75t_L g4459 ( 
.A(n_4108),
.Y(n_4459)
);

AOI322xp5_ASAP7_75t_L g4460 ( 
.A1(n_4156),
.A2(n_351),
.A3(n_350),
.B1(n_348),
.B2(n_346),
.C1(n_347),
.C2(n_349),
.Y(n_4460)
);

OAI321xp33_ASAP7_75t_L g4461 ( 
.A1(n_4156),
.A2(n_349),
.A3(n_351),
.B1(n_347),
.B2(n_348),
.C(n_350),
.Y(n_4461)
);

NAND2xp5_ASAP7_75t_L g4462 ( 
.A(n_4222),
.B(n_352),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_4155),
.Y(n_4463)
);

AOI22xp33_ASAP7_75t_L g4464 ( 
.A1(n_4402),
.A2(n_355),
.B1(n_352),
.B2(n_353),
.Y(n_4464)
);

AND2x2_ASAP7_75t_L g4465 ( 
.A(n_4427),
.B(n_353),
.Y(n_4465)
);

AO21x2_ASAP7_75t_L g4466 ( 
.A1(n_4284),
.A2(n_356),
.B(n_357),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4270),
.Y(n_4467)
);

AOI22xp33_ASAP7_75t_L g4468 ( 
.A1(n_4404),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.Y(n_4468)
);

NAND2xp5_ASAP7_75t_SL g4469 ( 
.A(n_4290),
.B(n_360),
.Y(n_4469)
);

OR2x2_ASAP7_75t_L g4470 ( 
.A(n_4396),
.B(n_360),
.Y(n_4470)
);

INVx1_ASAP7_75t_L g4471 ( 
.A(n_4299),
.Y(n_4471)
);

NOR3xp33_ASAP7_75t_L g4472 ( 
.A(n_4461),
.B(n_361),
.C(n_362),
.Y(n_4472)
);

OAI21xp5_ASAP7_75t_L g4473 ( 
.A1(n_4431),
.A2(n_361),
.B(n_362),
.Y(n_4473)
);

NOR3xp33_ASAP7_75t_L g4474 ( 
.A(n_4445),
.B(n_4439),
.C(n_4314),
.Y(n_4474)
);

AND2x2_ASAP7_75t_L g4475 ( 
.A(n_4444),
.B(n_363),
.Y(n_4475)
);

NAND3xp33_ASAP7_75t_L g4476 ( 
.A(n_4347),
.B(n_363),
.C(n_364),
.Y(n_4476)
);

NOR2x1_ASAP7_75t_SL g4477 ( 
.A(n_4371),
.B(n_4328),
.Y(n_4477)
);

AOI22xp33_ASAP7_75t_L g4478 ( 
.A1(n_4403),
.A2(n_369),
.B1(n_364),
.B2(n_365),
.Y(n_4478)
);

NAND4xp75_ASAP7_75t_L g4479 ( 
.A(n_4398),
.B(n_373),
.C(n_370),
.D(n_371),
.Y(n_4479)
);

AND2x2_ASAP7_75t_L g4480 ( 
.A(n_4380),
.B(n_370),
.Y(n_4480)
);

NOR3xp33_ASAP7_75t_L g4481 ( 
.A(n_4432),
.B(n_371),
.C(n_373),
.Y(n_4481)
);

OR2x2_ASAP7_75t_L g4482 ( 
.A(n_4394),
.B(n_374),
.Y(n_4482)
);

INVx1_ASAP7_75t_L g4483 ( 
.A(n_4351),
.Y(n_4483)
);

NAND4xp75_ASAP7_75t_L g4484 ( 
.A(n_4294),
.B(n_377),
.C(n_374),
.D(n_376),
.Y(n_4484)
);

OAI211xp5_ASAP7_75t_L g4485 ( 
.A1(n_4448),
.A2(n_380),
.B(n_378),
.C(n_379),
.Y(n_4485)
);

AND2x2_ASAP7_75t_L g4486 ( 
.A(n_4457),
.B(n_378),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_4357),
.Y(n_4487)
);

INVx1_ASAP7_75t_L g4488 ( 
.A(n_4395),
.Y(n_4488)
);

AOI22xp33_ASAP7_75t_SL g4489 ( 
.A1(n_4295),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_4489)
);

AND2x2_ASAP7_75t_L g4490 ( 
.A(n_4311),
.B(n_381),
.Y(n_4490)
);

INVx2_ASAP7_75t_L g4491 ( 
.A(n_4446),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4292),
.B(n_382),
.Y(n_4492)
);

AO21x2_ASAP7_75t_L g4493 ( 
.A1(n_4272),
.A2(n_382),
.B(n_384),
.Y(n_4493)
);

AOI22xp33_ASAP7_75t_L g4494 ( 
.A1(n_4410),
.A2(n_388),
.B1(n_385),
.B2(n_387),
.Y(n_4494)
);

OR2x2_ASAP7_75t_L g4495 ( 
.A(n_4319),
.B(n_385),
.Y(n_4495)
);

OR2x2_ASAP7_75t_L g4496 ( 
.A(n_4276),
.B(n_387),
.Y(n_4496)
);

AO21x2_ASAP7_75t_L g4497 ( 
.A1(n_4434),
.A2(n_389),
.B(n_390),
.Y(n_4497)
);

NOR2xp33_ASAP7_75t_L g4498 ( 
.A(n_4281),
.B(n_390),
.Y(n_4498)
);

AND2x2_ASAP7_75t_L g4499 ( 
.A(n_4372),
.B(n_391),
.Y(n_4499)
);

OR2x2_ASAP7_75t_L g4500 ( 
.A(n_4421),
.B(n_4428),
.Y(n_4500)
);

AND2x2_ASAP7_75t_L g4501 ( 
.A(n_4429),
.B(n_391),
.Y(n_4501)
);

AO21x2_ASAP7_75t_L g4502 ( 
.A1(n_4462),
.A2(n_392),
.B(n_393),
.Y(n_4502)
);

INVx1_ASAP7_75t_L g4503 ( 
.A(n_4397),
.Y(n_4503)
);

AOI221xp5_ASAP7_75t_L g4504 ( 
.A1(n_4376),
.A2(n_394),
.B1(n_392),
.B2(n_393),
.C(n_395),
.Y(n_4504)
);

AND2x2_ASAP7_75t_L g4505 ( 
.A(n_4456),
.B(n_394),
.Y(n_4505)
);

NAND4xp75_ASAP7_75t_L g4506 ( 
.A(n_4287),
.B(n_397),
.C(n_395),
.D(n_396),
.Y(n_4506)
);

NOR2xp33_ASAP7_75t_L g4507 ( 
.A(n_4381),
.B(n_4362),
.Y(n_4507)
);

NAND2xp5_ASAP7_75t_L g4508 ( 
.A(n_4360),
.B(n_396),
.Y(n_4508)
);

NAND4xp75_ASAP7_75t_L g4509 ( 
.A(n_4441),
.B(n_399),
.C(n_397),
.D(n_398),
.Y(n_4509)
);

AND2x4_ASAP7_75t_L g4510 ( 
.A(n_4341),
.B(n_4358),
.Y(n_4510)
);

AO22x2_ASAP7_75t_L g4511 ( 
.A1(n_4411),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.Y(n_4511)
);

NAND3xp33_ASAP7_75t_L g4512 ( 
.A(n_4442),
.B(n_400),
.C(n_402),
.Y(n_4512)
);

NAND3xp33_ASAP7_75t_L g4513 ( 
.A(n_4424),
.B(n_403),
.C(n_404),
.Y(n_4513)
);

AND2x2_ASAP7_75t_L g4514 ( 
.A(n_4463),
.B(n_405),
.Y(n_4514)
);

NAND4xp75_ASAP7_75t_L g4515 ( 
.A(n_4430),
.B(n_4435),
.C(n_4443),
.D(n_4345),
.Y(n_4515)
);

CKINVDCx5p33_ASAP7_75t_R g4516 ( 
.A(n_4310),
.Y(n_4516)
);

AOI22xp5_ASAP7_75t_L g4517 ( 
.A1(n_4370),
.A2(n_407),
.B1(n_405),
.B2(n_406),
.Y(n_4517)
);

OR2x2_ASAP7_75t_L g4518 ( 
.A(n_4366),
.B(n_406),
.Y(n_4518)
);

NAND3xp33_ASAP7_75t_L g4519 ( 
.A(n_4343),
.B(n_408),
.C(n_409),
.Y(n_4519)
);

NAND2xp5_ASAP7_75t_L g4520 ( 
.A(n_4273),
.B(n_4449),
.Y(n_4520)
);

NAND3xp33_ASAP7_75t_L g4521 ( 
.A(n_4271),
.B(n_408),
.C(n_409),
.Y(n_4521)
);

AND2x2_ASAP7_75t_L g4522 ( 
.A(n_4304),
.B(n_410),
.Y(n_4522)
);

OR2x2_ASAP7_75t_L g4523 ( 
.A(n_4378),
.B(n_410),
.Y(n_4523)
);

OAI211xp5_ASAP7_75t_SL g4524 ( 
.A1(n_4460),
.A2(n_413),
.B(n_411),
.C(n_412),
.Y(n_4524)
);

AND2x2_ASAP7_75t_L g4525 ( 
.A(n_4320),
.B(n_411),
.Y(n_4525)
);

AND2x2_ASAP7_75t_L g4526 ( 
.A(n_4440),
.B(n_413),
.Y(n_4526)
);

INVx1_ASAP7_75t_L g4527 ( 
.A(n_4329),
.Y(n_4527)
);

AND2x2_ASAP7_75t_L g4528 ( 
.A(n_4277),
.B(n_415),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4269),
.Y(n_4529)
);

AND2x2_ASAP7_75t_L g4530 ( 
.A(n_4278),
.B(n_416),
.Y(n_4530)
);

NOR3xp33_ASAP7_75t_SL g4531 ( 
.A(n_4275),
.B(n_416),
.C(n_417),
.Y(n_4531)
);

AND2x2_ASAP7_75t_L g4532 ( 
.A(n_4283),
.B(n_417),
.Y(n_4532)
);

INVx2_ASAP7_75t_L g4533 ( 
.A(n_4298),
.Y(n_4533)
);

AOI22xp33_ASAP7_75t_L g4534 ( 
.A1(n_4413),
.A2(n_420),
.B1(n_418),
.B2(n_419),
.Y(n_4534)
);

AO21x2_ASAP7_75t_L g4535 ( 
.A1(n_4291),
.A2(n_418),
.B(n_419),
.Y(n_4535)
);

AOI22xp5_ASAP7_75t_SL g4536 ( 
.A1(n_4322),
.A2(n_423),
.B1(n_420),
.B2(n_421),
.Y(n_4536)
);

NOR3xp33_ASAP7_75t_L g4537 ( 
.A(n_4303),
.B(n_423),
.C(n_424),
.Y(n_4537)
);

AND2x4_ASAP7_75t_L g4538 ( 
.A(n_4455),
.B(n_424),
.Y(n_4538)
);

OR2x2_ASAP7_75t_L g4539 ( 
.A(n_4323),
.B(n_425),
.Y(n_4539)
);

AND2x2_ASAP7_75t_L g4540 ( 
.A(n_4315),
.B(n_425),
.Y(n_4540)
);

AOI22xp5_ASAP7_75t_L g4541 ( 
.A1(n_4450),
.A2(n_428),
.B1(n_426),
.B2(n_427),
.Y(n_4541)
);

NOR3xp33_ASAP7_75t_L g4542 ( 
.A(n_4326),
.B(n_426),
.C(n_427),
.Y(n_4542)
);

NAND4xp75_ASAP7_75t_L g4543 ( 
.A(n_4433),
.B(n_430),
.C(n_428),
.D(n_429),
.Y(n_4543)
);

AND2x2_ASAP7_75t_L g4544 ( 
.A(n_4327),
.B(n_430),
.Y(n_4544)
);

INVx1_ASAP7_75t_L g4545 ( 
.A(n_4285),
.Y(n_4545)
);

INVx1_ASAP7_75t_L g4546 ( 
.A(n_4296),
.Y(n_4546)
);

NAND3xp33_ASAP7_75t_SL g4547 ( 
.A(n_4452),
.B(n_431),
.C(n_432),
.Y(n_4547)
);

AOI21xp33_ASAP7_75t_L g4548 ( 
.A1(n_4368),
.A2(n_433),
.B(n_432),
.Y(n_4548)
);

NAND3xp33_ASAP7_75t_L g4549 ( 
.A(n_4340),
.B(n_431),
.C(n_433),
.Y(n_4549)
);

AND2x2_ASAP7_75t_L g4550 ( 
.A(n_4425),
.B(n_434),
.Y(n_4550)
);

NAND2xp5_ASAP7_75t_L g4551 ( 
.A(n_4422),
.B(n_434),
.Y(n_4551)
);

INVxp67_ASAP7_75t_SL g4552 ( 
.A(n_4406),
.Y(n_4552)
);

BUFx3_ASAP7_75t_L g4553 ( 
.A(n_4363),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_SL g4554 ( 
.A(n_4391),
.B(n_435),
.Y(n_4554)
);

AND2x2_ASAP7_75t_L g4555 ( 
.A(n_4325),
.B(n_436),
.Y(n_4555)
);

NOR2xp33_ASAP7_75t_L g4556 ( 
.A(n_4436),
.B(n_436),
.Y(n_4556)
);

OA211x2_ASAP7_75t_L g4557 ( 
.A1(n_4302),
.A2(n_439),
.B(n_437),
.C(n_438),
.Y(n_4557)
);

NAND4xp75_ASAP7_75t_L g4558 ( 
.A(n_4344),
.B(n_439),
.C(n_437),
.D(n_438),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4379),
.Y(n_4559)
);

AND2x2_ASAP7_75t_L g4560 ( 
.A(n_4350),
.B(n_440),
.Y(n_4560)
);

AND2x4_ASAP7_75t_L g4561 ( 
.A(n_4328),
.B(n_4355),
.Y(n_4561)
);

INVx1_ASAP7_75t_L g4562 ( 
.A(n_4300),
.Y(n_4562)
);

AOI22xp5_ASAP7_75t_L g4563 ( 
.A1(n_4417),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_4563)
);

AND2x2_ASAP7_75t_L g4564 ( 
.A(n_4330),
.B(n_443),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_4301),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_SL g4566 ( 
.A(n_4274),
.B(n_4337),
.Y(n_4566)
);

HB1xp67_ASAP7_75t_L g4567 ( 
.A(n_4339),
.Y(n_4567)
);

OR2x2_ASAP7_75t_L g4568 ( 
.A(n_4349),
.B(n_444),
.Y(n_4568)
);

NOR2xp33_ASAP7_75t_L g4569 ( 
.A(n_4392),
.B(n_444),
.Y(n_4569)
);

NAND3xp33_ASAP7_75t_L g4570 ( 
.A(n_4399),
.B(n_445),
.C(n_446),
.Y(n_4570)
);

AND2x2_ASAP7_75t_L g4571 ( 
.A(n_4331),
.B(n_445),
.Y(n_4571)
);

NAND2xp5_ASAP7_75t_L g4572 ( 
.A(n_4359),
.B(n_447),
.Y(n_4572)
);

INVx1_ASAP7_75t_SL g4573 ( 
.A(n_4282),
.Y(n_4573)
);

AOI22xp33_ASAP7_75t_L g4574 ( 
.A1(n_4377),
.A2(n_449),
.B1(n_447),
.B2(n_448),
.Y(n_4574)
);

AO21x2_ASAP7_75t_L g4575 ( 
.A1(n_4293),
.A2(n_448),
.B(n_450),
.Y(n_4575)
);

NAND3xp33_ASAP7_75t_L g4576 ( 
.A(n_4453),
.B(n_450),
.C(n_451),
.Y(n_4576)
);

OR2x2_ASAP7_75t_L g4577 ( 
.A(n_4383),
.B(n_452),
.Y(n_4577)
);

NOR3xp33_ASAP7_75t_L g4578 ( 
.A(n_4361),
.B(n_452),
.C(n_453),
.Y(n_4578)
);

OR2x2_ASAP7_75t_L g4579 ( 
.A(n_4307),
.B(n_454),
.Y(n_4579)
);

NAND3xp33_ASAP7_75t_L g4580 ( 
.A(n_4280),
.B(n_454),
.C(n_456),
.Y(n_4580)
);

NOR3xp33_ASAP7_75t_L g4581 ( 
.A(n_4342),
.B(n_458),
.C(n_460),
.Y(n_4581)
);

INVx1_ASAP7_75t_L g4582 ( 
.A(n_4308),
.Y(n_4582)
);

NOR3xp33_ASAP7_75t_L g4583 ( 
.A(n_4288),
.B(n_461),
.C(n_462),
.Y(n_4583)
);

NOR3xp33_ASAP7_75t_L g4584 ( 
.A(n_4306),
.B(n_463),
.C(n_464),
.Y(n_4584)
);

OR2x2_ASAP7_75t_L g4585 ( 
.A(n_4317),
.B(n_463),
.Y(n_4585)
);

NAND2xp5_ASAP7_75t_L g4586 ( 
.A(n_4408),
.B(n_465),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_4348),
.B(n_467),
.Y(n_4587)
);

NAND2xp5_ASAP7_75t_L g4588 ( 
.A(n_4401),
.B(n_468),
.Y(n_4588)
);

INVx1_ASAP7_75t_L g4589 ( 
.A(n_4318),
.Y(n_4589)
);

OAI211xp5_ASAP7_75t_L g4590 ( 
.A1(n_4409),
.A2(n_470),
.B(n_468),
.C(n_469),
.Y(n_4590)
);

NAND2xp5_ASAP7_75t_L g4591 ( 
.A(n_4374),
.B(n_469),
.Y(n_4591)
);

NAND4xp75_ASAP7_75t_L g4592 ( 
.A(n_4419),
.B(n_4451),
.C(n_4305),
.D(n_4384),
.Y(n_4592)
);

AND2x2_ASAP7_75t_L g4593 ( 
.A(n_4354),
.B(n_470),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_4423),
.Y(n_4594)
);

AND2x2_ASAP7_75t_L g4595 ( 
.A(n_4346),
.B(n_472),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_4334),
.B(n_472),
.Y(n_4596)
);

NOR3xp33_ASAP7_75t_L g4597 ( 
.A(n_4316),
.B(n_4373),
.C(n_4365),
.Y(n_4597)
);

NOR2xp33_ASAP7_75t_L g4598 ( 
.A(n_4309),
.B(n_473),
.Y(n_4598)
);

AND2x2_ASAP7_75t_L g4599 ( 
.A(n_4438),
.B(n_473),
.Y(n_4599)
);

NAND2xp5_ASAP7_75t_L g4600 ( 
.A(n_4335),
.B(n_474),
.Y(n_4600)
);

NAND2xp5_ASAP7_75t_L g4601 ( 
.A(n_4338),
.B(n_474),
.Y(n_4601)
);

HB1xp67_ASAP7_75t_L g4602 ( 
.A(n_4487),
.Y(n_4602)
);

AND2x2_ASAP7_75t_L g4603 ( 
.A(n_4477),
.B(n_4510),
.Y(n_4603)
);

INVx1_ASAP7_75t_L g4604 ( 
.A(n_4567),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4467),
.B(n_4458),
.Y(n_4605)
);

AND2x2_ASAP7_75t_L g4606 ( 
.A(n_4474),
.B(n_4459),
.Y(n_4606)
);

AND2x2_ASAP7_75t_L g4607 ( 
.A(n_4490),
.B(n_4289),
.Y(n_4607)
);

INVx1_ASAP7_75t_L g4608 ( 
.A(n_4470),
.Y(n_4608)
);

INVx2_ASAP7_75t_L g4609 ( 
.A(n_4553),
.Y(n_4609)
);

INVx1_ASAP7_75t_L g4610 ( 
.A(n_4471),
.Y(n_4610)
);

INVx1_ASAP7_75t_L g4611 ( 
.A(n_4511),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4511),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4480),
.Y(n_4613)
);

OR2x2_ASAP7_75t_L g4614 ( 
.A(n_4495),
.B(n_4382),
.Y(n_4614)
);

OR2x2_ASAP7_75t_L g4615 ( 
.A(n_4500),
.B(n_4333),
.Y(n_4615)
);

AND2x2_ASAP7_75t_L g4616 ( 
.A(n_4573),
.B(n_4416),
.Y(n_4616)
);

INVx2_ASAP7_75t_L g4617 ( 
.A(n_4491),
.Y(n_4617)
);

INVx1_ASAP7_75t_L g4618 ( 
.A(n_4482),
.Y(n_4618)
);

INVx1_ASAP7_75t_L g4619 ( 
.A(n_4508),
.Y(n_4619)
);

HB1xp67_ASAP7_75t_L g4620 ( 
.A(n_4466),
.Y(n_4620)
);

OAI33xp33_ASAP7_75t_L g4621 ( 
.A1(n_4483),
.A2(n_4352),
.A3(n_4387),
.B1(n_4385),
.B2(n_4412),
.B3(n_4286),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_4568),
.Y(n_4622)
);

INVx1_ASAP7_75t_L g4623 ( 
.A(n_4600),
.Y(n_4623)
);

AND2x2_ASAP7_75t_L g4624 ( 
.A(n_4507),
.B(n_4388),
.Y(n_4624)
);

HB1xp67_ASAP7_75t_L g4625 ( 
.A(n_4496),
.Y(n_4625)
);

INVx1_ASAP7_75t_L g4626 ( 
.A(n_4601),
.Y(n_4626)
);

INVx6_ASAP7_75t_L g4627 ( 
.A(n_4538),
.Y(n_4627)
);

INVx1_ASAP7_75t_L g4628 ( 
.A(n_4503),
.Y(n_4628)
);

INVx2_ASAP7_75t_L g4629 ( 
.A(n_4561),
.Y(n_4629)
);

INVx1_ASAP7_75t_L g4630 ( 
.A(n_4579),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4585),
.Y(n_4631)
);

OAI31xp33_ASAP7_75t_L g4632 ( 
.A1(n_4520),
.A2(n_4390),
.A3(n_4297),
.B(n_4312),
.Y(n_4632)
);

BUFx2_ASAP7_75t_L g4633 ( 
.A(n_4473),
.Y(n_4633)
);

AND2x2_ASAP7_75t_L g4634 ( 
.A(n_4465),
.B(n_4389),
.Y(n_4634)
);

INVx3_ASAP7_75t_L g4635 ( 
.A(n_4525),
.Y(n_4635)
);

INVx1_ASAP7_75t_L g4636 ( 
.A(n_4527),
.Y(n_4636)
);

NAND2xp5_ASAP7_75t_L g4637 ( 
.A(n_4533),
.B(n_4353),
.Y(n_4637)
);

INVxp67_ASAP7_75t_SL g4638 ( 
.A(n_4556),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4597),
.B(n_4420),
.Y(n_4639)
);

BUFx3_ASAP7_75t_L g4640 ( 
.A(n_4544),
.Y(n_4640)
);

NAND2xp5_ASAP7_75t_L g4641 ( 
.A(n_4584),
.B(n_4472),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4539),
.Y(n_4642)
);

INVx1_ASAP7_75t_L g4643 ( 
.A(n_4577),
.Y(n_4643)
);

BUFx4f_ASAP7_75t_SL g4644 ( 
.A(n_4475),
.Y(n_4644)
);

INVx2_ASAP7_75t_L g4645 ( 
.A(n_4516),
.Y(n_4645)
);

BUFx12f_ASAP7_75t_L g4646 ( 
.A(n_4486),
.Y(n_4646)
);

OAI31xp33_ASAP7_75t_L g4647 ( 
.A1(n_4590),
.A2(n_4476),
.A3(n_4519),
.B(n_4570),
.Y(n_4647)
);

INVx2_ASAP7_75t_L g4648 ( 
.A(n_4599),
.Y(n_4648)
);

OR2x2_ASAP7_75t_L g4649 ( 
.A(n_4518),
.B(n_4405),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4542),
.B(n_4426),
.Y(n_4650)
);

INVx1_ASAP7_75t_L g4651 ( 
.A(n_4488),
.Y(n_4651)
);

AND2x2_ASAP7_75t_L g4652 ( 
.A(n_4501),
.B(n_4418),
.Y(n_4652)
);

INVx1_ASAP7_75t_L g4653 ( 
.A(n_4529),
.Y(n_4653)
);

NAND2xp5_ASAP7_75t_L g4654 ( 
.A(n_4493),
.B(n_4497),
.Y(n_4654)
);

INVx2_ASAP7_75t_L g4655 ( 
.A(n_4505),
.Y(n_4655)
);

INVx2_ASAP7_75t_L g4656 ( 
.A(n_4514),
.Y(n_4656)
);

INVx2_ASAP7_75t_L g4657 ( 
.A(n_4555),
.Y(n_4657)
);

OAI21xp5_ASAP7_75t_L g4658 ( 
.A1(n_4489),
.A2(n_4321),
.B(n_4356),
.Y(n_4658)
);

AOI21xp33_ASAP7_75t_L g4659 ( 
.A1(n_4552),
.A2(n_4324),
.B(n_4367),
.Y(n_4659)
);

INVx1_ASAP7_75t_SL g4660 ( 
.A(n_4528),
.Y(n_4660)
);

INVx2_ASAP7_75t_L g4661 ( 
.A(n_4560),
.Y(n_4661)
);

INVx2_ASAP7_75t_L g4662 ( 
.A(n_4523),
.Y(n_4662)
);

INVx4_ASAP7_75t_L g4663 ( 
.A(n_4522),
.Y(n_4663)
);

BUFx3_ASAP7_75t_L g4664 ( 
.A(n_4564),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4499),
.Y(n_4665)
);

XOR2xp5_ASAP7_75t_L g4666 ( 
.A(n_4515),
.B(n_4364),
.Y(n_4666)
);

OR2x2_ASAP7_75t_L g4667 ( 
.A(n_4566),
.B(n_4407),
.Y(n_4667)
);

OR2x2_ASAP7_75t_L g4668 ( 
.A(n_4572),
.B(n_4279),
.Y(n_4668)
);

AND2x2_ASAP7_75t_L g4669 ( 
.A(n_4469),
.B(n_4498),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4502),
.B(n_4437),
.Y(n_4670)
);

AND2x4_ASAP7_75t_L g4671 ( 
.A(n_4571),
.B(n_4447),
.Y(n_4671)
);

OR2x2_ASAP7_75t_L g4672 ( 
.A(n_4545),
.B(n_4336),
.Y(n_4672)
);

NOR2xp33_ASAP7_75t_L g4673 ( 
.A(n_4586),
.B(n_4332),
.Y(n_4673)
);

INVx2_ASAP7_75t_L g4674 ( 
.A(n_4558),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4546),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_4526),
.B(n_4454),
.Y(n_4676)
);

OAI32xp33_ASAP7_75t_L g4677 ( 
.A1(n_4481),
.A2(n_4375),
.A3(n_4369),
.B1(n_4414),
.B2(n_4400),
.Y(n_4677)
);

AND2x2_ASAP7_75t_L g4678 ( 
.A(n_4540),
.B(n_4393),
.Y(n_4678)
);

INVx1_ASAP7_75t_SL g4679 ( 
.A(n_4587),
.Y(n_4679)
);

INVx2_ASAP7_75t_L g4680 ( 
.A(n_4593),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4535),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4562),
.Y(n_4682)
);

AOI221xp5_ASAP7_75t_L g4683 ( 
.A1(n_4537),
.A2(n_4313),
.B1(n_4386),
.B2(n_4415),
.C(n_477),
.Y(n_4683)
);

AND2x2_ASAP7_75t_L g4684 ( 
.A(n_4532),
.B(n_475),
.Y(n_4684)
);

BUFx3_ASAP7_75t_L g4685 ( 
.A(n_4530),
.Y(n_4685)
);

AND2x2_ASAP7_75t_SL g4686 ( 
.A(n_4583),
.B(n_475),
.Y(n_4686)
);

AOI221xp5_ASAP7_75t_L g4687 ( 
.A1(n_4524),
.A2(n_478),
.B1(n_476),
.B2(n_477),
.C(n_479),
.Y(n_4687)
);

NAND4xp25_ASAP7_75t_L g4688 ( 
.A(n_4565),
.B(n_479),
.C(n_476),
.D(n_478),
.Y(n_4688)
);

INVx4_ASAP7_75t_L g4689 ( 
.A(n_4595),
.Y(n_4689)
);

BUFx3_ASAP7_75t_L g4690 ( 
.A(n_4550),
.Y(n_4690)
);

INVx2_ASAP7_75t_L g4691 ( 
.A(n_4575),
.Y(n_4691)
);

AND2x2_ASAP7_75t_SL g4692 ( 
.A(n_4578),
.B(n_480),
.Y(n_4692)
);

INVx2_ASAP7_75t_L g4693 ( 
.A(n_4559),
.Y(n_4693)
);

AND2x2_ASAP7_75t_L g4694 ( 
.A(n_4582),
.B(n_481),
.Y(n_4694)
);

AND2x2_ASAP7_75t_SL g4695 ( 
.A(n_4581),
.B(n_481),
.Y(n_4695)
);

AND3x1_ASAP7_75t_SL g4696 ( 
.A(n_4613),
.B(n_4594),
.C(n_4589),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4602),
.Y(n_4697)
);

CKINVDCx16_ASAP7_75t_R g4698 ( 
.A(n_4646),
.Y(n_4698)
);

NOR2xp33_ASAP7_75t_L g4699 ( 
.A(n_4644),
.B(n_4554),
.Y(n_4699)
);

OAI33xp33_ASAP7_75t_L g4700 ( 
.A1(n_4639),
.A2(n_4576),
.A3(n_4549),
.B1(n_4551),
.B2(n_4596),
.B3(n_4521),
.Y(n_4700)
);

INVx3_ASAP7_75t_L g4701 ( 
.A(n_4689),
.Y(n_4701)
);

OAI21xp33_ASAP7_75t_L g4702 ( 
.A1(n_4629),
.A2(n_4598),
.B(n_4563),
.Y(n_4702)
);

AOI22xp33_ASAP7_75t_SL g4703 ( 
.A1(n_4620),
.A2(n_4536),
.B1(n_4580),
.B2(n_4512),
.Y(n_4703)
);

OR2x2_ASAP7_75t_L g4704 ( 
.A(n_4679),
.B(n_4492),
.Y(n_4704)
);

OAI32xp33_ASAP7_75t_L g4705 ( 
.A1(n_4641),
.A2(n_4513),
.A3(n_4548),
.B1(n_4591),
.B2(n_4588),
.Y(n_4705)
);

NOR2x1p5_ASAP7_75t_SL g4706 ( 
.A(n_4617),
.B(n_4592),
.Y(n_4706)
);

INVx1_ASAP7_75t_L g4707 ( 
.A(n_4625),
.Y(n_4707)
);

OAI32xp33_ASAP7_75t_L g4708 ( 
.A1(n_4637),
.A2(n_4478),
.A3(n_4494),
.B1(n_4534),
.B2(n_4468),
.Y(n_4708)
);

INVx3_ASAP7_75t_L g4709 ( 
.A(n_4663),
.Y(n_4709)
);

NAND2xp5_ASAP7_75t_L g4710 ( 
.A(n_4660),
.B(n_4541),
.Y(n_4710)
);

AND2x2_ASAP7_75t_L g4711 ( 
.A(n_4603),
.B(n_4531),
.Y(n_4711)
);

NAND4xp75_ASAP7_75t_L g4712 ( 
.A(n_4647),
.B(n_4557),
.C(n_4517),
.D(n_4504),
.Y(n_4712)
);

OR2x2_ASAP7_75t_L g4713 ( 
.A(n_4604),
.B(n_4615),
.Y(n_4713)
);

INVx1_ASAP7_75t_L g4714 ( 
.A(n_4667),
.Y(n_4714)
);

AND2x2_ASAP7_75t_L g4715 ( 
.A(n_4609),
.B(n_4569),
.Y(n_4715)
);

AND2x4_ASAP7_75t_SL g4716 ( 
.A(n_4645),
.B(n_4624),
.Y(n_4716)
);

INVx1_ASAP7_75t_L g4717 ( 
.A(n_4622),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4685),
.B(n_4485),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_SL g4719 ( 
.A(n_4690),
.B(n_4464),
.Y(n_4719)
);

AOI22xp5_ASAP7_75t_L g4720 ( 
.A1(n_4692),
.A2(n_4547),
.B1(n_4506),
.B2(n_4543),
.Y(n_4720)
);

AOI211xp5_ASAP7_75t_SL g4721 ( 
.A1(n_4610),
.A2(n_4479),
.B(n_4484),
.C(n_4509),
.Y(n_4721)
);

INVx1_ASAP7_75t_L g4722 ( 
.A(n_4608),
.Y(n_4722)
);

OAI21xp33_ASAP7_75t_L g4723 ( 
.A1(n_4616),
.A2(n_4574),
.B(n_482),
.Y(n_4723)
);

OAI22xp33_ASAP7_75t_SL g4724 ( 
.A1(n_4654),
.A2(n_485),
.B1(n_483),
.B2(n_484),
.Y(n_4724)
);

AOI33xp33_ASAP7_75t_L g4725 ( 
.A1(n_4606),
.A2(n_487),
.A3(n_491),
.B1(n_485),
.B2(n_486),
.B3(n_490),
.Y(n_4725)
);

OR2x2_ASAP7_75t_L g4726 ( 
.A(n_4640),
.B(n_486),
.Y(n_4726)
);

INVx1_ASAP7_75t_L g4727 ( 
.A(n_4693),
.Y(n_4727)
);

INVx2_ASAP7_75t_L g4728 ( 
.A(n_4664),
.Y(n_4728)
);

NAND2x2_ASAP7_75t_L g4729 ( 
.A(n_4668),
.B(n_487),
.Y(n_4729)
);

HB1xp67_ASAP7_75t_L g4730 ( 
.A(n_4607),
.Y(n_4730)
);

INVx1_ASAP7_75t_L g4731 ( 
.A(n_4618),
.Y(n_4731)
);

INVx2_ASAP7_75t_L g4732 ( 
.A(n_4627),
.Y(n_4732)
);

AND2x2_ASAP7_75t_L g4733 ( 
.A(n_4605),
.B(n_490),
.Y(n_4733)
);

AOI22xp33_ASAP7_75t_L g4734 ( 
.A1(n_4619),
.A2(n_494),
.B1(n_491),
.B2(n_493),
.Y(n_4734)
);

AND2x2_ASAP7_75t_L g4735 ( 
.A(n_4676),
.B(n_495),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4627),
.Y(n_4736)
);

BUFx2_ASAP7_75t_L g4737 ( 
.A(n_4669),
.Y(n_4737)
);

AOI322xp5_ASAP7_75t_L g4738 ( 
.A1(n_4638),
.A2(n_500),
.A3(n_499),
.B1(n_497),
.B2(n_495),
.C1(n_496),
.C2(n_498),
.Y(n_4738)
);

INVx1_ASAP7_75t_L g4739 ( 
.A(n_4694),
.Y(n_4739)
);

INVx1_ASAP7_75t_L g4740 ( 
.A(n_4630),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4631),
.Y(n_4741)
);

OAI32xp33_ASAP7_75t_L g4742 ( 
.A1(n_4650),
.A2(n_498),
.A3(n_496),
.B1(n_497),
.B2(n_499),
.Y(n_4742)
);

AND2x4_ASAP7_75t_L g4743 ( 
.A(n_4680),
.B(n_500),
.Y(n_4743)
);

OAI32xp33_ASAP7_75t_L g4744 ( 
.A1(n_4670),
.A2(n_503),
.A3(n_501),
.B1(n_502),
.B2(n_504),
.Y(n_4744)
);

INVx1_ASAP7_75t_L g4745 ( 
.A(n_4642),
.Y(n_4745)
);

AND2x2_ASAP7_75t_L g4746 ( 
.A(n_4628),
.B(n_501),
.Y(n_4746)
);

AOI22xp33_ASAP7_75t_SL g4747 ( 
.A1(n_4633),
.A2(n_505),
.B1(n_503),
.B2(n_504),
.Y(n_4747)
);

INVx1_ASAP7_75t_L g4748 ( 
.A(n_4643),
.Y(n_4748)
);

INVx1_ASAP7_75t_L g4749 ( 
.A(n_4614),
.Y(n_4749)
);

INVx1_ASAP7_75t_L g4750 ( 
.A(n_4649),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4652),
.Y(n_4751)
);

INVx3_ASAP7_75t_L g4752 ( 
.A(n_4684),
.Y(n_4752)
);

NOR2xp33_ASAP7_75t_L g4753 ( 
.A(n_4635),
.B(n_4621),
.Y(n_4753)
);

INVx1_ASAP7_75t_L g4754 ( 
.A(n_4662),
.Y(n_4754)
);

BUFx2_ASAP7_75t_L g4755 ( 
.A(n_4634),
.Y(n_4755)
);

AOI211xp5_ASAP7_75t_L g4756 ( 
.A1(n_4677),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_4756)
);

NAND4xp75_ASAP7_75t_SL g4757 ( 
.A(n_4632),
.B(n_509),
.C(n_507),
.D(n_508),
.Y(n_4757)
);

NOR2xp33_ASAP7_75t_L g4758 ( 
.A(n_4698),
.B(n_4666),
.Y(n_4758)
);

INVx1_ASAP7_75t_L g4759 ( 
.A(n_4730),
.Y(n_4759)
);

INVx2_ASAP7_75t_L g4760 ( 
.A(n_4752),
.Y(n_4760)
);

INVx1_ASAP7_75t_L g4761 ( 
.A(n_4755),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4737),
.B(n_4678),
.Y(n_4762)
);

AOI22xp33_ASAP7_75t_L g4763 ( 
.A1(n_4700),
.A2(n_4612),
.B1(n_4611),
.B2(n_4681),
.Y(n_4763)
);

OR2x2_ASAP7_75t_L g4764 ( 
.A(n_4713),
.B(n_4636),
.Y(n_4764)
);

NAND3xp33_ASAP7_75t_L g4765 ( 
.A(n_4756),
.B(n_4683),
.C(n_4687),
.Y(n_4765)
);

OR2x2_ASAP7_75t_L g4766 ( 
.A(n_4697),
.B(n_4648),
.Y(n_4766)
);

NAND2xp5_ASAP7_75t_L g4767 ( 
.A(n_4733),
.B(n_4655),
.Y(n_4767)
);

OR2x2_ASAP7_75t_L g4768 ( 
.A(n_4751),
.B(n_4657),
.Y(n_4768)
);

INVx1_ASAP7_75t_L g4769 ( 
.A(n_4704),
.Y(n_4769)
);

INVx2_ASAP7_75t_L g4770 ( 
.A(n_4716),
.Y(n_4770)
);

OR2x2_ASAP7_75t_L g4771 ( 
.A(n_4714),
.B(n_4661),
.Y(n_4771)
);

NAND2xp5_ASAP7_75t_L g4772 ( 
.A(n_4743),
.B(n_4656),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4735),
.B(n_4695),
.Y(n_4773)
);

NAND2xp5_ASAP7_75t_L g4774 ( 
.A(n_4747),
.B(n_4673),
.Y(n_4774)
);

NAND2xp5_ASAP7_75t_L g4775 ( 
.A(n_4746),
.B(n_4665),
.Y(n_4775)
);

INVxp67_ASAP7_75t_L g4776 ( 
.A(n_4699),
.Y(n_4776)
);

AND2x2_ASAP7_75t_L g4777 ( 
.A(n_4711),
.B(n_4653),
.Y(n_4777)
);

INVx1_ASAP7_75t_L g4778 ( 
.A(n_4750),
.Y(n_4778)
);

OAI21xp33_ASAP7_75t_SL g4779 ( 
.A1(n_4753),
.A2(n_4682),
.B(n_4675),
.Y(n_4779)
);

AND2x2_ASAP7_75t_L g4780 ( 
.A(n_4701),
.B(n_4658),
.Y(n_4780)
);

HB1xp67_ASAP7_75t_L g4781 ( 
.A(n_4732),
.Y(n_4781)
);

INVx3_ASAP7_75t_L g4782 ( 
.A(n_4709),
.Y(n_4782)
);

INVx1_ASAP7_75t_SL g4783 ( 
.A(n_4757),
.Y(n_4783)
);

AOI22xp33_ASAP7_75t_L g4784 ( 
.A1(n_4703),
.A2(n_4691),
.B1(n_4686),
.B2(n_4674),
.Y(n_4784)
);

OR2x2_ASAP7_75t_L g4785 ( 
.A(n_4707),
.B(n_4749),
.Y(n_4785)
);

INVx2_ASAP7_75t_L g4786 ( 
.A(n_4726),
.Y(n_4786)
);

AND2x2_ASAP7_75t_L g4787 ( 
.A(n_4728),
.B(n_4671),
.Y(n_4787)
);

OR2x2_ASAP7_75t_L g4788 ( 
.A(n_4722),
.B(n_4651),
.Y(n_4788)
);

NAND2xp5_ASAP7_75t_L g4789 ( 
.A(n_4739),
.B(n_4623),
.Y(n_4789)
);

INVx1_ASAP7_75t_L g4790 ( 
.A(n_4725),
.Y(n_4790)
);

INVx1_ASAP7_75t_L g4791 ( 
.A(n_4729),
.Y(n_4791)
);

NOR2xp33_ASAP7_75t_L g4792 ( 
.A(n_4724),
.B(n_4626),
.Y(n_4792)
);

INVx2_ASAP7_75t_L g4793 ( 
.A(n_4736),
.Y(n_4793)
);

OR2x2_ASAP7_75t_L g4794 ( 
.A(n_4717),
.B(n_4672),
.Y(n_4794)
);

NAND2xp5_ASAP7_75t_L g4795 ( 
.A(n_4721),
.B(n_4688),
.Y(n_4795)
);

AND2x2_ASAP7_75t_L g4796 ( 
.A(n_4715),
.B(n_4659),
.Y(n_4796)
);

INVx2_ASAP7_75t_L g4797 ( 
.A(n_4754),
.Y(n_4797)
);

NAND5xp2_ASAP7_75t_SL g4798 ( 
.A(n_4706),
.B(n_512),
.C(n_510),
.D(n_511),
.E(n_513),
.Y(n_4798)
);

INVx2_ASAP7_75t_L g4799 ( 
.A(n_4712),
.Y(n_4799)
);

NOR4xp25_ASAP7_75t_SL g4800 ( 
.A(n_4719),
.B(n_514),
.C(n_510),
.D(n_511),
.Y(n_4800)
);

INVx3_ASAP7_75t_L g4801 ( 
.A(n_4731),
.Y(n_4801)
);

NAND2x1p5_ASAP7_75t_L g4802 ( 
.A(n_4740),
.B(n_515),
.Y(n_4802)
);

HB1xp67_ASAP7_75t_L g4803 ( 
.A(n_4718),
.Y(n_4803)
);

INVxp67_ASAP7_75t_L g4804 ( 
.A(n_4710),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4734),
.B(n_515),
.Y(n_4805)
);

INVx1_ASAP7_75t_L g4806 ( 
.A(n_4781),
.Y(n_4806)
);

NOR2xp33_ASAP7_75t_L g4807 ( 
.A(n_4783),
.B(n_4744),
.Y(n_4807)
);

OR2x2_ASAP7_75t_L g4808 ( 
.A(n_4762),
.B(n_4741),
.Y(n_4808)
);

OR2x6_ASAP7_75t_L g4809 ( 
.A(n_4793),
.B(n_4745),
.Y(n_4809)
);

INVx1_ASAP7_75t_SL g4810 ( 
.A(n_4796),
.Y(n_4810)
);

NOR2xp33_ASAP7_75t_L g4811 ( 
.A(n_4770),
.B(n_4705),
.Y(n_4811)
);

OAI221xp5_ASAP7_75t_L g4812 ( 
.A1(n_4763),
.A2(n_4720),
.B1(n_4702),
.B2(n_4727),
.C(n_4723),
.Y(n_4812)
);

AND2x2_ASAP7_75t_L g4813 ( 
.A(n_4761),
.B(n_4748),
.Y(n_4813)
);

NAND2xp5_ASAP7_75t_L g4814 ( 
.A(n_4787),
.B(n_4769),
.Y(n_4814)
);

INVx1_ASAP7_75t_L g4815 ( 
.A(n_4764),
.Y(n_4815)
);

NOR2xp33_ASAP7_75t_L g4816 ( 
.A(n_4773),
.B(n_4742),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4802),
.Y(n_4817)
);

NAND2xp5_ASAP7_75t_L g4818 ( 
.A(n_4777),
.B(n_4738),
.Y(n_4818)
);

INVx2_ASAP7_75t_L g4819 ( 
.A(n_4786),
.Y(n_4819)
);

AOI221xp5_ASAP7_75t_L g4820 ( 
.A1(n_4779),
.A2(n_4708),
.B1(n_4696),
.B2(n_519),
.C(n_516),
.Y(n_4820)
);

AOI211xp5_ASAP7_75t_L g4821 ( 
.A1(n_4758),
.A2(n_521),
.B(n_518),
.C(n_520),
.Y(n_4821)
);

INVx3_ASAP7_75t_L g4822 ( 
.A(n_4782),
.Y(n_4822)
);

INVx1_ASAP7_75t_L g4823 ( 
.A(n_4771),
.Y(n_4823)
);

NAND2xp5_ASAP7_75t_SL g4824 ( 
.A(n_4799),
.B(n_521),
.Y(n_4824)
);

NOR2xp33_ASAP7_75t_L g4825 ( 
.A(n_4774),
.B(n_4767),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4768),
.Y(n_4826)
);

INVx2_ASAP7_75t_L g4827 ( 
.A(n_4791),
.Y(n_4827)
);

AOI211xp5_ASAP7_75t_L g4828 ( 
.A1(n_4795),
.A2(n_524),
.B(n_522),
.C(n_523),
.Y(n_4828)
);

INVx1_ASAP7_75t_L g4829 ( 
.A(n_4759),
.Y(n_4829)
);

OR2x2_ASAP7_75t_L g4830 ( 
.A(n_4785),
.B(n_4766),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4794),
.Y(n_4831)
);

OAI21xp5_ASAP7_75t_L g4832 ( 
.A1(n_4765),
.A2(n_522),
.B(n_523),
.Y(n_4832)
);

INVx3_ASAP7_75t_L g4833 ( 
.A(n_4760),
.Y(n_4833)
);

OAI222xp33_ASAP7_75t_L g4834 ( 
.A1(n_4784),
.A2(n_527),
.B1(n_529),
.B2(n_525),
.C1(n_526),
.C2(n_528),
.Y(n_4834)
);

AND2x2_ASAP7_75t_L g4835 ( 
.A(n_4780),
.B(n_526),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_4792),
.B(n_528),
.Y(n_4836)
);

INVx1_ASAP7_75t_L g4837 ( 
.A(n_4775),
.Y(n_4837)
);

INVxp67_ASAP7_75t_SL g4838 ( 
.A(n_4801),
.Y(n_4838)
);

NAND2x1_ASAP7_75t_L g4839 ( 
.A(n_4778),
.B(n_529),
.Y(n_4839)
);

NAND2xp5_ASAP7_75t_L g4840 ( 
.A(n_4797),
.B(n_530),
.Y(n_4840)
);

NOR2x1_ASAP7_75t_L g4841 ( 
.A(n_4788),
.B(n_531),
.Y(n_4841)
);

OR2x2_ASAP7_75t_L g4842 ( 
.A(n_4789),
.B(n_531),
.Y(n_4842)
);

INVx1_ASAP7_75t_SL g4843 ( 
.A(n_4772),
.Y(n_4843)
);

INVx3_ASAP7_75t_L g4844 ( 
.A(n_4790),
.Y(n_4844)
);

INVx1_ASAP7_75t_SL g4845 ( 
.A(n_4803),
.Y(n_4845)
);

INVx1_ASAP7_75t_L g4846 ( 
.A(n_4804),
.Y(n_4846)
);

INVxp67_ASAP7_75t_SL g4847 ( 
.A(n_4776),
.Y(n_4847)
);

NAND2x1p5_ASAP7_75t_L g4848 ( 
.A(n_4805),
.B(n_533),
.Y(n_4848)
);

INVx1_ASAP7_75t_L g4849 ( 
.A(n_4798),
.Y(n_4849)
);

AND2x2_ASAP7_75t_L g4850 ( 
.A(n_4800),
.B(n_532),
.Y(n_4850)
);

OAI31xp33_ASAP7_75t_SL g4851 ( 
.A1(n_4758),
.A2(n_534),
.A3(n_532),
.B(n_533),
.Y(n_4851)
);

AOI22xp5_ASAP7_75t_L g4852 ( 
.A1(n_4791),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4781),
.B(n_535),
.Y(n_4853)
);

A2O1A1Ixp33_ASAP7_75t_L g4854 ( 
.A1(n_4779),
.A2(n_539),
.B(n_537),
.C(n_538),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4781),
.Y(n_4855)
);

OR2x2_ASAP7_75t_L g4856 ( 
.A(n_4830),
.B(n_539),
.Y(n_4856)
);

INVx1_ASAP7_75t_L g4857 ( 
.A(n_4814),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_4847),
.Y(n_4858)
);

AOI22xp5_ASAP7_75t_L g4859 ( 
.A1(n_4807),
.A2(n_550),
.B1(n_558),
.B2(n_540),
.Y(n_4859)
);

O2A1O1Ixp33_ASAP7_75t_L g4860 ( 
.A1(n_4854),
.A2(n_543),
.B(n_541),
.C(n_542),
.Y(n_4860)
);

INVx1_ASAP7_75t_L g4861 ( 
.A(n_4809),
.Y(n_4861)
);

INVx2_ASAP7_75t_L g4862 ( 
.A(n_4850),
.Y(n_4862)
);

AOI21xp33_ASAP7_75t_SL g4863 ( 
.A1(n_4831),
.A2(n_541),
.B(n_542),
.Y(n_4863)
);

OAI22xp5_ASAP7_75t_L g4864 ( 
.A1(n_4845),
.A2(n_548),
.B1(n_545),
.B2(n_546),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4851),
.B(n_545),
.Y(n_4865)
);

NAND2xp5_ASAP7_75t_L g4866 ( 
.A(n_4835),
.B(n_548),
.Y(n_4866)
);

INVx1_ASAP7_75t_SL g4867 ( 
.A(n_4810),
.Y(n_4867)
);

AOI22xp5_ASAP7_75t_L g4868 ( 
.A1(n_4827),
.A2(n_557),
.B1(n_565),
.B2(n_549),
.Y(n_4868)
);

INVx1_ASAP7_75t_L g4869 ( 
.A(n_4809),
.Y(n_4869)
);

NAND2xp5_ASAP7_75t_L g4870 ( 
.A(n_4841),
.B(n_549),
.Y(n_4870)
);

HB1xp67_ASAP7_75t_L g4871 ( 
.A(n_4839),
.Y(n_4871)
);

OAI22xp33_ASAP7_75t_SL g4872 ( 
.A1(n_4849),
.A2(n_552),
.B1(n_550),
.B2(n_551),
.Y(n_4872)
);

INVx2_ASAP7_75t_L g4873 ( 
.A(n_4848),
.Y(n_4873)
);

OAI22xp33_ASAP7_75t_L g4874 ( 
.A1(n_4818),
.A2(n_553),
.B1(n_551),
.B2(n_552),
.Y(n_4874)
);

BUFx2_ASAP7_75t_L g4875 ( 
.A(n_4806),
.Y(n_4875)
);

INVx1_ASAP7_75t_SL g4876 ( 
.A(n_4808),
.Y(n_4876)
);

O2A1O1Ixp5_ASAP7_75t_L g4877 ( 
.A1(n_4838),
.A2(n_556),
.B(n_554),
.C(n_555),
.Y(n_4877)
);

OAI22xp5_ASAP7_75t_L g4878 ( 
.A1(n_4855),
.A2(n_557),
.B1(n_554),
.B2(n_555),
.Y(n_4878)
);

NAND2xp5_ASAP7_75t_L g4879 ( 
.A(n_4825),
.B(n_558),
.Y(n_4879)
);

AND2x4_ASAP7_75t_L g4880 ( 
.A(n_4833),
.B(n_559),
.Y(n_4880)
);

INVx1_ASAP7_75t_L g4881 ( 
.A(n_4826),
.Y(n_4881)
);

AOI22xp5_ASAP7_75t_L g4882 ( 
.A1(n_4816),
.A2(n_4843),
.B1(n_4846),
.B2(n_4820),
.Y(n_4882)
);

INVx1_ASAP7_75t_L g4883 ( 
.A(n_4823),
.Y(n_4883)
);

INVx1_ASAP7_75t_L g4884 ( 
.A(n_4853),
.Y(n_4884)
);

OAI221xp5_ASAP7_75t_SL g4885 ( 
.A1(n_4812),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.C(n_563),
.Y(n_4885)
);

NAND2xp5_ASAP7_75t_L g4886 ( 
.A(n_4821),
.B(n_560),
.Y(n_4886)
);

NAND2xp5_ASAP7_75t_L g4887 ( 
.A(n_4828),
.B(n_4817),
.Y(n_4887)
);

NAND2xp5_ASAP7_75t_SL g4888 ( 
.A(n_4815),
.B(n_561),
.Y(n_4888)
);

INVx1_ASAP7_75t_L g4889 ( 
.A(n_4842),
.Y(n_4889)
);

OAI22xp5_ASAP7_75t_L g4890 ( 
.A1(n_4837),
.A2(n_565),
.B1(n_562),
.B2(n_564),
.Y(n_4890)
);

NAND3xp33_ASAP7_75t_L g4891 ( 
.A(n_4811),
.B(n_4832),
.C(n_4819),
.Y(n_4891)
);

INVx1_ASAP7_75t_SL g4892 ( 
.A(n_4813),
.Y(n_4892)
);

NAND2xp5_ASAP7_75t_L g4893 ( 
.A(n_4822),
.B(n_566),
.Y(n_4893)
);

INVx1_ASAP7_75t_L g4894 ( 
.A(n_4836),
.Y(n_4894)
);

INVx2_ASAP7_75t_SL g4895 ( 
.A(n_4829),
.Y(n_4895)
);

AND2x4_ASAP7_75t_L g4896 ( 
.A(n_4840),
.B(n_566),
.Y(n_4896)
);

INVx1_ASAP7_75t_L g4897 ( 
.A(n_4844),
.Y(n_4897)
);

OAI322xp33_ASAP7_75t_L g4898 ( 
.A1(n_4824),
.A2(n_572),
.A3(n_571),
.B1(n_569),
.B2(n_567),
.C1(n_568),
.C2(n_570),
.Y(n_4898)
);

BUFx2_ASAP7_75t_L g4899 ( 
.A(n_4852),
.Y(n_4899)
);

O2A1O1Ixp5_ASAP7_75t_L g4900 ( 
.A1(n_4834),
.A2(n_570),
.B(n_567),
.C(n_568),
.Y(n_4900)
);

AND2x2_ASAP7_75t_L g4901 ( 
.A(n_4845),
.B(n_571),
.Y(n_4901)
);

AOI222xp33_ASAP7_75t_L g4902 ( 
.A1(n_4820),
.A2(n_575),
.B1(n_577),
.B2(n_573),
.C1(n_574),
.C2(n_576),
.Y(n_4902)
);

OAI221xp5_ASAP7_75t_L g4903 ( 
.A1(n_4820),
.A2(n_576),
.B1(n_573),
.B2(n_575),
.C(n_577),
.Y(n_4903)
);

INVx1_ASAP7_75t_L g4904 ( 
.A(n_4830),
.Y(n_4904)
);

AOI22xp5_ASAP7_75t_L g4905 ( 
.A1(n_4807),
.A2(n_586),
.B1(n_595),
.B2(n_578),
.Y(n_4905)
);

AOI22xp5_ASAP7_75t_L g4906 ( 
.A1(n_4807),
.A2(n_587),
.B1(n_596),
.B2(n_579),
.Y(n_4906)
);

OAI22xp5_ASAP7_75t_L g4907 ( 
.A1(n_4845),
.A2(n_581),
.B1(n_579),
.B2(n_580),
.Y(n_4907)
);

INVx3_ASAP7_75t_L g4908 ( 
.A(n_4839),
.Y(n_4908)
);

NAND2xp5_ASAP7_75t_L g4909 ( 
.A(n_4851),
.B(n_581),
.Y(n_4909)
);

INVx1_ASAP7_75t_SL g4910 ( 
.A(n_4830),
.Y(n_4910)
);

AND2x2_ASAP7_75t_L g4911 ( 
.A(n_4845),
.B(n_582),
.Y(n_4911)
);

AOI221xp5_ASAP7_75t_L g4912 ( 
.A1(n_4820),
.A2(n_601),
.B1(n_612),
.B2(n_593),
.C(n_583),
.Y(n_4912)
);

INVx1_ASAP7_75t_L g4913 ( 
.A(n_4830),
.Y(n_4913)
);

INVx1_ASAP7_75t_L g4914 ( 
.A(n_4856),
.Y(n_4914)
);

INVx1_ASAP7_75t_L g4915 ( 
.A(n_4904),
.Y(n_4915)
);

OAI32xp33_ASAP7_75t_L g4916 ( 
.A1(n_4910),
.A2(n_585),
.A3(n_583),
.B1(n_584),
.B2(n_586),
.Y(n_4916)
);

INVx1_ASAP7_75t_SL g4917 ( 
.A(n_4892),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4913),
.Y(n_4918)
);

AND2x2_ASAP7_75t_L g4919 ( 
.A(n_4867),
.B(n_4876),
.Y(n_4919)
);

INVx1_ASAP7_75t_L g4920 ( 
.A(n_4866),
.Y(n_4920)
);

OAI32xp33_ASAP7_75t_L g4921 ( 
.A1(n_4871),
.A2(n_588),
.A3(n_584),
.B1(n_585),
.B2(n_589),
.Y(n_4921)
);

INVxp67_ASAP7_75t_L g4922 ( 
.A(n_4908),
.Y(n_4922)
);

AOI211x1_ASAP7_75t_L g4923 ( 
.A1(n_4891),
.A2(n_590),
.B(n_588),
.C(n_589),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4880),
.B(n_590),
.Y(n_4924)
);

HB1xp67_ASAP7_75t_L g4925 ( 
.A(n_4880),
.Y(n_4925)
);

OR2x2_ASAP7_75t_L g4926 ( 
.A(n_4875),
.B(n_591),
.Y(n_4926)
);

OAI221xp5_ASAP7_75t_L g4927 ( 
.A1(n_4882),
.A2(n_594),
.B1(n_591),
.B2(n_593),
.C(n_595),
.Y(n_4927)
);

AND2x2_ASAP7_75t_L g4928 ( 
.A(n_4901),
.B(n_594),
.Y(n_4928)
);

INVxp67_ASAP7_75t_SL g4929 ( 
.A(n_4865),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_4870),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4911),
.Y(n_4931)
);

XOR2x2_ASAP7_75t_L g4932 ( 
.A(n_4885),
.B(n_596),
.Y(n_4932)
);

NAND2xp5_ASAP7_75t_L g4933 ( 
.A(n_4862),
.B(n_597),
.Y(n_4933)
);

INVxp67_ASAP7_75t_L g4934 ( 
.A(n_4909),
.Y(n_4934)
);

NAND2xp5_ASAP7_75t_L g4935 ( 
.A(n_4896),
.B(n_597),
.Y(n_4935)
);

INVx1_ASAP7_75t_L g4936 ( 
.A(n_4879),
.Y(n_4936)
);

INVx2_ASAP7_75t_L g4937 ( 
.A(n_4900),
.Y(n_4937)
);

AOI21xp5_ASAP7_75t_L g4938 ( 
.A1(n_4888),
.A2(n_598),
.B(n_599),
.Y(n_4938)
);

INVx1_ASAP7_75t_L g4939 ( 
.A(n_4896),
.Y(n_4939)
);

INVx2_ASAP7_75t_SL g4940 ( 
.A(n_4861),
.Y(n_4940)
);

INVx1_ASAP7_75t_L g4941 ( 
.A(n_4889),
.Y(n_4941)
);

AOI221xp5_ASAP7_75t_L g4942 ( 
.A1(n_4903),
.A2(n_602),
.B1(n_598),
.B2(n_600),
.C(n_603),
.Y(n_4942)
);

AO22x2_ASAP7_75t_L g4943 ( 
.A1(n_4869),
.A2(n_603),
.B1(n_600),
.B2(n_602),
.Y(n_4943)
);

XNOR2x2_ASAP7_75t_L g4944 ( 
.A(n_4893),
.B(n_606),
.Y(n_4944)
);

INVx1_ASAP7_75t_L g4945 ( 
.A(n_4858),
.Y(n_4945)
);

INVx1_ASAP7_75t_L g4946 ( 
.A(n_4877),
.Y(n_4946)
);

INVx1_ASAP7_75t_L g4947 ( 
.A(n_4886),
.Y(n_4947)
);

AOI31xp33_ASAP7_75t_L g4948 ( 
.A1(n_4857),
.A2(n_609),
.A3(n_606),
.B(n_608),
.Y(n_4948)
);

NAND2xp5_ASAP7_75t_L g4949 ( 
.A(n_4863),
.B(n_610),
.Y(n_4949)
);

INVx1_ASAP7_75t_L g4950 ( 
.A(n_4898),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_4873),
.B(n_611),
.Y(n_4951)
);

OAI332xp33_ASAP7_75t_L g4952 ( 
.A1(n_4887),
.A2(n_617),
.A3(n_616),
.B1(n_614),
.B2(n_618),
.B3(n_611),
.C1(n_613),
.C2(n_615),
.Y(n_4952)
);

AOI211xp5_ASAP7_75t_L g4953 ( 
.A1(n_4912),
.A2(n_616),
.B(n_613),
.C(n_614),
.Y(n_4953)
);

NAND2xp5_ASAP7_75t_L g4954 ( 
.A(n_4872),
.B(n_617),
.Y(n_4954)
);

XNOR2x2_ASAP7_75t_L g4955 ( 
.A(n_4864),
.B(n_618),
.Y(n_4955)
);

INVx1_ASAP7_75t_L g4956 ( 
.A(n_4881),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4894),
.B(n_619),
.Y(n_4957)
);

INVx1_ASAP7_75t_L g4958 ( 
.A(n_4883),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4899),
.Y(n_4959)
);

INVx1_ASAP7_75t_L g4960 ( 
.A(n_4895),
.Y(n_4960)
);

INVx2_ASAP7_75t_L g4961 ( 
.A(n_4884),
.Y(n_4961)
);

INVx1_ASAP7_75t_L g4962 ( 
.A(n_4897),
.Y(n_4962)
);

NAND2xp33_ASAP7_75t_SL g4963 ( 
.A(n_4907),
.B(n_620),
.Y(n_4963)
);

INVx1_ASAP7_75t_L g4964 ( 
.A(n_4859),
.Y(n_4964)
);

OAI21xp33_ASAP7_75t_L g4965 ( 
.A1(n_4902),
.A2(n_620),
.B(n_621),
.Y(n_4965)
);

AOI222xp33_ASAP7_75t_L g4966 ( 
.A1(n_4874),
.A2(n_623),
.B1(n_625),
.B2(n_621),
.C1(n_622),
.C2(n_624),
.Y(n_4966)
);

INVx2_ASAP7_75t_L g4967 ( 
.A(n_4905),
.Y(n_4967)
);

INVxp67_ASAP7_75t_L g4968 ( 
.A(n_4890),
.Y(n_4968)
);

INVx2_ASAP7_75t_L g4969 ( 
.A(n_4906),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4878),
.Y(n_4970)
);

INVx2_ASAP7_75t_L g4971 ( 
.A(n_4868),
.Y(n_4971)
);

NAND2xp5_ASAP7_75t_L g4972 ( 
.A(n_4860),
.B(n_622),
.Y(n_4972)
);

AND2x2_ASAP7_75t_L g4973 ( 
.A(n_4910),
.B(n_626),
.Y(n_4973)
);

INVx1_ASAP7_75t_L g4974 ( 
.A(n_4856),
.Y(n_4974)
);

INVx1_ASAP7_75t_L g4975 ( 
.A(n_4856),
.Y(n_4975)
);

INVx2_ASAP7_75t_L g4976 ( 
.A(n_4908),
.Y(n_4976)
);

OAI221xp5_ASAP7_75t_L g4977 ( 
.A1(n_4882),
.A2(n_628),
.B1(n_626),
.B2(n_627),
.C(n_629),
.Y(n_4977)
);

NAND2xp5_ASAP7_75t_L g4978 ( 
.A(n_4910),
.B(n_629),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4910),
.B(n_630),
.Y(n_4979)
);

INVx1_ASAP7_75t_L g4980 ( 
.A(n_4856),
.Y(n_4980)
);

NAND2xp5_ASAP7_75t_L g4981 ( 
.A(n_4910),
.B(n_631),
.Y(n_4981)
);

NAND4xp75_ASAP7_75t_L g4982 ( 
.A(n_4882),
.B(n_634),
.C(n_631),
.D(n_632),
.Y(n_4982)
);

AND2x2_ASAP7_75t_L g4983 ( 
.A(n_4910),
.B(n_634),
.Y(n_4983)
);

INVx2_ASAP7_75t_L g4984 ( 
.A(n_4908),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4856),
.Y(n_4985)
);

AND2x2_ASAP7_75t_L g4986 ( 
.A(n_4910),
.B(n_635),
.Y(n_4986)
);

INVx1_ASAP7_75t_L g4987 ( 
.A(n_4856),
.Y(n_4987)
);

HB1xp67_ASAP7_75t_L g4988 ( 
.A(n_4871),
.Y(n_4988)
);

OR2x2_ASAP7_75t_L g4989 ( 
.A(n_4910),
.B(n_635),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4910),
.B(n_636),
.Y(n_4990)
);

INVx1_ASAP7_75t_SL g4991 ( 
.A(n_4910),
.Y(n_4991)
);

INVx1_ASAP7_75t_L g4992 ( 
.A(n_4856),
.Y(n_4992)
);

NAND3xp33_ASAP7_75t_SL g4993 ( 
.A(n_4910),
.B(n_637),
.C(n_638),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4910),
.A2(n_637),
.B(n_638),
.Y(n_4994)
);

INVx2_ASAP7_75t_L g4995 ( 
.A(n_4908),
.Y(n_4995)
);

INVx1_ASAP7_75t_L g4996 ( 
.A(n_4856),
.Y(n_4996)
);

NAND2xp5_ASAP7_75t_L g4997 ( 
.A(n_4910),
.B(n_639),
.Y(n_4997)
);

INVx1_ASAP7_75t_L g4998 ( 
.A(n_4856),
.Y(n_4998)
);

INVx1_ASAP7_75t_L g4999 ( 
.A(n_4856),
.Y(n_4999)
);

OAI22xp5_ASAP7_75t_L g5000 ( 
.A1(n_4910),
.A2(n_642),
.B1(n_640),
.B2(n_641),
.Y(n_5000)
);

INVxp67_ASAP7_75t_L g5001 ( 
.A(n_4871),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4856),
.Y(n_5002)
);

NAND2xp5_ASAP7_75t_L g5003 ( 
.A(n_4991),
.B(n_640),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4919),
.A2(n_641),
.B(n_642),
.Y(n_5004)
);

NAND4xp25_ASAP7_75t_L g5005 ( 
.A(n_4917),
.B(n_646),
.C(n_647),
.D(n_645),
.Y(n_5005)
);

OAI21xp33_ASAP7_75t_L g5006 ( 
.A1(n_4940),
.A2(n_643),
.B(n_646),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_L g5007 ( 
.A(n_4923),
.B(n_647),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4925),
.Y(n_5008)
);

INVx1_ASAP7_75t_L g5009 ( 
.A(n_4943),
.Y(n_5009)
);

INVx1_ASAP7_75t_L g5010 ( 
.A(n_4943),
.Y(n_5010)
);

INVx1_ASAP7_75t_L g5011 ( 
.A(n_4988),
.Y(n_5011)
);

AOI21xp33_ASAP7_75t_SL g5012 ( 
.A1(n_4946),
.A2(n_4926),
.B(n_4948),
.Y(n_5012)
);

INVxp67_ASAP7_75t_L g5013 ( 
.A(n_4928),
.Y(n_5013)
);

BUFx3_ASAP7_75t_L g5014 ( 
.A(n_4976),
.Y(n_5014)
);

NAND2xp5_ASAP7_75t_L g5015 ( 
.A(n_4937),
.B(n_648),
.Y(n_5015)
);

INVx1_ASAP7_75t_L g5016 ( 
.A(n_4944),
.Y(n_5016)
);

INVx1_ASAP7_75t_L g5017 ( 
.A(n_4959),
.Y(n_5017)
);

AO21x1_ASAP7_75t_L g5018 ( 
.A1(n_4978),
.A2(n_648),
.B(n_650),
.Y(n_5018)
);

INVx1_ASAP7_75t_L g5019 ( 
.A(n_4973),
.Y(n_5019)
);

INVxp67_ASAP7_75t_L g5020 ( 
.A(n_4983),
.Y(n_5020)
);

INVx1_ASAP7_75t_L g5021 ( 
.A(n_4986),
.Y(n_5021)
);

AOI32xp33_ASAP7_75t_L g5022 ( 
.A1(n_4915),
.A2(n_652),
.A3(n_650),
.B1(n_651),
.B2(n_653),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_L g5023 ( 
.A(n_4952),
.B(n_651),
.Y(n_5023)
);

INVx1_ASAP7_75t_SL g5024 ( 
.A(n_4989),
.Y(n_5024)
);

INVx2_ASAP7_75t_L g5025 ( 
.A(n_4955),
.Y(n_5025)
);

NOR2x1_ASAP7_75t_L g5026 ( 
.A(n_4984),
.B(n_652),
.Y(n_5026)
);

NAND4xp25_ASAP7_75t_L g5027 ( 
.A(n_4960),
.B(n_4918),
.C(n_4922),
.D(n_4995),
.Y(n_5027)
);

AOI211xp5_ASAP7_75t_L g5028 ( 
.A1(n_5001),
.A2(n_655),
.B(n_653),
.C(n_654),
.Y(n_5028)
);

INVx1_ASAP7_75t_L g5029 ( 
.A(n_4935),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_4914),
.B(n_658),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4939),
.Y(n_5031)
);

INVx1_ASAP7_75t_L g5032 ( 
.A(n_4924),
.Y(n_5032)
);

HB1xp67_ASAP7_75t_L g5033 ( 
.A(n_4982),
.Y(n_5033)
);

NAND2xp5_ASAP7_75t_SL g5034 ( 
.A(n_4966),
.B(n_659),
.Y(n_5034)
);

INVx1_ASAP7_75t_L g5035 ( 
.A(n_4954),
.Y(n_5035)
);

INVx2_ASAP7_75t_L g5036 ( 
.A(n_4932),
.Y(n_5036)
);

INVx1_ASAP7_75t_SL g5037 ( 
.A(n_4963),
.Y(n_5037)
);

INVx1_ASAP7_75t_L g5038 ( 
.A(n_4974),
.Y(n_5038)
);

INVx2_ASAP7_75t_SL g5039 ( 
.A(n_4961),
.Y(n_5039)
);

BUFx2_ASAP7_75t_L g5040 ( 
.A(n_4979),
.Y(n_5040)
);

INVx1_ASAP7_75t_L g5041 ( 
.A(n_4975),
.Y(n_5041)
);

NAND2xp5_ASAP7_75t_L g5042 ( 
.A(n_4980),
.B(n_659),
.Y(n_5042)
);

OR2x2_ASAP7_75t_L g5043 ( 
.A(n_4981),
.B(n_4990),
.Y(n_5043)
);

NAND2xp5_ASAP7_75t_L g5044 ( 
.A(n_4985),
.B(n_660),
.Y(n_5044)
);

NAND2xp5_ASAP7_75t_SL g5045 ( 
.A(n_4931),
.B(n_661),
.Y(n_5045)
);

NAND2xp5_ASAP7_75t_L g5046 ( 
.A(n_4987),
.B(n_663),
.Y(n_5046)
);

O2A1O1Ixp33_ASAP7_75t_L g5047 ( 
.A1(n_4927),
.A2(n_666),
.B(n_664),
.C(n_665),
.Y(n_5047)
);

INVxp67_ASAP7_75t_SL g5048 ( 
.A(n_4997),
.Y(n_5048)
);

INVx2_ASAP7_75t_L g5049 ( 
.A(n_4992),
.Y(n_5049)
);

XNOR2xp5_ASAP7_75t_L g5050 ( 
.A(n_4993),
.B(n_666),
.Y(n_5050)
);

INVx1_ASAP7_75t_L g5051 ( 
.A(n_4996),
.Y(n_5051)
);

NOR3xp33_ASAP7_75t_L g5052 ( 
.A(n_4977),
.B(n_665),
.C(n_667),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4998),
.B(n_667),
.Y(n_5053)
);

AOI22xp33_ASAP7_75t_L g5054 ( 
.A1(n_4930),
.A2(n_670),
.B1(n_668),
.B2(n_669),
.Y(n_5054)
);

OR2x2_ASAP7_75t_L g5055 ( 
.A(n_4941),
.B(n_670),
.Y(n_5055)
);

AND2x2_ASAP7_75t_L g5056 ( 
.A(n_4962),
.B(n_671),
.Y(n_5056)
);

NAND2xp33_ASAP7_75t_L g5057 ( 
.A(n_4956),
.B(n_671),
.Y(n_5057)
);

AND2x2_ASAP7_75t_L g5058 ( 
.A(n_4958),
.B(n_672),
.Y(n_5058)
);

NOR2xp33_ASAP7_75t_L g5059 ( 
.A(n_4921),
.B(n_672),
.Y(n_5059)
);

OAI21x1_ASAP7_75t_L g5060 ( 
.A1(n_4994),
.A2(n_673),
.B(n_674),
.Y(n_5060)
);

BUFx2_ASAP7_75t_L g5061 ( 
.A(n_4934),
.Y(n_5061)
);

OR2x2_ASAP7_75t_L g5062 ( 
.A(n_4945),
.B(n_674),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_4999),
.B(n_675),
.Y(n_5063)
);

INVx2_ASAP7_75t_L g5064 ( 
.A(n_5002),
.Y(n_5064)
);

NAND2xp5_ASAP7_75t_L g5065 ( 
.A(n_4929),
.B(n_676),
.Y(n_5065)
);

XNOR2xp5_ASAP7_75t_L g5066 ( 
.A(n_4950),
.B(n_677),
.Y(n_5066)
);

AOI31xp33_ASAP7_75t_R g5067 ( 
.A1(n_4965),
.A2(n_679),
.A3(n_676),
.B(n_678),
.Y(n_5067)
);

NAND2xp33_ASAP7_75t_SL g5068 ( 
.A(n_5000),
.B(n_678),
.Y(n_5068)
);

OA21x2_ASAP7_75t_SL g5069 ( 
.A1(n_4933),
.A2(n_681),
.B(n_680),
.Y(n_5069)
);

AND2x2_ASAP7_75t_L g5070 ( 
.A(n_4970),
.B(n_679),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4949),
.Y(n_5071)
);

AND2x2_ASAP7_75t_L g5072 ( 
.A(n_4936),
.B(n_680),
.Y(n_5072)
);

INVx1_ASAP7_75t_L g5073 ( 
.A(n_4972),
.Y(n_5073)
);

INVx2_ASAP7_75t_L g5074 ( 
.A(n_4920),
.Y(n_5074)
);

NAND2xp33_ASAP7_75t_R g5075 ( 
.A(n_4951),
.B(n_4957),
.Y(n_5075)
);

XNOR2x2_ASAP7_75t_L g5076 ( 
.A(n_4938),
.B(n_681),
.Y(n_5076)
);

NAND2xp5_ASAP7_75t_L g5077 ( 
.A(n_4953),
.B(n_682),
.Y(n_5077)
);

INVx1_ASAP7_75t_L g5078 ( 
.A(n_4916),
.Y(n_5078)
);

NAND2xp5_ASAP7_75t_L g5079 ( 
.A(n_4968),
.B(n_683),
.Y(n_5079)
);

NAND2xp5_ASAP7_75t_L g5080 ( 
.A(n_4964),
.B(n_683),
.Y(n_5080)
);

INVx1_ASAP7_75t_L g5081 ( 
.A(n_4967),
.Y(n_5081)
);

NAND3xp33_ASAP7_75t_L g5082 ( 
.A(n_4942),
.B(n_4947),
.C(n_4969),
.Y(n_5082)
);

AOI22xp33_ASAP7_75t_L g5083 ( 
.A1(n_4971),
.A2(n_686),
.B1(n_684),
.B2(n_685),
.Y(n_5083)
);

NOR2xp33_ASAP7_75t_SL g5084 ( 
.A(n_4991),
.B(n_684),
.Y(n_5084)
);

INVx1_ASAP7_75t_L g5085 ( 
.A(n_4925),
.Y(n_5085)
);

INVx1_ASAP7_75t_SL g5086 ( 
.A(n_4991),
.Y(n_5086)
);

AND2x2_ASAP7_75t_L g5087 ( 
.A(n_4919),
.B(n_686),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4925),
.Y(n_5088)
);

AND4x1_ASAP7_75t_L g5089 ( 
.A(n_5084),
.B(n_689),
.C(n_687),
.D(n_688),
.Y(n_5089)
);

AO22x2_ASAP7_75t_L g5090 ( 
.A1(n_5009),
.A2(n_690),
.B1(n_687),
.B2(n_688),
.Y(n_5090)
);

AOI211xp5_ASAP7_75t_SL g5091 ( 
.A1(n_5017),
.A2(n_692),
.B(n_690),
.C(n_691),
.Y(n_5091)
);

OAI21xp33_ASAP7_75t_SL g5092 ( 
.A1(n_5086),
.A2(n_692),
.B(n_693),
.Y(n_5092)
);

NOR2x1_ASAP7_75t_L g5093 ( 
.A(n_5014),
.B(n_693),
.Y(n_5093)
);

AOI22xp5_ASAP7_75t_L g5094 ( 
.A1(n_5061),
.A2(n_696),
.B1(n_694),
.B2(n_695),
.Y(n_5094)
);

OAI21xp33_ASAP7_75t_L g5095 ( 
.A1(n_5027),
.A2(n_5039),
.B(n_5008),
.Y(n_5095)
);

OAI21x1_ASAP7_75t_L g5096 ( 
.A1(n_5026),
.A2(n_5060),
.B(n_5004),
.Y(n_5096)
);

AOI211xp5_ASAP7_75t_L g5097 ( 
.A1(n_5012),
.A2(n_698),
.B(n_695),
.C(n_697),
.Y(n_5097)
);

OAI211xp5_ASAP7_75t_L g5098 ( 
.A1(n_5011),
.A2(n_700),
.B(n_697),
.C(n_699),
.Y(n_5098)
);

NOR3xp33_ASAP7_75t_L g5099 ( 
.A(n_5016),
.B(n_699),
.C(n_701),
.Y(n_5099)
);

AOI22xp5_ASAP7_75t_L g5100 ( 
.A1(n_5035),
.A2(n_704),
.B1(n_702),
.B2(n_703),
.Y(n_5100)
);

NOR3x1_ASAP7_75t_L g5101 ( 
.A(n_5003),
.B(n_705),
.C(n_706),
.Y(n_5101)
);

AO22x2_ASAP7_75t_L g5102 ( 
.A1(n_5010),
.A2(n_707),
.B1(n_705),
.B2(n_706),
.Y(n_5102)
);

AOI211x1_ASAP7_75t_L g5103 ( 
.A1(n_5085),
.A2(n_709),
.B(n_707),
.C(n_708),
.Y(n_5103)
);

INVx2_ASAP7_75t_L g5104 ( 
.A(n_5076),
.Y(n_5104)
);

NAND2xp5_ASAP7_75t_L g5105 ( 
.A(n_5087),
.B(n_709),
.Y(n_5105)
);

NOR2x1_ASAP7_75t_L g5106 ( 
.A(n_5088),
.B(n_710),
.Y(n_5106)
);

NOR2x1_ASAP7_75t_L g5107 ( 
.A(n_5038),
.B(n_711),
.Y(n_5107)
);

AND2x2_ASAP7_75t_L g5108 ( 
.A(n_5041),
.B(n_712),
.Y(n_5108)
);

AOI211x1_ASAP7_75t_L g5109 ( 
.A1(n_5018),
.A2(n_714),
.B(n_712),
.C(n_713),
.Y(n_5109)
);

AO22x2_ASAP7_75t_L g5110 ( 
.A1(n_5025),
.A2(n_717),
.B1(n_713),
.B2(n_716),
.Y(n_5110)
);

INVx1_ASAP7_75t_L g5111 ( 
.A(n_5050),
.Y(n_5111)
);

INVx2_ASAP7_75t_SL g5112 ( 
.A(n_5056),
.Y(n_5112)
);

AOI21xp5_ASAP7_75t_L g5113 ( 
.A1(n_5023),
.A2(n_717),
.B(n_718),
.Y(n_5113)
);

NOR3x1_ASAP7_75t_L g5114 ( 
.A(n_5045),
.B(n_718),
.C(n_719),
.Y(n_5114)
);

NOR3xp33_ASAP7_75t_L g5115 ( 
.A(n_5015),
.B(n_719),
.C(n_720),
.Y(n_5115)
);

INVx1_ASAP7_75t_L g5116 ( 
.A(n_5007),
.Y(n_5116)
);

AOI22xp5_ASAP7_75t_L g5117 ( 
.A1(n_5073),
.A2(n_723),
.B1(n_721),
.B2(n_722),
.Y(n_5117)
);

AOI21xp5_ASAP7_75t_L g5118 ( 
.A1(n_5057),
.A2(n_721),
.B(n_722),
.Y(n_5118)
);

AOI21xp5_ASAP7_75t_L g5119 ( 
.A1(n_5006),
.A2(n_723),
.B(n_724),
.Y(n_5119)
);

NOR2xp33_ASAP7_75t_L g5120 ( 
.A(n_5005),
.B(n_724),
.Y(n_5120)
);

AOI211xp5_ASAP7_75t_L g5121 ( 
.A1(n_5051),
.A2(n_727),
.B(n_725),
.C(n_726),
.Y(n_5121)
);

AOI22xp5_ASAP7_75t_L g5122 ( 
.A1(n_5075),
.A2(n_727),
.B1(n_725),
.B2(n_726),
.Y(n_5122)
);

OR2x2_ASAP7_75t_L g5123 ( 
.A(n_5049),
.B(n_728),
.Y(n_5123)
);

AOI21xp5_ASAP7_75t_L g5124 ( 
.A1(n_5068),
.A2(n_729),
.B(n_730),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_5024),
.B(n_730),
.Y(n_5125)
);

AOI21xp5_ASAP7_75t_L g5126 ( 
.A1(n_5064),
.A2(n_731),
.B(n_733),
.Y(n_5126)
);

INVx1_ASAP7_75t_L g5127 ( 
.A(n_5072),
.Y(n_5127)
);

NOR3xp33_ASAP7_75t_L g5128 ( 
.A(n_5065),
.B(n_733),
.C(n_734),
.Y(n_5128)
);

HB1xp67_ASAP7_75t_L g5129 ( 
.A(n_5013),
.Y(n_5129)
);

AOI22xp5_ASAP7_75t_L g5130 ( 
.A1(n_5071),
.A2(n_736),
.B1(n_734),
.B2(n_735),
.Y(n_5130)
);

NOR3xp33_ASAP7_75t_L g5131 ( 
.A(n_5080),
.B(n_735),
.C(n_736),
.Y(n_5131)
);

OAI21xp33_ASAP7_75t_L g5132 ( 
.A1(n_5031),
.A2(n_737),
.B(n_738),
.Y(n_5132)
);

INVx1_ASAP7_75t_L g5133 ( 
.A(n_5058),
.Y(n_5133)
);

OR2x2_ASAP7_75t_L g5134 ( 
.A(n_5062),
.B(n_738),
.Y(n_5134)
);

INVx2_ASAP7_75t_L g5135 ( 
.A(n_5055),
.Y(n_5135)
);

OAI21xp33_ASAP7_75t_SL g5136 ( 
.A1(n_5037),
.A2(n_739),
.B(n_740),
.Y(n_5136)
);

AOI211xp5_ASAP7_75t_L g5137 ( 
.A1(n_5059),
.A2(n_5074),
.B(n_5066),
.C(n_5078),
.Y(n_5137)
);

AOI22xp5_ASAP7_75t_L g5138 ( 
.A1(n_5048),
.A2(n_742),
.B1(n_740),
.B2(n_741),
.Y(n_5138)
);

NAND2xp5_ASAP7_75t_L g5139 ( 
.A(n_5020),
.B(n_741),
.Y(n_5139)
);

NOR2x1_ASAP7_75t_L g5140 ( 
.A(n_5030),
.B(n_742),
.Y(n_5140)
);

AOI22xp5_ASAP7_75t_L g5141 ( 
.A1(n_5019),
.A2(n_745),
.B1(n_743),
.B2(n_744),
.Y(n_5141)
);

NAND2xp5_ASAP7_75t_L g5142 ( 
.A(n_5021),
.B(n_743),
.Y(n_5142)
);

AOI221xp5_ASAP7_75t_L g5143 ( 
.A1(n_5029),
.A2(n_747),
.B1(n_744),
.B2(n_746),
.C(n_748),
.Y(n_5143)
);

INVx1_ASAP7_75t_L g5144 ( 
.A(n_5040),
.Y(n_5144)
);

INVx1_ASAP7_75t_L g5145 ( 
.A(n_5070),
.Y(n_5145)
);

OAI211xp5_ASAP7_75t_SL g5146 ( 
.A1(n_5036),
.A2(n_749),
.B(n_746),
.C(n_747),
.Y(n_5146)
);

NOR2xp33_ASAP7_75t_L g5147 ( 
.A(n_5033),
.B(n_749),
.Y(n_5147)
);

OAI21xp5_ASAP7_75t_L g5148 ( 
.A1(n_5079),
.A2(n_750),
.B(n_751),
.Y(n_5148)
);

AOI22xp5_ASAP7_75t_L g5149 ( 
.A1(n_5032),
.A2(n_752),
.B1(n_750),
.B2(n_751),
.Y(n_5149)
);

XOR2x2_ASAP7_75t_L g5150 ( 
.A(n_5082),
.B(n_752),
.Y(n_5150)
);

NOR2xp67_ASAP7_75t_L g5151 ( 
.A(n_5042),
.B(n_753),
.Y(n_5151)
);

AOI22xp5_ASAP7_75t_L g5152 ( 
.A1(n_5034),
.A2(n_758),
.B1(n_754),
.B2(n_757),
.Y(n_5152)
);

INVx1_ASAP7_75t_L g5153 ( 
.A(n_5043),
.Y(n_5153)
);

OAI22xp5_ASAP7_75t_L g5154 ( 
.A1(n_5083),
.A2(n_760),
.B1(n_757),
.B2(n_759),
.Y(n_5154)
);

OAI22x1_ASAP7_75t_L g5155 ( 
.A1(n_5081),
.A2(n_762),
.B1(n_760),
.B2(n_761),
.Y(n_5155)
);

AOI21xp5_ASAP7_75t_L g5156 ( 
.A1(n_5044),
.A2(n_5053),
.B(n_5046),
.Y(n_5156)
);

AO22x2_ASAP7_75t_L g5157 ( 
.A1(n_5063),
.A2(n_764),
.B1(n_762),
.B2(n_763),
.Y(n_5157)
);

NAND2xp5_ASAP7_75t_L g5158 ( 
.A(n_5028),
.B(n_763),
.Y(n_5158)
);

OR2x2_ASAP7_75t_L g5159 ( 
.A(n_5077),
.B(n_764),
.Y(n_5159)
);

AOI211xp5_ASAP7_75t_L g5160 ( 
.A1(n_5052),
.A2(n_5047),
.B(n_5067),
.C(n_5069),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_5022),
.B(n_765),
.Y(n_5161)
);

NOR3x1_ASAP7_75t_L g5162 ( 
.A(n_5054),
.B(n_765),
.C(n_766),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_5086),
.B(n_767),
.Y(n_5163)
);

AOI21xp5_ASAP7_75t_L g5164 ( 
.A1(n_5086),
.A2(n_767),
.B(n_768),
.Y(n_5164)
);

NAND2xp5_ASAP7_75t_L g5165 ( 
.A(n_5086),
.B(n_768),
.Y(n_5165)
);

NOR3xp33_ASAP7_75t_SL g5166 ( 
.A(n_5027),
.B(n_769),
.C(n_770),
.Y(n_5166)
);

AOI22xp5_ASAP7_75t_L g5167 ( 
.A1(n_5061),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.Y(n_5167)
);

INVxp67_ASAP7_75t_L g5168 ( 
.A(n_5084),
.Y(n_5168)
);

INVx1_ASAP7_75t_L g5169 ( 
.A(n_5018),
.Y(n_5169)
);

INVx2_ASAP7_75t_L g5170 ( 
.A(n_5014),
.Y(n_5170)
);

AOI211x1_ASAP7_75t_L g5171 ( 
.A1(n_5027),
.A2(n_774),
.B(n_772),
.C(n_773),
.Y(n_5171)
);

INVx2_ASAP7_75t_SL g5172 ( 
.A(n_5014),
.Y(n_5172)
);

AOI211xp5_ASAP7_75t_L g5173 ( 
.A1(n_5012),
.A2(n_776),
.B(n_773),
.C(n_775),
.Y(n_5173)
);

NOR3xp33_ASAP7_75t_SL g5174 ( 
.A(n_5027),
.B(n_775),
.C(n_776),
.Y(n_5174)
);

AOI211xp5_ASAP7_75t_L g5175 ( 
.A1(n_5012),
.A2(n_780),
.B(n_778),
.C(n_779),
.Y(n_5175)
);

NOR2xp33_ASAP7_75t_L g5176 ( 
.A(n_5084),
.B(n_779),
.Y(n_5176)
);

INVx1_ASAP7_75t_L g5177 ( 
.A(n_5090),
.Y(n_5177)
);

NOR2x1_ASAP7_75t_L g5178 ( 
.A(n_5170),
.B(n_780),
.Y(n_5178)
);

INVx1_ASAP7_75t_L g5179 ( 
.A(n_5090),
.Y(n_5179)
);

INVx1_ASAP7_75t_L g5180 ( 
.A(n_5102),
.Y(n_5180)
);

INVx1_ASAP7_75t_L g5181 ( 
.A(n_5102),
.Y(n_5181)
);

INVx1_ASAP7_75t_L g5182 ( 
.A(n_5110),
.Y(n_5182)
);

INVx2_ASAP7_75t_L g5183 ( 
.A(n_5157),
.Y(n_5183)
);

AND2x2_ASAP7_75t_L g5184 ( 
.A(n_5172),
.B(n_781),
.Y(n_5184)
);

INVxp67_ASAP7_75t_L g5185 ( 
.A(n_5093),
.Y(n_5185)
);

OAI22xp5_ASAP7_75t_L g5186 ( 
.A1(n_5163),
.A2(n_785),
.B1(n_783),
.B2(n_784),
.Y(n_5186)
);

NAND2xp5_ASAP7_75t_L g5187 ( 
.A(n_5109),
.B(n_786),
.Y(n_5187)
);

OAI22xp33_ASAP7_75t_L g5188 ( 
.A1(n_5104),
.A2(n_788),
.B1(n_785),
.B2(n_787),
.Y(n_5188)
);

OAI21xp5_ASAP7_75t_SL g5189 ( 
.A1(n_5129),
.A2(n_787),
.B(n_788),
.Y(n_5189)
);

NAND2x1p5_ASAP7_75t_L g5190 ( 
.A(n_5144),
.B(n_789),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_5171),
.B(n_5103),
.Y(n_5191)
);

NAND2xp5_ASAP7_75t_L g5192 ( 
.A(n_5091),
.B(n_790),
.Y(n_5192)
);

AOI31xp33_ASAP7_75t_L g5193 ( 
.A1(n_5095),
.A2(n_791),
.A3(n_789),
.B(n_790),
.Y(n_5193)
);

A2O1A1Ixp33_ASAP7_75t_L g5194 ( 
.A1(n_5113),
.A2(n_794),
.B(n_792),
.C(n_793),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5110),
.Y(n_5195)
);

AOI22xp33_ASAP7_75t_L g5196 ( 
.A1(n_5116),
.A2(n_5135),
.B1(n_5151),
.B2(n_5140),
.Y(n_5196)
);

OAI21xp5_ASAP7_75t_SL g5197 ( 
.A1(n_5168),
.A2(n_792),
.B(n_793),
.Y(n_5197)
);

NAND2x1_ASAP7_75t_L g5198 ( 
.A(n_5106),
.B(n_794),
.Y(n_5198)
);

OAI22xp33_ASAP7_75t_SL g5199 ( 
.A1(n_5169),
.A2(n_5134),
.B1(n_5123),
.B2(n_5153),
.Y(n_5199)
);

INVx2_ASAP7_75t_SL g5200 ( 
.A(n_5108),
.Y(n_5200)
);

NOR2xp33_ASAP7_75t_L g5201 ( 
.A(n_5089),
.B(n_796),
.Y(n_5201)
);

OAI211xp5_ASAP7_75t_L g5202 ( 
.A1(n_5092),
.A2(n_798),
.B(n_796),
.C(n_797),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_SL g5203 ( 
.A(n_5136),
.B(n_799),
.Y(n_5203)
);

INVx1_ASAP7_75t_L g5204 ( 
.A(n_5157),
.Y(n_5204)
);

INVx1_ASAP7_75t_L g5205 ( 
.A(n_5107),
.Y(n_5205)
);

INVxp67_ASAP7_75t_L g5206 ( 
.A(n_5176),
.Y(n_5206)
);

INVx2_ASAP7_75t_L g5207 ( 
.A(n_5101),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_SL g5208 ( 
.A(n_5166),
.B(n_5174),
.Y(n_5208)
);

OAI21xp33_ASAP7_75t_SL g5209 ( 
.A1(n_5165),
.A2(n_800),
.B(n_801),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_5114),
.B(n_5120),
.Y(n_5210)
);

XNOR2xp5_ASAP7_75t_L g5211 ( 
.A(n_5150),
.B(n_803),
.Y(n_5211)
);

OA22x2_ASAP7_75t_L g5212 ( 
.A1(n_5152),
.A2(n_806),
.B1(n_804),
.B2(n_805),
.Y(n_5212)
);

INVx1_ASAP7_75t_L g5213 ( 
.A(n_5105),
.Y(n_5213)
);

OAI21xp33_ASAP7_75t_L g5214 ( 
.A1(n_5147),
.A2(n_805),
.B(n_806),
.Y(n_5214)
);

AND2x2_ASAP7_75t_L g5215 ( 
.A(n_5099),
.B(n_807),
.Y(n_5215)
);

INVx1_ASAP7_75t_L g5216 ( 
.A(n_5155),
.Y(n_5216)
);

INVx1_ASAP7_75t_SL g5217 ( 
.A(n_5159),
.Y(n_5217)
);

AOI21xp5_ASAP7_75t_L g5218 ( 
.A1(n_5164),
.A2(n_807),
.B(n_808),
.Y(n_5218)
);

INVx2_ASAP7_75t_L g5219 ( 
.A(n_5096),
.Y(n_5219)
);

A2O1A1Ixp33_ASAP7_75t_L g5220 ( 
.A1(n_5119),
.A2(n_811),
.B(n_809),
.C(n_810),
.Y(n_5220)
);

INVx1_ASAP7_75t_L g5221 ( 
.A(n_5112),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_5125),
.Y(n_5222)
);

XNOR2xp5_ASAP7_75t_L g5223 ( 
.A(n_5137),
.B(n_809),
.Y(n_5223)
);

AND2x2_ASAP7_75t_L g5224 ( 
.A(n_5097),
.B(n_810),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_5160),
.B(n_813),
.Y(n_5225)
);

AOI22xp33_ASAP7_75t_L g5226 ( 
.A1(n_5127),
.A2(n_5133),
.B1(n_5145),
.B2(n_5156),
.Y(n_5226)
);

AND3x4_ASAP7_75t_L g5227 ( 
.A(n_5128),
.B(n_5131),
.C(n_5115),
.Y(n_5227)
);

INVx1_ASAP7_75t_L g5228 ( 
.A(n_5146),
.Y(n_5228)
);

OAI21xp33_ASAP7_75t_SL g5229 ( 
.A1(n_5161),
.A2(n_812),
.B(n_813),
.Y(n_5229)
);

HB1xp67_ASAP7_75t_L g5230 ( 
.A(n_5162),
.Y(n_5230)
);

INVx1_ASAP7_75t_L g5231 ( 
.A(n_5142),
.Y(n_5231)
);

AOI22xp5_ASAP7_75t_L g5232 ( 
.A1(n_5111),
.A2(n_815),
.B1(n_812),
.B2(n_814),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5158),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_5139),
.Y(n_5234)
);

AND2x4_ASAP7_75t_L g5235 ( 
.A(n_5148),
.B(n_816),
.Y(n_5235)
);

XOR2x2_ASAP7_75t_L g5236 ( 
.A(n_5173),
.B(n_5175),
.Y(n_5236)
);

NOR2x1p5_ASAP7_75t_L g5237 ( 
.A(n_5098),
.B(n_5132),
.Y(n_5237)
);

AOI322xp5_ASAP7_75t_L g5238 ( 
.A1(n_5122),
.A2(n_823),
.A3(n_820),
.B1(n_818),
.B2(n_816),
.C1(n_817),
.C2(n_819),
.Y(n_5238)
);

INVx1_ASAP7_75t_L g5239 ( 
.A(n_5138),
.Y(n_5239)
);

OAI21xp33_ASAP7_75t_SL g5240 ( 
.A1(n_5124),
.A2(n_819),
.B(n_820),
.Y(n_5240)
);

NAND2xp5_ASAP7_75t_SL g5241 ( 
.A(n_5121),
.B(n_823),
.Y(n_5241)
);

AOI211xp5_ASAP7_75t_SL g5242 ( 
.A1(n_5126),
.A2(n_826),
.B(n_824),
.C(n_825),
.Y(n_5242)
);

INVx1_ASAP7_75t_L g5243 ( 
.A(n_5141),
.Y(n_5243)
);

AOI221xp5_ASAP7_75t_L g5244 ( 
.A1(n_5118),
.A2(n_826),
.B1(n_824),
.B2(n_825),
.C(n_827),
.Y(n_5244)
);

OAI22xp33_ASAP7_75t_L g5245 ( 
.A1(n_5100),
.A2(n_829),
.B1(n_827),
.B2(n_828),
.Y(n_5245)
);

NOR2xp33_ASAP7_75t_L g5246 ( 
.A(n_5154),
.B(n_829),
.Y(n_5246)
);

OAI22xp5_ASAP7_75t_L g5247 ( 
.A1(n_5117),
.A2(n_5167),
.B1(n_5094),
.B2(n_5130),
.Y(n_5247)
);

XOR2x2_ASAP7_75t_L g5248 ( 
.A(n_5149),
.B(n_830),
.Y(n_5248)
);

CKINVDCx20_ASAP7_75t_R g5249 ( 
.A(n_5143),
.Y(n_5249)
);

INVx1_ASAP7_75t_L g5250 ( 
.A(n_5090),
.Y(n_5250)
);

OAI221xp5_ASAP7_75t_L g5251 ( 
.A1(n_5129),
.A2(n_832),
.B1(n_830),
.B2(n_831),
.C(n_833),
.Y(n_5251)
);

AOI21xp5_ASAP7_75t_L g5252 ( 
.A1(n_5095),
.A2(n_831),
.B(n_833),
.Y(n_5252)
);

NOR3xp33_ASAP7_75t_L g5253 ( 
.A(n_5144),
.B(n_834),
.C(n_835),
.Y(n_5253)
);

NAND2xp5_ASAP7_75t_L g5254 ( 
.A(n_5185),
.B(n_834),
.Y(n_5254)
);

HB1xp67_ASAP7_75t_L g5255 ( 
.A(n_5198),
.Y(n_5255)
);

INVxp67_ASAP7_75t_SL g5256 ( 
.A(n_5178),
.Y(n_5256)
);

OA22x2_ASAP7_75t_L g5257 ( 
.A1(n_5197),
.A2(n_838),
.B1(n_835),
.B2(n_836),
.Y(n_5257)
);

AOI22xp5_ASAP7_75t_L g5258 ( 
.A1(n_5219),
.A2(n_839),
.B1(n_836),
.B2(n_838),
.Y(n_5258)
);

NOR2xp67_ASAP7_75t_L g5259 ( 
.A(n_5221),
.B(n_839),
.Y(n_5259)
);

NAND4xp25_ASAP7_75t_SL g5260 ( 
.A(n_5252),
.B(n_842),
.C(n_840),
.D(n_841),
.Y(n_5260)
);

INVx1_ASAP7_75t_L g5261 ( 
.A(n_5190),
.Y(n_5261)
);

AO22x2_ASAP7_75t_L g5262 ( 
.A1(n_5177),
.A2(n_842),
.B1(n_840),
.B2(n_841),
.Y(n_5262)
);

AO22x1_ASAP7_75t_L g5263 ( 
.A1(n_5253),
.A2(n_845),
.B1(n_843),
.B2(n_844),
.Y(n_5263)
);

AO22x1_ASAP7_75t_L g5264 ( 
.A1(n_5216),
.A2(n_846),
.B1(n_843),
.B2(n_845),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_5205),
.B(n_847),
.Y(n_5265)
);

NOR4xp25_ASAP7_75t_L g5266 ( 
.A(n_5229),
.B(n_849),
.C(n_847),
.D(n_848),
.Y(n_5266)
);

AOI22xp5_ASAP7_75t_L g5267 ( 
.A1(n_5247),
.A2(n_5233),
.B1(n_5231),
.B2(n_5200),
.Y(n_5267)
);

AOI22xp5_ASAP7_75t_L g5268 ( 
.A1(n_5210),
.A2(n_851),
.B1(n_849),
.B2(n_850),
.Y(n_5268)
);

NOR2x1_ASAP7_75t_L g5269 ( 
.A(n_5184),
.B(n_850),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5191),
.Y(n_5270)
);

AOI22xp5_ASAP7_75t_L g5271 ( 
.A1(n_5203),
.A2(n_854),
.B1(n_852),
.B2(n_853),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_L g5272 ( 
.A(n_5207),
.B(n_852),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_SL g5273 ( 
.A(n_5199),
.B(n_853),
.Y(n_5273)
);

AOI22xp5_ASAP7_75t_L g5274 ( 
.A1(n_5234),
.A2(n_857),
.B1(n_855),
.B2(n_856),
.Y(n_5274)
);

AO22x2_ASAP7_75t_L g5275 ( 
.A1(n_5179),
.A2(n_859),
.B1(n_857),
.B2(n_858),
.Y(n_5275)
);

HB1xp67_ASAP7_75t_L g5276 ( 
.A(n_5180),
.Y(n_5276)
);

INVxp67_ASAP7_75t_SL g5277 ( 
.A(n_5192),
.Y(n_5277)
);

NAND2xp5_ASAP7_75t_L g5278 ( 
.A(n_5182),
.B(n_859),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5181),
.Y(n_5279)
);

HB1xp67_ASAP7_75t_L g5280 ( 
.A(n_5250),
.Y(n_5280)
);

AOI22xp5_ASAP7_75t_L g5281 ( 
.A1(n_5201),
.A2(n_863),
.B1(n_861),
.B2(n_862),
.Y(n_5281)
);

NOR2x1_ASAP7_75t_L g5282 ( 
.A(n_5189),
.B(n_863),
.Y(n_5282)
);

AOI22xp5_ASAP7_75t_L g5283 ( 
.A1(n_5228),
.A2(n_866),
.B1(n_864),
.B2(n_865),
.Y(n_5283)
);

INVx2_ASAP7_75t_L g5284 ( 
.A(n_5183),
.Y(n_5284)
);

AOI221xp5_ASAP7_75t_L g5285 ( 
.A1(n_5218),
.A2(n_867),
.B1(n_865),
.B2(n_866),
.C(n_868),
.Y(n_5285)
);

NAND2xp5_ASAP7_75t_L g5286 ( 
.A(n_5195),
.B(n_869),
.Y(n_5286)
);

INVx1_ASAP7_75t_L g5287 ( 
.A(n_5187),
.Y(n_5287)
);

AO22x1_ASAP7_75t_L g5288 ( 
.A1(n_5204),
.A2(n_872),
.B1(n_870),
.B2(n_871),
.Y(n_5288)
);

AOI22xp5_ASAP7_75t_L g5289 ( 
.A1(n_5213),
.A2(n_872),
.B1(n_870),
.B2(n_871),
.Y(n_5289)
);

NOR2x1p5_ASAP7_75t_L g5290 ( 
.A(n_5225),
.B(n_873),
.Y(n_5290)
);

NOR2x1_ASAP7_75t_L g5291 ( 
.A(n_5188),
.B(n_874),
.Y(n_5291)
);

NOR2x1_ASAP7_75t_L g5292 ( 
.A(n_5251),
.B(n_874),
.Y(n_5292)
);

INVx1_ASAP7_75t_L g5293 ( 
.A(n_5212),
.Y(n_5293)
);

INVx3_ASAP7_75t_L g5294 ( 
.A(n_5235),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5230),
.Y(n_5295)
);

AOI22xp5_ASAP7_75t_L g5296 ( 
.A1(n_5222),
.A2(n_877),
.B1(n_875),
.B2(n_876),
.Y(n_5296)
);

INVx2_ASAP7_75t_L g5297 ( 
.A(n_5236),
.Y(n_5297)
);

INVx2_ASAP7_75t_L g5298 ( 
.A(n_5235),
.Y(n_5298)
);

NOR2x1_ASAP7_75t_L g5299 ( 
.A(n_5193),
.B(n_875),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_5211),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_SL g5301 ( 
.A(n_5226),
.B(n_877),
.Y(n_5301)
);

OAI22xp5_ASAP7_75t_SL g5302 ( 
.A1(n_5227),
.A2(n_880),
.B1(n_878),
.B2(n_879),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_5242),
.B(n_878),
.Y(n_5303)
);

NOR2xp67_ASAP7_75t_L g5304 ( 
.A(n_5202),
.B(n_880),
.Y(n_5304)
);

NAND2xp5_ASAP7_75t_SL g5305 ( 
.A(n_5244),
.B(n_881),
.Y(n_5305)
);

AOI22xp5_ASAP7_75t_L g5306 ( 
.A1(n_5217),
.A2(n_884),
.B1(n_882),
.B2(n_883),
.Y(n_5306)
);

NOR3xp33_ASAP7_75t_L g5307 ( 
.A(n_5206),
.B(n_884),
.C(n_885),
.Y(n_5307)
);

NOR2x1_ASAP7_75t_L g5308 ( 
.A(n_5186),
.B(n_885),
.Y(n_5308)
);

NOR4xp25_ASAP7_75t_L g5309 ( 
.A(n_5196),
.B(n_5208),
.C(n_5239),
.D(n_5209),
.Y(n_5309)
);

INVx1_ASAP7_75t_L g5310 ( 
.A(n_5262),
.Y(n_5310)
);

AOI221xp5_ASAP7_75t_L g5311 ( 
.A1(n_5295),
.A2(n_5240),
.B1(n_5246),
.B2(n_5241),
.C(n_5243),
.Y(n_5311)
);

INVx1_ASAP7_75t_L g5312 ( 
.A(n_5262),
.Y(n_5312)
);

INVx2_ASAP7_75t_L g5313 ( 
.A(n_5275),
.Y(n_5313)
);

CKINVDCx5p33_ASAP7_75t_R g5314 ( 
.A(n_5267),
.Y(n_5314)
);

OAI211xp5_ASAP7_75t_SL g5315 ( 
.A1(n_5273),
.A2(n_5214),
.B(n_5194),
.C(n_5238),
.Y(n_5315)
);

INVx1_ASAP7_75t_L g5316 ( 
.A(n_5275),
.Y(n_5316)
);

A2O1A1Ixp33_ASAP7_75t_SL g5317 ( 
.A1(n_5270),
.A2(n_5215),
.B(n_5224),
.C(n_5223),
.Y(n_5317)
);

A2O1A1Ixp33_ASAP7_75t_L g5318 ( 
.A1(n_5259),
.A2(n_5220),
.B(n_5232),
.C(n_5237),
.Y(n_5318)
);

AOI22x1_ASAP7_75t_L g5319 ( 
.A1(n_5261),
.A2(n_5249),
.B1(n_5248),
.B2(n_5245),
.Y(n_5319)
);

AO22x2_ASAP7_75t_L g5320 ( 
.A1(n_5256),
.A2(n_889),
.B1(n_886),
.B2(n_887),
.Y(n_5320)
);

OAI21xp5_ASAP7_75t_SL g5321 ( 
.A1(n_5281),
.A2(n_886),
.B(n_887),
.Y(n_5321)
);

INVx2_ASAP7_75t_SL g5322 ( 
.A(n_5269),
.Y(n_5322)
);

INVx1_ASAP7_75t_L g5323 ( 
.A(n_5255),
.Y(n_5323)
);

NAND4xp75_ASAP7_75t_L g5324 ( 
.A(n_5279),
.B(n_892),
.C(n_890),
.D(n_891),
.Y(n_5324)
);

NOR2x1_ASAP7_75t_L g5325 ( 
.A(n_5265),
.B(n_893),
.Y(n_5325)
);

OAI21xp5_ASAP7_75t_L g5326 ( 
.A1(n_5299),
.A2(n_895),
.B(n_896),
.Y(n_5326)
);

BUFx2_ASAP7_75t_L g5327 ( 
.A(n_5282),
.Y(n_5327)
);

INVx1_ASAP7_75t_L g5328 ( 
.A(n_5302),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_L g5329 ( 
.A(n_5266),
.B(n_895),
.Y(n_5329)
);

CKINVDCx16_ASAP7_75t_R g5330 ( 
.A(n_5309),
.Y(n_5330)
);

NOR2xp33_ASAP7_75t_R g5331 ( 
.A(n_5260),
.B(n_896),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_5288),
.B(n_897),
.Y(n_5332)
);

NOR2x1_ASAP7_75t_L g5333 ( 
.A(n_5254),
.B(n_898),
.Y(n_5333)
);

OAI22xp5_ASAP7_75t_L g5334 ( 
.A1(n_5258),
.A2(n_5268),
.B1(n_5271),
.B2(n_5293),
.Y(n_5334)
);

AOI221xp5_ASAP7_75t_L g5335 ( 
.A1(n_5287),
.A2(n_5276),
.B1(n_5280),
.B2(n_5297),
.C(n_5301),
.Y(n_5335)
);

AOI22xp5_ASAP7_75t_L g5336 ( 
.A1(n_5284),
.A2(n_901),
.B1(n_898),
.B2(n_899),
.Y(n_5336)
);

AOI311xp33_ASAP7_75t_L g5337 ( 
.A1(n_5300),
.A2(n_903),
.A3(n_901),
.B(n_902),
.C(n_904),
.Y(n_5337)
);

XNOR2x2_ASAP7_75t_SL g5338 ( 
.A(n_5306),
.B(n_902),
.Y(n_5338)
);

NOR2xp33_ASAP7_75t_L g5339 ( 
.A(n_5294),
.B(n_5303),
.Y(n_5339)
);

AOI22xp5_ASAP7_75t_L g5340 ( 
.A1(n_5277),
.A2(n_906),
.B1(n_903),
.B2(n_905),
.Y(n_5340)
);

BUFx2_ASAP7_75t_L g5341 ( 
.A(n_5294),
.Y(n_5341)
);

CKINVDCx5p33_ASAP7_75t_R g5342 ( 
.A(n_5298),
.Y(n_5342)
);

NOR2x1p5_ASAP7_75t_L g5343 ( 
.A(n_5272),
.B(n_905),
.Y(n_5343)
);

NAND2xp5_ASAP7_75t_L g5344 ( 
.A(n_5304),
.B(n_906),
.Y(n_5344)
);

INVx2_ASAP7_75t_L g5345 ( 
.A(n_5320),
.Y(n_5345)
);

NOR2x1_ASAP7_75t_L g5346 ( 
.A(n_5323),
.B(n_5278),
.Y(n_5346)
);

AND2x4_ASAP7_75t_L g5347 ( 
.A(n_5341),
.B(n_5308),
.Y(n_5347)
);

NOR2xp33_ASAP7_75t_L g5348 ( 
.A(n_5330),
.B(n_5286),
.Y(n_5348)
);

AOI22xp5_ASAP7_75t_L g5349 ( 
.A1(n_5335),
.A2(n_5290),
.B1(n_5292),
.B2(n_5291),
.Y(n_5349)
);

INVx1_ASAP7_75t_L g5350 ( 
.A(n_5320),
.Y(n_5350)
);

INVx1_ASAP7_75t_L g5351 ( 
.A(n_5314),
.Y(n_5351)
);

NOR2x1_ASAP7_75t_L g5352 ( 
.A(n_5324),
.B(n_5305),
.Y(n_5352)
);

NOR2xp67_ASAP7_75t_L g5353 ( 
.A(n_5340),
.B(n_5336),
.Y(n_5353)
);

INVx1_ASAP7_75t_L g5354 ( 
.A(n_5310),
.Y(n_5354)
);

AND2x2_ASAP7_75t_L g5355 ( 
.A(n_5337),
.B(n_5257),
.Y(n_5355)
);

NOR2x1_ASAP7_75t_L g5356 ( 
.A(n_5329),
.B(n_5264),
.Y(n_5356)
);

NAND4xp75_ASAP7_75t_L g5357 ( 
.A(n_5325),
.B(n_5285),
.C(n_5296),
.D(n_5283),
.Y(n_5357)
);

NOR2xp33_ASAP7_75t_L g5358 ( 
.A(n_5313),
.B(n_5263),
.Y(n_5358)
);

NAND4xp75_ASAP7_75t_L g5359 ( 
.A(n_5339),
.B(n_5333),
.C(n_5311),
.D(n_5326),
.Y(n_5359)
);

AOI22xp5_ASAP7_75t_L g5360 ( 
.A1(n_5334),
.A2(n_5307),
.B1(n_5289),
.B2(n_5274),
.Y(n_5360)
);

OAI211xp5_ASAP7_75t_L g5361 ( 
.A1(n_5332),
.A2(n_910),
.B(n_908),
.C(n_909),
.Y(n_5361)
);

HB1xp67_ASAP7_75t_L g5362 ( 
.A(n_5347),
.Y(n_5362)
);

NAND2xp5_ASAP7_75t_L g5363 ( 
.A(n_5347),
.B(n_5322),
.Y(n_5363)
);

AND2x2_ASAP7_75t_L g5364 ( 
.A(n_5355),
.B(n_5327),
.Y(n_5364)
);

HB1xp67_ASAP7_75t_L g5365 ( 
.A(n_5350),
.Y(n_5365)
);

AO22x2_ASAP7_75t_L g5366 ( 
.A1(n_5345),
.A2(n_5316),
.B1(n_5312),
.B2(n_5344),
.Y(n_5366)
);

OAI22xp5_ASAP7_75t_L g5367 ( 
.A1(n_5349),
.A2(n_5342),
.B1(n_5318),
.B2(n_5328),
.Y(n_5367)
);

O2A1O1Ixp33_ASAP7_75t_L g5368 ( 
.A1(n_5354),
.A2(n_5317),
.B(n_5321),
.C(n_5315),
.Y(n_5368)
);

INVx1_ASAP7_75t_L g5369 ( 
.A(n_5351),
.Y(n_5369)
);

AOI211xp5_ASAP7_75t_SL g5370 ( 
.A1(n_5348),
.A2(n_5338),
.B(n_5319),
.C(n_5331),
.Y(n_5370)
);

NOR4xp25_ASAP7_75t_L g5371 ( 
.A(n_5358),
.B(n_5343),
.C(n_910),
.D(n_908),
.Y(n_5371)
);

OAI221xp5_ASAP7_75t_SL g5372 ( 
.A1(n_5360),
.A2(n_5361),
.B1(n_5359),
.B2(n_5356),
.C(n_5346),
.Y(n_5372)
);

OR2x2_ASAP7_75t_L g5373 ( 
.A(n_5362),
.B(n_5357),
.Y(n_5373)
);

AND2x2_ASAP7_75t_L g5374 ( 
.A(n_5364),
.B(n_5352),
.Y(n_5374)
);

NOR2x1_ASAP7_75t_L g5375 ( 
.A(n_5363),
.B(n_5353),
.Y(n_5375)
);

NAND3xp33_ASAP7_75t_L g5376 ( 
.A(n_5370),
.B(n_909),
.C(n_911),
.Y(n_5376)
);

INVx1_ASAP7_75t_L g5377 ( 
.A(n_5365),
.Y(n_5377)
);

OAI21xp5_ASAP7_75t_L g5378 ( 
.A1(n_5369),
.A2(n_912),
.B(n_913),
.Y(n_5378)
);

XOR2x1_ASAP7_75t_SL g5379 ( 
.A(n_5366),
.B(n_912),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_5374),
.Y(n_5380)
);

CKINVDCx5p33_ASAP7_75t_R g5381 ( 
.A(n_5377),
.Y(n_5381)
);

OAI322xp33_ASAP7_75t_L g5382 ( 
.A1(n_5373),
.A2(n_5367),
.A3(n_5368),
.B1(n_5372),
.B2(n_5366),
.C1(n_5371),
.C2(n_916),
.Y(n_5382)
);

CKINVDCx20_ASAP7_75t_R g5383 ( 
.A(n_5379),
.Y(n_5383)
);

HB1xp67_ASAP7_75t_L g5384 ( 
.A(n_5375),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5384),
.Y(n_5385)
);

HB1xp67_ASAP7_75t_L g5386 ( 
.A(n_5380),
.Y(n_5386)
);

OR2x2_ASAP7_75t_L g5387 ( 
.A(n_5385),
.B(n_5381),
.Y(n_5387)
);

OAI22xp5_ASAP7_75t_L g5388 ( 
.A1(n_5387),
.A2(n_5386),
.B1(n_5383),
.B2(n_5376),
.Y(n_5388)
);

AND2x4_ASAP7_75t_L g5389 ( 
.A(n_5388),
.B(n_5378),
.Y(n_5389)
);

NAND2xp5_ASAP7_75t_L g5390 ( 
.A(n_5389),
.B(n_5382),
.Y(n_5390)
);

INVx4_ASAP7_75t_L g5391 ( 
.A(n_5390),
.Y(n_5391)
);

OAI21xp5_ASAP7_75t_SL g5392 ( 
.A1(n_5391),
.A2(n_914),
.B(n_915),
.Y(n_5392)
);

OAI22xp33_ASAP7_75t_L g5393 ( 
.A1(n_5392),
.A2(n_916),
.B1(n_914),
.B2(n_915),
.Y(n_5393)
);

NAND2xp5_ASAP7_75t_L g5394 ( 
.A(n_5393),
.B(n_917),
.Y(n_5394)
);

AOI21xp33_ASAP7_75t_L g5395 ( 
.A1(n_5394),
.A2(n_918),
.B(n_919),
.Y(n_5395)
);

AOI211xp5_ASAP7_75t_L g5396 ( 
.A1(n_5395),
.A2(n_920),
.B(n_918),
.C(n_919),
.Y(n_5396)
);


endmodule