module fake_jpeg_17884_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx6_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_39),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_15),
.B1(n_26),
.B2(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_53),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_15),
.B1(n_26),
.B2(n_23),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_26),
.B1(n_29),
.B2(n_23),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_59),
.B1(n_18),
.B2(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_37),
.A2(n_27),
.B1(n_24),
.B2(n_22),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_42),
.C(n_40),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_61),
.B(n_72),
.Y(n_114)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_63),
.B(n_71),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_69),
.B1(n_87),
.B2(n_16),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_66),
.B(n_68),
.Y(n_117)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_45),
.B(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_37),
.B1(n_17),
.B2(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_49),
.B(n_19),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_70),
.B(n_75),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_31),
.Y(n_72)
);

XNOR2x1_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_31),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_16),
.C(n_25),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_33),
.B1(n_24),
.B2(n_22),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_2),
.B(n_3),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_56),
.A2(n_50),
.B1(n_44),
.B2(n_54),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_33),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_83),
.B(n_96),
.Y(n_105)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_77),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_21),
.B1(n_19),
.B2(n_17),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_78),
.B(n_81),
.Y(n_111)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_89),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_31),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_57),
.B(n_21),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_88),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_86),
.Y(n_113)
);

OAI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_50),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_58),
.B(n_25),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_90),
.B(n_94),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_51),
.B(n_1),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_43),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_95),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_102),
.A2(n_91),
.B1(n_77),
.B2(n_28),
.Y(n_148)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_63),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_81),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_109),
.B(n_115),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_66),
.B(n_76),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_76),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_116),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_118),
.B(n_96),
.Y(n_126)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_119),
.Y(n_125)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_120),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_1),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_123),
.B(n_2),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_124),
.B(n_137),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_126),
.A2(n_133),
.B(n_144),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_141),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_128),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_61),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_129),
.B(n_132),
.C(n_143),
.Y(n_173)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_109),
.A2(n_68),
.A3(n_60),
.B1(n_83),
.B2(n_67),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_131),
.B(n_145),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_117),
.C(n_105),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_83),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_136),
.B(n_131),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_99),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_149),
.Y(n_160)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_85),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_65),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_142),
.B(n_146),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_65),
.C(n_60),
.Y(n_143)
);

AOI211xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_75),
.B(n_86),
.C(n_16),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_91),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_28),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_147),
.A2(n_110),
.B(n_112),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_148),
.A2(n_102),
.B1(n_104),
.B2(n_113),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_101),
.B(n_25),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_134),
.B(n_111),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_140),
.A2(n_107),
.B1(n_123),
.B2(n_113),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_155),
.B(n_170),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_159),
.A2(n_20),
.B(n_103),
.Y(n_185)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_168),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_121),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_166),
.B(n_167),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_100),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_100),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_171),
.Y(n_189)
);

NOR4xp25_ASAP7_75t_L g170 ( 
.A(n_136),
.B(n_120),
.C(n_119),
.D(n_106),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_143),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_106),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_145),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_144),
.A2(n_148),
.B1(n_126),
.B2(n_129),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_175),
.A2(n_28),
.B1(n_20),
.B2(n_92),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_178),
.B(n_155),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_175),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_163),
.B1(n_152),
.B2(n_158),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_147),
.C(n_103),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_181),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_135),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_156),
.Y(n_203)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_195),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_20),
.B1(n_4),
.B2(n_6),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_190),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_3),
.B1(n_6),
.B2(n_8),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_8),
.C(n_9),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_191),
.B(n_193),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_8),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_165),
.B(n_10),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_161),
.Y(n_195)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_150),
.CI(n_157),
.CON(n_198),
.SN(n_198)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_198),
.B(n_199),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_183),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_203),
.Y(n_214)
);

OAI322xp33_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_157),
.A3(n_164),
.B1(n_153),
.B2(n_152),
.C1(n_151),
.C2(n_169),
.Y(n_202)
);

OA21x2_ASAP7_75t_SL g215 ( 
.A1(n_202),
.A2(n_205),
.B(n_187),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_164),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_176),
.Y(n_225)
);

OAI21x1_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_156),
.B(n_163),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_194),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_209),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_215),
.A2(n_217),
.B(n_226),
.Y(n_234)
);

NOR2xp67_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_177),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_188),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_222),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_187),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_207),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_224),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_190),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_228),
.C(n_197),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_210),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_210),
.A2(n_177),
.B(n_176),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_182),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_197),
.B(n_180),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_232),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_220),
.A2(n_222),
.B(n_218),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_235),
.B(n_237),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_201),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_226),
.A2(n_210),
.B1(n_227),
.B2(n_216),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_233),
.A2(n_216),
.B1(n_185),
.B2(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_193),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_231),
.B(n_234),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_198),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_198),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_239),
.B(n_191),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_219),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_246),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_200),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_235),
.B(n_229),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_200),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_247),
.B(n_237),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_248),
.A2(n_242),
.B1(n_245),
.B2(n_240),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_240),
.C(n_11),
.Y(n_255)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_247),
.B(n_181),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_251),
.B(n_10),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_254),
.B(n_256),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_257),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_10),
.C(n_11),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_252),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_259),
.B(n_11),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_260),
.B(n_248),
.C(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_262),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_263),
.A2(n_258),
.B(n_13),
.Y(n_264)
);


endmodule