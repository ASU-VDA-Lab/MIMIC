module real_jpeg_2142_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_216;
wire n_167;
wire n_179;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_1),
.A2(n_53),
.B1(n_54),
.B2(n_65),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_1),
.A2(n_39),
.B1(n_46),
.B2(n_65),
.Y(n_159)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_34),
.Y(n_33)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_3),
.A2(n_33),
.B(n_34),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_3),
.B(n_100),
.Y(n_137)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_3),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_3),
.B(n_52),
.Y(n_170)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_3),
.A2(n_26),
.B(n_178),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_39),
.C(n_90),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_3),
.A2(n_53),
.B1(n_54),
.B2(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_3),
.B(n_42),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_3),
.B(n_94),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_4),
.A2(n_26),
.B1(n_27),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_4),
.A2(n_31),
.B1(n_34),
.B2(n_61),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_4),
.A2(n_53),
.B1(n_54),
.B2(n_61),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_4),
.A2(n_39),
.B1(n_46),
.B2(n_61),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_39),
.B1(n_46),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_6),
.A2(n_39),
.B1(n_46),
.B2(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_6),
.Y(n_84)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_9),
.A2(n_31),
.B1(n_34),
.B2(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_9),
.A2(n_26),
.B1(n_27),
.B2(n_72),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_72),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_9),
.A2(n_39),
.B1(n_46),
.B2(n_72),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_39),
.B1(n_46),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_11),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_11),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_93)
);

BUFx16f_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_13),
.A2(n_26),
.B1(n_27),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_13),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_104),
.Y(n_107)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_13),
.A2(n_39),
.B1(n_46),
.B2(n_104),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_14),
.A2(n_31),
.B1(n_34),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_14),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_14),
.A2(n_26),
.B1(n_27),
.B2(n_75),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_75),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_14),
.A2(n_39),
.B1(n_46),
.B2(n_75),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_39),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_16),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_16),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_124),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_111),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_111),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_76),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_50),
.C(n_66),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_24),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_25),
.B(n_37),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_29),
.A3(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_26),
.A2(n_27),
.B1(n_56),
.B2(n_58),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g70 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_36),
.Y(n_70)
);

OAI32xp33_ASAP7_75t_L g153 ( 
.A1(n_26),
.A2(n_54),
.A3(n_56),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_27),
.B(n_155),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_29),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_36),
.Y(n_69)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_38),
.A2(n_42),
.B1(n_80),
.B2(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_38),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_38),
.A2(n_42),
.B1(n_44),
.B2(n_140),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_38),
.A2(n_42),
.B1(n_159),
.B2(n_172),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_38),
.A2(n_42),
.B1(n_155),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_38),
.A2(n_42),
.B1(n_198),
.B2(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_39),
.A2(n_46),
.B1(n_90),
.B2(n_91),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_39),
.B(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_41),
.A2(n_48),
.B1(n_81),
.B2(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_41),
.A2(n_110),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_41),
.A2(n_110),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_50),
.B(n_66),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_50)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_51),
.A2(n_60),
.B1(n_62),
.B2(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_51),
.A2(n_62),
.B1(n_121),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_51),
.A2(n_62),
.B1(n_135),
.B2(n_177),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_59),
.Y(n_51)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_52),
.A2(n_64),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AO22x2_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_54),
.B1(n_90),
.B2(n_91),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_53),
.B(n_58),
.Y(n_156)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_54),
.B(n_186),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_73),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_67),
.A2(n_70),
.B1(n_71),
.B2(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_68),
.A2(n_74),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_96),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_85),
.B2(n_95),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_88),
.B1(n_93),
.B2(n_94),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_92),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_94),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_88),
.A2(n_94),
.B1(n_118),
.B2(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_88),
.A2(n_94),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_88),
.A2(n_94),
.B1(n_168),
.B2(n_189),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_92),
.A2(n_108),
.B1(n_151),
.B2(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_105),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_109),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.C(n_115),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_112),
.B(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_115),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_120),
.C(n_122),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_120),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_143),
.B(n_218),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_141),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_128),
.B(n_141),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_132),
.B(n_133),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.C(n_138),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_140),
.Y(n_160)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_163),
.B(n_217),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_161),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_146),
.B(n_161),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_152),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_147),
.B(n_214),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_152),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_153),
.B(n_157),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_154),
.Y(n_178)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_212),
.B(n_216),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_181),
.B(n_211),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_173),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_170),
.C(n_171),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_167),
.B(n_170),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_169),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_172),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_174),
.B(n_176),
.C(n_179),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_179),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_192),
.B(n_210),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_188),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_204),
.B(n_209),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_199),
.B(n_203),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_201),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_205),
.B(n_208),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_215),
.Y(n_216)
);


endmodule