module fake_jpeg_13103_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_13),
.Y(n_45)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_19),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

OA22x2_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_49)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_17),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_52),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_23),
.B1(n_28),
.B2(n_26),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_34),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_49),
.A2(n_36),
.B1(n_37),
.B2(n_35),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_56),
.B1(n_24),
.B2(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_58),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_62),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_43),
.B(n_22),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_65),
.B(n_68),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_52),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_29),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_45),
.B1(n_37),
.B2(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_67),
.A2(n_60),
.B1(n_53),
.B2(n_33),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_17),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_50),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_75),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_71),
.B(n_51),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_28),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_72),
.B(n_79),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_58),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_56),
.A2(n_32),
.B1(n_47),
.B2(n_29),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_77),
.B1(n_30),
.B2(n_69),
.Y(n_86)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_84),
.Y(n_94)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_20),
.A3(n_16),
.B1(n_14),
.B2(n_42),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g87 ( 
.A(n_83),
.B(n_59),
.CI(n_19),
.CON(n_87),
.SN(n_87)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_24),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_87),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_55),
.B(n_64),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_88),
.A2(n_90),
.B(n_91),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_84),
.A2(n_61),
.B1(n_18),
.B2(n_57),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_78),
.A2(n_63),
.B(n_16),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_72),
.C(n_77),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_14),
.Y(n_95)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_70),
.A2(n_32),
.B1(n_57),
.B2(n_20),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_97),
.A2(n_79),
.B1(n_74),
.B2(n_44),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_59),
.B(n_30),
.C(n_50),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_51),
.B(n_74),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_80),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_106),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_87),
.B(n_75),
.CON(n_101),
.SN(n_101)
);

NOR2x1_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_92),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_9),
.C(n_8),
.Y(n_102)
);

FAx1_ASAP7_75t_SL g110 ( 
.A(n_102),
.B(n_104),
.CI(n_7),
.CON(n_110),
.SN(n_110)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_89),
.Y(n_103)
);

INVxp67_ASAP7_75t_SL g111 ( 
.A(n_103),
.Y(n_111)
);

NOR4xp25_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_85),
.C(n_59),
.D(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_108),
.B(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_110),
.B(n_109),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_116),
.Y(n_118)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_106),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_114),
.A2(n_115),
.B1(n_117),
.B2(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_96),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_107),
.A2(n_90),
.B1(n_92),
.B2(n_98),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_116),
.B(n_99),
.C(n_105),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_122),
.C(n_123),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_110),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_99),
.C(n_105),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_101),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_119),
.B(n_113),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_124),
.A2(n_122),
.B(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_129),
.C(n_2),
.Y(n_133)
);

OAI31xp33_ASAP7_75t_L g129 ( 
.A1(n_126),
.A2(n_112),
.A3(n_118),
.B(n_110),
.Y(n_129)
);

CKINVDCx5p33_ASAP7_75t_R g131 ( 
.A(n_127),
.Y(n_131)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_131),
.A2(n_117),
.A3(n_98),
.B1(n_114),
.B2(n_115),
.C1(n_1),
.C2(n_4),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_133),
.C(n_130),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_135),
.C(n_3),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_3),
.C(n_4),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_5),
.Y(n_137)
);


endmodule