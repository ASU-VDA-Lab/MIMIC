module real_aes_9917_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_2036, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_2036;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_2003;
wire n_1279;
wire n_1314;
wire n_2014;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_2029;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_2006;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_2031;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1994;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1284;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_2004;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_1945;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_2012;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_1499;
wire n_700;
wire n_948;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_2033;
wire n_1769;
wire n_1812;
wire n_1985;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_2023;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_1409;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_2019;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1078;
wire n_1638;
wire n_495;
wire n_1072;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1986;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_2032;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_2027;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_2034;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_2028;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_1457;
wire n_719;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_2011;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_2030;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1049;
wire n_559;
wire n_1277;
wire n_1584;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_1916;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_2010;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_1430;
wire n_907;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1390 ( .A1(n_0), .A2(n_188), .B1(n_1391), .B2(n_1392), .C(n_1393), .Y(n_1390) );
AOI221xp5_ASAP7_75t_L g1424 ( .A1(n_0), .A2(n_372), .B1(n_676), .B2(n_678), .C(n_1425), .Y(n_1424) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_1), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_1), .A2(n_360), .B1(n_640), .B2(n_790), .Y(n_789) );
OA22x2_ASAP7_75t_L g1123 ( .A1(n_2), .A2(n_1124), .B1(n_1186), .B2(n_1187), .Y(n_1123) );
INVxp67_ASAP7_75t_SL g1187 ( .A(n_2), .Y(n_1187) );
AOI22xp5_ASAP7_75t_L g1714 ( .A1(n_3), .A2(n_364), .B1(n_1700), .B2(n_1703), .Y(n_1714) );
CKINVDCx5p33_ASAP7_75t_R g841 ( .A(n_4), .Y(n_841) );
INVx1_ASAP7_75t_L g842 ( .A(n_5), .Y(n_842) );
INVx1_ASAP7_75t_L g1574 ( .A(n_6), .Y(n_1574) );
INVxp33_ASAP7_75t_L g781 ( .A(n_7), .Y(n_781) );
AOI21xp33_ASAP7_75t_L g799 ( .A1(n_7), .A2(n_800), .B(n_801), .Y(n_799) );
INVx1_ASAP7_75t_L g1345 ( .A(n_8), .Y(n_1345) );
AOI221xp5_ASAP7_75t_SL g1365 ( .A1(n_8), .A2(n_145), .B1(n_635), .B2(n_1160), .C(n_1366), .Y(n_1365) );
INVx1_ASAP7_75t_L g764 ( .A(n_9), .Y(n_764) );
INVx1_ASAP7_75t_L g1339 ( .A(n_10), .Y(n_1339) );
AOI221xp5_ASAP7_75t_L g1373 ( .A1(n_10), .A2(n_250), .B1(n_1156), .B2(n_1374), .C(n_1375), .Y(n_1373) );
AOI221xp5_ASAP7_75t_L g821 ( .A1(n_11), .A2(n_106), .B1(n_822), .B2(n_823), .C(n_824), .Y(n_821) );
INVx1_ASAP7_75t_L g848 ( .A(n_11), .Y(n_848) );
AOI22xp33_ASAP7_75t_SL g1293 ( .A1(n_12), .A2(n_170), .B1(n_463), .B2(n_1294), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_12), .A2(n_65), .B1(n_623), .B2(n_925), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_13), .A2(n_316), .B1(n_593), .B2(n_595), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_13), .A2(n_346), .B1(n_638), .B2(n_640), .Y(n_637) );
XNOR2x2_ASAP7_75t_L g1286 ( .A(n_14), .B(n_1287), .Y(n_1286) );
INVxp33_ASAP7_75t_L g779 ( .A(n_15), .Y(n_779) );
NAND2xp33_ASAP7_75t_SL g797 ( .A(n_15), .B(n_798), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g1500 ( .A(n_16), .Y(n_1500) );
CKINVDCx20_ASAP7_75t_R g1935 ( .A(n_17), .Y(n_1935) );
AOI22xp5_ASAP7_75t_L g1715 ( .A1(n_18), .A2(n_310), .B1(n_1693), .B2(n_1711), .Y(n_1715) );
AOI22xp33_ASAP7_75t_SL g1296 ( .A1(n_19), .A2(n_65), .B1(n_1115), .B2(n_1297), .Y(n_1296) );
AOI21xp33_ASAP7_75t_L g1318 ( .A1(n_19), .A2(n_554), .B(n_1099), .Y(n_1318) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_20), .A2(n_262), .B1(n_1127), .B2(n_1128), .Y(n_1126) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_20), .Y(n_1181) );
CKINVDCx5p33_ASAP7_75t_R g1083 ( .A(n_21), .Y(n_1083) );
INVxp67_ASAP7_75t_L g1451 ( .A(n_22), .Y(n_1451) );
AOI221xp5_ASAP7_75t_L g1472 ( .A1(n_22), .A2(n_69), .B1(n_635), .B2(n_675), .C(n_788), .Y(n_1472) );
CKINVDCx16_ASAP7_75t_R g1691 ( .A(n_23), .Y(n_1691) );
XNOR2xp5_ASAP7_75t_L g1906 ( .A(n_23), .B(n_1907), .Y(n_1906) );
AOI22xp33_ASAP7_75t_L g1974 ( .A1(n_23), .A2(n_1975), .B1(n_1978), .B2(n_2029), .Y(n_1974) );
INVxp33_ASAP7_75t_L g1582 ( .A(n_24), .Y(n_1582) );
AOI221xp5_ASAP7_75t_L g1629 ( .A1(n_24), .A2(n_89), .B1(n_474), .B2(n_1630), .C(n_1631), .Y(n_1629) );
OAI221xp5_ASAP7_75t_L g1024 ( .A1(n_25), .A2(n_78), .B1(n_1025), .B2(n_1027), .C(n_1028), .Y(n_1024) );
INVx1_ASAP7_75t_L g1062 ( .A(n_25), .Y(n_1062) );
INVx1_ASAP7_75t_L g1310 ( .A(n_26), .Y(n_1310) );
AOI22xp33_ASAP7_75t_L g1320 ( .A1(n_26), .A2(n_325), .B1(n_925), .B2(n_1099), .Y(n_1320) );
OAI221xp5_ASAP7_75t_L g774 ( .A1(n_27), .A2(n_340), .B1(n_722), .B2(n_731), .C(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g802 ( .A(n_27), .Y(n_802) );
OAI22xp5_ASAP7_75t_L g1987 ( .A1(n_28), .A2(n_362), .B1(n_511), .B2(n_659), .Y(n_1987) );
INVxp67_ASAP7_75t_SL g2028 ( .A(n_28), .Y(n_2028) );
INVx1_ASAP7_75t_L g895 ( .A(n_29), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_29), .A2(n_63), .B1(n_945), .B2(n_947), .Y(n_944) );
OAI221xp5_ASAP7_75t_L g1448 ( .A1(n_30), .A2(n_132), .B1(n_722), .B2(n_775), .C(n_855), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1469 ( .A1(n_30), .A2(n_132), .B1(n_615), .B2(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g646 ( .A(n_31), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_32), .A2(n_182), .B1(n_595), .B2(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g628 ( .A(n_32), .Y(n_628) );
INVxp33_ASAP7_75t_L g884 ( .A(n_33), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g923 ( .A1(n_33), .A2(n_91), .B1(n_924), .B2(n_925), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1603 ( .A1(n_34), .A2(n_359), .B1(n_795), .B2(n_1604), .Y(n_1603) );
INVxp67_ASAP7_75t_SL g1642 ( .A(n_34), .Y(n_1642) );
AOI221xp5_ASAP7_75t_L g833 ( .A1(n_35), .A2(n_252), .B1(n_635), .B2(n_788), .C(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g862 ( .A(n_35), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g1481 ( .A(n_36), .Y(n_1481) );
INVx1_ASAP7_75t_L g1043 ( .A(n_37), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1340 ( .A1(n_38), .A2(n_329), .B1(n_722), .B2(n_727), .C(n_731), .Y(n_1340) );
OAI22xp5_ASAP7_75t_L g1372 ( .A1(n_38), .A2(n_329), .B1(n_1166), .B2(n_1167), .Y(n_1372) );
INVx1_ASAP7_75t_L g381 ( .A(n_39), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g1699 ( .A1(n_40), .A2(n_176), .B1(n_1700), .B2(n_1703), .Y(n_1699) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_41), .A2(n_333), .B1(n_466), .B2(n_468), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g546 ( .A1(n_41), .A2(n_166), .B1(n_547), .B2(n_549), .C(n_554), .Y(n_546) );
OAI221xp5_ASAP7_75t_L g890 ( .A1(n_42), .A2(n_215), .B1(n_727), .B2(n_732), .C(n_891), .Y(n_890) );
OAI33xp33_ASAP7_75t_L g932 ( .A1(n_42), .A2(n_215), .A3(n_566), .B1(n_933), .B2(n_934), .B3(n_2036), .Y(n_932) );
INVx1_ASAP7_75t_L g1484 ( .A(n_43), .Y(n_1484) );
AOI221xp5_ASAP7_75t_L g1506 ( .A1(n_43), .A2(n_200), .B1(n_662), .B2(n_1507), .C(n_1509), .Y(n_1506) );
OAI221xp5_ASAP7_75t_L g1132 ( .A1(n_44), .A2(n_79), .B1(n_727), .B2(n_731), .C(n_891), .Y(n_1132) );
OAI222xp33_ASAP7_75t_L g1165 ( .A1(n_44), .A2(n_79), .B1(n_246), .B2(n_1042), .C1(n_1166), .C2(n_1167), .Y(n_1165) );
INVx1_ASAP7_75t_L g771 ( .A(n_45), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g1795 ( .A1(n_46), .A2(n_243), .B1(n_1687), .B2(n_1754), .Y(n_1795) );
AOI21xp33_ASAP7_75t_L g1093 ( .A1(n_47), .A2(n_547), .B(n_941), .Y(n_1093) );
AOI221xp5_ASAP7_75t_L g1117 ( .A1(n_47), .A2(n_98), .B1(n_449), .B2(n_470), .C(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1991 ( .A(n_48), .Y(n_1991) );
OAI221xp5_ASAP7_75t_L g2008 ( .A1(n_48), .A2(n_319), .B1(n_1391), .B2(n_2009), .C(n_2010), .Y(n_2008) );
INVx1_ASAP7_75t_L g1589 ( .A(n_49), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_50), .A2(n_356), .B1(n_444), .B2(n_1544), .Y(n_1543) );
OAI22xp5_ASAP7_75t_L g1563 ( .A1(n_50), .A2(n_270), .B1(n_1078), .B2(n_1564), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g1358 ( .A(n_51), .Y(n_1358) );
INVxp33_ASAP7_75t_SL g588 ( .A(n_52), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_52), .A2(n_167), .B1(n_620), .B2(n_621), .Y(n_619) );
OAI222xp33_ASAP7_75t_L g1257 ( .A1(n_53), .A2(n_191), .B1(n_296), .B2(n_1258), .C1(n_1260), .C2(n_1261), .Y(n_1257) );
AOI221xp5_ASAP7_75t_L g1281 ( .A1(n_53), .A2(n_191), .B1(n_1282), .B2(n_1283), .C(n_1284), .Y(n_1281) );
AOI22xp5_ASAP7_75t_L g1709 ( .A1(n_54), .A2(n_140), .B1(n_1700), .B2(n_1703), .Y(n_1709) );
AO221x2_ASAP7_75t_L g1717 ( .A1(n_55), .A2(n_272), .B1(n_1693), .B2(n_1711), .C(n_1718), .Y(n_1717) );
CKINVDCx16_ASAP7_75t_R g1694 ( .A(n_56), .Y(n_1694) );
INVx1_ASAP7_75t_L g500 ( .A(n_57), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_58), .A2(n_346), .B1(n_472), .B2(n_597), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_58), .A2(n_316), .B1(n_630), .B2(n_632), .C(n_635), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g674 ( .A1(n_59), .A2(n_187), .B1(n_635), .B2(n_675), .C(n_676), .Y(n_674) );
INVxp33_ASAP7_75t_SL g706 ( .A(n_59), .Y(n_706) );
CKINVDCx5p33_ASAP7_75t_R g1291 ( .A(n_60), .Y(n_1291) );
INVx1_ASAP7_75t_L g656 ( .A(n_61), .Y(n_656) );
AOI22xp5_ASAP7_75t_SL g1731 ( .A1(n_62), .A2(n_259), .B1(n_1687), .B2(n_1693), .Y(n_1731) );
INVx1_ASAP7_75t_L g899 ( .A(n_63), .Y(n_899) );
OAI221xp5_ASAP7_75t_L g1397 ( .A1(n_64), .A2(n_122), .B1(n_732), .B2(n_891), .C(n_1398), .Y(n_1397) );
OAI221xp5_ASAP7_75t_SL g1421 ( .A1(n_64), .A2(n_122), .B1(n_1166), .B2(n_1167), .C(n_1422), .Y(n_1421) );
INVx1_ASAP7_75t_L g908 ( .A(n_66), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g1144 ( .A(n_67), .Y(n_1144) );
XOR2xp5_ASAP7_75t_L g650 ( .A(n_68), .B(n_651), .Y(n_650) );
INVxp33_ASAP7_75t_L g1455 ( .A(n_69), .Y(n_1455) );
AOI22xp33_ASAP7_75t_L g1606 ( .A1(n_70), .A2(n_227), .B1(n_1251), .B2(n_1607), .Y(n_1606) );
OAI22xp5_ASAP7_75t_L g1654 ( .A1(n_70), .A2(n_227), .B1(n_1655), .B2(n_1657), .Y(n_1654) );
INVx1_ASAP7_75t_L g1536 ( .A(n_71), .Y(n_1536) );
INVx1_ASAP7_75t_L g1953 ( .A(n_72), .Y(n_1953) );
OAI22xp33_ASAP7_75t_L g1962 ( .A1(n_72), .A2(n_135), .B1(n_1586), .B2(n_1963), .Y(n_1962) );
AOI22xp33_ASAP7_75t_L g1919 ( .A1(n_73), .A2(n_373), .B1(n_1920), .B2(n_1921), .Y(n_1919) );
INVx1_ASAP7_75t_L g1940 ( .A(n_73), .Y(n_1940) );
AOI22xp33_ASAP7_75t_L g1538 ( .A1(n_74), .A2(n_169), .B1(n_1054), .B2(n_1539), .Y(n_1538) );
AOI221xp5_ASAP7_75t_L g1547 ( .A1(n_74), .A2(n_239), .B1(n_521), .B2(n_1548), .C(n_1550), .Y(n_1547) );
CKINVDCx14_ASAP7_75t_R g1759 ( .A(n_75), .Y(n_1759) );
AOI22xp33_ASAP7_75t_L g2000 ( .A1(n_76), .A2(n_231), .B1(n_1433), .B2(n_1989), .Y(n_2000) );
AOI22xp33_ASAP7_75t_L g2017 ( .A1(n_76), .A2(n_231), .B1(n_2018), .B2(n_2020), .Y(n_2017) );
OAI221xp5_ASAP7_75t_L g1085 ( .A1(n_77), .A2(n_150), .B1(n_934), .B2(n_1081), .C(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1122 ( .A(n_77), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1057 ( .A1(n_78), .A2(n_232), .B1(n_1058), .B2(n_1060), .C(n_1061), .Y(n_1057) );
INVx1_ASAP7_75t_L g879 ( .A(n_80), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g1497 ( .A(n_81), .Y(n_1497) );
CKINVDCx5p33_ASAP7_75t_R g1141 ( .A(n_82), .Y(n_1141) );
AOI21xp33_ASAP7_75t_L g971 ( .A1(n_83), .A2(n_972), .B(n_973), .Y(n_971) );
INVxp33_ASAP7_75t_L g999 ( .A(n_83), .Y(n_999) );
AOI22xp33_ASAP7_75t_L g1211 ( .A1(n_84), .A2(n_226), .B1(n_1212), .B2(n_1214), .Y(n_1211) );
INVxp67_ASAP7_75t_SL g1232 ( .A(n_84), .Y(n_1232) );
XOR2x2_ASAP7_75t_L g1569 ( .A(n_85), .B(n_1570), .Y(n_1569) );
OAI22xp33_ASAP7_75t_L g829 ( .A1(n_86), .A2(n_237), .B1(n_830), .B2(n_831), .Y(n_829) );
OAI221xp5_ASAP7_75t_L g853 ( .A1(n_86), .A2(n_237), .B1(n_727), .B2(n_854), .C(n_855), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1793 ( .A1(n_87), .A2(n_236), .B1(n_1700), .B2(n_1794), .Y(n_1793) );
INVxp33_ASAP7_75t_L g887 ( .A(n_88), .Y(n_887) );
AOI21xp33_ASAP7_75t_L g926 ( .A1(n_88), .A2(n_824), .B(n_927), .Y(n_926) );
INVxp33_ASAP7_75t_L g1584 ( .A(n_89), .Y(n_1584) );
INVx1_ASAP7_75t_L g1217 ( .A(n_90), .Y(n_1217) );
INVxp33_ASAP7_75t_L g888 ( .A(n_91), .Y(n_888) );
INVx1_ASAP7_75t_L g1531 ( .A(n_92), .Y(n_1531) );
CKINVDCx20_ASAP7_75t_R g966 ( .A(n_93), .Y(n_966) );
CKINVDCx5p33_ASAP7_75t_R g1308 ( .A(n_94), .Y(n_1308) );
INVxp33_ASAP7_75t_L g1447 ( .A(n_95), .Y(n_1447) );
AOI22xp33_ASAP7_75t_L g1467 ( .A1(n_95), .A2(n_374), .B1(n_640), .B2(n_1468), .Y(n_1467) );
CKINVDCx5p33_ASAP7_75t_R g1917 ( .A(n_96), .Y(n_1917) );
AOI22xp33_ASAP7_75t_L g1299 ( .A1(n_97), .A2(n_195), .B1(n_467), .B2(n_470), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g1326 ( .A1(n_97), .A2(n_195), .B1(n_561), .B2(n_1327), .Y(n_1326) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_98), .A2(n_257), .B1(n_925), .B2(n_946), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_99), .A2(n_194), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1069 ( .A(n_99), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g471 ( .A1(n_100), .A2(n_111), .B1(n_466), .B2(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g572 ( .A(n_100), .Y(n_572) );
INVxp33_ASAP7_75t_SL g2004 ( .A(n_101), .Y(n_2004) );
AOI22xp33_ASAP7_75t_L g2024 ( .A1(n_101), .A2(n_361), .B1(n_2020), .B2(n_2022), .Y(n_2024) );
OAI221xp5_ASAP7_75t_L g1485 ( .A1(n_102), .A2(n_178), .B1(n_775), .B2(n_891), .C(n_1002), .Y(n_1485) );
OAI22xp33_ASAP7_75t_L g1505 ( .A1(n_102), .A2(n_178), .B1(n_511), .B2(n_516), .Y(n_1505) );
CKINVDCx14_ASAP7_75t_R g1719 ( .A(n_103), .Y(n_1719) );
CKINVDCx5p33_ASAP7_75t_R g1360 ( .A(n_104), .Y(n_1360) );
OR2x2_ASAP7_75t_L g414 ( .A(n_105), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g435 ( .A(n_105), .Y(n_435) );
BUFx2_ASAP7_75t_L g458 ( .A(n_105), .Y(n_458) );
BUFx2_ASAP7_75t_L g488 ( .A(n_105), .Y(n_488) );
INVx1_ASAP7_75t_L g850 ( .A(n_106), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g1300 ( .A1(n_107), .A2(n_120), .B1(n_463), .B2(n_1294), .Y(n_1300) );
INVx1_ASAP7_75t_L g1325 ( .A(n_107), .Y(n_1325) );
CKINVDCx5p33_ASAP7_75t_R g963 ( .A(n_108), .Y(n_963) );
AOI221xp5_ASAP7_75t_L g977 ( .A1(n_109), .A2(n_248), .B1(n_978), .B2(n_980), .C(n_983), .Y(n_977) );
INVxp67_ASAP7_75t_SL g1010 ( .A(n_109), .Y(n_1010) );
INVx1_ASAP7_75t_L g1349 ( .A(n_110), .Y(n_1349) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_110), .A2(n_298), .B1(n_1369), .B2(n_1370), .Y(n_1368) );
INVx1_ASAP7_75t_L g509 ( .A(n_111), .Y(n_509) );
AOI221xp5_ASAP7_75t_SL g1034 ( .A1(n_112), .A2(n_117), .B1(n_630), .B2(n_800), .C(n_973), .Y(n_1034) );
INVx1_ASAP7_75t_L g1053 ( .A(n_112), .Y(n_1053) );
INVx1_ASAP7_75t_L g1030 ( .A(n_113), .Y(n_1030) );
AOI221xp5_ASAP7_75t_L g1199 ( .A1(n_114), .A2(n_138), .B1(n_560), .B2(n_1200), .C(n_1201), .Y(n_1199) );
INVxp33_ASAP7_75t_L g1222 ( .A(n_114), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1475 ( .A1(n_115), .A2(n_1476), .B1(n_1517), .B2(n_1518), .Y(n_1475) );
INVx1_ASAP7_75t_L g1517 ( .A(n_115), .Y(n_1517) );
INVx1_ASAP7_75t_L g1408 ( .A(n_116), .Y(n_1408) );
INVx1_ASAP7_75t_L g1052 ( .A(n_117), .Y(n_1052) );
XOR2x2_ASAP7_75t_L g1073 ( .A(n_118), .B(n_1074), .Y(n_1073) );
INVxp67_ASAP7_75t_SL g902 ( .A(n_119), .Y(n_902) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_119), .A2(n_327), .B1(n_937), .B2(n_939), .C(n_941), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g1313 ( .A(n_120), .B(n_571), .Y(n_1313) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_121), .A2(n_246), .B1(n_485), .B2(n_1130), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g1179 ( .A(n_121), .Y(n_1179) );
OA22x2_ASAP7_75t_L g1190 ( .A1(n_123), .A2(n_1191), .B1(n_1192), .B2(n_1241), .Y(n_1190) );
CKINVDCx16_ASAP7_75t_R g1241 ( .A(n_123), .Y(n_1241) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_124), .Y(n_1356) );
CKINVDCx5p33_ASAP7_75t_R g1418 ( .A(n_125), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g1098 ( .A1(n_126), .A2(n_286), .B1(n_621), .B2(n_1099), .Y(n_1098) );
OAI211xp5_ASAP7_75t_L g1101 ( .A1(n_126), .A2(n_1102), .B(n_1104), .C(n_1106), .Y(n_1101) );
OAI22xp33_ASAP7_75t_L g1932 ( .A1(n_127), .A2(n_225), .B1(n_1597), .B2(n_1933), .Y(n_1932) );
INVx1_ASAP7_75t_L g1960 ( .A(n_127), .Y(n_1960) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_128), .A2(n_199), .B1(n_658), .B2(n_659), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g721 ( .A1(n_128), .A2(n_199), .B1(n_722), .B2(n_727), .C(n_731), .Y(n_721) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_129), .Y(n_820) );
AOI221xp5_ASAP7_75t_L g1037 ( .A1(n_130), .A2(n_204), .B1(n_635), .B2(n_675), .C(n_676), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g1064 ( .A1(n_130), .A2(n_194), .B1(n_1065), .B2(n_1067), .C(n_1068), .Y(n_1064) );
XNOR2x1_ASAP7_75t_L g1438 ( .A(n_131), .B(n_1439), .Y(n_1438) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_133), .A2(n_357), .B1(n_597), .B2(n_599), .Y(n_598) );
INVxp33_ASAP7_75t_L g645 ( .A(n_133), .Y(n_645) );
INVx1_ASAP7_75t_L g1561 ( .A(n_134), .Y(n_1561) );
AOI221xp5_ASAP7_75t_L g1954 ( .A1(n_135), .A2(n_315), .B1(n_474), .B2(n_1955), .C(n_1956), .Y(n_1954) );
CKINVDCx5p33_ASAP7_75t_R g1362 ( .A(n_136), .Y(n_1362) );
CKINVDCx5p33_ASAP7_75t_R g1499 ( .A(n_137), .Y(n_1499) );
INVxp33_ASAP7_75t_L g1224 ( .A(n_138), .Y(n_1224) );
OAI222xp33_ASAP7_75t_L g1262 ( .A1(n_139), .A2(n_218), .B1(n_354), .B2(n_831), .C1(n_1042), .C2(n_1263), .Y(n_1262) );
INVx1_ASAP7_75t_L g1274 ( .A(n_139), .Y(n_1274) );
OAI22xp33_ASAP7_75t_L g1080 ( .A1(n_141), .A2(n_337), .B1(n_682), .B2(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1116 ( .A1(n_141), .A2(n_203), .B1(n_475), .B2(n_594), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1100 ( .A1(n_142), .A2(n_824), .B(n_927), .Y(n_1100) );
INVx1_ASAP7_75t_L g1107 ( .A(n_142), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1077 ( .A1(n_143), .A2(n_203), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_143), .A2(n_337), .B1(n_431), .B2(n_1115), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_144), .Y(n_816) );
INVx1_ASAP7_75t_L g1348 ( .A(n_145), .Y(n_1348) );
AOI221xp5_ASAP7_75t_L g1997 ( .A1(n_146), .A2(n_328), .B1(n_675), .B2(n_1998), .C(n_1999), .Y(n_1997) );
AOI22xp33_ASAP7_75t_L g2021 ( .A1(n_146), .A2(n_328), .B1(n_2022), .B2(n_2023), .Y(n_2021) );
INVx1_ASAP7_75t_L g1533 ( .A(n_147), .Y(n_1533) );
INVx1_ASAP7_75t_L g1948 ( .A(n_148), .Y(n_1948) );
OAI22xp33_ASAP7_75t_L g1964 ( .A1(n_148), .A2(n_315), .B1(n_1965), .B2(n_1967), .Y(n_1964) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_149), .Y(n_1089) );
INVx1_ASAP7_75t_L g1105 ( .A(n_150), .Y(n_1105) );
INVx1_ASAP7_75t_L g1032 ( .A(n_151), .Y(n_1032) );
INVx1_ASAP7_75t_L g669 ( .A(n_152), .Y(n_669) );
AOI22xp5_ASAP7_75t_SL g1730 ( .A1(n_153), .A2(n_184), .B1(n_1700), .B2(n_1703), .Y(n_1730) );
CKINVDCx5p33_ASAP7_75t_R g1150 ( .A(n_154), .Y(n_1150) );
AOI221xp5_ASAP7_75t_L g1252 ( .A1(n_155), .A2(n_326), .B1(n_554), .B2(n_788), .C(n_1253), .Y(n_1252) );
INVx1_ASAP7_75t_L g1280 ( .A(n_155), .Y(n_1280) );
INVx1_ASAP7_75t_L g1387 ( .A(n_156), .Y(n_1387) );
CKINVDCx5p33_ASAP7_75t_R g1502 ( .A(n_157), .Y(n_1502) );
INVx1_ASAP7_75t_L g1458 ( .A(n_158), .Y(n_1458) );
INVx1_ASAP7_75t_L g1677 ( .A(n_159), .Y(n_1677) );
INVxp33_ASAP7_75t_SL g2003 ( .A(n_160), .Y(n_2003) );
AOI22xp33_ASAP7_75t_L g2025 ( .A1(n_160), .A2(n_306), .B1(n_2018), .B2(n_2023), .Y(n_2025) );
INVx1_ASAP7_75t_L g420 ( .A(n_161), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_161), .A2(n_283), .B1(n_511), .B2(n_516), .Y(n_510) );
XNOR2x1_ASAP7_75t_L g576 ( .A(n_162), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g1208 ( .A(n_163), .Y(n_1208) );
INVx1_ASAP7_75t_L g685 ( .A(n_164), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g916 ( .A(n_165), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_166), .A2(n_331), .B1(n_461), .B2(n_463), .Y(n_460) );
INVxp33_ASAP7_75t_SL g583 ( .A(n_167), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g1209 ( .A1(n_168), .A2(n_242), .B1(n_547), .B2(n_939), .C(n_1210), .Y(n_1209) );
INVxp67_ASAP7_75t_SL g1237 ( .A(n_168), .Y(n_1237) );
INVx1_ASAP7_75t_L g1552 ( .A(n_169), .Y(n_1552) );
INVx1_ASAP7_75t_L g1316 ( .A(n_170), .Y(n_1316) );
XOR2x1_ASAP7_75t_L g403 ( .A(n_171), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g885 ( .A(n_172), .Y(n_885) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_172), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g1411 ( .A(n_173), .Y(n_1411) );
CKINVDCx16_ASAP7_75t_R g1684 ( .A(n_174), .Y(n_1684) );
INVx1_ASAP7_75t_L g1595 ( .A(n_175), .Y(n_1595) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_177), .A2(n_219), .B1(n_662), .B2(n_664), .C(n_666), .Y(n_661) );
INVxp33_ASAP7_75t_L g735 ( .A(n_177), .Y(n_735) );
INVx1_ASAP7_75t_L g1460 ( .A(n_179), .Y(n_1460) );
INVx1_ASAP7_75t_L g1678 ( .A(n_180), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1683 ( .A(n_180), .B(n_1676), .Y(n_1683) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_181), .A2(n_266), .B1(n_525), .B2(n_662), .Y(n_1035) );
OAI221xp5_ASAP7_75t_L g1048 ( .A1(n_181), .A2(n_266), .B1(n_1049), .B2(n_1050), .C(n_1051), .Y(n_1048) );
INVxp33_ASAP7_75t_L g644 ( .A(n_182), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g1601 ( .A1(n_183), .A2(n_213), .B1(n_1200), .B2(n_1602), .Y(n_1601) );
INVxp67_ASAP7_75t_SL g1641 ( .A(n_183), .Y(n_1641) );
INVx1_ASAP7_75t_L g773 ( .A(n_185), .Y(n_773) );
INVx2_ASAP7_75t_L g393 ( .A(n_186), .Y(n_393) );
INVxp67_ASAP7_75t_L g693 ( .A(n_187), .Y(n_693) );
INVx1_ASAP7_75t_L g1423 ( .A(n_188), .Y(n_1423) );
AOI22xp33_ASAP7_75t_L g1929 ( .A1(n_189), .A2(n_370), .B1(n_640), .B2(n_1930), .Y(n_1929) );
OAI22xp5_ASAP7_75t_L g1937 ( .A1(n_189), .A2(n_370), .B1(n_1655), .B2(n_1657), .Y(n_1937) );
BUFx3_ASAP7_75t_L g497 ( .A(n_190), .Y(n_497) );
INVx1_ASAP7_75t_L g524 ( .A(n_190), .Y(n_524) );
INVx1_ASAP7_75t_L g1488 ( .A(n_192), .Y(n_1488) );
AOI22xp33_ASAP7_75t_L g1514 ( .A1(n_192), .A2(n_309), .B1(n_795), .B2(n_945), .Y(n_1514) );
INVx1_ASAP7_75t_L g1578 ( .A(n_193), .Y(n_1578) );
INVx1_ASAP7_75t_L g910 ( .A(n_196), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g1338 ( .A(n_197), .Y(n_1338) );
INVxp33_ASAP7_75t_L g782 ( .A(n_198), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_198), .A2(n_317), .B1(n_794), .B2(n_795), .Y(n_793) );
INVx1_ASAP7_75t_L g1480 ( .A(n_200), .Y(n_1480) );
INVx1_ASAP7_75t_L g585 ( .A(n_201), .Y(n_585) );
INVx1_ASAP7_75t_L g684 ( .A(n_202), .Y(n_684) );
INVx1_ASAP7_75t_L g1070 ( .A(n_204), .Y(n_1070) );
INVxp67_ASAP7_75t_L g1401 ( .A(n_205), .Y(n_1401) );
AOI22xp33_ASAP7_75t_L g1432 ( .A1(n_205), .A2(n_345), .B1(n_795), .B2(n_1433), .Y(n_1432) );
OAI22xp33_ASAP7_75t_R g1206 ( .A1(n_206), .A2(n_368), .B1(n_659), .B2(n_1166), .Y(n_1206) );
OAI221xp5_ASAP7_75t_L g1226 ( .A1(n_206), .A2(n_368), .B1(n_855), .B2(n_891), .C(n_1227), .Y(n_1226) );
OAI221xp5_ASAP7_75t_SL g967 ( .A1(n_207), .A2(n_363), .B1(n_613), .B2(n_659), .C(n_968), .Y(n_967) );
OAI221xp5_ASAP7_75t_L g1001 ( .A1(n_207), .A2(n_363), .B1(n_728), .B2(n_891), .C(n_1002), .Y(n_1001) );
CKINVDCx5p33_ASAP7_75t_R g1336 ( .A(n_208), .Y(n_1336) );
INVx1_ASAP7_75t_L g1216 ( .A(n_209), .Y(n_1216) );
INVx1_ASAP7_75t_L g1395 ( .A(n_210), .Y(n_1395) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_211), .A2(n_350), .B1(n_678), .B2(n_681), .Y(n_677) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_211), .Y(n_699) );
INVx1_ASAP7_75t_L g1031 ( .A(n_212), .Y(n_1031) );
INVxp67_ASAP7_75t_SL g1646 ( .A(n_213), .Y(n_1646) );
INVx1_ASAP7_75t_L g673 ( .A(n_214), .Y(n_673) );
CKINVDCx5p33_ASAP7_75t_R g1148 ( .A(n_216), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g1615 ( .A(n_217), .Y(n_1615) );
INVx1_ASAP7_75t_L g1267 ( .A(n_218), .Y(n_1267) );
INVxp33_ASAP7_75t_L g738 ( .A(n_219), .Y(n_738) );
INVx1_ASAP7_75t_L g653 ( .A(n_220), .Y(n_653) );
INVxp33_ASAP7_75t_SL g1527 ( .A(n_221), .Y(n_1527) );
AOI221xp5_ASAP7_75t_L g1553 ( .A1(n_221), .A2(n_273), .B1(n_521), .B2(n_1554), .C(n_1555), .Y(n_1553) );
AOI22xp33_ASAP7_75t_L g1250 ( .A1(n_222), .A2(n_313), .B1(n_681), .B2(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1272 ( .A(n_222), .Y(n_1272) );
INVx1_ASAP7_75t_L g806 ( .A(n_223), .Y(n_806) );
INVx1_ASAP7_75t_L g447 ( .A(n_224), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g520 ( .A1(n_224), .A2(n_318), .B1(n_521), .B2(n_525), .C(n_526), .Y(n_520) );
INVx1_ASAP7_75t_L g1958 ( .A(n_225), .Y(n_1958) );
INVxp67_ASAP7_75t_SL g1238 ( .A(n_226), .Y(n_1238) );
INVxp67_ASAP7_75t_L g1454 ( .A(n_228), .Y(n_1454) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_228), .A2(n_285), .B1(n_640), .B2(n_836), .Y(n_1473) );
INVx1_ASAP7_75t_L g990 ( .A(n_229), .Y(n_990) );
INVx1_ASAP7_75t_L g492 ( .A(n_230), .Y(n_492) );
INVx1_ASAP7_75t_L g538 ( .A(n_230), .Y(n_538) );
INVx1_ASAP7_75t_L g1029 ( .A(n_232), .Y(n_1029) );
INVxp33_ASAP7_75t_SL g587 ( .A(n_233), .Y(n_587) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_233), .A2(n_536), .B(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g906 ( .A(n_234), .Y(n_906) );
CKINVDCx20_ASAP7_75t_R g1757 ( .A(n_235), .Y(n_1757) );
CKINVDCx5p33_ASAP7_75t_R g1095 ( .A(n_238), .Y(n_1095) );
INVx1_ASAP7_75t_L g1537 ( .A(n_239), .Y(n_1537) );
INVx1_ASAP7_75t_L g1457 ( .A(n_240), .Y(n_1457) );
AOI22xp33_ASAP7_75t_SL g1605 ( .A1(n_241), .A2(n_300), .B1(n_1212), .B2(n_1602), .Y(n_1605) );
OAI211xp5_ASAP7_75t_SL g1623 ( .A1(n_241), .A2(n_1624), .B(n_1628), .C(n_1632), .Y(n_1623) );
INVxp67_ASAP7_75t_SL g1233 ( .A(n_242), .Y(n_1233) );
XNOR2x1_ASAP7_75t_L g1329 ( .A(n_243), .B(n_1330), .Y(n_1329) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_244), .A2(n_335), .B1(n_630), .B2(n_800), .C(n_973), .Y(n_1249) );
INVx1_ASAP7_75t_L g1270 ( .A(n_244), .Y(n_1270) );
CKINVDCx14_ASAP7_75t_R g1720 ( .A(n_245), .Y(n_1720) );
INVx1_ASAP7_75t_L g1461 ( .A(n_247), .Y(n_1461) );
INVx1_ASAP7_75t_L g1008 ( .A(n_248), .Y(n_1008) );
CKINVDCx5p33_ASAP7_75t_R g1290 ( .A(n_249), .Y(n_1290) );
INVx1_ASAP7_75t_L g1334 ( .A(n_250), .Y(n_1334) );
AOI22xp33_ASAP7_75t_L g825 ( .A1(n_251), .A2(n_258), .B1(n_826), .B2(n_828), .Y(n_825) );
INVx1_ASAP7_75t_L g847 ( .A(n_251), .Y(n_847) );
INVx1_ASAP7_75t_L g864 ( .A(n_252), .Y(n_864) );
INVxp33_ASAP7_75t_L g756 ( .A(n_253), .Y(n_756) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_253), .A2(n_290), .B1(n_635), .B2(n_787), .C(n_788), .Y(n_786) );
INVx1_ASAP7_75t_L g1205 ( .A(n_254), .Y(n_1205) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_255), .A2(n_320), .B1(n_986), .B2(n_987), .Y(n_985) );
INVx1_ASAP7_75t_L g1007 ( .A(n_255), .Y(n_1007) );
INVx1_ASAP7_75t_L g1197 ( .A(n_256), .Y(n_1197) );
INVx1_ASAP7_75t_L g1119 ( .A(n_257), .Y(n_1119) );
INVx1_ASAP7_75t_L g851 ( .A(n_258), .Y(n_851) );
XNOR2xp5_ASAP7_75t_L g811 ( .A(n_259), .B(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g1928 ( .A(n_260), .Y(n_1928) );
OAI211xp5_ASAP7_75t_SL g1946 ( .A1(n_260), .A2(n_1624), .B(n_1947), .C(n_1957), .Y(n_1946) );
INVx1_ASAP7_75t_L g1311 ( .A(n_261), .Y(n_1311) );
OAI211xp5_ASAP7_75t_L g1323 ( .A1(n_261), .A2(n_1042), .B(n_1324), .C(n_1328), .Y(n_1323) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_262), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_263), .Y(n_1151) );
INVx1_ASAP7_75t_L g1925 ( .A(n_264), .Y(n_1925) );
OAI221xp5_ASAP7_75t_L g1938 ( .A1(n_264), .A2(n_1638), .B1(n_1939), .B2(n_1943), .C(n_1945), .Y(n_1938) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_265), .A2(n_303), .B1(n_461), .B2(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g569 ( .A(n_265), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g1916 ( .A(n_267), .Y(n_1916) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_268), .A2(n_279), .B1(n_621), .B2(n_634), .Y(n_970) );
INVxp33_ASAP7_75t_L g1000 ( .A(n_268), .Y(n_1000) );
INVx1_ASAP7_75t_L g1492 ( .A(n_269), .Y(n_1492) );
AOI221xp5_ASAP7_75t_L g1512 ( .A1(n_269), .A2(n_291), .B1(n_547), .B2(n_549), .C(n_1513), .Y(n_1512) );
INVxp67_ASAP7_75t_SL g1542 ( .A(n_270), .Y(n_1542) );
CKINVDCx5p33_ASAP7_75t_R g1463 ( .A(n_271), .Y(n_1463) );
XNOR2x1_ASAP7_75t_L g1245 ( .A(n_272), .B(n_1246), .Y(n_1245) );
INVxp33_ASAP7_75t_SL g1530 ( .A(n_273), .Y(n_1530) );
INVx1_ASAP7_75t_L g1409 ( .A(n_274), .Y(n_1409) );
CKINVDCx20_ASAP7_75t_R g1679 ( .A(n_275), .Y(n_1679) );
BUFx3_ASAP7_75t_L g499 ( .A(n_276), .Y(n_499) );
INVx1_ASAP7_75t_L g506 ( .A(n_276), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g1139 ( .A(n_277), .Y(n_1139) );
AO221x2_ASAP7_75t_L g1753 ( .A1(n_278), .A2(n_349), .B1(n_1754), .B2(n_1755), .C(n_1756), .Y(n_1753) );
INVxp33_ASAP7_75t_L g996 ( .A(n_279), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g1710 ( .A1(n_280), .A2(n_281), .B1(n_1693), .B2(n_1711), .Y(n_1710) );
INVx1_ASAP7_75t_L g1015 ( .A(n_281), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_282), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_282), .B(n_353), .Y(n_415) );
AND2x2_ASAP7_75t_L g436 ( .A(n_282), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g481 ( .A(n_282), .Y(n_481) );
INVx1_ASAP7_75t_L g416 ( .A(n_283), .Y(n_416) );
CKINVDCx5p33_ASAP7_75t_R g1353 ( .A(n_284), .Y(n_1353) );
INVxp67_ASAP7_75t_L g1452 ( .A(n_285), .Y(n_1452) );
INVx1_ASAP7_75t_L g1110 ( .A(n_286), .Y(n_1110) );
AOI21xp5_ASAP7_75t_L g1992 ( .A1(n_287), .A2(n_801), .B(n_929), .Y(n_1992) );
INVx1_ASAP7_75t_L g2012 ( .A(n_287), .Y(n_2012) );
OAI332xp33_ASAP7_75t_L g1133 ( .A1(n_288), .A2(n_477), .A3(n_689), .B1(n_1134), .B2(n_1138), .B3(n_1143), .C1(n_1149), .C2(n_1152), .Y(n_1133) );
INVx1_ASAP7_75t_L g1183 ( .A(n_288), .Y(n_1183) );
INVx1_ASAP7_75t_L g668 ( .A(n_289), .Y(n_668) );
INVxp67_ASAP7_75t_L g746 ( .A(n_290), .Y(n_746) );
INVx1_ASAP7_75t_L g1490 ( .A(n_291), .Y(n_1490) );
INVx1_ASAP7_75t_L g1560 ( .A(n_292), .Y(n_1560) );
INVx2_ASAP7_75t_L g494 ( .A(n_293), .Y(n_494) );
OR2x2_ASAP7_75t_L g508 ( .A(n_293), .B(n_492), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g1136 ( .A(n_294), .Y(n_1136) );
INVxp67_ASAP7_75t_L g1405 ( .A(n_295), .Y(n_1405) );
AOI221xp5_ASAP7_75t_L g1429 ( .A1(n_295), .A2(n_343), .B1(n_1210), .B2(n_1430), .C(n_1431), .Y(n_1429) );
INVx1_ASAP7_75t_L g1285 ( .A(n_296), .Y(n_1285) );
CKINVDCx16_ASAP7_75t_R g1020 ( .A(n_297), .Y(n_1020) );
INVx1_ASAP7_75t_L g1343 ( .A(n_298), .Y(n_1343) );
INVx1_ASAP7_75t_L g976 ( .A(n_299), .Y(n_976) );
OAI221xp5_ASAP7_75t_L g1637 ( .A1(n_300), .A2(n_1638), .B1(n_1640), .B2(n_1645), .C(n_1653), .Y(n_1637) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_301), .A2(n_332), .B1(n_638), .B2(n_640), .Y(n_1254) );
INVx1_ASAP7_75t_L g1279 ( .A(n_301), .Y(n_1279) );
AOI22xp5_ASAP7_75t_SL g1705 ( .A1(n_302), .A2(n_307), .B1(n_1687), .B2(n_1693), .Y(n_1705) );
INVx1_ASAP7_75t_L g545 ( .A(n_303), .Y(n_545) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_304), .Y(n_442) );
INVx1_ASAP7_75t_L g1412 ( .A(n_305), .Y(n_1412) );
INVxp67_ASAP7_75t_SL g1996 ( .A(n_306), .Y(n_1996) );
AOI221xp5_ASAP7_75t_L g1988 ( .A1(n_308), .A2(n_319), .B1(n_675), .B2(n_1989), .C(n_1990), .Y(n_1988) );
INVxp33_ASAP7_75t_L g2011 ( .A(n_308), .Y(n_2011) );
INVx1_ASAP7_75t_L g1493 ( .A(n_309), .Y(n_1493) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_311), .Y(n_1194) );
INVx1_ASAP7_75t_L g1304 ( .A(n_312), .Y(n_1304) );
AOI21xp5_ASAP7_75t_L g1321 ( .A1(n_312), .A2(n_671), .B(n_946), .Y(n_1321) );
INVx1_ASAP7_75t_L g1269 ( .A(n_313), .Y(n_1269) );
CKINVDCx5p33_ASAP7_75t_R g1483 ( .A(n_314), .Y(n_1483) );
INVxp33_ASAP7_75t_L g778 ( .A(n_317), .Y(n_778) );
INVx1_ASAP7_75t_L g428 ( .A(n_318), .Y(n_428) );
INVx1_ASAP7_75t_L g1011 ( .A(n_320), .Y(n_1011) );
INVx1_ASAP7_75t_L g767 ( .A(n_321), .Y(n_767) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_322), .Y(n_580) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_322), .A2(n_348), .B1(n_613), .B2(n_615), .C(n_617), .Y(n_612) );
INVx1_ASAP7_75t_L g913 ( .A(n_323), .Y(n_913) );
CKINVDCx5p33_ASAP7_75t_R g1495 ( .A(n_324), .Y(n_1495) );
INVx1_ASAP7_75t_L g1307 ( .A(n_325), .Y(n_1307) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_326), .A2(n_332), .B1(n_868), .B2(n_1058), .C(n_1278), .Y(n_1277) );
INVxp33_ASAP7_75t_L g897 ( .A(n_327), .Y(n_897) );
XNOR2xp5_ASAP7_75t_L g1979 ( .A(n_330), .B(n_1980), .Y(n_1979) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_331), .A2(n_333), .B1(n_557), .B2(n_560), .Y(n_556) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_334), .A2(n_365), .B1(n_836), .B2(n_838), .Y(n_835) );
INVx1_ASAP7_75t_L g866 ( .A(n_334), .Y(n_866) );
INVx1_ASAP7_75t_L g1276 ( .A(n_335), .Y(n_1276) );
CKINVDCx5p33_ASAP7_75t_R g1256 ( .A(n_336), .Y(n_1256) );
INVx1_ASAP7_75t_L g969 ( .A(n_338), .Y(n_969) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g1674 ( .A(n_339), .B(n_381), .Y(n_1674) );
AND3x2_ASAP7_75t_L g1690 ( .A(n_339), .B(n_381), .C(n_1677), .Y(n_1690) );
INVx1_ASAP7_75t_L g803 ( .A(n_340), .Y(n_803) );
INVx2_ASAP7_75t_L g394 ( .A(n_341), .Y(n_394) );
XNOR2x2_ASAP7_75t_L g1523 ( .A(n_342), .B(n_1524), .Y(n_1523) );
INVxp67_ASAP7_75t_SL g1406 ( .A(n_343), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_344), .Y(n_438) );
INVxp33_ASAP7_75t_SL g1403 ( .A(n_345), .Y(n_1403) );
INVx1_ASAP7_75t_L g1528 ( .A(n_347), .Y(n_1528) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_348), .Y(n_581) );
AOI22x1_ASAP7_75t_L g740 ( .A1(n_349), .A2(n_741), .B1(n_742), .B2(n_807), .Y(n_740) );
INVx1_ASAP7_75t_L g807 ( .A(n_349), .Y(n_807) );
INVxp33_ASAP7_75t_L g703 ( .A(n_350), .Y(n_703) );
CKINVDCx5p33_ASAP7_75t_R g1135 ( .A(n_351), .Y(n_1135) );
INVx1_ASAP7_75t_L g1203 ( .A(n_352), .Y(n_1203) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
INVx2_ASAP7_75t_L g437 ( .A(n_353), .Y(n_437) );
INVx1_ASAP7_75t_L g1266 ( .A(n_354), .Y(n_1266) );
INVxp33_ASAP7_75t_L g1446 ( .A(n_355), .Y(n_1446) );
AOI221xp5_ASAP7_75t_L g1466 ( .A1(n_355), .A2(n_358), .B1(n_800), .B2(n_940), .C(n_973), .Y(n_1466) );
OAI22xp33_ASAP7_75t_L g1565 ( .A1(n_356), .A2(n_369), .B1(n_633), .B2(n_1081), .Y(n_1565) );
INVxp67_ASAP7_75t_L g611 ( .A(n_357), .Y(n_611) );
INVxp33_ASAP7_75t_L g1444 ( .A(n_358), .Y(n_1444) );
INVxp67_ASAP7_75t_SL g1652 ( .A(n_359), .Y(n_1652) );
INVxp33_ASAP7_75t_L g753 ( .A(n_360), .Y(n_753) );
INVxp67_ASAP7_75t_SL g1986 ( .A(n_361), .Y(n_1986) );
INVxp67_ASAP7_75t_SL g2027 ( .A(n_362), .Y(n_2027) );
INVx1_ASAP7_75t_L g861 ( .A(n_365), .Y(n_861) );
CKINVDCx5p33_ASAP7_75t_R g1983 ( .A(n_366), .Y(n_1983) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_367), .Y(n_817) );
INVxp67_ASAP7_75t_SL g1541 ( .A(n_369), .Y(n_1541) );
INVx1_ASAP7_75t_L g989 ( .A(n_371), .Y(n_989) );
INVxp33_ASAP7_75t_SL g1394 ( .A(n_372), .Y(n_1394) );
INVx1_ASAP7_75t_L g1942 ( .A(n_373), .Y(n_1942) );
INVxp33_ASAP7_75t_L g1443 ( .A(n_374), .Y(n_1443) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_397), .B(n_1664), .Y(n_375) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_384), .Y(n_378) );
AND2x4_ASAP7_75t_L g1973 ( .A(n_379), .B(n_385), .Y(n_1973) );
NOR2xp33_ASAP7_75t_SL g379 ( .A(n_380), .B(n_382), .Y(n_379) );
INVx1_ASAP7_75t_SL g1977 ( .A(n_380), .Y(n_1977) );
NAND2xp5_ASAP7_75t_L g2034 ( .A(n_380), .B(n_382), .Y(n_2034) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g1976 ( .A(n_382), .B(n_1977), .Y(n_1976) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_386), .B(n_390), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g459 ( .A(n_388), .B(n_396), .Y(n_459) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OR2x2_ASAP7_75t_L g690 ( .A(n_389), .B(n_691), .Y(n_690) );
OR2x6_ASAP7_75t_L g390 ( .A(n_391), .B(n_395), .Y(n_390) );
OR2x2_ASAP7_75t_L g485 ( .A(n_391), .B(n_414), .Y(n_485) );
BUFx6f_ASAP7_75t_L g705 ( .A(n_391), .Y(n_705) );
INVx2_ASAP7_75t_SL g717 ( .A(n_391), .Y(n_717) );
BUFx2_ASAP7_75t_L g860 ( .A(n_391), .Y(n_860) );
INVx1_ASAP7_75t_L g1006 ( .A(n_391), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1118 ( .A1(n_391), .A2(n_759), .B1(n_1089), .B2(n_1119), .Y(n_1118) );
INVx2_ASAP7_75t_SL g1231 ( .A(n_391), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g1284 ( .A1(n_391), .A2(n_759), .B1(n_1256), .B2(n_1285), .Y(n_1284) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g412 ( .A(n_393), .Y(n_412) );
INVx1_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
AND2x4_ASAP7_75t_L g433 ( .A(n_393), .B(n_426), .Y(n_433) );
AND2x2_ASAP7_75t_L g446 ( .A(n_393), .B(n_394), .Y(n_446) );
INVx2_ASAP7_75t_L g451 ( .A(n_393), .Y(n_451) );
INVx1_ASAP7_75t_L g419 ( .A(n_394), .Y(n_419) );
INVx2_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
INVx1_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_394), .B(n_451), .Y(n_698) );
INVx1_ASAP7_75t_L g711 ( .A(n_394), .Y(n_711) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
XOR2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_952), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_808), .B2(n_809), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AO22x2_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_648), .B2(n_649), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_576), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_482), .Y(n_404) );
AND4x1_ASAP7_75t_L g405 ( .A(n_406), .B(n_427), .C(n_441), .D(n_454), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_416), .B1(n_417), .B2(n_420), .C(n_421), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g1566 ( .A1(n_407), .A2(n_422), .B1(n_1560), .B2(n_1561), .C(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_409), .A2(n_417), .B1(n_422), .B2(n_580), .C(n_581), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g1072 ( .A1(n_409), .A2(n_417), .B1(n_422), .B2(n_1031), .C(n_1032), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_409), .A2(n_1071), .B1(n_1083), .B2(n_1105), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1265 ( .A1(n_409), .A2(n_417), .B1(n_422), .B2(n_1266), .C(n_1267), .Y(n_1265) );
AOI221xp5_ASAP7_75t_L g1289 ( .A1(n_409), .A2(n_417), .B1(n_422), .B2(n_1290), .C(n_1291), .Y(n_1289) );
AOI221xp5_ASAP7_75t_L g2026 ( .A1(n_409), .A2(n_417), .B1(n_422), .B2(n_2027), .C(n_2028), .Y(n_2026) );
AND2x4_ASAP7_75t_L g409 ( .A(n_410), .B(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
AND2x2_ASAP7_75t_L g710 ( .A(n_412), .B(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_412), .B(n_711), .Y(n_760) );
AND2x4_ASAP7_75t_L g417 ( .A(n_413), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_L g422 ( .A(n_413), .B(n_423), .Y(n_422) );
NAND2x1_ASAP7_75t_SL g724 ( .A(n_413), .B(n_725), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g728 ( .A(n_413), .B(n_729), .Y(n_728) );
NAND2x1p5_ASAP7_75t_L g732 ( .A(n_413), .B(n_440), .Y(n_732) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g1621 ( .A(n_415), .Y(n_1621) );
AOI21xp5_ASAP7_75t_L g1121 ( .A1(n_417), .A2(n_422), .B(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1568 ( .A(n_417), .Y(n_1568) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_418), .B(n_1619), .Y(n_1634) );
AND2x2_ASAP7_75t_L g1959 ( .A(n_418), .B(n_1619), .Y(n_1959) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g726 ( .A(n_419), .Y(n_726) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
HB1xp67_ASAP7_75t_L g2023 ( .A(n_423), .Y(n_2023) );
BUFx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
BUFx3_ASAP7_75t_L g440 ( .A(n_424), .Y(n_440) );
INVx1_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
BUFx6f_ASAP7_75t_L g1056 ( .A(n_424), .Y(n_1056) );
BUFx3_ASAP7_75t_L g1545 ( .A(n_424), .Y(n_1545) );
AND2x4_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_429), .B1(n_438), .B2(n_439), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_429), .A2(n_439), .B1(n_884), .B2(n_885), .Y(n_883) );
HB1xp67_ASAP7_75t_L g1396 ( .A(n_429), .Y(n_1396) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
BUFx2_ASAP7_75t_L g584 ( .A(n_430), .Y(n_584) );
BUFx2_ASAP7_75t_L g736 ( .A(n_430), .Y(n_736) );
BUFx2_ASAP7_75t_L g997 ( .A(n_430), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_430), .A2(n_1203), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
BUFx2_ASAP7_75t_L g1273 ( .A(n_430), .Y(n_1273) );
BUFx2_ASAP7_75t_L g1335 ( .A(n_430), .Y(n_1335) );
AOI22xp33_ASAP7_75t_L g1442 ( .A1(n_430), .A2(n_439), .B1(n_1443), .B2(n_1444), .Y(n_1442) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_434), .Y(n_430) );
BUFx3_ASAP7_75t_L g701 ( .A(n_431), .Y(n_701) );
INVx1_ASAP7_75t_L g714 ( .A(n_431), .Y(n_714) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g601 ( .A(n_432), .Y(n_601) );
BUFx6f_ASAP7_75t_L g1298 ( .A(n_432), .Y(n_1298) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_433), .Y(n_470) );
INVx1_ASAP7_75t_L g1651 ( .A(n_433), .Y(n_1651) );
AND2x6_ASAP7_75t_L g439 ( .A(n_434), .B(n_440), .Y(n_439) );
AND2x4_ASAP7_75t_L g443 ( .A(n_434), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g448 ( .A(n_434), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g739 ( .A(n_434), .B(n_449), .Y(n_739) );
AND2x2_ASAP7_75t_L g852 ( .A(n_434), .B(n_449), .Y(n_852) );
AND2x2_ASAP7_75t_L g889 ( .A(n_434), .B(n_449), .Y(n_889) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_434), .A2(n_476), .B1(n_1048), .B2(n_1057), .Y(n_1047) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_434), .B(n_449), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_434), .B(n_1109), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1111 ( .A(n_434), .B(n_601), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1120 ( .A(n_434), .B(n_475), .Y(n_1120) );
AND2x4_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx1_ASAP7_75t_L g478 ( .A(n_435), .Y(n_478) );
OR2x2_ASAP7_75t_L g1577 ( .A(n_435), .B(n_508), .Y(n_1577) );
INVx2_ASAP7_75t_L g1627 ( .A(n_436), .Y(n_1627) );
AND2x4_ASAP7_75t_L g1639 ( .A(n_436), .B(n_462), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1656 ( .A(n_436), .B(n_450), .Y(n_1656) );
INVx1_ASAP7_75t_L g480 ( .A(n_437), .Y(n_480) );
INVx1_ASAP7_75t_L g691 ( .A(n_437), .Y(n_691) );
OAI221xp5_ASAP7_75t_L g526 ( .A1(n_438), .A2(n_442), .B1(n_527), .B2(n_532), .C(n_535), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_439), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_439), .A2(n_668), .B1(n_735), .B2(n_736), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_439), .A2(n_584), .B1(n_778), .B2(n_779), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_439), .A2(n_736), .B1(n_847), .B2(n_848), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_439), .A2(n_969), .B1(n_996), .B2(n_997), .Y(n_995) );
INVx1_ASAP7_75t_SL g1128 ( .A(n_439), .Y(n_1128) );
BUFx2_ASAP7_75t_L g1225 ( .A(n_439), .Y(n_1225) );
AOI22xp5_ASAP7_75t_L g1268 ( .A1(n_439), .A2(n_739), .B1(n_1269), .B2(n_1270), .Y(n_1268) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_439), .A2(n_1103), .B1(n_1307), .B2(n_1308), .Y(n_1306) );
AOI22xp33_ASAP7_75t_L g1333 ( .A1(n_439), .A2(n_1334), .B1(n_1335), .B2(n_1336), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_439), .A2(n_1273), .B1(n_1480), .B2(n_1481), .Y(n_1479) );
AOI22xp33_ASAP7_75t_L g1526 ( .A1(n_439), .A2(n_1335), .B1(n_1527), .B2(n_1528), .Y(n_1526) );
BUFx2_ASAP7_75t_L g595 ( .A(n_440), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_443), .B1(n_447), .B2(n_448), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_443), .A2(n_448), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_443), .A2(n_669), .B1(n_738), .B2(n_739), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_443), .A2(n_739), .B1(n_781), .B2(n_782), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g849 ( .A1(n_443), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_849) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_443), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_443), .A2(n_448), .B1(n_999), .B2(n_1000), .Y(n_998) );
BUFx2_ASAP7_75t_L g1221 ( .A(n_443), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1303 ( .A(n_443), .B(n_1304), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_443), .A2(n_852), .B1(n_1338), .B2(n_1339), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_443), .A2(n_852), .B1(n_1446), .B2(n_1447), .Y(n_1445) );
AOI22xp33_ASAP7_75t_L g1482 ( .A1(n_443), .A2(n_889), .B1(n_1483), .B2(n_1484), .Y(n_1482) );
AOI21xp5_ASAP7_75t_L g1532 ( .A1(n_443), .A2(n_1533), .B(n_1534), .Y(n_1532) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_SL g1109 ( .A(n_445), .Y(n_1109) );
INVx2_ASAP7_75t_L g2019 ( .A(n_445), .Y(n_2019) );
INVx3_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_446), .Y(n_462) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
BUFx2_ASAP7_75t_L g597 ( .A(n_450), .Y(n_597) );
INVx1_ASAP7_75t_L g1059 ( .A(n_450), .Y(n_1059) );
INVx1_ASAP7_75t_L g1066 ( .A(n_450), .Y(n_1066) );
BUFx6f_ASAP7_75t_L g1115 ( .A(n_450), .Y(n_1115) );
AND2x4_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx1_ASAP7_75t_L g730 ( .A(n_451), .Y(n_730) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI33xp33_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_460), .A3(n_465), .B1(n_471), .B2(n_473), .B3(n_476), .Y(n_454) );
BUFx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g2016 ( .A(n_456), .Y(n_2016) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_459), .Y(n_456) );
BUFx2_ASAP7_75t_L g575 ( .A(n_457), .Y(n_575) );
AND2x4_ASAP7_75t_L g591 ( .A(n_457), .B(n_459), .Y(n_591) );
AOI31xp33_ASAP7_75t_L g917 ( .A1(n_457), .A2(n_918), .A3(n_935), .B(n_949), .Y(n_917) );
INVx2_ASAP7_75t_L g1045 ( .A(n_457), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_457), .B(n_1302), .Y(n_1301) );
OR2x6_ASAP7_75t_L g1600 ( .A(n_457), .B(n_943), .Y(n_1600) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_L g608 ( .A(n_458), .Y(n_608) );
OR2x6_ASAP7_75t_L g689 ( .A(n_458), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g1644 ( .A(n_459), .Y(n_1644) );
BUFx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_462), .Y(n_594) );
INVx3_ASAP7_75t_L g1295 ( .A(n_462), .Y(n_1295) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx3_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g472 ( .A(n_470), .Y(n_472) );
INVx2_ASAP7_75t_SL g896 ( .A(n_470), .Y(n_896) );
INVx2_ASAP7_75t_SL g907 ( .A(n_470), .Y(n_907) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_470), .Y(n_1050) );
INVx4_ASAP7_75t_L g1137 ( .A(n_470), .Y(n_1137) );
INVx1_ASAP7_75t_L g772 ( .A(n_472), .Y(n_772) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI33xp33_ASAP7_75t_L g589 ( .A1(n_476), .A2(n_590), .A3(n_592), .B1(n_596), .B2(n_598), .B3(n_602), .Y(n_589) );
INVx1_ASAP7_75t_L g914 ( .A(n_476), .Y(n_914) );
AOI322xp5_ASAP7_75t_L g1113 ( .A1(n_476), .A2(n_591), .A3(n_1095), .B1(n_1114), .B2(n_1116), .C1(n_1117), .C2(n_1120), .Y(n_1113) );
AOI222xp33_ASAP7_75t_L g1275 ( .A1(n_476), .A2(n_591), .B1(n_1108), .B2(n_1276), .C1(n_1277), .C2(n_1281), .Y(n_1275) );
INVx6_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx5_ASAP7_75t_L g720 ( .A(n_477), .Y(n_720) );
OR2x6_ASAP7_75t_L g477 ( .A(n_478), .B(n_479), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g1594 ( .A(n_478), .B(n_490), .Y(n_1594) );
INVx2_ASAP7_75t_L g1302 ( .A(n_479), .Y(n_1302) );
BUFx2_ASAP7_75t_L g1956 ( .A(n_479), .Y(n_1956) );
NAND2x1p5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
AOI21xp33_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_500), .B(n_501), .Y(n_482) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_483), .A2(n_916), .B(n_917), .Y(n_915) );
AOI21xp5_ASAP7_75t_L g1361 ( .A1(n_483), .A2(n_1362), .B(n_1363), .Y(n_1361) );
AOI21xp5_ASAP7_75t_L g1501 ( .A1(n_483), .A2(n_1502), .B(n_1503), .Y(n_1501) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx5_ASAP7_75t_L g647 ( .A(n_484), .Y(n_647) );
INVx2_ASAP7_75t_L g843 ( .A(n_484), .Y(n_843) );
INVx1_ASAP7_75t_L g1982 ( .A(n_484), .Y(n_1982) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
INVx2_ASAP7_75t_L g1071 ( .A(n_485), .Y(n_1071) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x6_ASAP7_75t_L g1616 ( .A(n_487), .B(n_1617), .Y(n_1616) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x4_ASAP7_75t_L g1609 ( .A(n_488), .B(n_537), .Y(n_1609) );
INVx2_ASAP7_75t_L g1042 ( .A(n_489), .Y(n_1042) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_495), .Y(n_489) );
AND2x4_ASAP7_75t_L g512 ( .A(n_490), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g517 ( .A(n_490), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g566 ( .A(n_490), .Y(n_566) );
AND2x4_ASAP7_75t_L g614 ( .A(n_490), .B(n_513), .Y(n_614) );
AND2x4_ASAP7_75t_L g616 ( .A(n_490), .B(n_518), .Y(n_616) );
BUFx2_ASAP7_75t_L g642 ( .A(n_490), .Y(n_642) );
AND2x2_ASAP7_75t_L g660 ( .A(n_490), .B(n_518), .Y(n_660) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_493), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x4_ASAP7_75t_L g537 ( .A(n_493), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g555 ( .A(n_494), .B(n_538), .Y(n_555) );
INVx2_ASAP7_75t_L g559 ( .A(n_495), .Y(n_559) );
INVx6_ASAP7_75t_L g624 ( .A(n_495), .Y(n_624) );
BUFx2_ASAP7_75t_L g927 ( .A(n_495), .Y(n_927) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
INVx1_ASAP7_75t_L g519 ( .A(n_496), .Y(n_519) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g505 ( .A(n_497), .B(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g544 ( .A(n_497), .B(n_499), .Y(n_544) );
INVx1_ASAP7_75t_L g515 ( .A(n_498), .Y(n_515) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x4_ASAP7_75t_L g523 ( .A(n_499), .B(n_524), .Y(n_523) );
AOI31xp33_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_539), .A3(n_568), .B(n_575), .Y(n_501) );
AOI211xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_509), .B(n_510), .C(n_520), .Y(n_502) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_503), .A2(n_611), .B(n_612), .Y(n_610) );
AOI211xp5_ASAP7_75t_L g655 ( .A1(n_503), .A2(n_656), .B(n_657), .C(n_661), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_503), .A2(n_570), .B1(n_764), .B2(n_771), .Y(n_804) );
INVx1_ASAP7_75t_L g920 ( .A(n_503), .Y(n_920) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_503), .A2(n_966), .B(n_967), .Y(n_965) );
HB1xp67_ASAP7_75t_L g1198 ( .A(n_503), .Y(n_1198) );
AOI211xp5_ASAP7_75t_L g1371 ( .A1(n_503), .A2(n_1353), .B(n_1372), .C(n_1373), .Y(n_1371) );
AOI221xp5_ASAP7_75t_L g1465 ( .A1(n_503), .A2(n_1457), .B1(n_1466), .B2(n_1467), .C(n_1469), .Y(n_1465) );
AOI211xp5_ASAP7_75t_L g1504 ( .A1(n_503), .A2(n_1497), .B(n_1505), .C(n_1506), .Y(n_1504) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
BUFx3_ASAP7_75t_L g525 ( .A(n_504), .Y(n_525) );
INVx2_ASAP7_75t_SL g938 ( .A(n_504), .Y(n_938) );
INVx1_ASAP7_75t_L g1508 ( .A(n_504), .Y(n_1508) );
BUFx6f_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g548 ( .A(n_505), .Y(n_548) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_505), .Y(n_620) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_505), .Y(n_634) );
BUFx2_ASAP7_75t_L g675 ( .A(n_505), .Y(n_675) );
BUFx6f_ASAP7_75t_L g787 ( .A(n_505), .Y(n_787) );
BUFx2_ASAP7_75t_L g924 ( .A(n_505), .Y(n_924) );
BUFx3_ASAP7_75t_L g1099 ( .A(n_505), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g1253 ( .A(n_505), .Y(n_1253) );
INVx1_ASAP7_75t_L g531 ( .A(n_506), .Y(n_531) );
AND2x4_ASAP7_75t_L g542 ( .A(n_507), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g818 ( .A(n_507), .B(n_787), .Y(n_818) );
AOI222xp33_ASAP7_75t_L g1023 ( .A1(n_507), .A2(n_512), .B1(n_660), .B2(n_1024), .C1(n_1031), .C2(n_1032), .Y(n_1023) );
OAI21xp5_ASAP7_75t_L g1076 ( .A1(n_507), .A2(n_1077), .B(n_1080), .Y(n_1076) );
AOI221xp5_ASAP7_75t_L g1255 ( .A1(n_507), .A2(n_570), .B1(n_1256), .B2(n_1257), .C(n_1262), .Y(n_1255) );
A2O1A1Ixp33_ASAP7_75t_L g1324 ( .A1(n_507), .A2(n_940), .B(n_1325), .C(n_1326), .Y(n_1324) );
OAI21xp5_ASAP7_75t_L g1562 ( .A1(n_507), .A2(n_1563), .B(n_1565), .Y(n_1562) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g571 ( .A(n_508), .B(n_534), .Y(n_571) );
OR2x2_ASAP7_75t_L g574 ( .A(n_508), .B(n_563), .Y(n_574) );
A2O1A1Ixp33_ASAP7_75t_SL g1154 ( .A1(n_508), .A2(n_1155), .B(n_1159), .C(n_1164), .Y(n_1154) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g658 ( .A(n_512), .Y(n_658) );
AOI322xp5_ASAP7_75t_L g792 ( .A1(n_512), .A2(n_517), .A3(n_793), .B1(n_797), .B2(n_799), .C1(n_802), .C2(n_803), .Y(n_792) );
INVx2_ASAP7_75t_SL g1166 ( .A(n_512), .Y(n_1166) );
INVx2_ASAP7_75t_SL g1470 ( .A(n_512), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_512), .A2(n_660), .B1(n_1560), .B2(n_1561), .Y(n_1559) );
INVxp67_ASAP7_75t_L g934 ( .A(n_513), .Y(n_934) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g1592 ( .A(n_514), .Y(n_1592) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_SL g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g933 ( .A(n_518), .Y(n_933) );
INVx1_ASAP7_75t_L g1086 ( .A(n_518), .Y(n_1086) );
BUFx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
HB1xp67_ASAP7_75t_L g1370 ( .A(n_521), .Y(n_1370) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g682 ( .A(n_522), .Y(n_682) );
INVx1_ASAP7_75t_L g796 ( .A(n_522), .Y(n_796) );
INVx1_ASAP7_75t_L g948 ( .A(n_522), .Y(n_948) );
BUFx6f_ASAP7_75t_L g987 ( .A(n_522), .Y(n_987) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g563 ( .A(n_523), .Y(n_563) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_523), .Y(n_621) );
INVx1_ASAP7_75t_L g663 ( .A(n_523), .Y(n_663) );
INVx1_ASAP7_75t_L g1158 ( .A(n_523), .Y(n_1158) );
INVx1_ASAP7_75t_L g530 ( .A(n_524), .Y(n_530) );
INVxp67_ASAP7_75t_L g1178 ( .A(n_525), .Y(n_1178) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g618 ( .A(n_528), .Y(n_618) );
INVx2_ASAP7_75t_SL g1081 ( .A(n_528), .Y(n_1081) );
INVx1_ASAP7_75t_L g1202 ( .A(n_528), .Y(n_1202) );
BUFx4f_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g667 ( .A(n_529), .Y(n_667) );
INVx1_ASAP7_75t_L g931 ( .A(n_529), .Y(n_931) );
INVx2_ASAP7_75t_L g1091 ( .A(n_529), .Y(n_1091) );
INVx1_ASAP7_75t_L g1259 ( .A(n_529), .Y(n_1259) );
BUFx2_ASAP7_75t_L g1377 ( .A(n_529), .Y(n_1377) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
OR2x2_ASAP7_75t_L g534 ( .A(n_530), .B(n_531), .Y(n_534) );
OAI221xp5_ASAP7_75t_L g666 ( .A1(n_532), .A2(n_667), .B1(n_668), .B2(n_669), .C(n_670), .Y(n_666) );
OAI221xp5_ASAP7_75t_L g1509 ( .A1(n_532), .A2(n_535), .B1(n_1481), .B2(n_1483), .C(n_1510), .Y(n_1509) );
OAI221xp5_ASAP7_75t_L g1555 ( .A1(n_532), .A2(n_618), .B1(n_1528), .B2(n_1533), .C(n_1556), .Y(n_1555) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g1026 ( .A(n_534), .Y(n_1026) );
BUFx2_ASAP7_75t_L g1204 ( .A(n_534), .Y(n_1204) );
INVx1_ASAP7_75t_L g1915 ( .A(n_534), .Y(n_1915) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_535), .A2(n_1202), .B1(n_1203), .B2(n_1204), .C(n_1205), .Y(n_1201) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g801 ( .A(n_536), .Y(n_801) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g671 ( .A(n_537), .Y(n_671) );
INVx1_ASAP7_75t_L g824 ( .A(n_537), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g973 ( .A(n_537), .Y(n_973) );
HB1xp67_ASAP7_75t_L g1556 ( .A(n_537), .Y(n_1556) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_545), .B1(n_546), .B2(n_556), .C(n_564), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_540), .A2(n_564), .B1(n_913), .B2(n_936), .C(n_944), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g1511 ( .A1(n_540), .A2(n_564), .B1(n_1500), .B2(n_1512), .C(n_1514), .Y(n_1511) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g627 ( .A(n_542), .Y(n_627) );
INVx2_ASAP7_75t_SL g840 ( .A(n_542), .Y(n_840) );
BUFx6f_ASAP7_75t_L g975 ( .A(n_542), .Y(n_975) );
INVx1_ASAP7_75t_L g1995 ( .A(n_542), .Y(n_1995) );
INVx2_ASAP7_75t_SL g631 ( .A(n_543), .Y(n_631) );
AND2x4_ASAP7_75t_L g641 ( .A(n_543), .B(n_642), .Y(n_641) );
BUFx3_ASAP7_75t_L g676 ( .A(n_543), .Y(n_676) );
BUFx4f_ASAP7_75t_L g940 ( .A(n_543), .Y(n_940) );
BUFx6f_ASAP7_75t_L g1163 ( .A(n_543), .Y(n_1163) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_544), .Y(n_553) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g794 ( .A(n_548), .Y(n_794) );
INVx1_ASAP7_75t_L g834 ( .A(n_548), .Y(n_834) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g1431 ( .A(n_550), .Y(n_1431) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_L g567 ( .A(n_553), .Y(n_567) );
INVx1_ASAP7_75t_L g982 ( .A(n_553), .Y(n_982) );
INVx1_ASAP7_75t_L g984 ( .A(n_554), .Y(n_984) );
BUFx2_ASAP7_75t_L g1210 ( .A(n_554), .Y(n_1210) );
INVx2_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
BUFx3_ASAP7_75t_L g636 ( .A(n_555), .Y(n_636) );
INVx2_ASAP7_75t_L g943 ( .A(n_555), .Y(n_943) );
INVx1_ASAP7_75t_L g1513 ( .A(n_555), .Y(n_1513) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g1583 ( .A(n_558), .B(n_1576), .Y(n_1583) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g822 ( .A(n_559), .Y(n_822) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
BUFx2_ASAP7_75t_L g925 ( .A(n_562), .Y(n_925) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g838 ( .A(n_563), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_564), .A2(n_626), .B1(n_673), .B2(n_674), .C(n_677), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g785 ( .A1(n_564), .A2(n_626), .B1(n_767), .B2(n_786), .C(n_789), .Y(n_785) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_564), .A2(n_975), .B1(n_976), .B2(n_977), .C(n_985), .Y(n_974) );
AOI21xp33_ASAP7_75t_L g1033 ( .A1(n_564), .A2(n_1034), .B(n_1035), .Y(n_1033) );
INVx1_ASAP7_75t_L g1164 ( .A(n_564), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g1207 ( .A1(n_564), .A2(n_626), .B1(n_1208), .B2(n_1209), .C(n_1211), .Y(n_1207) );
AOI221xp5_ASAP7_75t_L g1364 ( .A1(n_564), .A2(n_975), .B1(n_1360), .B2(n_1365), .C(n_1368), .Y(n_1364) );
INVx1_ASAP7_75t_L g1435 ( .A(n_564), .Y(n_1435) );
AOI221xp5_ASAP7_75t_L g1471 ( .A1(n_564), .A2(n_975), .B1(n_1461), .B2(n_1472), .C(n_1473), .Y(n_1471) );
HB1xp67_ASAP7_75t_L g2001 ( .A(n_564), .Y(n_2001) );
AND2x4_ASAP7_75t_L g564 ( .A(n_565), .B(n_567), .Y(n_564) );
INVx1_ASAP7_75t_SL g565 ( .A(n_566), .Y(n_565) );
OR2x2_ASAP7_75t_L g1167 ( .A(n_566), .B(n_933), .Y(n_1167) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_567), .Y(n_788) );
AOI22xp5_ASAP7_75t_L g1028 ( .A1(n_567), .A2(n_787), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
INVx1_ASAP7_75t_L g1367 ( .A(n_567), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_572), .B2(n_573), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_570), .A2(n_573), .B1(n_644), .B2(n_645), .Y(n_643) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_570), .A2(n_573), .B1(n_684), .B2(n_685), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g815 ( .A1(n_570), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_815) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_570), .A2(n_573), .B1(n_908), .B2(n_910), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_570), .A2(n_573), .B1(n_989), .B2(n_990), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1215 ( .A1(n_570), .A2(n_573), .B1(n_1216), .B2(n_1217), .Y(n_1215) );
AOI22xp33_ASAP7_75t_SL g1379 ( .A1(n_570), .A2(n_573), .B1(n_1356), .B2(n_1358), .Y(n_1379) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_570), .A2(n_573), .B1(n_1409), .B2(n_1411), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1474 ( .A1(n_570), .A2(n_573), .B1(n_1458), .B2(n_1460), .Y(n_1474) );
AOI22xp33_ASAP7_75t_L g1515 ( .A1(n_570), .A2(n_573), .B1(n_1495), .B2(n_1499), .Y(n_1515) );
AOI22xp33_ASAP7_75t_L g2002 ( .A1(n_570), .A2(n_573), .B1(n_2003), .B2(n_2004), .Y(n_2002) );
INVx6_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_573), .B(n_773), .Y(n_805) );
AOI221xp5_ASAP7_75t_L g819 ( .A1(n_573), .A2(n_820), .B1(n_821), .B2(n_825), .C(n_829), .Y(n_819) );
INVx4_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
CKINVDCx8_ASAP7_75t_R g1185 ( .A(n_575), .Y(n_1185) );
OAI31xp33_ASAP7_75t_SL g1936 ( .A1(n_575), .A2(n_1937), .A3(n_1938), .B(n_1946), .Y(n_1936) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_605), .Y(n_577) );
AND4x1_ASAP7_75t_L g578 ( .A(n_579), .B(n_582), .C(n_586), .D(n_589), .Y(n_578) );
OAI211xp5_ASAP7_75t_L g617 ( .A1(n_585), .A2(n_618), .B(n_619), .C(n_622), .Y(n_617) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g1063 ( .A1(n_591), .A2(n_1043), .B1(n_1064), .B2(n_1071), .Y(n_1063) );
AOI33xp33_ASAP7_75t_L g1292 ( .A1(n_591), .A2(n_1293), .A3(n_1296), .B1(n_1299), .B2(n_1300), .B3(n_1301), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g604 ( .A(n_594), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g1051 ( .A1(n_594), .A2(n_1052), .B1(n_1053), .B2(n_1054), .Y(n_1051) );
HB1xp67_ASAP7_75t_L g2022 ( .A(n_597), .Y(n_2022) );
INVx2_ASAP7_75t_SL g1350 ( .A(n_599), .Y(n_1350) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g1060 ( .A(n_600), .Y(n_1060) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g751 ( .A(n_601), .Y(n_751) );
INVx2_ASAP7_75t_L g869 ( .A(n_601), .Y(n_869) );
INVx2_ASAP7_75t_L g871 ( .A(n_601), .Y(n_871) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_606), .A2(n_609), .B1(n_646), .B2(n_647), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_606), .A2(n_647), .B1(n_784), .B2(n_806), .Y(n_783) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_606), .A2(n_814), .B1(n_842), .B2(n_843), .Y(n_813) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
BUFx8_ASAP7_75t_SL g686 ( .A(n_607), .Y(n_686) );
AOI31xp33_ASAP7_75t_L g1195 ( .A1(n_607), .A2(n_1196), .A3(n_1207), .B(n_1215), .Y(n_1195) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
BUFx2_ASAP7_75t_L g992 ( .A(n_608), .Y(n_992) );
NAND3xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_625), .C(n_643), .Y(n_609) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx4_ASAP7_75t_L g830 ( .A(n_614), .Y(n_830) );
INVx1_ASAP7_75t_SL g1263 ( .A(n_614), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1328 ( .A1(n_614), .A2(n_616), .B1(n_1290), .B2(n_1291), .Y(n_1328) );
INVx2_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g831 ( .A(n_616), .Y(n_831) );
OAI211xp5_ASAP7_75t_L g968 ( .A1(n_618), .A2(n_969), .B(n_970), .C(n_971), .Y(n_968) );
INVx2_ASAP7_75t_L g665 ( .A(n_620), .Y(n_665) );
INVx2_ASAP7_75t_SL g827 ( .A(n_620), .Y(n_827) );
BUFx3_ASAP7_75t_L g1175 ( .A(n_620), .Y(n_1175) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_621), .Y(n_640) );
BUFx3_ASAP7_75t_L g828 ( .A(n_621), .Y(n_828) );
INVx1_ASAP7_75t_L g1608 ( .A(n_621), .Y(n_1608) );
INVx1_ASAP7_75t_L g1922 ( .A(n_621), .Y(n_1922) );
INVx1_ASAP7_75t_L g791 ( .A(n_623), .Y(n_791) );
INVx2_ASAP7_75t_SL g623 ( .A(n_624), .Y(n_623) );
HB1xp67_ASAP7_75t_L g639 ( .A(n_624), .Y(n_639) );
INVx2_ASAP7_75t_L g680 ( .A(n_624), .Y(n_680) );
BUFx6f_ASAP7_75t_L g837 ( .A(n_624), .Y(n_837) );
INVx1_ASAP7_75t_L g946 ( .A(n_624), .Y(n_946) );
INVx2_ASAP7_75t_L g972 ( .A(n_624), .Y(n_972) );
INVx1_ASAP7_75t_L g1039 ( .A(n_624), .Y(n_1039) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_628), .B1(n_629), .B2(n_637), .C(n_641), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g798 ( .A(n_631), .Y(n_798) );
INVx1_ASAP7_75t_L g823 ( .A(n_631), .Y(n_823) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx3_ASAP7_75t_L g1251 ( .A(n_634), .Y(n_1251) );
INVx1_ASAP7_75t_L g1327 ( .A(n_634), .Y(n_1327) );
BUFx2_ASAP7_75t_L g1430 ( .A(n_634), .Y(n_1430) );
INVx1_ASAP7_75t_L g1931 ( .A(n_634), .Y(n_1931) );
INVx3_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g1173 ( .A1(n_636), .A2(n_930), .B1(n_1135), .B2(n_1141), .C(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1999 ( .A(n_636), .Y(n_1999) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g1172 ( .A(n_640), .Y(n_1172) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_641), .A2(n_833), .B1(n_835), .B2(n_839), .C(n_841), .Y(n_832) );
AOI221xp5_ASAP7_75t_L g1248 ( .A1(n_641), .A2(n_1249), .B1(n_1250), .B2(n_1252), .C(n_1254), .Y(n_1248) );
INVx1_ASAP7_75t_L g1322 ( .A(n_641), .Y(n_1322) );
BUFx3_ASAP7_75t_L g1087 ( .A(n_642), .Y(n_1087) );
AOI21xp33_ASAP7_75t_L g652 ( .A1(n_647), .A2(n_653), .B(n_654), .Y(n_652) );
AOI21xp33_ASAP7_75t_SL g962 ( .A1(n_647), .A2(n_963), .B(n_964), .Y(n_962) );
INVx1_ASAP7_75t_L g1417 ( .A(n_647), .Y(n_1417) );
AOI21xp33_ASAP7_75t_SL g1462 ( .A1(n_647), .A2(n_1463), .B(n_1464), .Y(n_1462) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
XOR2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_740), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_687), .Y(n_651) );
AOI31xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_672), .A3(n_683), .B(n_686), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_656), .A2(n_685), .B1(n_713), .B2(n_714), .Y(n_712) );
INVx3_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g1040 ( .A(n_663), .Y(n_1040) );
INVx1_ASAP7_75t_L g1214 ( .A(n_663), .Y(n_1214) );
INVx2_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g1378 ( .A(n_671), .Y(n_1378) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_673), .A2(n_684), .B1(n_716), .B2(n_718), .Y(n_715) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx6f_ASAP7_75t_L g800 ( .A(n_680), .Y(n_800) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g1176 ( .A1(n_682), .A2(n_1177), .B1(n_1178), .B2(n_1179), .Y(n_1176) );
OAI221xp5_ASAP7_75t_L g1422 ( .A1(n_682), .A2(n_938), .B1(n_1395), .B2(n_1423), .C(n_1424), .Y(n_1422) );
INVx1_ASAP7_75t_L g1989 ( .A(n_682), .Y(n_1989) );
AOI31xp33_ASAP7_75t_L g1419 ( .A1(n_686), .A2(n_1420), .A3(n_1426), .B(n_1436), .Y(n_1419) );
AOI31xp33_ASAP7_75t_L g1464 ( .A1(n_686), .A2(n_1465), .A3(n_1471), .B(n_1474), .Y(n_1464) );
OAI31xp33_ASAP7_75t_L g1622 ( .A1(n_686), .A2(n_1623), .A3(n_1637), .B(n_1654), .Y(n_1622) );
INVx5_ASAP7_75t_L g2006 ( .A(n_686), .Y(n_2006) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_688), .B(n_721), .C(n_733), .Y(n_687) );
OAI33xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_692), .A3(n_702), .B1(n_712), .B2(n_715), .B3(n_719), .Y(n_688) );
OAI33xp33_ASAP7_75t_L g744 ( .A1(n_689), .A2(n_719), .A3(n_745), .B1(n_752), .B2(n_761), .B3(n_768), .Y(n_744) );
OAI33xp33_ASAP7_75t_L g856 ( .A1(n_689), .A2(n_719), .A3(n_857), .B1(n_863), .B2(n_870), .B3(n_872), .Y(n_856) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_689), .Y(n_893) );
OAI33xp33_ASAP7_75t_L g1003 ( .A1(n_689), .A2(n_719), .A3(n_1004), .B1(n_1009), .B2(n_1012), .B3(n_1014), .Y(n_1003) );
OAI33xp33_ASAP7_75t_L g1228 ( .A1(n_689), .A2(n_914), .A3(n_1229), .B1(n_1234), .B2(n_1239), .B3(n_1240), .Y(n_1228) );
OAI33xp33_ASAP7_75t_L g1341 ( .A1(n_689), .A2(n_719), .A3(n_1342), .B1(n_1347), .B2(n_1351), .B3(n_1357), .Y(n_1341) );
OAI33xp33_ASAP7_75t_L g1449 ( .A1(n_689), .A2(n_719), .A3(n_1450), .B1(n_1453), .B2(n_1456), .B3(n_1459), .Y(n_1449) );
OAI33xp33_ASAP7_75t_L g1486 ( .A1(n_689), .A2(n_719), .A3(n_1487), .B1(n_1491), .B2(n_1494), .B3(n_1498), .Y(n_1486) );
OAI22xp5_ASAP7_75t_L g1534 ( .A1(n_689), .A2(n_719), .B1(n_1535), .B2(n_1540), .Y(n_1534) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_699), .B2(n_700), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g1450 ( .A1(n_694), .A2(n_1137), .B1(n_1451), .B2(n_1452), .Y(n_1450) );
OAI22xp5_ASAP7_75t_L g1456 ( .A1(n_694), .A2(n_751), .B1(n_1457), .B2(n_1458), .Y(n_1456) );
OAI22xp5_ASAP7_75t_L g1939 ( .A1(n_694), .A2(n_1940), .B1(n_1941), .B2(n_1942), .Y(n_1939) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g713 ( .A(n_695), .Y(n_713) );
INVx2_ASAP7_75t_L g865 ( .A(n_695), .Y(n_865) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx2_ASAP7_75t_L g1496 ( .A(n_696), .Y(n_1496) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
BUFx3_ASAP7_75t_L g770 ( .A(n_697), .Y(n_770) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g749 ( .A(n_698), .Y(n_749) );
BUFx2_ASAP7_75t_L g1147 ( .A(n_698), .Y(n_1147) );
OAI22xp33_ASAP7_75t_L g1498 ( .A1(n_700), .A2(n_1489), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
CKINVDCx5p33_ASAP7_75t_R g700 ( .A(n_701), .Y(n_700) );
OAI22xp33_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_706), .B2(n_707), .Y(n_702) );
OAI221xp5_ASAP7_75t_L g1943 ( .A1(n_704), .A2(n_1643), .B1(n_1916), .B2(n_1917), .C(n_1944), .Y(n_1943) );
BUFx2_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g755 ( .A(n_705), .Y(n_755) );
INVx1_ASAP7_75t_L g763 ( .A(n_705), .Y(n_763) );
OAI22xp33_ASAP7_75t_L g909 ( .A1(n_705), .A2(n_910), .B1(n_911), .B2(n_913), .Y(n_909) );
OAI22xp33_ASAP7_75t_L g1061 ( .A1(n_705), .A2(n_709), .B1(n_1030), .B2(n_1062), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1068 ( .A1(n_705), .A2(n_709), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
OAI22xp5_ASAP7_75t_SL g1149 ( .A1(n_705), .A2(n_873), .B1(n_1150), .B2(n_1151), .Y(n_1149) );
OAI22xp33_ASAP7_75t_L g1494 ( .A1(n_705), .A2(n_1495), .B1(n_1496), .B2(n_1497), .Y(n_1494) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g1489 ( .A(n_708), .Y(n_1489) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g718 ( .A(n_709), .Y(n_718) );
INVx3_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
BUFx2_ASAP7_75t_L g766 ( .A(n_710), .Y(n_766) );
INVx2_ASAP7_75t_L g912 ( .A(n_710), .Y(n_912) );
INVx2_ASAP7_75t_L g1944 ( .A(n_710), .Y(n_1944) );
OAI22xp33_ASAP7_75t_SL g898 ( .A1(n_716), .A2(n_899), .B1(n_900), .B2(n_902), .Y(n_898) );
OAI22xp33_ASAP7_75t_L g1459 ( .A1(n_716), .A2(n_718), .B1(n_1460), .B2(n_1461), .Y(n_1459) );
OAI22xp33_ASAP7_75t_L g1487 ( .A1(n_716), .A2(n_1488), .B1(n_1489), .B2(n_1490), .Y(n_1487) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g1014 ( .A1(n_718), .A2(n_754), .B1(n_976), .B2(n_989), .Y(n_1014) );
INVx1_ASAP7_75t_L g1414 ( .A(n_719), .Y(n_1414) );
CKINVDCx8_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g891 ( .A(n_723), .Y(n_891) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_724), .Y(n_854) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g1227 ( .A(n_727), .Y(n_1227) );
HB1xp67_ASAP7_75t_L g1398 ( .A(n_727), .Y(n_1398) );
BUFx4f_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
BUFx4f_ASAP7_75t_L g775 ( .A(n_728), .Y(n_775) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x6_ASAP7_75t_L g1636 ( .A(n_730), .B(n_1620), .Y(n_1636) );
BUFx3_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g855 ( .A(n_732), .Y(n_855) );
BUFx2_ASAP7_75t_L g1002 ( .A(n_732), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_737), .Y(n_733) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_743), .B(n_783), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_774), .C(n_776), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_750), .B2(n_751), .Y(n_745) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_748), .A2(n_772), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
HB1xp67_ASAP7_75t_L g1236 ( .A(n_749), .Y(n_1236) );
OAI22xp5_ASAP7_75t_L g1143 ( .A1(n_751), .A2(n_1144), .B1(n_1145), .B2(n_1148), .Y(n_1143) );
INVx2_ASAP7_75t_L g1283 ( .A(n_751), .Y(n_1283) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_756), .B2(n_757), .Y(n_752) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g1453 ( .A1(n_757), .A2(n_1230), .B1(n_1454), .B2(n_1455), .Y(n_1453) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx2_ASAP7_75t_L g873 ( .A(n_758), .Y(n_873) );
INVx2_ASAP7_75t_L g1359 ( .A(n_758), .Y(n_1359) );
INVx2_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
BUFx3_ASAP7_75t_L g1142 ( .A(n_759), .Y(n_1142) );
OAI22xp5_ASAP7_75t_L g1278 ( .A1(n_759), .A2(n_860), .B1(n_1279), .B2(n_1280), .Y(n_1278) );
BUFx6f_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_764), .B1(n_765), .B2(n_767), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g857 ( .A1(n_765), .A2(n_858), .B1(n_861), .B2(n_862), .Y(n_857) );
OAI22xp33_ASAP7_75t_L g1004 ( .A1(n_765), .A2(n_1005), .B1(n_1007), .B2(n_1008), .Y(n_1004) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
OAI22xp5_ASAP7_75t_L g768 ( .A1(n_769), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_768) );
INVx2_ASAP7_75t_L g901 ( .A(n_769), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_769), .A2(n_966), .B1(n_990), .B2(n_1013), .Y(n_1012) );
OAI22xp5_ASAP7_75t_L g1134 ( .A1(n_769), .A2(n_1135), .B1(n_1136), .B2(n_1137), .Y(n_1134) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
INVx2_ASAP7_75t_SL g905 ( .A(n_770), .Y(n_905) );
INVx2_ASAP7_75t_L g1049 ( .A(n_770), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_780), .Y(n_776) );
NAND4xp25_ASAP7_75t_L g784 ( .A(n_785), .B(n_792), .C(n_804), .D(n_805), .Y(n_784) );
INVx1_ASAP7_75t_L g979 ( .A(n_787), .Y(n_979) );
INVx1_ASAP7_75t_L g1079 ( .A(n_787), .Y(n_1079) );
BUFx2_ASAP7_75t_L g1920 ( .A(n_787), .Y(n_1920) );
A2O1A1Ixp33_ASAP7_75t_L g1558 ( .A1(n_788), .A2(n_927), .B(n_1087), .C(n_1531), .Y(n_1558) );
HB1xp67_ASAP7_75t_L g1998 ( .A(n_788), .Y(n_1998) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_794), .B(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
HB1xp67_ASAP7_75t_L g1433 ( .A(n_800), .Y(n_1433) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
AOI22xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_874), .B1(n_950), .B2(n_951), .Y(n_809) );
INVx1_ASAP7_75t_L g950 ( .A(n_810), .Y(n_950) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_813), .B(n_844), .Y(n_812) );
NAND3xp33_ASAP7_75t_SL g814 ( .A(n_815), .B(n_819), .C(n_832), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g872 ( .A1(n_816), .A2(n_841), .B1(n_858), .B2(n_873), .Y(n_872) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_817), .A2(n_820), .B1(n_865), .B2(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g1184 ( .A(n_824), .Y(n_1184) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
OAI221xp5_ASAP7_75t_L g1550 ( .A1(n_827), .A2(n_984), .B1(n_1536), .B2(n_1551), .C(n_1552), .Y(n_1550) );
AOI22xp33_ASAP7_75t_L g1155 ( .A1(n_836), .A2(n_1148), .B1(n_1150), .B2(n_1156), .Y(n_1155) );
INVx4_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g1084 ( .A(n_837), .Y(n_1084) );
INVx2_ASAP7_75t_L g1213 ( .A(n_837), .Y(n_1213) );
INVx1_ASAP7_75t_L g1564 ( .A(n_838), .Y(n_1564) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
AOI21xp5_ASAP7_75t_L g1193 ( .A1(n_843), .A2(n_1194), .B(n_1195), .Y(n_1193) );
NOR3xp33_ASAP7_75t_L g844 ( .A(n_845), .B(n_853), .C(n_856), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_846), .B(n_849), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_852), .A2(n_1205), .B1(n_1221), .B2(n_1222), .Y(n_1220) );
INVx1_ASAP7_75t_L g1391 ( .A(n_852), .Y(n_1391) );
INVx2_ASAP7_75t_SL g858 ( .A(n_859), .Y(n_858) );
INVx2_ASAP7_75t_SL g859 ( .A(n_860), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B1(n_866), .B2(n_867), .Y(n_863) );
OAI221xp5_ASAP7_75t_L g1947 ( .A1(n_865), .A2(n_1948), .B1(n_1949), .B2(n_1953), .C(n_1954), .Y(n_1947) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
HB1xp67_ASAP7_75t_L g1013 ( .A(n_869), .Y(n_1013) );
OAI22xp33_ASAP7_75t_L g894 ( .A1(n_873), .A2(n_895), .B1(n_896), .B2(n_897), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g1229 ( .A1(n_873), .A2(n_1230), .B1(n_1232), .B2(n_1233), .Y(n_1229) );
OAI22xp33_ASAP7_75t_L g1240 ( .A1(n_873), .A2(n_907), .B1(n_1208), .B2(n_1217), .Y(n_1240) );
OAI22xp5_ASAP7_75t_L g1404 ( .A1(n_873), .A2(n_900), .B1(n_1405), .B2(n_1406), .Y(n_1404) );
INVx1_ASAP7_75t_L g951 ( .A(n_874), .Y(n_951) );
HB1xp67_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
XNOR2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g880 ( .A(n_881), .B(n_915), .Y(n_880) );
NOR3xp33_ASAP7_75t_SL g881 ( .A(n_882), .B(n_890), .C(n_892), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g882 ( .A(n_883), .B(n_886), .Y(n_882) );
AOI22xp33_ASAP7_75t_SL g1529 ( .A1(n_889), .A2(n_1071), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
OAI33xp33_ASAP7_75t_L g892 ( .A1(n_893), .A2(n_894), .A3(n_898), .B1(n_903), .B2(n_909), .B3(n_914), .Y(n_892) );
OAI33xp33_ASAP7_75t_L g1399 ( .A1(n_893), .A2(n_1400), .A3(n_1404), .B1(n_1407), .B2(n_1410), .B3(n_1413), .Y(n_1399) );
INVxp67_ASAP7_75t_L g1067 ( .A(n_896), .Y(n_1067) );
OAI221xp5_ASAP7_75t_L g1628 ( .A1(n_896), .A2(n_1049), .B1(n_1574), .B2(n_1578), .C(n_1629), .Y(n_1628) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_900), .A2(n_1050), .B1(n_1408), .B2(n_1409), .Y(n_1407) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_906), .B1(n_907), .B2(n_908), .Y(n_903) );
OAI22xp33_ASAP7_75t_L g1239 ( .A1(n_904), .A2(n_1197), .B1(n_1216), .B2(n_1230), .Y(n_1239) );
BUFx2_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI221xp5_ASAP7_75t_L g1540 ( .A1(n_905), .A2(n_907), .B1(n_1541), .B2(n_1542), .C(n_1543), .Y(n_1540) );
AOI21xp5_ASAP7_75t_L g918 ( .A1(n_906), .A2(n_919), .B(n_921), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_907), .A2(n_1235), .B1(n_1237), .B2(n_1238), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
OR2x2_ASAP7_75t_L g1653 ( .A(n_912), .B(n_1620), .Y(n_1653) );
OR2x6_ASAP7_75t_L g1945 ( .A(n_912), .B(n_1620), .Y(n_1945) );
AOI211xp5_ASAP7_75t_SL g1985 ( .A1(n_919), .A2(n_1986), .B(n_1987), .C(n_1988), .Y(n_1985) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI31xp33_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_926), .A3(n_928), .B(n_932), .Y(n_922) );
INVx1_ASAP7_75t_L g1260 ( .A(n_924), .Y(n_1260) );
INVx1_ASAP7_75t_L g1027 ( .A(n_925), .Y(n_1027) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
OAI221xp5_ASAP7_75t_L g1180 ( .A1(n_930), .A2(n_1181), .B1(n_1182), .B2(n_1183), .C(n_1184), .Y(n_1180) );
BUFx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g1927 ( .A(n_931), .Y(n_1927) );
OR2x6_ASAP7_75t_L g1597 ( .A(n_933), .B(n_1594), .Y(n_1597) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx1_ASAP7_75t_L g1468 ( .A(n_938), .Y(n_1468) );
BUFx2_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
HB1xp67_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g1549 ( .A(n_946), .Y(n_1549) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_953), .B(n_1661), .Y(n_952) );
INVxp67_ASAP7_75t_SL g953 ( .A(n_954), .Y(n_953) );
NOR2xp33_ASAP7_75t_L g954 ( .A(n_955), .B(n_1382), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx2_ASAP7_75t_L g1663 ( .A(n_956), .Y(n_1663) );
AO22x2_ASAP7_75t_L g956 ( .A1(n_957), .A2(n_958), .B1(n_1189), .B2(n_1381), .Y(n_956) );
INVx2_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
XNOR2x1_ASAP7_75t_L g958 ( .A(n_959), .B(n_1016), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
XNOR2x1_ASAP7_75t_L g960 ( .A(n_961), .B(n_1015), .Y(n_960) );
AND2x2_ASAP7_75t_L g961 ( .A(n_962), .B(n_993), .Y(n_961) );
AOI31xp33_ASAP7_75t_L g964 ( .A1(n_965), .A2(n_974), .A3(n_988), .B(n_991), .Y(n_964) );
BUFx3_ASAP7_75t_L g986 ( .A(n_972), .Y(n_986) );
HB1xp67_ASAP7_75t_L g1369 ( .A(n_972), .Y(n_1369) );
INVx1_ASAP7_75t_L g1428 ( .A(n_975), .Y(n_1428) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
OR2x2_ASAP7_75t_L g1967 ( .A(n_979), .B(n_1577), .Y(n_1967) );
HB1xp67_ASAP7_75t_L g980 ( .A(n_981), .Y(n_980) );
AND2x2_ASAP7_75t_L g1910 ( .A(n_981), .B(n_1613), .Y(n_1910) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx1_ASAP7_75t_L g983 ( .A(n_984), .Y(n_983) );
INVx2_ASAP7_75t_SL g1261 ( .A(n_987), .Y(n_1261) );
AOI21xp5_ASAP7_75t_L g1247 ( .A1(n_991), .A2(n_1248), .B(n_1255), .Y(n_1247) );
AOI31xp33_ASAP7_75t_L g1363 ( .A1(n_991), .A2(n_1364), .A3(n_1371), .B(n_1379), .Y(n_1363) );
INVx2_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
OAI31xp33_ASAP7_75t_L g1312 ( .A1(n_992), .A2(n_1313), .A3(n_1314), .B(n_1323), .Y(n_1312) );
NOR3xp33_ASAP7_75t_SL g993 ( .A(n_994), .B(n_1001), .C(n_1003), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_998), .Y(n_994) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1006), .Y(n_1140) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1006), .Y(n_1402) );
OAI22x1_ASAP7_75t_L g1016 ( .A1(n_1017), .A2(n_1018), .B1(n_1123), .B2(n_1188), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
XNOR2x1_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1073), .Y(n_1018) );
XNOR2x1_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1021), .Y(n_1019) );
OR2x2_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1046), .Y(n_1021) );
AOI31xp33_ASAP7_75t_SL g1022 ( .A1(n_1023), .A2(n_1033), .A3(n_1036), .B(n_1044), .Y(n_1022) );
OAI221xp5_ASAP7_75t_L g1375 ( .A1(n_1025), .A2(n_1336), .B1(n_1338), .B2(n_1376), .C(n_1378), .Y(n_1375) );
OAI221xp5_ASAP7_75t_L g1924 ( .A1(n_1025), .A2(n_1925), .B1(n_1926), .B2(n_1928), .C(n_1929), .Y(n_1924) );
INVx2_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
INVx2_ASAP7_75t_L g1078 ( .A(n_1026), .Y(n_1078) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_1026), .Y(n_1171) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1026), .Y(n_1182) );
INVx1_ASAP7_75t_L g1966 ( .A(n_1026), .Y(n_1966) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1038), .B1(n_1041), .B2(n_1043), .Y(n_1036) );
BUFx2_ASAP7_75t_L g1604 ( .A(n_1039), .Y(n_1604) );
INVx2_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx2_ASAP7_75t_L g1044 ( .A(n_1045), .Y(n_1044) );
AOI211xp5_ASAP7_75t_L g1074 ( .A1(n_1045), .A2(n_1075), .B(n_1101), .C(n_1112), .Y(n_1074) );
NOR2xp67_ASAP7_75t_L g1617 ( .A(n_1045), .B(n_1618), .Y(n_1617) );
NAND3xp33_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1063), .C(n_1072), .Y(n_1046) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_1049), .A2(n_1348), .B1(n_1349), .B2(n_1350), .Y(n_1347) );
OAI22xp5_ASAP7_75t_L g1400 ( .A1(n_1050), .A2(n_1401), .B1(n_1402), .B2(n_1403), .Y(n_1400) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx2_ASAP7_75t_SL g1055 ( .A(n_1056), .Y(n_1055) );
INVx2_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g1941 ( .A(n_1060), .Y(n_1941) );
INVx1_ASAP7_75t_L g1065 ( .A(n_1066), .Y(n_1065) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1066), .Y(n_1282) );
AOI22xp5_ASAP7_75t_L g1271 ( .A1(n_1071), .A2(n_1272), .B1(n_1273), .B2(n_1274), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_1071), .A2(n_1111), .B1(n_1310), .B2(n_1311), .Y(n_1309) );
NAND4xp25_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1082), .C(n_1088), .D(n_1094), .Y(n_1075) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1079), .Y(n_1374) );
A2O1A1Ixp33_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1084), .B(n_1085), .C(n_1087), .Y(n_1082) );
OAI211xp5_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1090), .B(n_1092), .C(n_1093), .Y(n_1088) );
OAI211xp5_ASAP7_75t_L g1319 ( .A1(n_1090), .A2(n_1308), .B(n_1320), .C(n_1321), .Y(n_1319) );
BUFx3_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
INVx1_ASAP7_75t_L g1097 ( .A(n_1091), .Y(n_1097) );
OR2x6_ASAP7_75t_L g1586 ( .A(n_1091), .B(n_1577), .Y(n_1586) );
OAI211xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1096), .B(n_1098), .C(n_1100), .Y(n_1094) );
INVx2_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_1099), .Y(n_1161) );
BUFx3_ASAP7_75t_L g1200 ( .A(n_1099), .Y(n_1200) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1127 ( .A(n_1103), .Y(n_1127) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_1107), .A2(n_1108), .B1(n_1110), .B2(n_1111), .Y(n_1106) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1108), .Y(n_1152) );
NAND2xp5_ASAP7_75t_L g1618 ( .A(n_1109), .B(n_1619), .Y(n_1618) );
BUFx2_ASAP7_75t_L g1955 ( .A(n_1109), .Y(n_1955) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1111), .Y(n_1130) );
NAND2xp5_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1121), .Y(n_1112) );
INVx2_ASAP7_75t_L g1188 ( .A(n_1123), .Y(n_1188) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1124), .Y(n_1186) );
NAND3xp33_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1131), .C(n_1153), .Y(n_1124) );
NOR2xp33_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1129), .Y(n_1125) );
NOR2xp33_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1133), .Y(n_1131) );
OAI22xp5_ASAP7_75t_L g1169 ( .A1(n_1136), .A2(n_1139), .B1(n_1170), .B2(n_1172), .Y(n_1169) );
INVx2_ASAP7_75t_L g2020 ( .A(n_1137), .Y(n_2020) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1140), .B1(n_1141), .B2(n_1142), .Y(n_1138) );
BUFx3_ASAP7_75t_L g1346 ( .A(n_1142), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_1144), .A2(n_1151), .B1(n_1160), .B2(n_1162), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1491 ( .A1(n_1145), .A2(n_1350), .B1(n_1492), .B2(n_1493), .Y(n_1491) );
OAI221xp5_ASAP7_75t_L g1535 ( .A1(n_1145), .A2(n_1354), .B1(n_1536), .B2(n_1537), .C(n_1538), .Y(n_1535) );
INVx2_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx2_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
BUFx2_ASAP7_75t_L g1352 ( .A(n_1147), .Y(n_1352) );
OAI31xp33_ASAP7_75t_L g1153 ( .A1(n_1154), .A2(n_1165), .A3(n_1168), .B(n_1185), .Y(n_1153) );
BUFx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx2_ASAP7_75t_L g1157 ( .A(n_1158), .Y(n_1157) );
OR2x6_ASAP7_75t_L g1580 ( .A(n_1158), .B(n_1577), .Y(n_1580) );
OR2x2_ASAP7_75t_L g1963 ( .A(n_1158), .B(n_1577), .Y(n_1963) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
BUFx2_ASAP7_75t_SL g1162 ( .A(n_1163), .Y(n_1162) );
HB1xp67_ASAP7_75t_L g1602 ( .A(n_1163), .Y(n_1602) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1163), .B(n_1613), .Y(n_1612) );
OAI22xp5_ASAP7_75t_L g1168 ( .A1(n_1169), .A2(n_1173), .B1(n_1176), .B2(n_1180), .Y(n_1168) );
OAI21xp5_ASAP7_75t_SL g1990 ( .A1(n_1170), .A2(n_1991), .B(n_1992), .Y(n_1990) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g1516 ( .A(n_1185), .Y(n_1516) );
OAI31xp33_ASAP7_75t_SL g1546 ( .A1(n_1185), .A2(n_1547), .A3(n_1553), .B(n_1557), .Y(n_1546) );
INVx1_ASAP7_75t_SL g1381 ( .A(n_1189), .Y(n_1381) );
XNOR2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1242), .Y(n_1189) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1218), .Y(n_1192) );
AOI211xp5_ASAP7_75t_L g1196 ( .A1(n_1197), .A2(n_1198), .B(n_1199), .C(n_1206), .Y(n_1196) );
AOI21xp5_ASAP7_75t_L g1420 ( .A1(n_1198), .A2(n_1408), .B(n_1421), .Y(n_1420) );
OAI211xp5_ASAP7_75t_L g1315 ( .A1(n_1202), .A2(n_1316), .B(n_1317), .C(n_1318), .Y(n_1315) );
BUFx2_ASAP7_75t_L g1918 ( .A(n_1202), .Y(n_1918) );
HB1xp67_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
NOR3xp33_ASAP7_75t_L g1218 ( .A(n_1219), .B(n_1226), .C(n_1228), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1223), .Y(n_1219) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_1221), .A2(n_1394), .B1(n_1395), .B2(n_1396), .Y(n_1393) );
INVx1_ASAP7_75t_L g2009 ( .A(n_1221), .Y(n_2009) );
INVxp67_ASAP7_75t_SL g1392 ( .A(n_1225), .Y(n_1392) );
AOI22xp33_ASAP7_75t_L g2010 ( .A1(n_1225), .A2(n_1273), .B1(n_2011), .B2(n_2012), .Y(n_2010) );
BUFx2_ASAP7_75t_L g1344 ( .A(n_1230), .Y(n_1344) );
OAI221xp5_ASAP7_75t_L g1640 ( .A1(n_1230), .A2(n_1346), .B1(n_1641), .B2(n_1642), .C(n_1643), .Y(n_1640) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1645 ( .A1(n_1235), .A2(n_1646), .B1(n_1647), .B2(n_1652), .Y(n_1645) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1236), .Y(n_1235) );
AOI22xp5_ASAP7_75t_L g1242 ( .A1(n_1243), .A2(n_1244), .B1(n_1329), .B2(n_1380), .Y(n_1242) );
INVx1_ASAP7_75t_SL g1243 ( .A(n_1244), .Y(n_1243) );
XNOR2x1_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1286), .Y(n_1244) );
NOR2x1_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1264), .Y(n_1246) );
HB1xp67_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
NAND4xp25_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1268), .C(n_1271), .D(n_1275), .Y(n_1264) );
NAND3xp33_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1305), .C(n_1312), .Y(n_1287) );
AND3x1_ASAP7_75t_L g1288 ( .A(n_1289), .B(n_1292), .C(n_1303), .Y(n_1288) );
INVx2_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx2_ASAP7_75t_L g1539 ( .A(n_1295), .Y(n_1539) );
INVx2_ASAP7_75t_SL g1630 ( .A(n_1295), .Y(n_1630) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
INVx2_ASAP7_75t_L g1355 ( .A(n_1298), .Y(n_1355) );
INVx2_ASAP7_75t_SL g1631 ( .A(n_1302), .Y(n_1631) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1309), .Y(n_1305) );
NAND3xp33_ASAP7_75t_L g1314 ( .A(n_1315), .B(n_1319), .C(n_1322), .Y(n_1314) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1327), .Y(n_1554) );
INVx2_ASAP7_75t_L g1380 ( .A(n_1329), .Y(n_1380) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1361), .Y(n_1330) );
NOR3xp33_ASAP7_75t_SL g1331 ( .A(n_1332), .B(n_1340), .C(n_1341), .Y(n_1331) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1337), .Y(n_1332) );
OAI22xp33_ASAP7_75t_L g1342 ( .A1(n_1343), .A2(n_1344), .B1(n_1345), .B2(n_1346), .Y(n_1342) );
OAI22xp33_ASAP7_75t_L g1357 ( .A1(n_1344), .A2(n_1358), .B1(n_1359), .B2(n_1360), .Y(n_1357) );
OAI22xp33_ASAP7_75t_L g1410 ( .A1(n_1346), .A2(n_1402), .B1(n_1411), .B2(n_1412), .Y(n_1410) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_1352), .A2(n_1353), .B1(n_1354), .B2(n_1356), .Y(n_1351) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1377), .Y(n_1510) );
INVx2_ASAP7_75t_SL g1551 ( .A(n_1377), .Y(n_1551) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1378), .Y(n_1425) );
AND2x2_ASAP7_75t_L g1662 ( .A(n_1382), .B(n_1663), .Y(n_1662) );
AO22x1_ASAP7_75t_L g1382 ( .A1(n_1383), .A2(n_1384), .B1(n_1519), .B2(n_1660), .Y(n_1382) );
INVx2_ASAP7_75t_L g1383 ( .A(n_1384), .Y(n_1383) );
XNOR2x1_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1437), .Y(n_1384) );
INVx2_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
XNOR2x1_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1388), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1415), .Y(n_1388) );
NOR3xp33_ASAP7_75t_SL g1389 ( .A(n_1390), .B(n_1397), .C(n_1399), .Y(n_1389) );
AOI221xp5_ASAP7_75t_L g1426 ( .A1(n_1412), .A2(n_1427), .B1(n_1429), .B2(n_1432), .C(n_1434), .Y(n_1426) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1414), .Y(n_1413) );
AOI33xp33_ASAP7_75t_L g2014 ( .A1(n_1414), .A2(n_2015), .A3(n_2017), .B1(n_2021), .B2(n_2024), .B3(n_2025), .Y(n_2014) );
AOI21xp5_ASAP7_75t_L g1415 ( .A1(n_1416), .A2(n_1418), .B(n_1419), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1417), .Y(n_1416) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
XOR2x2_ASAP7_75t_L g1437 ( .A(n_1438), .B(n_1475), .Y(n_1437) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1462), .Y(n_1439) );
NOR3xp33_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1448), .C(n_1449), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1445), .Y(n_1441) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1476), .Y(n_1518) );
AND2x2_ASAP7_75t_L g1476 ( .A(n_1477), .B(n_1501), .Y(n_1476) );
NOR3xp33_ASAP7_75t_L g1477 ( .A(n_1478), .B(n_1485), .C(n_1486), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1482), .Y(n_1478) );
AOI31xp33_ASAP7_75t_L g1503 ( .A1(n_1504), .A2(n_1511), .A3(n_1515), .B(n_1516), .Y(n_1503) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1508), .Y(n_1507) );
INVxp67_ASAP7_75t_SL g1660 ( .A(n_1519), .Y(n_1660) );
AOI22xp33_ASAP7_75t_L g1519 ( .A1(n_1520), .A2(n_1521), .B1(n_1569), .B2(n_1659), .Y(n_1519) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
HB1xp67_ASAP7_75t_L g1522 ( .A(n_1523), .Y(n_1522) );
NAND4xp25_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1532), .C(n_1546), .D(n_1566), .Y(n_1524) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1529), .Y(n_1525) );
BUFx6f_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
AND2x4_ASAP7_75t_L g1625 ( .A(n_1545), .B(n_1626), .Y(n_1625) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
NAND3xp33_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1559), .C(n_1562), .Y(n_1557) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1569), .Y(n_1659) );
NAND3xp33_ASAP7_75t_L g1570 ( .A(n_1571), .B(n_1614), .C(n_1622), .Y(n_1570) );
NOR2xp33_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1587), .Y(n_1571) );
NAND2xp5_ASAP7_75t_L g1572 ( .A(n_1573), .B(n_1581), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1573 ( .A1(n_1574), .A2(n_1575), .B1(n_1578), .B2(n_1579), .Y(n_1573) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1577), .Y(n_1576) );
OR2x2_ASAP7_75t_L g1965 ( .A(n_1577), .B(n_1966), .Y(n_1965) );
CKINVDCx6p67_ASAP7_75t_R g1579 ( .A(n_1580), .Y(n_1579) );
AOI22xp33_ASAP7_75t_L g1581 ( .A1(n_1582), .A2(n_1583), .B1(n_1584), .B2(n_1585), .Y(n_1581) );
CKINVDCx6p67_ASAP7_75t_R g1585 ( .A(n_1586), .Y(n_1585) );
NAND3xp33_ASAP7_75t_SL g1587 ( .A(n_1588), .B(n_1598), .C(n_1610), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1588 ( .A1(n_1589), .A2(n_1590), .B1(n_1595), .B2(n_1596), .Y(n_1588) );
AOI22xp33_ASAP7_75t_L g1632 ( .A1(n_1589), .A2(n_1595), .B1(n_1633), .B2(n_1635), .Y(n_1632) );
INVx2_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
HB1xp67_ASAP7_75t_L g1933 ( .A(n_1591), .Y(n_1933) );
NAND2x1p5_ASAP7_75t_L g1591 ( .A(n_1592), .B(n_1593), .Y(n_1591) );
INVx2_ASAP7_75t_SL g1593 ( .A(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1594), .Y(n_1613) );
INVx2_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
AOI33xp33_ASAP7_75t_L g1598 ( .A1(n_1599), .A2(n_1601), .A3(n_1603), .B1(n_1605), .B2(n_1606), .B3(n_1609), .Y(n_1598) );
CKINVDCx5p33_ASAP7_75t_R g1599 ( .A(n_1600), .Y(n_1599) );
OAI22xp5_ASAP7_75t_SL g1911 ( .A1(n_1600), .A2(n_1912), .B1(n_1923), .B2(n_1924), .Y(n_1911) );
INVx1_ASAP7_75t_L g1607 ( .A(n_1608), .Y(n_1607) );
INVx4_ASAP7_75t_L g1923 ( .A(n_1609), .Y(n_1923) );
INVx1_ASAP7_75t_L g1610 ( .A(n_1611), .Y(n_1610) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_1615), .B(n_1616), .Y(n_1614) );
NAND2xp5_ASAP7_75t_L g1934 ( .A(n_1616), .B(n_1935), .Y(n_1934) );
INVx1_ASAP7_75t_L g1619 ( .A(n_1620), .Y(n_1619) );
INVx2_ASAP7_75t_L g1620 ( .A(n_1621), .Y(n_1620) );
INVx8_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
AND2x4_ASAP7_75t_L g1658 ( .A(n_1626), .B(n_1650), .Y(n_1658) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1627), .Y(n_1626) );
HB1xp67_ASAP7_75t_L g1633 ( .A(n_1634), .Y(n_1633) );
AOI22xp33_ASAP7_75t_L g1957 ( .A1(n_1635), .A2(n_1958), .B1(n_1959), .B2(n_1960), .Y(n_1957) );
CKINVDCx11_ASAP7_75t_R g1635 ( .A(n_1636), .Y(n_1635) );
CKINVDCx6p67_ASAP7_75t_R g1638 ( .A(n_1639), .Y(n_1638) );
INVx2_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1648), .Y(n_1647) );
INVx1_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
INVx1_ASAP7_75t_L g1649 ( .A(n_1650), .Y(n_1649) );
INVx2_ASAP7_75t_L g1650 ( .A(n_1651), .Y(n_1650) );
INVx1_ASAP7_75t_L g1952 ( .A(n_1651), .Y(n_1952) );
INVx3_ASAP7_75t_L g1655 ( .A(n_1656), .Y(n_1655) );
INVx3_ASAP7_75t_L g1657 ( .A(n_1658), .Y(n_1657) );
INVx1_ASAP7_75t_L g1661 ( .A(n_1662), .Y(n_1661) );
OAI221xp5_ASAP7_75t_L g1664 ( .A1(n_1665), .A2(n_1902), .B1(n_1903), .B2(n_1968), .C(n_1974), .Y(n_1664) );
AOI311xp33_ASAP7_75t_L g1665 ( .A1(n_1666), .A2(n_1761), .A3(n_1789), .B(n_1796), .C(n_1868), .Y(n_1665) );
OAI211xp5_ASAP7_75t_L g1666 ( .A1(n_1667), .A2(n_1695), .B(n_1721), .C(n_1747), .Y(n_1666) );
A2O1A1Ixp33_ASAP7_75t_L g1721 ( .A1(n_1667), .A2(n_1722), .B(n_1726), .C(n_1732), .Y(n_1721) );
INVx1_ASAP7_75t_L g1667 ( .A(n_1668), .Y(n_1667) );
NAND2xp5_ASAP7_75t_L g1813 ( .A(n_1668), .B(n_1814), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1895 ( .A(n_1668), .B(n_1790), .Y(n_1895) );
INVx1_ASAP7_75t_L g1668 ( .A(n_1669), .Y(n_1668) );
INVx2_ASAP7_75t_SL g1737 ( .A(n_1669), .Y(n_1737) );
AND2x2_ASAP7_75t_L g1772 ( .A(n_1669), .B(n_1729), .Y(n_1772) );
AND2x4_ASAP7_75t_L g1786 ( .A(n_1669), .B(n_1728), .Y(n_1786) );
NAND2xp5_ASAP7_75t_L g1811 ( .A(n_1669), .B(n_1790), .Y(n_1811) );
AND2x2_ASAP7_75t_L g1817 ( .A(n_1669), .B(n_1818), .Y(n_1817) );
NOR2xp33_ASAP7_75t_L g1859 ( .A(n_1669), .B(n_1818), .Y(n_1859) );
HB1xp67_ASAP7_75t_L g1886 ( .A(n_1669), .Y(n_1886) );
CKINVDCx5p33_ASAP7_75t_R g1669 ( .A(n_1670), .Y(n_1669) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1670), .B(n_1729), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1824 ( .A(n_1670), .B(n_1728), .Y(n_1824) );
OR2x2_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1685), .Y(n_1670) );
OAI22xp5_ASAP7_75t_L g1671 ( .A1(n_1672), .A2(n_1679), .B1(n_1680), .B2(n_1684), .Y(n_1671) );
BUFx3_ASAP7_75t_L g1758 ( .A(n_1672), .Y(n_1758) );
BUFx6f_ASAP7_75t_L g1672 ( .A(n_1673), .Y(n_1672) );
OAI22xp5_ASAP7_75t_L g1718 ( .A1(n_1673), .A2(n_1682), .B1(n_1719), .B2(n_1720), .Y(n_1718) );
OR2x2_ASAP7_75t_L g1673 ( .A(n_1674), .B(n_1675), .Y(n_1673) );
OR2x2_ASAP7_75t_L g1682 ( .A(n_1674), .B(n_1683), .Y(n_1682) );
INVx1_ASAP7_75t_L g1702 ( .A(n_1674), .Y(n_1702) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1675), .Y(n_1701) );
NAND2xp5_ASAP7_75t_L g1675 ( .A(n_1676), .B(n_1678), .Y(n_1675) );
HB1xp67_ASAP7_75t_L g2032 ( .A(n_1676), .Y(n_2032) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1678), .Y(n_1689) );
HB1xp67_ASAP7_75t_L g1760 ( .A(n_1680), .Y(n_1760) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
INVx1_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1683), .Y(n_1704) );
OAI22xp5_ASAP7_75t_L g1685 ( .A1(n_1686), .A2(n_1691), .B1(n_1692), .B2(n_1694), .Y(n_1685) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
BUFx3_ASAP7_75t_L g1755 ( .A(n_1687), .Y(n_1755) );
AND2x4_ASAP7_75t_L g1687 ( .A(n_1688), .B(n_1690), .Y(n_1687) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1688), .B(n_1690), .Y(n_1711) );
HB1xp67_ASAP7_75t_L g2033 ( .A(n_1688), .Y(n_2033) );
INVx1_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
AND2x4_ASAP7_75t_L g1693 ( .A(n_1689), .B(n_1690), .Y(n_1693) );
INVx2_ASAP7_75t_L g1754 ( .A(n_1692), .Y(n_1754) );
INVx2_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1706), .Y(n_1695) );
NAND2xp5_ASAP7_75t_L g1723 ( .A(n_1696), .B(n_1724), .Y(n_1723) );
OAI321xp33_ASAP7_75t_SL g1809 ( .A1(n_1696), .A2(n_1810), .A3(n_1811), .B1(n_1812), .B2(n_1813), .C(n_1815), .Y(n_1809) );
NAND2xp5_ASAP7_75t_L g1821 ( .A(n_1696), .B(n_1739), .Y(n_1821) );
INVx2_ASAP7_75t_L g1696 ( .A(n_1697), .Y(n_1696) );
NAND2xp5_ASAP7_75t_L g1808 ( .A(n_1697), .B(n_1712), .Y(n_1808) );
NAND2xp5_ASAP7_75t_SL g1843 ( .A(n_1697), .B(n_1844), .Y(n_1843) );
AND2x2_ASAP7_75t_L g1874 ( .A(n_1697), .B(n_1772), .Y(n_1874) );
BUFx2_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1698), .B(n_1736), .Y(n_1735) );
INVx2_ASAP7_75t_L g1743 ( .A(n_1698), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1764 ( .A(n_1698), .B(n_1765), .Y(n_1764) );
OR2x2_ASAP7_75t_L g1782 ( .A(n_1698), .B(n_1770), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1698), .B(n_1725), .Y(n_1801) );
INVx2_ASAP7_75t_L g1818 ( .A(n_1698), .Y(n_1818) );
AND2x2_ASAP7_75t_L g1698 ( .A(n_1699), .B(n_1705), .Y(n_1698) );
AND2x4_ASAP7_75t_L g1700 ( .A(n_1701), .B(n_1702), .Y(n_1700) );
AND2x4_ASAP7_75t_L g1703 ( .A(n_1702), .B(n_1704), .Y(n_1703) );
BUFx2_ASAP7_75t_L g1794 ( .A(n_1703), .Y(n_1794) );
INVx2_ASAP7_75t_L g1748 ( .A(n_1706), .Y(n_1748) );
NAND2xp5_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1712), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1707), .B(n_1735), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1707), .B(n_1745), .Y(n_1744) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1707), .B(n_1740), .Y(n_1765) );
AND2x2_ASAP7_75t_L g1771 ( .A(n_1707), .B(n_1750), .Y(n_1771) );
INVxp67_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
BUFx2_ASAP7_75t_L g1725 ( .A(n_1708), .Y(n_1725) );
BUFx3_ASAP7_75t_L g1770 ( .A(n_1708), .Y(n_1770) );
OR2x2_ASAP7_75t_L g1854 ( .A(n_1708), .B(n_1717), .Y(n_1854) );
AND2x2_ASAP7_75t_L g1708 ( .A(n_1709), .B(n_1710), .Y(n_1708) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1712), .B(n_1770), .Y(n_1769) );
NOR2xp33_ASAP7_75t_L g1852 ( .A(n_1712), .B(n_1853), .Y(n_1852) );
INVx1_ASAP7_75t_L g1863 ( .A(n_1712), .Y(n_1863) );
NAND3xp33_ASAP7_75t_SL g1881 ( .A(n_1712), .B(n_1742), .C(n_1805), .Y(n_1881) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1713), .B(n_1716), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1736 ( .A(n_1713), .B(n_1717), .Y(n_1736) );
INVx2_ASAP7_75t_L g1741 ( .A(n_1713), .Y(n_1741) );
OR2x2_ASAP7_75t_L g1746 ( .A(n_1713), .B(n_1717), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_1713), .B(n_1770), .Y(n_1816) );
NOR2xp33_ASAP7_75t_L g1844 ( .A(n_1713), .B(n_1770), .Y(n_1844) );
AND2x2_ASAP7_75t_L g1713 ( .A(n_1714), .B(n_1715), .Y(n_1713) );
NOR2x1_ASAP7_75t_L g1724 ( .A(n_1716), .B(n_1725), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1867 ( .A(n_1716), .B(n_1770), .Y(n_1867) );
INVx2_ASAP7_75t_SL g1716 ( .A(n_1717), .Y(n_1716) );
AND2x2_ASAP7_75t_L g1740 ( .A(n_1717), .B(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
NOR2xp33_ASAP7_75t_L g1879 ( .A(n_1723), .B(n_1826), .Y(n_1879) );
INVx1_ASAP7_75t_L g1865 ( .A(n_1724), .Y(n_1865) );
AND2x2_ASAP7_75t_L g1739 ( .A(n_1725), .B(n_1740), .Y(n_1739) );
AND2x2_ASAP7_75t_L g1788 ( .A(n_1725), .B(n_1736), .Y(n_1788) );
A2O1A1Ixp33_ASAP7_75t_L g1732 ( .A1(n_1726), .A2(n_1733), .B(n_1737), .C(n_1738), .Y(n_1732) );
OAI221xp5_ASAP7_75t_L g1773 ( .A1(n_1726), .A2(n_1727), .B1(n_1774), .B2(n_1776), .C(n_1778), .Y(n_1773) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
AOI22xp33_ASAP7_75t_L g1883 ( .A1(n_1727), .A2(n_1762), .B1(n_1824), .B2(n_1884), .Y(n_1883) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1728), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1814 ( .A(n_1728), .B(n_1792), .Y(n_1814) );
OR2x2_ASAP7_75t_L g1826 ( .A(n_1728), .B(n_1827), .Y(n_1826) );
INVx3_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
OR2x2_ASAP7_75t_L g1850 ( .A(n_1729), .B(n_1792), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1891 ( .A(n_1729), .B(n_1791), .Y(n_1891) );
AND2x2_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1731), .Y(n_1729) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1735), .Y(n_1812) );
O2A1O1Ixp33_ASAP7_75t_L g1869 ( .A1(n_1735), .A2(n_1870), .B(n_1871), .C(n_1872), .Y(n_1869) );
INVx1_ASAP7_75t_L g1775 ( .A(n_1736), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1736), .B(n_1743), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1742 ( .A(n_1737), .B(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1763 ( .A(n_1737), .Y(n_1763) );
NOR2xp33_ASAP7_75t_L g1780 ( .A(n_1737), .B(n_1781), .Y(n_1780) );
NOR2xp33_ASAP7_75t_L g1840 ( .A(n_1737), .B(n_1826), .Y(n_1840) );
INVx2_ASAP7_75t_L g1848 ( .A(n_1737), .Y(n_1848) );
AOI21xp33_ASAP7_75t_SL g1738 ( .A1(n_1739), .A2(n_1742), .B(n_1744), .Y(n_1738) );
OAI211xp5_ASAP7_75t_L g1837 ( .A1(n_1739), .A2(n_1818), .B(n_1824), .C(n_1838), .Y(n_1837) );
A2O1A1Ixp33_ASAP7_75t_SL g1882 ( .A1(n_1739), .A2(n_1856), .B(n_1883), .C(n_1888), .Y(n_1882) );
AND2x2_ASAP7_75t_L g1800 ( .A(n_1740), .B(n_1801), .Y(n_1800) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1740), .Y(n_1832) );
NAND2xp5_ASAP7_75t_L g1810 ( .A(n_1741), .B(n_1770), .Y(n_1810) );
OAI321xp33_ASAP7_75t_L g1872 ( .A1(n_1741), .A2(n_1861), .A3(n_1873), .B1(n_1875), .B2(n_1876), .C(n_1878), .Y(n_1872) );
NOR2xp33_ASAP7_75t_L g1745 ( .A(n_1743), .B(n_1746), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1743), .B(n_1750), .Y(n_1749) );
AND2x2_ASAP7_75t_L g1877 ( .A(n_1743), .B(n_1816), .Y(n_1877) );
INVx1_ASAP7_75t_L g1887 ( .A(n_1744), .Y(n_1887) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1746), .Y(n_1750) );
OR2x2_ASAP7_75t_L g1781 ( .A(n_1746), .B(n_1782), .Y(n_1781) );
NOR2xp33_ASAP7_75t_L g1822 ( .A(n_1746), .B(n_1823), .Y(n_1822) );
O2A1O1Ixp33_ASAP7_75t_L g1747 ( .A1(n_1748), .A2(n_1749), .B(n_1751), .C(n_1752), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1870 ( .A(n_1749), .B(n_1770), .Y(n_1870) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1750), .B(n_1801), .Y(n_1849) );
CKINVDCx5p33_ASAP7_75t_R g1806 ( .A(n_1751), .Y(n_1806) );
AOI211xp5_ASAP7_75t_SL g1819 ( .A1(n_1751), .A2(n_1820), .B(n_1822), .C(n_1825), .Y(n_1819) );
NAND4xp25_ASAP7_75t_L g1899 ( .A(n_1751), .B(n_1801), .C(n_1838), .D(n_1900), .Y(n_1899) );
INVx3_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
INVx3_ASAP7_75t_L g1778 ( .A(n_1753), .Y(n_1778) );
A2O1A1Ixp33_ASAP7_75t_SL g1796 ( .A1(n_1753), .A2(n_1797), .B(n_1819), .C(n_1835), .Y(n_1796) );
AND2x2_ASAP7_75t_L g1856 ( .A(n_1753), .B(n_1857), .Y(n_1856) );
CKINVDCx5p33_ASAP7_75t_R g1902 ( .A(n_1755), .Y(n_1902) );
OAI22xp33_ASAP7_75t_L g1756 ( .A1(n_1757), .A2(n_1758), .B1(n_1759), .B2(n_1760), .Y(n_1756) );
NAND4xp25_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1766), .C(n_1779), .D(n_1783), .Y(n_1761) );
OR2x2_ASAP7_75t_L g1762 ( .A(n_1763), .B(n_1764), .Y(n_1762) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1764), .Y(n_1890) );
AOI21xp33_ASAP7_75t_L g1766 ( .A1(n_1767), .A2(n_1772), .B(n_1773), .Y(n_1766) );
INVx1_ASAP7_75t_L g1767 ( .A(n_1768), .Y(n_1767) );
NOR2xp33_ASAP7_75t_L g1768 ( .A(n_1769), .B(n_1771), .Y(n_1768) );
OR2x2_ASAP7_75t_L g1774 ( .A(n_1770), .B(n_1775), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1829 ( .A(n_1770), .B(n_1777), .Y(n_1829) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1771), .Y(n_1860) );
AOI221xp5_ASAP7_75t_L g1797 ( .A1(n_1772), .A2(n_1798), .B1(n_1802), .B2(n_1807), .C(n_1809), .Y(n_1797) );
AOI21xp5_ASAP7_75t_L g1888 ( .A1(n_1772), .A2(n_1786), .B(n_1828), .Y(n_1888) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1774), .Y(n_1845) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1778), .B(n_1790), .Y(n_1789) );
O2A1O1Ixp33_ASAP7_75t_L g1846 ( .A1(n_1778), .A2(n_1808), .B(n_1847), .C(n_1850), .Y(n_1846) );
OAI211xp5_ASAP7_75t_L g1868 ( .A1(n_1778), .A2(n_1869), .B(n_1882), .C(n_1889), .Y(n_1868) );
INVxp67_ASAP7_75t_SL g1779 ( .A(n_1780), .Y(n_1779) );
O2A1O1Ixp33_ASAP7_75t_L g1889 ( .A1(n_1780), .A2(n_1890), .B(n_1891), .C(n_1892), .Y(n_1889) );
NAND2xp5_ASAP7_75t_L g1798 ( .A(n_1781), .B(n_1799), .Y(n_1798) );
NOR2xp33_ASAP7_75t_L g1898 ( .A(n_1781), .B(n_1886), .Y(n_1898) );
OR2x2_ASAP7_75t_L g1862 ( .A(n_1782), .B(n_1863), .Y(n_1862) );
INVxp67_ASAP7_75t_L g1783 ( .A(n_1784), .Y(n_1783) );
NOR2xp33_ASAP7_75t_L g1784 ( .A(n_1785), .B(n_1787), .Y(n_1784) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
AND2x2_ASAP7_75t_L g1834 ( .A(n_1786), .B(n_1790), .Y(n_1834) );
INVx1_ASAP7_75t_L g1787 ( .A(n_1788), .Y(n_1787) );
OAI332xp33_ASAP7_75t_L g1851 ( .A1(n_1789), .A2(n_1848), .A3(n_1852), .B1(n_1855), .B2(n_1858), .B3(n_1860), .C1(n_1861), .C2(n_1862), .Y(n_1851) );
INVx2_ASAP7_75t_L g1838 ( .A(n_1790), .Y(n_1838) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1791), .Y(n_1805) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1792), .Y(n_1791) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1792), .Y(n_1827) );
INVx1_ASAP7_75t_L g1875 ( .A(n_1792), .Y(n_1875) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1793), .B(n_1795), .Y(n_1792) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
NAND2xp5_ASAP7_75t_L g1839 ( .A(n_1800), .B(n_1840), .Y(n_1839) );
INVx1_ASAP7_75t_L g1802 ( .A(n_1803), .Y(n_1802) );
OR2x2_ASAP7_75t_L g1803 ( .A(n_1804), .B(n_1806), .Y(n_1803) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1805), .Y(n_1804) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1805), .Y(n_1857) );
AOI211xp5_ASAP7_75t_L g1864 ( .A1(n_1805), .A2(n_1823), .B(n_1865), .C(n_1866), .Y(n_1864) );
INVx1_ASAP7_75t_L g1807 ( .A(n_1808), .Y(n_1807) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1811), .Y(n_1871) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1814), .Y(n_1861) );
NAND2xp5_ASAP7_75t_L g1815 ( .A(n_1816), .B(n_1817), .Y(n_1815) );
NAND2xp5_ASAP7_75t_L g1823 ( .A(n_1818), .B(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1820 ( .A(n_1821), .Y(n_1820) );
OAI21xp33_ASAP7_75t_L g1825 ( .A1(n_1826), .A2(n_1828), .B(n_1830), .Y(n_1825) );
INVx1_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
INVxp33_ASAP7_75t_L g1830 ( .A(n_1831), .Y(n_1830) );
NOR2xp33_ASAP7_75t_L g1831 ( .A(n_1832), .B(n_1833), .Y(n_1831) );
NAND2xp5_ASAP7_75t_L g1901 ( .A(n_1832), .B(n_1863), .Y(n_1901) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1834), .Y(n_1833) );
OAI21xp5_ASAP7_75t_L g1841 ( .A1(n_1834), .A2(n_1842), .B(n_1845), .Y(n_1841) );
NOR4xp25_ASAP7_75t_L g1835 ( .A(n_1836), .B(n_1846), .C(n_1851), .D(n_1864), .Y(n_1835) );
NAND3xp33_ASAP7_75t_L g1836 ( .A(n_1837), .B(n_1839), .C(n_1841), .Y(n_1836) );
A2O1A1Ixp33_ASAP7_75t_L g1892 ( .A1(n_1838), .A2(n_1893), .B(n_1897), .C(n_1899), .Y(n_1892) );
INVx1_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
NAND2xp5_ASAP7_75t_L g1847 ( .A(n_1848), .B(n_1849), .Y(n_1847) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1854), .Y(n_1853) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1859), .Y(n_1858) );
INVxp67_ASAP7_75t_L g1896 ( .A(n_1862), .Y(n_1896) );
INVx1_ASAP7_75t_L g1866 ( .A(n_1867), .Y(n_1866) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1874), .Y(n_1873) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1877), .Y(n_1876) );
NOR2xp33_ASAP7_75t_L g1878 ( .A(n_1879), .B(n_1880), .Y(n_1878) );
INVx1_ASAP7_75t_L g1880 ( .A(n_1881), .Y(n_1880) );
INVxp33_ASAP7_75t_L g1884 ( .A(n_1885), .Y(n_1884) );
NOR2xp33_ASAP7_75t_L g1885 ( .A(n_1886), .B(n_1887), .Y(n_1885) );
NAND2xp5_ASAP7_75t_L g1893 ( .A(n_1894), .B(n_1896), .Y(n_1893) );
INVx1_ASAP7_75t_L g1894 ( .A(n_1895), .Y(n_1894) );
INVx1_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
INVx1_ASAP7_75t_L g1900 ( .A(n_1901), .Y(n_1900) );
CKINVDCx14_ASAP7_75t_R g1903 ( .A(n_1904), .Y(n_1903) );
HB1xp67_ASAP7_75t_L g1904 ( .A(n_1905), .Y(n_1904) );
INVx1_ASAP7_75t_L g1905 ( .A(n_1906), .Y(n_1905) );
AND4x1_ASAP7_75t_L g1907 ( .A(n_1908), .B(n_1934), .C(n_1936), .D(n_1961), .Y(n_1907) );
NOR3xp33_ASAP7_75t_SL g1908 ( .A(n_1909), .B(n_1911), .C(n_1932), .Y(n_1908) );
BUFx2_ASAP7_75t_L g1909 ( .A(n_1910), .Y(n_1909) );
OAI221xp5_ASAP7_75t_L g1912 ( .A1(n_1913), .A2(n_1916), .B1(n_1917), .B2(n_1918), .C(n_1919), .Y(n_1912) );
BUFx2_ASAP7_75t_L g1913 ( .A(n_1914), .Y(n_1913) );
INVx2_ASAP7_75t_L g1914 ( .A(n_1915), .Y(n_1914) );
INVx1_ASAP7_75t_L g1921 ( .A(n_1922), .Y(n_1921) );
INVx2_ASAP7_75t_L g1926 ( .A(n_1927), .Y(n_1926) );
INVx1_ASAP7_75t_L g1930 ( .A(n_1931), .Y(n_1930) );
INVx1_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
INVx1_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
INVx1_ASAP7_75t_L g1951 ( .A(n_1952), .Y(n_1951) );
NOR2xp33_ASAP7_75t_L g1961 ( .A(n_1962), .B(n_1964), .Y(n_1961) );
CKINVDCx14_ASAP7_75t_R g1968 ( .A(n_1969), .Y(n_1968) );
INVx4_ASAP7_75t_L g1969 ( .A(n_1970), .Y(n_1969) );
INVx1_ASAP7_75t_L g1970 ( .A(n_1971), .Y(n_1970) );
INVx1_ASAP7_75t_L g1971 ( .A(n_1972), .Y(n_1971) );
INVx1_ASAP7_75t_L g1972 ( .A(n_1973), .Y(n_1972) );
HB1xp67_ASAP7_75t_SL g1975 ( .A(n_1976), .Y(n_1975) );
A2O1A1Ixp33_ASAP7_75t_L g2030 ( .A1(n_1977), .A2(n_2031), .B(n_2033), .C(n_2034), .Y(n_2030) );
INVxp33_ASAP7_75t_SL g1978 ( .A(n_1979), .Y(n_1978) );
AND2x2_ASAP7_75t_L g1980 ( .A(n_1981), .B(n_2007), .Y(n_1980) );
AOI21xp5_ASAP7_75t_L g1981 ( .A1(n_1982), .A2(n_1983), .B(n_1984), .Y(n_1981) );
AOI31xp33_ASAP7_75t_L g1984 ( .A1(n_1985), .A2(n_1993), .A3(n_2002), .B(n_2005), .Y(n_1984) );
AOI221xp5_ASAP7_75t_L g1993 ( .A1(n_1994), .A2(n_1996), .B1(n_1997), .B2(n_2000), .C(n_2001), .Y(n_1993) );
CKINVDCx5p33_ASAP7_75t_R g1994 ( .A(n_1995), .Y(n_1994) );
INVx1_ASAP7_75t_SL g2005 ( .A(n_2006), .Y(n_2005) );
NOR2xp33_ASAP7_75t_L g2007 ( .A(n_2008), .B(n_2013), .Y(n_2007) );
NAND2xp5_ASAP7_75t_SL g2013 ( .A(n_2014), .B(n_2026), .Y(n_2013) );
INVx2_ASAP7_75t_L g2015 ( .A(n_2016), .Y(n_2015) );
BUFx3_ASAP7_75t_L g2018 ( .A(n_2019), .Y(n_2018) );
HB1xp67_ASAP7_75t_L g2029 ( .A(n_2030), .Y(n_2029) );
INVx1_ASAP7_75t_L g2031 ( .A(n_2032), .Y(n_2031) );
endmodule