module fake_netlist_6_1007_n_2357 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_223, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_2357);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_223;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_2357;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_813;
wire n_395;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1950;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_320;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_231;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2348;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_1098;
wire n_391;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_400;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_1147;
wire n_763;
wire n_1848;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_2334;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_973;
wire n_359;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_202),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_14),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_77),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_68),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_138),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_118),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_147),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_155),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_51),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_58),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_193),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_29),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_129),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_46),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_51),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_150),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_198),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_84),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_160),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_15),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_71),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_199),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_66),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_112),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_41),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_2),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_68),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_151),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_38),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_48),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_223),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_132),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_157),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_22),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_12),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_97),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_115),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_152),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_90),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_15),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_67),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_48),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_12),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_26),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_124),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_34),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_71),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_173),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_117),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_25),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_75),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_65),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_166),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g284 ( 
.A(n_209),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_196),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_161),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_125),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_63),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_172),
.Y(n_289)
);

BUFx2_ASAP7_75t_L g290 ( 
.A(n_18),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_81),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_22),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_76),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_76),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_34),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_11),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_18),
.Y(n_297)
);

BUFx5_ASAP7_75t_L g298 ( 
.A(n_136),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_159),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_17),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_119),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_66),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_98),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_218),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_75),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_21),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_2),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_144),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_146),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_87),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_116),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_85),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_94),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_106),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_142),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_73),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_108),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_201),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_16),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_53),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_14),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_133),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_195),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_194),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_130),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_145),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_82),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_73),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_11),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_176),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_189),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_217),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_61),
.Y(n_333)
);

BUFx10_ASAP7_75t_L g334 ( 
.A(n_111),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_38),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_113),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_50),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_36),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_204),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_171),
.Y(n_340)
);

INVx2_ASAP7_75t_SL g341 ( 
.A(n_184),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_92),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_21),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_190),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_37),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_186),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_65),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_121),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_91),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_137),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_17),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_27),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_91),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_175),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_180),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_41),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_102),
.Y(n_357)
);

CKINVDCx12_ASAP7_75t_R g358 ( 
.A(n_78),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_214),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_86),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_182),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_140),
.Y(n_362)
);

BUFx10_ASAP7_75t_L g363 ( 
.A(n_135),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_77),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_163),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_87),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_79),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_148),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_126),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_85),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_220),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_131),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_60),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_170),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_59),
.Y(n_375)
);

BUFx10_ASAP7_75t_L g376 ( 
.A(n_191),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_26),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_165),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_183),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_74),
.Y(n_380)
);

BUFx3_ASAP7_75t_L g381 ( 
.A(n_162),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_86),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_95),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_70),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_79),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_120),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_134),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_25),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_62),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_127),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_4),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_4),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_221),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_141),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_36),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_53),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_89),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_31),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_30),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_30),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_212),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_60),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_107),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_174),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_46),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_19),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_169),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_35),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_16),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_24),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_222),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_197),
.Y(n_412)
);

BUFx2_ASAP7_75t_SL g413 ( 
.A(n_225),
.Y(n_413)
);

INVx2_ASAP7_75t_SL g414 ( 
.A(n_64),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_96),
.Y(n_415)
);

BUFx8_ASAP7_75t_SL g416 ( 
.A(n_188),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_52),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_37),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_82),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_158),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_49),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_59),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_3),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_23),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_7),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_208),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_84),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_5),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_216),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_43),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_61),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_27),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_78),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_88),
.Y(n_434)
);

INVx2_ASAP7_75t_SL g435 ( 
.A(n_90),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_57),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_177),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_207),
.Y(n_438)
);

INVxp67_ASAP7_75t_SL g439 ( 
.A(n_8),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_139),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_6),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_211),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_29),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_49),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_358),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_232),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_261),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_302),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_302),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_275),
.Y(n_450)
);

INVxp67_ASAP7_75t_SL g451 ( 
.A(n_258),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_373),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_284),
.B(n_0),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_226),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_389),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_226),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_227),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_227),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_313),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_373),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_380),
.Y(n_461)
);

BUFx6f_ASAP7_75t_SL g462 ( 
.A(n_334),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_380),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_315),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_396),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_229),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_396),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_229),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_326),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_370),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_336),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_244),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_416),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_370),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_230),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_251),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_237),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_251),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_263),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_238),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_284),
.B(n_0),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_263),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_234),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_234),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_243),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_233),
.Y(n_488)
);

NOR2xp67_ASAP7_75t_L g489 ( 
.A(n_389),
.B(n_1),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_236),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_245),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_249),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_246),
.Y(n_493)
);

INVxp33_ASAP7_75t_L g494 ( 
.A(n_290),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_239),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_239),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_241),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_370),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_252),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_241),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_253),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_262),
.Y(n_502)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_290),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_370),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_266),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_255),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_312),
.B(n_1),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_248),
.Y(n_508)
);

NOR2xp67_ASAP7_75t_L g509 ( 
.A(n_312),
.B(n_3),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_256),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_267),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_341),
.B(n_5),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_248),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_259),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_264),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g516 ( 
.A(n_414),
.B(n_6),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_268),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_279),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_341),
.B(n_7),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_278),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_283),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_285),
.Y(n_522)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_334),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_278),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_270),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_299),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_299),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_370),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_271),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_414),
.B(n_8),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_377),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_358),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_286),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_272),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_274),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_276),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_317),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_254),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_277),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_317),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_390),
.B(n_9),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_287),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_435),
.B(n_9),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_348),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_289),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_377),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_348),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_308),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_280),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_309),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_254),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_282),
.Y(n_552)
);

NOR2xp67_ASAP7_75t_L g553 ( 
.A(n_435),
.B(n_10),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_355),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_355),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_311),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_357),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_390),
.B(n_10),
.Y(n_558)
);

CKINVDCx14_ASAP7_75t_R g559 ( 
.A(n_431),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_357),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_368),
.Y(n_561)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_288),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_368),
.B(n_13),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_559),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_472),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_473),
.Y(n_567)
);

NAND2xp33_ASAP7_75t_SL g568 ( 
.A(n_494),
.B(n_441),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_488),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_472),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_490),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_448),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_472),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_491),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_538),
.B(n_254),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_504),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_470),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_470),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_474),
.Y(n_579)
);

BUFx2_ASAP7_75t_L g580 ( 
.A(n_448),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_474),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_498),
.B(n_301),
.Y(n_582)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_546),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_498),
.A2(n_242),
.B(n_300),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_504),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g586 ( 
.A(n_531),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_528),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_455),
.B(n_303),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_528),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_455),
.Y(n_590)
);

INVx6_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_R g592 ( 
.A(n_475),
.B(n_314),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_472),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_478),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_493),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_512),
.B(n_370),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_478),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_501),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_502),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_558),
.B(n_318),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_483),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_505),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_483),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_454),
.Y(n_604)
);

INVx6_ASAP7_75t_L g605 ( 
.A(n_551),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_476),
.A2(n_265),
.B1(n_294),
.B2(n_228),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_456),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_457),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_458),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_511),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_445),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_466),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_468),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_485),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_551),
.B(n_303),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_486),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_446),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_449),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_449),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_452),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_503),
.A2(n_441),
.B1(n_384),
.B2(n_392),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_479),
.Y(n_623)
);

INVxp67_ASAP7_75t_SL g624 ( 
.A(n_496),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_497),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_500),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_508),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_SL g628 ( 
.A(n_453),
.B(n_247),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_513),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_520),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_524),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_452),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_526),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_527),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_517),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_537),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_540),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_544),
.B(n_303),
.Y(n_638)
);

OA21x2_ASAP7_75t_L g639 ( 
.A1(n_547),
.A2(n_242),
.B(n_300),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_554),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_482),
.B(n_334),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_555),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_518),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_557),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_521),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_560),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_522),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_460),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_561),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_489),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_451),
.B(n_564),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_519),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_541),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_507),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_533),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_542),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_545),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_509),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_601),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_601),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_588),
.B(n_381),
.Y(n_661)
);

INVxp67_ASAP7_75t_SL g662 ( 
.A(n_570),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_652),
.A2(n_242),
.B1(n_424),
.B2(n_250),
.Y(n_663)
);

INVx8_ASAP7_75t_L g664 ( 
.A(n_651),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_601),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_628),
.B(n_475),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_565),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_628),
.B(n_477),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_607),
.Y(n_669)
);

AO22x2_ASAP7_75t_L g670 ( 
.A1(n_621),
.A2(n_562),
.B1(n_250),
.B2(n_257),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_605),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_652),
.B(n_477),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_605),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_653),
.B(n_481),
.Y(n_674)
);

NAND3x1_ASAP7_75t_L g675 ( 
.A(n_651),
.B(n_257),
.C(n_231),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_586),
.B(n_523),
.Y(n_676)
);

INVx2_ASAP7_75t_SL g677 ( 
.A(n_605),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_576),
.Y(n_678)
);

BUFx4f_ASAP7_75t_L g679 ( 
.A(n_639),
.Y(n_679)
);

BUFx10_ASAP7_75t_L g680 ( 
.A(n_565),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_600),
.B(n_481),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_617),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_601),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_576),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_607),
.Y(n_685)
);

NOR2xp33_ASAP7_75t_L g686 ( 
.A(n_600),
.B(n_487),
.Y(n_686)
);

INVx5_ASAP7_75t_L g687 ( 
.A(n_629),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_608),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_588),
.B(n_381),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_653),
.B(n_301),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_601),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_605),
.B(n_487),
.Y(n_692)
);

AND3x2_ASAP7_75t_L g693 ( 
.A(n_580),
.B(n_439),
.C(n_424),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_576),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_586),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_588),
.B(n_381),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_605),
.Y(n_697)
);

INVx4_ASAP7_75t_L g698 ( 
.A(n_629),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_654),
.B(n_492),
.Y(n_699)
);

AND2x6_ASAP7_75t_L g700 ( 
.A(n_575),
.B(n_378),
.Y(n_700)
);

INVx4_ASAP7_75t_SL g701 ( 
.A(n_591),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_605),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_585),
.Y(n_703)
);

OR2x6_ASAP7_75t_L g704 ( 
.A(n_580),
.B(n_532),
.Y(n_704)
);

INVxp67_ASAP7_75t_SL g705 ( 
.A(n_570),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_575),
.B(n_378),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_641),
.B(n_492),
.Y(n_707)
);

AND2x6_ASAP7_75t_L g708 ( 
.A(n_575),
.B(n_383),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_641),
.B(n_244),
.Y(n_709)
);

CKINVDCx14_ASAP7_75t_R g710 ( 
.A(n_580),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_651),
.B(n_244),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_608),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_572),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_583),
.B(n_460),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_583),
.B(n_461),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_611),
.B(n_499),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_609),
.Y(n_717)
);

AND2x2_ASAP7_75t_SL g718 ( 
.A(n_639),
.B(n_596),
.Y(n_718)
);

INVx6_ASAP7_75t_L g719 ( 
.A(n_615),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_609),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_612),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_614),
.Y(n_722)
);

AND2x6_ASAP7_75t_L g723 ( 
.A(n_615),
.B(n_383),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_612),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_613),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_613),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_625),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_596),
.B(n_650),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_568),
.A2(n_550),
.B1(n_556),
.B2(n_548),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_625),
.Y(n_730)
);

INVx4_ASAP7_75t_L g731 ( 
.A(n_629),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_601),
.Y(n_732)
);

AND2x2_ASAP7_75t_SL g733 ( 
.A(n_639),
.B(n_393),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_572),
.Y(n_734)
);

NAND3xp33_ASAP7_75t_L g735 ( 
.A(n_650),
.B(n_506),
.C(n_499),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_627),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_654),
.B(n_244),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_627),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_630),
.Y(n_739)
);

BUFx10_ASAP7_75t_L g740 ( 
.A(n_567),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_569),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_630),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_601),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_658),
.B(n_506),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_640),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_571),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_615),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_624),
.B(n_644),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_629),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_574),
.Y(n_750)
);

OAI22xp33_ASAP7_75t_L g751 ( 
.A1(n_658),
.A2(n_269),
.B1(n_417),
.B2(n_260),
.Y(n_751)
);

OR2x2_ASAP7_75t_SL g752 ( 
.A(n_619),
.B(n_231),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_614),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_624),
.B(n_644),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_585),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_585),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_611),
.B(n_510),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_588),
.B(n_393),
.Y(n_758)
);

INVx3_ASAP7_75t_L g759 ( 
.A(n_601),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_640),
.Y(n_760)
);

OR2x2_ASAP7_75t_L g761 ( 
.A(n_618),
.B(n_461),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_638),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_623),
.Y(n_763)
);

AND2x6_ASAP7_75t_L g764 ( 
.A(n_638),
.B(n_404),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_646),
.Y(n_765)
);

INVx4_ASAP7_75t_SL g766 ( 
.A(n_591),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_646),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_614),
.B(n_510),
.Y(n_768)
);

AND2x6_ASAP7_75t_L g769 ( 
.A(n_638),
.B(n_404),
.Y(n_769)
);

AND2x2_ASAP7_75t_SL g770 ( 
.A(n_639),
.B(n_407),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_590),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_590),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_649),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_614),
.B(n_514),
.Y(n_774)
);

INVx1_ASAP7_75t_SL g775 ( 
.A(n_623),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_622),
.B(n_514),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_618),
.B(n_515),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_622),
.Y(n_778)
);

INVx4_ASAP7_75t_L g779 ( 
.A(n_629),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_622),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_590),
.Y(n_781)
);

BUFx3_ASAP7_75t_L g782 ( 
.A(n_639),
.Y(n_782)
);

NAND3xp33_ASAP7_75t_L g783 ( 
.A(n_568),
.B(n_525),
.C(n_515),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_588),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_590),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_617),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_622),
.B(n_525),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_622),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_639),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_637),
.B(n_529),
.Y(n_790)
);

INVx4_ASAP7_75t_SL g791 ( 
.A(n_591),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_637),
.Y(n_792)
);

INVx4_ASAP7_75t_L g793 ( 
.A(n_629),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_595),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_637),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_618),
.B(n_529),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_616),
.B(n_407),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_577),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_637),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_620),
.B(n_534),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_584),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_616),
.B(n_411),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_619),
.Y(n_803)
);

OR2x6_ASAP7_75t_L g804 ( 
.A(n_620),
.B(n_413),
.Y(n_804)
);

OR2x6_ASAP7_75t_L g805 ( 
.A(n_620),
.B(n_413),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_637),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_577),
.Y(n_807)
);

AND2x6_ASAP7_75t_L g808 ( 
.A(n_594),
.B(n_411),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_578),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_578),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_584),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_579),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_632),
.B(n_463),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_632),
.Y(n_814)
);

BUFx10_ASAP7_75t_L g815 ( 
.A(n_657),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_632),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_672),
.B(n_534),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_681),
.B(n_629),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_679),
.B(n_592),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_681),
.B(n_629),
.Y(n_820)
);

INVx8_ASAP7_75t_L g821 ( 
.A(n_664),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_686),
.B(n_642),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_798),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_798),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_784),
.Y(n_825)
);

AOI22xp5_ASAP7_75t_L g826 ( 
.A1(n_686),
.A2(n_484),
.B1(n_480),
.B2(n_648),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_719),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_776),
.B(n_642),
.Y(n_828)
);

INVxp67_ASAP7_75t_L g829 ( 
.A(n_695),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_679),
.B(n_592),
.Y(n_830)
);

BUFx4f_ASAP7_75t_L g831 ( 
.A(n_804),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_776),
.B(n_642),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_676),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_733),
.A2(n_584),
.B1(n_281),
.B2(n_295),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_787),
.B(n_642),
.Y(n_835)
);

OAI22xp5_ASAP7_75t_L g836 ( 
.A1(n_762),
.A2(n_450),
.B1(n_459),
.B2(n_447),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_733),
.A2(n_584),
.B1(n_281),
.B2(n_295),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_807),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_770),
.B(n_244),
.Y(n_839)
);

INVxp67_ASAP7_75t_SL g840 ( 
.A(n_789),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_784),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_787),
.B(n_642),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_790),
.B(n_642),
.Y(n_843)
);

INVxp67_ASAP7_75t_L g844 ( 
.A(n_716),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_762),
.B(n_648),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_669),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_747),
.A2(n_469),
.B1(n_471),
.B2(n_464),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_685),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_678),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_777),
.B(n_648),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_790),
.B(n_642),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_747),
.B(n_642),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_716),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_807),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_728),
.B(n_604),
.Y(n_855)
);

NOR2x1p5_ASAP7_75t_L g856 ( 
.A(n_674),
.B(n_463),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_688),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_712),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_717),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_678),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_781),
.B(n_719),
.Y(n_861)
);

AOI22xp5_ASAP7_75t_L g862 ( 
.A1(n_707),
.A2(n_664),
.B1(n_668),
.B2(n_666),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_781),
.B(n_604),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_720),
.Y(n_864)
);

BUFx8_ASAP7_75t_L g865 ( 
.A(n_796),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_748),
.B(n_535),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_719),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_721),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_693),
.Y(n_869)
);

AOI22xp33_ASAP7_75t_L g870 ( 
.A1(n_770),
.A2(n_584),
.B1(n_297),
.B2(n_310),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_724),
.Y(n_871)
);

OR2x6_ASAP7_75t_L g872 ( 
.A(n_704),
.B(n_606),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_725),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_781),
.B(n_604),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_809),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_664),
.B(n_700),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_726),
.Y(n_877)
);

A2O1A1Ixp33_ASAP7_75t_L g878 ( 
.A1(n_707),
.A2(n_530),
.B(n_543),
.C(n_516),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_684),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_727),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_664),
.B(n_604),
.Y(n_881)
);

AND2x4_ASAP7_75t_L g882 ( 
.A(n_722),
.B(n_616),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_730),
.Y(n_883)
);

OAI22xp33_ASAP7_75t_L g884 ( 
.A1(n_754),
.A2(n_621),
.B1(n_553),
.B2(n_240),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_699),
.B(n_535),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_700),
.B(n_626),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_700),
.B(n_626),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_736),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_789),
.B(n_244),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_700),
.B(n_626),
.Y(n_890)
);

AND2x2_ASAP7_75t_SL g891 ( 
.A(n_666),
.B(n_438),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_789),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_738),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_700),
.B(n_626),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_809),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_744),
.B(n_536),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_SL g897 ( 
.A1(n_668),
.A2(n_606),
.B1(n_462),
.B2(n_467),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_722),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_663),
.A2(n_297),
.B(n_310),
.C(n_273),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_706),
.B(n_631),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_714),
.B(n_465),
.Y(n_901)
);

NAND2x1p5_ASAP7_75t_L g902 ( 
.A(n_782),
.B(n_584),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_706),
.B(n_631),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_706),
.B(n_631),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_SL g905 ( 
.A(n_741),
.B(n_598),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_718),
.A2(n_316),
.B1(n_327),
.B2(n_273),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_768),
.B(n_536),
.Y(n_907)
);

AND2x6_ASAP7_75t_SL g908 ( 
.A(n_704),
.B(n_316),
.Y(n_908)
);

OAI21xp33_ASAP7_75t_L g909 ( 
.A1(n_663),
.A2(n_549),
.B(n_539),
.Y(n_909)
);

NAND3xp33_ASAP7_75t_L g910 ( 
.A(n_735),
.B(n_549),
.C(n_539),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_739),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_718),
.A2(n_333),
.B1(n_345),
.B2(n_327),
.Y(n_912)
);

NOR2xp67_ASAP7_75t_L g913 ( 
.A(n_783),
.B(n_599),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_757),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_742),
.Y(n_915)
);

INVx4_ASAP7_75t_L g916 ( 
.A(n_753),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_745),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_708),
.B(n_633),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_684),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_741),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_708),
.A2(n_467),
.B1(n_465),
.B2(n_552),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_760),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_708),
.B(n_633),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_774),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_765),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_711),
.B(n_552),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_767),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_L g928 ( 
.A(n_800),
.B(n_563),
.C(n_602),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_711),
.B(n_563),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_708),
.B(n_633),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_708),
.B(n_634),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_789),
.B(n_634),
.Y(n_932)
);

NOR2x1_ASAP7_75t_L g933 ( 
.A(n_692),
.B(n_715),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_SL g934 ( 
.A1(n_670),
.A2(n_462),
.B1(n_635),
.B2(n_610),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_752),
.B(n_462),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_811),
.B(n_634),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_782),
.A2(n_382),
.B1(n_430),
.B2(n_432),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_773),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_761),
.B(n_656),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_812),
.B(n_235),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_694),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_694),
.Y(n_942)
);

AND2x6_ASAP7_75t_L g943 ( 
.A(n_801),
.B(n_420),
.Y(n_943)
);

OR2x2_ASAP7_75t_L g944 ( 
.A(n_813),
.B(n_814),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_811),
.B(n_438),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_811),
.B(n_753),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_810),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_734),
.B(n_816),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_661),
.B(n_636),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_764),
.A2(n_371),
.B1(n_304),
.B2(n_372),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_810),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_811),
.B(n_438),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_661),
.Y(n_953)
);

BUFx8_ASAP7_75t_L g954 ( 
.A(n_682),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_801),
.B(n_438),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_771),
.B(n_772),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_764),
.A2(n_769),
.B1(n_723),
.B2(n_689),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_778),
.B(n_438),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_804),
.A2(n_420),
.B1(n_429),
.B2(n_426),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_661),
.Y(n_960)
);

BUFx6f_ASAP7_75t_SL g961 ( 
.A(n_815),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_689),
.B(n_636),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_804),
.B(n_805),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_710),
.B(n_763),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_771),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_709),
.B(n_292),
.C(n_291),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_689),
.Y(n_967)
);

NOR2x1p5_ASAP7_75t_L g968 ( 
.A(n_746),
.B(n_643),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_696),
.Y(n_969)
);

INVx1_ASAP7_75t_SL g970 ( 
.A(n_775),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_780),
.B(n_438),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_696),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_696),
.Y(n_973)
);

AND2x6_ASAP7_75t_SL g974 ( 
.A(n_704),
.B(n_333),
.Y(n_974)
);

AOI22xp33_ASAP7_75t_L g975 ( 
.A1(n_764),
.A2(n_367),
.B1(n_430),
.B2(n_432),
.Y(n_975)
);

BUFx5_ASAP7_75t_L g976 ( 
.A(n_788),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_703),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_797),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_772),
.B(n_634),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_SL g980 ( 
.A1(n_670),
.A2(n_710),
.B1(n_805),
.B2(n_804),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_713),
.B(n_645),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_785),
.B(n_758),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_785),
.B(n_579),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_703),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_755),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_702),
.Y(n_986)
);

INVx1_ASAP7_75t_SL g987 ( 
.A(n_682),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_949),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_827),
.B(n_758),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_965),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_970),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_882),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_892),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_829),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_866),
.B(n_764),
.Y(n_995)
);

INVx4_ASAP7_75t_L g996 ( 
.A(n_892),
.Y(n_996)
);

HB1xp67_ASAP7_75t_L g997 ( 
.A(n_924),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_844),
.B(n_803),
.Y(n_998)
);

AND2x2_ASAP7_75t_L g999 ( 
.A(n_850),
.B(n_805),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_892),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_965),
.Y(n_1001)
);

AND2x4_ASAP7_75t_L g1002 ( 
.A(n_827),
.B(n_758),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_949),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_892),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_866),
.B(n_764),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_853),
.B(n_805),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_967),
.Y(n_1007)
);

INVx3_ASAP7_75t_L g1008 ( 
.A(n_967),
.Y(n_1008)
);

NAND3xp33_ASAP7_75t_L g1009 ( 
.A(n_926),
.B(n_729),
.C(n_655),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_914),
.B(n_833),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_920),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_962),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_867),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_823),
.Y(n_1014)
);

OAI21xp33_ASAP7_75t_L g1015 ( 
.A1(n_885),
.A2(n_670),
.B(n_690),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_891),
.B(n_769),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_821),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_817),
.B(n_647),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_962),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_891),
.A2(n_769),
.B1(n_709),
.B2(n_723),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_964),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_862),
.B(n_769),
.Y(n_1022)
);

INVx2_ASAP7_75t_SL g1023 ( 
.A(n_882),
.Y(n_1023)
);

OR2x6_ASAP7_75t_SL g1024 ( 
.A(n_836),
.B(n_746),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_840),
.B(n_769),
.Y(n_1025)
);

NOR2x1_ASAP7_75t_L g1026 ( 
.A(n_910),
.B(n_751),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_978),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_867),
.B(n_898),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_821),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_986),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_906),
.A2(n_675),
.B1(n_705),
.B2(n_662),
.Y(n_1031)
);

AND2x4_ASAP7_75t_L g1032 ( 
.A(n_898),
.B(n_702),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_823),
.Y(n_1033)
);

OR2x4_ASAP7_75t_L g1034 ( 
.A(n_885),
.B(n_345),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_817),
.B(n_750),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_824),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_916),
.B(n_797),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_834),
.B(n_792),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_821),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_845),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_SL g1041 ( 
.A(n_905),
.B(n_750),
.Y(n_1041)
);

INVx6_ASAP7_75t_L g1042 ( 
.A(n_865),
.Y(n_1042)
);

INVx5_ASAP7_75t_L g1043 ( 
.A(n_943),
.Y(n_1043)
);

BUFx3_ASAP7_75t_L g1044 ( 
.A(n_954),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_906),
.A2(n_723),
.B1(n_808),
.B2(n_802),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_824),
.Y(n_1046)
);

A2O1A1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_912),
.A2(n_690),
.B(n_802),
.C(n_797),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_SL g1048 ( 
.A(n_954),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_986),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_838),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_926),
.B(n_723),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_SL g1052 ( 
.A(n_826),
.B(n_897),
.C(n_921),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_986),
.Y(n_1053)
);

OR2x6_ASAP7_75t_L g1054 ( 
.A(n_924),
.B(n_675),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_838),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_929),
.B(n_723),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_929),
.B(n_795),
.Y(n_1057)
);

BUFx3_ASAP7_75t_L g1058 ( 
.A(n_865),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_854),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_907),
.B(n_799),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_944),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_834),
.B(n_806),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_854),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_SL g1064 ( 
.A(n_884),
.B(n_296),
.C(n_293),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_875),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_884),
.B(n_306),
.C(n_305),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_875),
.Y(n_1067)
);

INVx1_ASAP7_75t_SL g1068 ( 
.A(n_981),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_831),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_R g1070 ( 
.A(n_961),
.B(n_794),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_986),
.Y(n_1071)
);

OR2x2_ASAP7_75t_L g1072 ( 
.A(n_987),
.B(n_794),
.Y(n_1072)
);

INVx3_ASAP7_75t_L g1073 ( 
.A(n_895),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_895),
.Y(n_1074)
);

INVx1_ASAP7_75t_SL g1075 ( 
.A(n_901),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_869),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_896),
.B(n_815),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_943),
.Y(n_1078)
);

AND2x4_ASAP7_75t_L g1079 ( 
.A(n_916),
.B(n_802),
.Y(n_1079)
);

AND2x4_ASAP7_75t_L g1080 ( 
.A(n_953),
.B(n_671),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_839),
.A2(n_673),
.B(n_671),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_960),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_969),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_R g1084 ( 
.A(n_961),
.B(n_786),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_948),
.B(n_667),
.Y(n_1085)
);

INVx5_ASAP7_75t_L g1086 ( 
.A(n_943),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_972),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_907),
.B(n_673),
.Y(n_1088)
);

CKINVDCx11_ASAP7_75t_R g1089 ( 
.A(n_908),
.Y(n_1089)
);

AND2x2_ASAP7_75t_L g1090 ( 
.A(n_896),
.B(n_815),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_837),
.B(n_659),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_973),
.Y(n_1092)
);

HB1xp67_ASAP7_75t_L g1093 ( 
.A(n_847),
.Y(n_1093)
);

AND2x2_ASAP7_75t_SL g1094 ( 
.A(n_912),
.B(n_831),
.Y(n_1094)
);

A2O1A1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_937),
.A2(n_347),
.B(n_352),
.C(n_351),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_946),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_947),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_984),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_933),
.A2(n_808),
.B1(n_697),
.B2(n_677),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_837),
.B(n_677),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_870),
.B(n_940),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_951),
.Y(n_1102)
);

BUFx3_ASAP7_75t_L g1103 ( 
.A(n_846),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_968),
.Y(n_1104)
);

NOR2x1_ASAP7_75t_L g1105 ( 
.A(n_913),
.B(n_737),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_SL g1106 ( 
.A(n_909),
.B(n_319),
.C(n_307),
.Y(n_1106)
);

INVxp67_ASAP7_75t_SL g1107 ( 
.A(n_902),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_936),
.A2(n_697),
.B(n_698),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_870),
.B(n_808),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_940),
.B(n_808),
.Y(n_1110)
);

AND2x2_ASAP7_75t_SL g1111 ( 
.A(n_975),
.B(n_429),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_948),
.B(n_667),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_984),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_943),
.A2(n_808),
.B1(n_737),
.B2(n_683),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_848),
.B(n_667),
.Y(n_1115)
);

INVx4_ASAP7_75t_L g1116 ( 
.A(n_943),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_839),
.A2(n_660),
.B(n_659),
.Y(n_1117)
);

NOR2xp67_ASAP7_75t_L g1118 ( 
.A(n_939),
.B(n_636),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_818),
.B(n_820),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_825),
.Y(n_1120)
);

OR2x2_ASAP7_75t_L g1121 ( 
.A(n_928),
.B(n_786),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_822),
.B(n_659),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_855),
.B(n_857),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_974),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_858),
.B(n_660),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_849),
.Y(n_1126)
);

BUFx10_ASAP7_75t_L g1127 ( 
.A(n_963),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_841),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_902),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_859),
.B(n_701),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_976),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_864),
.B(n_701),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_872),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_868),
.B(n_871),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_861),
.Y(n_1135)
);

INVx4_ASAP7_75t_L g1136 ( 
.A(n_976),
.Y(n_1136)
);

HB1xp67_ASAP7_75t_L g1137 ( 
.A(n_873),
.Y(n_1137)
);

INVxp67_ASAP7_75t_SL g1138 ( 
.A(n_932),
.Y(n_1138)
);

AND2x4_ASAP7_75t_L g1139 ( 
.A(n_877),
.B(n_701),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_872),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_880),
.Y(n_1141)
);

BUFx2_ASAP7_75t_L g1142 ( 
.A(n_872),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_883),
.B(n_660),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_860),
.Y(n_1144)
);

HB1xp67_ASAP7_75t_L g1145 ( 
.A(n_888),
.Y(n_1145)
);

INVx5_ASAP7_75t_L g1146 ( 
.A(n_879),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_893),
.Y(n_1147)
);

INVx5_ASAP7_75t_L g1148 ( 
.A(n_919),
.Y(n_1148)
);

CKINVDCx20_ASAP7_75t_R g1149 ( 
.A(n_959),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_980),
.Y(n_1150)
);

XNOR2xp5_ASAP7_75t_L g1151 ( 
.A(n_856),
.B(n_740),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_941),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_911),
.B(n_766),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_915),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_942),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_917),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_922),
.B(n_665),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_925),
.B(n_665),
.Y(n_1158)
);

INVx3_ASAP7_75t_L g1159 ( 
.A(n_977),
.Y(n_1159)
);

HB1xp67_ASAP7_75t_L g1160 ( 
.A(n_927),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_876),
.Y(n_1161)
);

BUFx2_ASAP7_75t_L g1162 ( 
.A(n_963),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_935),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_937),
.A2(n_352),
.B(n_351),
.C(n_436),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_985),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_982),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_938),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_983),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_863),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_956),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_886),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_878),
.B(n_680),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_R g1173 ( 
.A(n_935),
.B(n_740),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_976),
.Y(n_1174)
);

INVx3_ASAP7_75t_SL g1175 ( 
.A(n_819),
.Y(n_1175)
);

BUFx8_ASAP7_75t_SL g1176 ( 
.A(n_934),
.Y(n_1176)
);

AO22x1_ASAP7_75t_L g1177 ( 
.A1(n_881),
.A2(n_408),
.B1(n_321),
.B2(n_398),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_966),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_852),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_976),
.Y(n_1180)
);

AOI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1057),
.A2(n_832),
.B(n_828),
.Y(n_1181)
);

OAI21x1_ASAP7_75t_L g1182 ( 
.A1(n_1108),
.A2(n_842),
.B(n_835),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1100),
.A2(n_955),
.B(n_952),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1141),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1122),
.A2(n_851),
.B(n_843),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_994),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1109),
.A2(n_955),
.B(n_952),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1147),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1117),
.A2(n_889),
.B(n_945),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_1017),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_SL g1191 ( 
.A1(n_1078),
.A2(n_957),
.B(n_890),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_990),
.Y(n_1192)
);

CKINVDCx8_ASAP7_75t_R g1193 ( 
.A(n_1104),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_990),
.Y(n_1194)
);

OA21x2_ASAP7_75t_L g1195 ( 
.A1(n_1119),
.A2(n_889),
.B(n_945),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1131),
.Y(n_1196)
);

OAI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1091),
.A2(n_830),
.B(n_819),
.Y(n_1197)
);

AOI221xp5_ASAP7_75t_L g1198 ( 
.A1(n_1035),
.A2(n_878),
.B1(n_975),
.B2(n_428),
.C(n_353),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1091),
.A2(n_830),
.B(n_887),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1156),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_991),
.Y(n_1201)
);

AOI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1022),
.A2(n_1056),
.B(n_1051),
.Y(n_1202)
);

BUFx6f_ASAP7_75t_L g1203 ( 
.A(n_1017),
.Y(n_1203)
);

AO21x1_ASAP7_75t_L g1204 ( 
.A1(n_1101),
.A2(n_900),
.B(n_894),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_L g1205 ( 
.A(n_1035),
.B(n_740),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1167),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_999),
.B(n_899),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1081),
.A2(n_1180),
.B(n_1174),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1027),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1180),
.A2(n_874),
.B(n_903),
.Y(n_1210)
);

INVx3_ASAP7_75t_L g1211 ( 
.A(n_1131),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1047),
.A2(n_918),
.A3(n_923),
.B(n_904),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1036),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_SL g1214 ( 
.A1(n_1131),
.A2(n_931),
.B(n_930),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1011),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1123),
.B(n_950),
.Y(n_1216)
);

BUFx3_ASAP7_75t_L g1217 ( 
.A(n_1011),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_L g1218 ( 
.A1(n_995),
.A2(n_979),
.B(n_971),
.Y(n_1218)
);

INVx3_ASAP7_75t_L g1219 ( 
.A(n_1136),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1038),
.A2(n_971),
.B(n_958),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1180),
.A2(n_958),
.B(n_683),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1168),
.B(n_899),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_SL g1223 ( 
.A1(n_1078),
.A2(n_367),
.B(n_347),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1174),
.A2(n_683),
.B(n_665),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_SL g1225 ( 
.A1(n_1136),
.A2(n_731),
.B(n_698),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1025),
.A2(n_732),
.B(n_691),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1018),
.B(n_680),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1136),
.A2(n_731),
.B(n_698),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1017),
.B(n_691),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1129),
.A2(n_732),
.B(n_691),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1047),
.A2(n_406),
.A3(n_397),
.B(n_436),
.Y(n_1231)
);

BUFx2_ASAP7_75t_SL g1232 ( 
.A(n_1017),
.Y(n_1232)
);

AOI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1005),
.A2(n_756),
.B(n_755),
.Y(n_1233)
);

OAI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1062),
.A2(n_743),
.B(n_732),
.Y(n_1234)
);

BUFx12f_ASAP7_75t_SL g1235 ( 
.A(n_1054),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1031),
.A2(n_1095),
.A3(n_1164),
.B(n_1172),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1129),
.A2(n_759),
.B(n_743),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1129),
.A2(n_759),
.B(n_743),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1062),
.A2(n_1016),
.B(n_1138),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1001),
.A2(n_759),
.B(n_756),
.Y(n_1240)
);

OAI21x1_ASAP7_75t_L g1241 ( 
.A1(n_1001),
.A2(n_976),
.B(n_587),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_996),
.A2(n_749),
.B(n_731),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_996),
.A2(n_779),
.B(n_749),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1073),
.A2(n_1033),
.B(n_1014),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1073),
.A2(n_1033),
.B(n_1014),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1179),
.B(n_976),
.Y(n_1246)
);

OAI21x1_ASAP7_75t_L g1247 ( 
.A1(n_1073),
.A2(n_587),
.B(n_581),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1050),
.A2(n_589),
.B(n_581),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1172),
.A2(n_793),
.A3(n_779),
.B(n_749),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1098),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_SL g1251 ( 
.A1(n_1110),
.A2(n_344),
.B(n_334),
.Y(n_1251)
);

OAI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1060),
.A2(n_793),
.B(n_779),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1018),
.B(n_359),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_996),
.A2(n_793),
.B(n_687),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1050),
.A2(n_589),
.B(n_594),
.Y(n_1255)
);

BUFx12f_ASAP7_75t_L g1256 ( 
.A(n_1042),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1061),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1170),
.B(n_603),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1085),
.B(n_680),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1020),
.A2(n_582),
.B(n_573),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_997),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1059),
.A2(n_603),
.B(n_597),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1042),
.Y(n_1263)
);

AOI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1009),
.A2(n_1068),
.B(n_1085),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1169),
.A2(n_582),
.B(n_573),
.Y(n_1265)
);

OAI21xp33_ASAP7_75t_L g1266 ( 
.A1(n_1041),
.A2(n_328),
.B(n_320),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1170),
.A2(n_573),
.B(n_566),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1040),
.B(n_597),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_1059),
.A2(n_597),
.B(n_573),
.Y(n_1269)
);

INVx4_ASAP7_75t_L g1270 ( 
.A(n_1029),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1094),
.B(n_322),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1094),
.B(n_323),
.Y(n_1272)
);

OAI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1114),
.A2(n_593),
.B(n_566),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1065),
.A2(n_597),
.B(n_593),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1045),
.A2(n_593),
.B(n_566),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1021),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1098),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_1070),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1065),
.A2(n_593),
.B(n_566),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1134),
.B(n_324),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1134),
.B(n_325),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1134),
.B(n_330),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1067),
.A2(n_570),
.B(n_397),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1077),
.B(n_240),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1046),
.Y(n_1285)
);

OAI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1107),
.A2(n_570),
.B(n_687),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1067),
.A2(n_570),
.B(n_406),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1088),
.A2(n_382),
.B(n_687),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1074),
.A2(n_791),
.B(n_766),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1053),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1074),
.A2(n_791),
.B(n_766),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1090),
.B(n_240),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1120),
.B(n_331),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1128),
.B(n_332),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1125),
.A2(n_791),
.B(n_687),
.Y(n_1295)
);

NOR4xp25_ASAP7_75t_L g1296 ( 
.A(n_1052),
.B(n_422),
.C(n_349),
.D(n_412),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_993),
.A2(n_374),
.B(n_442),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1111),
.B(n_339),
.Y(n_1298)
);

BUFx3_ASAP7_75t_L g1299 ( 
.A(n_1013),
.Y(n_1299)
);

BUFx2_ASAP7_75t_L g1300 ( 
.A(n_1162),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1075),
.B(n_349),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1006),
.A2(n_387),
.B1(n_340),
.B2(n_342),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1111),
.B(n_346),
.Y(n_1303)
);

AO21x2_ASAP7_75t_L g1304 ( 
.A1(n_1099),
.A2(n_298),
.B(n_344),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_993),
.A2(n_386),
.B(n_440),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1143),
.A2(n_1158),
.B(n_1157),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1113),
.A2(n_298),
.B(n_185),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1171),
.B(n_298),
.Y(n_1308)
);

INVx2_ASAP7_75t_L g1309 ( 
.A(n_1113),
.Y(n_1309)
);

NOR4xp25_ASAP7_75t_L g1310 ( 
.A(n_1015),
.B(n_422),
.C(n_349),
.D(n_376),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_993),
.A2(n_1004),
.B(n_1000),
.Y(n_1311)
);

A2O1A1Ixp33_ASAP7_75t_L g1312 ( 
.A1(n_1095),
.A2(n_422),
.B(n_366),
.C(n_364),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1007),
.A2(n_298),
.B(n_178),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1053),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1055),
.A2(n_1063),
.B(n_1006),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1137),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_993),
.A2(n_379),
.B(n_437),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1171),
.B(n_298),
.Y(n_1318)
);

BUFx2_ASAP7_75t_L g1319 ( 
.A(n_1054),
.Y(n_1319)
);

AOI221xp5_ASAP7_75t_L g1320 ( 
.A1(n_1149),
.A2(n_1093),
.B1(n_998),
.B2(n_1150),
.C(n_1010),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1164),
.A2(n_433),
.B(n_444),
.C(n_443),
.Y(n_1321)
);

AO31x2_ASAP7_75t_L g1322 ( 
.A1(n_1078),
.A2(n_298),
.A3(n_19),
.B(n_20),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1154),
.B(n_350),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1126),
.A2(n_354),
.B(n_361),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1010),
.B(n_362),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1000),
.A2(n_415),
.B(n_403),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1112),
.B(n_365),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1029),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1171),
.B(n_298),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1007),
.A2(n_298),
.B(n_149),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1000),
.A2(n_401),
.B(n_394),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_SL g1332 ( 
.A1(n_1116),
.A2(n_143),
.B(n_93),
.Y(n_1332)
);

AO21x1_ASAP7_75t_L g1333 ( 
.A1(n_1116),
.A2(n_298),
.B(n_344),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1126),
.A2(n_369),
.B(n_434),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1007),
.A2(n_123),
.B(n_224),
.Y(n_1335)
);

AO31x2_ASAP7_75t_L g1336 ( 
.A1(n_1116),
.A2(n_1102),
.A3(n_1097),
.B(n_1155),
.Y(n_1336)
);

INVx2_ASAP7_75t_SL g1337 ( 
.A(n_1053),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_1084),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1145),
.Y(n_1339)
);

OAI21xp5_ASAP7_75t_L g1340 ( 
.A1(n_1144),
.A2(n_395),
.B(n_427),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1029),
.B(n_591),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1160),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1008),
.A2(n_114),
.B(n_219),
.Y(n_1343)
);

A2O1A1Ixp33_ASAP7_75t_L g1344 ( 
.A1(n_1064),
.A2(n_338),
.B(n_337),
.C(n_335),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1144),
.A2(n_13),
.A3(n_20),
.B(n_23),
.Y(n_1345)
);

AND2x4_ASAP7_75t_L g1346 ( 
.A(n_989),
.B(n_99),
.Y(n_1346)
);

AOI22x1_ASAP7_75t_L g1347 ( 
.A1(n_1197),
.A2(n_1175),
.B1(n_1178),
.B2(n_1008),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1241),
.A2(n_1105),
.B(n_1008),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1192),
.Y(n_1349)
);

OAI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1216),
.A2(n_1026),
.B(n_1106),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1253),
.B(n_1112),
.Y(n_1351)
);

OAI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1199),
.A2(n_1083),
.B(n_1082),
.Y(n_1352)
);

OAI221xp5_ASAP7_75t_L g1353 ( 
.A1(n_1198),
.A2(n_1163),
.B1(n_1066),
.B2(n_1121),
.C(n_998),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1241),
.A2(n_1159),
.B(n_1155),
.Y(n_1354)
);

BUFx6f_ASAP7_75t_L g1355 ( 
.A(n_1190),
.Y(n_1355)
);

CKINVDCx8_ASAP7_75t_R g1356 ( 
.A(n_1278),
.Y(n_1356)
);

INVxp67_ASAP7_75t_SL g1357 ( 
.A(n_1186),
.Y(n_1357)
);

O2A1O1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1264),
.A2(n_1054),
.B(n_1115),
.C(n_1072),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1201),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1320),
.A2(n_1149),
.B1(n_1150),
.B2(n_1054),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1298),
.A2(n_1103),
.B1(n_1176),
.B2(n_1002),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_1346),
.B(n_1013),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1303),
.A2(n_1103),
.B1(n_1176),
.B2(n_1002),
.Y(n_1363)
);

AO21x2_ASAP7_75t_L g1364 ( 
.A1(n_1202),
.A2(n_1118),
.B(n_1092),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1283),
.A2(n_1159),
.B(n_1152),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1227),
.B(n_1096),
.Y(n_1366)
);

BUFx2_ASAP7_75t_SL g1367 ( 
.A(n_1215),
.Y(n_1367)
);

O2A1O1Ixp33_ASAP7_75t_L g1368 ( 
.A1(n_1205),
.A2(n_1115),
.B(n_1175),
.C(n_1076),
.Y(n_1368)
);

AO31x2_ASAP7_75t_L g1369 ( 
.A1(n_1204),
.A2(n_1165),
.A3(n_1152),
.B(n_1087),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1190),
.Y(n_1370)
);

AO21x2_ASAP7_75t_L g1371 ( 
.A1(n_1181),
.A2(n_1003),
.B(n_988),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1183),
.A2(n_1083),
.B(n_1023),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1338),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1283),
.A2(n_1159),
.B(n_1165),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1192),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1215),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1300),
.Y(n_1377)
);

OAI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1259),
.A2(n_1028),
.B1(n_1023),
.B2(n_992),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1194),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1287),
.A2(n_1049),
.B(n_1030),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1287),
.A2(n_1049),
.B(n_1030),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1325),
.B(n_1096),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1284),
.B(n_1096),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1225),
.A2(n_1043),
.B(n_1086),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1271),
.A2(n_1002),
.B1(n_989),
.B2(n_1012),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1284),
.B(n_1096),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1272),
.A2(n_989),
.B1(n_1019),
.B2(n_1140),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1279),
.A2(n_1030),
.B(n_1049),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1194),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1279),
.A2(n_1071),
.B(n_1161),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1250),
.Y(n_1391)
);

BUFx3_ASAP7_75t_L g1392 ( 
.A(n_1217),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1256),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1269),
.A2(n_1071),
.B(n_1161),
.Y(n_1394)
);

OAI21xp5_ASAP7_75t_L g1395 ( 
.A1(n_1187),
.A2(n_992),
.B(n_1080),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1296),
.A2(n_1037),
.B(n_1079),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_L g1397 ( 
.A1(n_1269),
.A2(n_1071),
.B(n_1161),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1250),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1344),
.A2(n_1069),
.B(n_1142),
.C(n_1133),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1190),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1277),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1277),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1309),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1185),
.A2(n_1080),
.B(n_1037),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1186),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1207),
.B(n_1166),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1309),
.Y(n_1407)
);

NAND2x1p5_ASAP7_75t_L g1408 ( 
.A(n_1196),
.B(n_1043),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1257),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1258),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1292),
.B(n_1166),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1217),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1327),
.A2(n_1028),
.B1(n_1069),
.B2(n_1043),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1213),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1225),
.A2(n_1043),
.B(n_1086),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1244),
.Y(n_1416)
);

NAND2x1p5_ASAP7_75t_L g1417 ( 
.A(n_1196),
.B(n_1043),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_SL g1418 ( 
.A1(n_1191),
.A2(n_1151),
.B(n_1127),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1274),
.A2(n_1245),
.B(n_1244),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1285),
.Y(n_1420)
);

AOI221xp5_ASAP7_75t_L g1421 ( 
.A1(n_1266),
.A2(n_1173),
.B1(n_329),
.B2(n_343),
.C(n_356),
.Y(n_1421)
);

AND2x4_ASAP7_75t_L g1422 ( 
.A(n_1346),
.B(n_1028),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1256),
.Y(n_1423)
);

BUFx2_ASAP7_75t_L g1424 ( 
.A(n_1276),
.Y(n_1424)
);

OA21x2_ASAP7_75t_L g1425 ( 
.A1(n_1185),
.A2(n_1080),
.B(n_1037),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1248),
.Y(n_1426)
);

AND2x4_ASAP7_75t_L g1427 ( 
.A(n_1346),
.B(n_1029),
.Y(n_1427)
);

NAND3xp33_ASAP7_75t_L g1428 ( 
.A(n_1344),
.B(n_1177),
.C(n_1104),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1245),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1262),
.Y(n_1430)
);

NAND2x1p5_ASAP7_75t_L g1431 ( 
.A(n_1196),
.B(n_1086),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1274),
.A2(n_1161),
.B(n_1148),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1321),
.A2(n_1124),
.B(n_1044),
.C(n_1058),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1261),
.B(n_1316),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1261),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1262),
.A2(n_1148),
.B(n_1146),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1240),
.A2(n_1226),
.B(n_1247),
.Y(n_1437)
);

OAI21x1_ASAP7_75t_SL g1438 ( 
.A1(n_1332),
.A2(n_1127),
.B(n_1034),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1240),
.A2(n_1226),
.B(n_1247),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1210),
.A2(n_1148),
.B(n_1146),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1182),
.A2(n_1079),
.B(n_1032),
.Y(n_1441)
);

NAND2xp33_ASAP7_75t_L g1442 ( 
.A(n_1211),
.B(n_1086),
.Y(n_1442)
);

INVx3_ASAP7_75t_L g1443 ( 
.A(n_1211),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1248),
.Y(n_1444)
);

OR2x6_ASAP7_75t_L g1445 ( 
.A(n_1319),
.B(n_1039),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1207),
.A2(n_1166),
.B1(n_1127),
.B2(n_1171),
.Y(n_1446)
);

OA21x2_ASAP7_75t_L g1447 ( 
.A1(n_1182),
.A2(n_1079),
.B(n_1032),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1211),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1301),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1255),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1184),
.Y(n_1451)
);

CKINVDCx11_ASAP7_75t_R g1452 ( 
.A(n_1193),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1210),
.A2(n_1148),
.B(n_1146),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1188),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1222),
.B(n_1166),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1255),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1224),
.Y(n_1457)
);

OAI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1323),
.A2(n_1034),
.B1(n_1024),
.B2(n_1042),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1224),
.Y(n_1459)
);

OAI21xp5_ASAP7_75t_L g1460 ( 
.A1(n_1239),
.A2(n_1032),
.B(n_1153),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1236),
.B(n_1135),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1200),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1301),
.Y(n_1463)
);

AO21x2_ASAP7_75t_L g1464 ( 
.A1(n_1204),
.A2(n_1173),
.B(n_1153),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1292),
.A2(n_1135),
.B1(n_363),
.B2(n_376),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1336),
.Y(n_1466)
);

OAI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1230),
.A2(n_1148),
.B(n_1146),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1206),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1219),
.A2(n_1000),
.B(n_1004),
.Y(n_1469)
);

AND2x4_ASAP7_75t_L g1470 ( 
.A(n_1299),
.B(n_1039),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1336),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1231),
.Y(n_1472)
);

OA21x2_ASAP7_75t_L g1473 ( 
.A1(n_1307),
.A2(n_421),
.B(n_391),
.Y(n_1473)
);

BUFx12f_ASAP7_75t_L g1474 ( 
.A(n_1263),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1235),
.A2(n_1135),
.B1(n_363),
.B2(n_344),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1299),
.B(n_1039),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1230),
.A2(n_1135),
.B(n_1053),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1338),
.A2(n_1084),
.B1(n_1070),
.B2(n_1044),
.Y(n_1478)
);

OAI21x1_ASAP7_75t_L g1479 ( 
.A1(n_1237),
.A2(n_1039),
.B(n_1004),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1268),
.B(n_1130),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1307),
.A2(n_409),
.B(n_375),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1219),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1190),
.Y(n_1483)
);

INVx2_ASAP7_75t_L g1484 ( 
.A(n_1336),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1222),
.B(n_1130),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1231),
.Y(n_1486)
);

AOI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1233),
.A2(n_1288),
.B(n_1218),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1231),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1270),
.B(n_1130),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1208),
.A2(n_405),
.B(n_385),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1270),
.B(n_1132),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1339),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1336),
.Y(n_1493)
);

OAI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1315),
.A2(n_1139),
.B(n_1132),
.Y(n_1494)
);

OAI21x1_ASAP7_75t_L g1495 ( 
.A1(n_1237),
.A2(n_1139),
.B(n_1132),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1238),
.A2(n_103),
.B(n_100),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1342),
.B(n_1293),
.Y(n_1497)
);

A2O1A1Ixp33_ASAP7_75t_L g1498 ( 
.A1(n_1340),
.A2(n_1058),
.B(n_360),
.C(n_410),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1236),
.B(n_388),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1236),
.B(n_363),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1235),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1268),
.B(n_399),
.Y(n_1502)
);

AND2x2_ASAP7_75t_SL g1503 ( 
.A(n_1310),
.B(n_1048),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1209),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1238),
.A2(n_168),
.B(n_104),
.Y(n_1505)
);

INVx1_ASAP7_75t_SL g1506 ( 
.A(n_1278),
.Y(n_1506)
);

OAI222xp33_ASAP7_75t_L g1507 ( 
.A1(n_1302),
.A2(n_402),
.B1(n_400),
.B2(n_418),
.C1(n_419),
.C2(n_423),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1231),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_1280),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1295),
.A2(n_179),
.B(n_109),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1295),
.A2(n_181),
.B(n_110),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1294),
.B(n_425),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1203),
.Y(n_1513)
);

AO31x2_ASAP7_75t_L g1514 ( 
.A1(n_1333),
.A2(n_24),
.A3(n_28),
.B(n_31),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1281),
.A2(n_1089),
.B1(n_412),
.B2(n_376),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_SL g1516 ( 
.A(n_1193),
.B(n_412),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1231),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_SL g1518 ( 
.A1(n_1223),
.A2(n_213),
.B(n_210),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_SL g1519 ( 
.A1(n_1282),
.A2(n_1089),
.B1(n_412),
.B2(n_376),
.Y(n_1519)
);

AOI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1219),
.A2(n_591),
.B(n_206),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1208),
.A2(n_591),
.B(n_32),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1221),
.A2(n_205),
.B(n_200),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1263),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1195),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_SL g1525 ( 
.A1(n_1519),
.A2(n_1353),
.B1(n_1351),
.B2(n_1503),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1360),
.A2(n_1246),
.B1(n_1334),
.B2(n_1232),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1406),
.B(n_1312),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1406),
.B(n_1312),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1350),
.A2(n_1308),
.B(n_1318),
.Y(n_1529)
);

OR2x6_ASAP7_75t_SL g1530 ( 
.A(n_1393),
.B(n_1251),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1485),
.B(n_1236),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1485),
.B(n_1236),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1361),
.A2(n_1286),
.B1(n_1324),
.B2(n_1270),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1455),
.B(n_1322),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1427),
.B(n_1290),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1451),
.Y(n_1536)
);

AND2x4_ASAP7_75t_L g1537 ( 
.A(n_1427),
.B(n_1290),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1455),
.B(n_1322),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1449),
.B(n_1322),
.Y(n_1539)
);

NAND2x1p5_ASAP7_75t_L g1540 ( 
.A(n_1443),
.B(n_1203),
.Y(n_1540)
);

NOR2xp33_ASAP7_75t_L g1541 ( 
.A(n_1509),
.B(n_1308),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1451),
.Y(n_1542)
);

BUFx3_ASAP7_75t_L g1543 ( 
.A(n_1376),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1500),
.A2(n_1333),
.B1(n_1304),
.B2(n_1220),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1463),
.A2(n_1515),
.B1(n_1410),
.B2(n_1366),
.Y(n_1545)
);

OAI21x1_ASAP7_75t_L g1546 ( 
.A1(n_1437),
.A2(n_1313),
.B(n_1330),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1377),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1497),
.B(n_1322),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1442),
.A2(n_1214),
.B(n_1252),
.Y(n_1549)
);

OAI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1363),
.A2(n_1387),
.B1(n_1446),
.B2(n_1368),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1362),
.A2(n_1357),
.B1(n_1385),
.B2(n_1358),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1500),
.A2(n_1304),
.B1(n_1318),
.B2(n_1329),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1452),
.Y(n_1553)
);

NOR2xp33_ASAP7_75t_R g1554 ( 
.A(n_1393),
.B(n_1203),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_SL g1555 ( 
.A1(n_1503),
.A2(n_1304),
.B1(n_1343),
.B2(n_1335),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1410),
.B(n_1329),
.Y(n_1556)
);

INVx3_ASAP7_75t_L g1557 ( 
.A(n_1489),
.Y(n_1557)
);

NAND2xp33_ASAP7_75t_SL g1558 ( 
.A(n_1422),
.B(n_1203),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1454),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1373),
.Y(n_1560)
);

NAND2x1p5_ASAP7_75t_L g1561 ( 
.A(n_1443),
.B(n_1328),
.Y(n_1561)
);

AOI21xp33_ASAP7_75t_L g1562 ( 
.A1(n_1399),
.A2(n_1265),
.B(n_1195),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1503),
.A2(n_1343),
.B1(n_1335),
.B2(n_1313),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1502),
.B(n_1322),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1362),
.B(n_1345),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1419),
.A2(n_1330),
.B(n_1306),
.Y(n_1566)
);

AO31x2_ASAP7_75t_L g1567 ( 
.A1(n_1472),
.A2(n_1228),
.A3(n_1243),
.B(n_1242),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1462),
.Y(n_1568)
);

CKINVDCx8_ASAP7_75t_R g1569 ( 
.A(n_1367),
.Y(n_1569)
);

AOI221xp5_ASAP7_75t_L g1570 ( 
.A1(n_1507),
.A2(n_1297),
.B1(n_1305),
.B2(n_1331),
.C(n_1317),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1437),
.A2(n_1306),
.B(n_1221),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1362),
.B(n_1345),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1349),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1424),
.B(n_1212),
.Y(n_1574)
);

AOI21xp5_ASAP7_75t_L g1575 ( 
.A1(n_1442),
.A2(n_1214),
.B(n_1195),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1349),
.Y(n_1576)
);

INVx3_ASAP7_75t_L g1577 ( 
.A(n_1489),
.Y(n_1577)
);

INVx3_ASAP7_75t_L g1578 ( 
.A(n_1489),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1384),
.A2(n_1189),
.B(n_1260),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1424),
.B(n_1377),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_L g1581 ( 
.A1(n_1499),
.A2(n_1234),
.B1(n_1189),
.B2(n_1275),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1491),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1359),
.B(n_1345),
.Y(n_1583)
);

INVxp33_ASAP7_75t_L g1584 ( 
.A(n_1409),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1499),
.A2(n_1273),
.B1(n_1267),
.B2(n_1337),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1461),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1480),
.B(n_1337),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1439),
.A2(n_1289),
.B(n_1291),
.Y(n_1589)
);

CKINVDCx8_ASAP7_75t_R g1590 ( 
.A(n_1367),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1468),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1375),
.Y(n_1592)
);

HB1xp67_ASAP7_75t_L g1593 ( 
.A(n_1461),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1422),
.A2(n_1328),
.B1(n_1326),
.B2(n_1314),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1411),
.B(n_1314),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1382),
.B(n_1212),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1414),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1512),
.B(n_1422),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1504),
.B(n_1501),
.Y(n_1599)
);

INVx6_ASAP7_75t_L g1600 ( 
.A(n_1474),
.Y(n_1600)
);

CKINVDCx20_ASAP7_75t_R g1601 ( 
.A(n_1373),
.Y(n_1601)
);

BUFx10_ASAP7_75t_L g1602 ( 
.A(n_1423),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1414),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1435),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1501),
.B(n_1345),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_SL g1606 ( 
.A(n_1427),
.B(n_1328),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1423),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1458),
.A2(n_1328),
.B1(n_1341),
.B2(n_1229),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1375),
.Y(n_1609)
);

NOR2xp33_ASAP7_75t_SL g1610 ( 
.A(n_1523),
.B(n_1229),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1379),
.Y(n_1611)
);

OAI22xp33_ASAP7_75t_L g1612 ( 
.A1(n_1492),
.A2(n_1341),
.B1(n_1311),
.B2(n_1212),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1376),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1440),
.A2(n_1291),
.B(n_1289),
.Y(n_1614)
);

AOI221xp5_ASAP7_75t_L g1615 ( 
.A1(n_1433),
.A2(n_1254),
.B1(n_1212),
.B2(n_33),
.C(n_35),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1392),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1405),
.B(n_1212),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1405),
.B(n_1341),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1491),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1379),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1428),
.A2(n_1341),
.B1(n_1249),
.B2(n_33),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1475),
.A2(n_1249),
.B1(n_32),
.B2(n_39),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1420),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1389),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1465),
.A2(n_1249),
.B1(n_39),
.B2(n_40),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1391),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1439),
.A2(n_1453),
.B(n_1440),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1391),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1516),
.A2(n_28),
.B1(n_40),
.B2(n_42),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1398),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1506),
.B(n_1249),
.Y(n_1631)
);

INVx2_ASAP7_75t_L g1632 ( 
.A(n_1398),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1392),
.B(n_42),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1347),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_1634)
);

INVxp33_ASAP7_75t_L g1635 ( 
.A(n_1434),
.Y(n_1635)
);

INVx2_ASAP7_75t_L g1636 ( 
.A(n_1401),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1419),
.A2(n_44),
.B(n_45),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1389),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1412),
.B(n_47),
.Y(n_1639)
);

AOI222xp33_ASAP7_75t_L g1640 ( 
.A1(n_1421),
.A2(n_47),
.B1(n_50),
.B2(n_52),
.C1(n_54),
.C2(n_55),
.Y(n_1640)
);

AOI22xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1418),
.A2(n_1347),
.B1(n_1474),
.B2(n_1378),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1412),
.B(n_54),
.Y(n_1642)
);

NAND2xp33_ASAP7_75t_R g1643 ( 
.A(n_1445),
.B(n_187),
.Y(n_1643)
);

CKINVDCx6p67_ASAP7_75t_R g1644 ( 
.A(n_1470),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1356),
.B(n_55),
.Y(n_1645)
);

A2O1A1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1498),
.A2(n_1352),
.B(n_1460),
.C(n_1395),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1470),
.Y(n_1647)
);

OAI22xp5_ASAP7_75t_L g1648 ( 
.A1(n_1478),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1648)
);

AOI22xp33_ASAP7_75t_L g1649 ( 
.A1(n_1418),
.A2(n_56),
.B1(n_62),
.B2(n_63),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1356),
.A2(n_64),
.B1(n_67),
.B2(n_69),
.Y(n_1650)
);

AOI22xp33_ASAP7_75t_L g1651 ( 
.A1(n_1472),
.A2(n_69),
.B1(n_70),
.B2(n_72),
.Y(n_1651)
);

AND2x4_ASAP7_75t_SL g1652 ( 
.A(n_1470),
.B(n_101),
.Y(n_1652)
);

NOR2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1523),
.B(n_167),
.Y(n_1653)
);

NOR3xp33_ASAP7_75t_SL g1654 ( 
.A(n_1413),
.B(n_72),
.C(n_74),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1401),
.B(n_1407),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1445),
.B(n_1402),
.Y(n_1656)
);

AOI22xp33_ASAP7_75t_L g1657 ( 
.A1(n_1486),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1491),
.B(n_122),
.Y(n_1658)
);

NOR2xp33_ASAP7_75t_SL g1659 ( 
.A(n_1476),
.B(n_128),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1355),
.Y(n_1660)
);

AOI22xp33_ASAP7_75t_SL g1661 ( 
.A1(n_1438),
.A2(n_80),
.B1(n_83),
.B2(n_88),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1407),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_R g1663 ( 
.A(n_1355),
.B(n_153),
.Y(n_1663)
);

INVx2_ASAP7_75t_SL g1664 ( 
.A(n_1476),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1494),
.A2(n_89),
.B1(n_154),
.B2(n_164),
.Y(n_1665)
);

INVx5_ASAP7_75t_L g1666 ( 
.A(n_1355),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1415),
.A2(n_1372),
.B(n_1447),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1476),
.B(n_1445),
.Y(n_1668)
);

INVx3_ASAP7_75t_L g1669 ( 
.A(n_1355),
.Y(n_1669)
);

BUFx6f_ASAP7_75t_SL g1670 ( 
.A(n_1445),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1403),
.B(n_1355),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_1370),
.Y(n_1673)
);

NOR2x1_ASAP7_75t_SL g1674 ( 
.A(n_1364),
.B(n_1396),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1370),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1466),
.Y(n_1676)
);

AOI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1441),
.A2(n_1447),
.B(n_1408),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1466),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_L g1679 ( 
.A1(n_1486),
.A2(n_1488),
.B1(n_1508),
.B2(n_1517),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1370),
.Y(n_1680)
);

HB1xp67_ASAP7_75t_L g1681 ( 
.A(n_1471),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1488),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1431),
.A2(n_1417),
.B1(n_1408),
.B2(n_1493),
.Y(n_1683)
);

OAI222xp33_ASAP7_75t_L g1684 ( 
.A1(n_1508),
.A2(n_1517),
.B1(n_1520),
.B2(n_1471),
.C1(n_1493),
.C2(n_1484),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1464),
.B(n_1369),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1370),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1370),
.B(n_1400),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1400),
.B(n_1483),
.Y(n_1688)
);

OAI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1431),
.A2(n_1408),
.B1(n_1417),
.B2(n_1484),
.Y(n_1689)
);

NOR2xp33_ASAP7_75t_L g1690 ( 
.A(n_1464),
.B(n_1396),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_SL g1691 ( 
.A(n_1400),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1416),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1438),
.A2(n_1518),
.B1(n_1371),
.B2(n_1364),
.Y(n_1693)
);

CKINVDCx5p33_ASAP7_75t_R g1694 ( 
.A(n_1400),
.Y(n_1694)
);

CKINVDCx14_ASAP7_75t_R g1695 ( 
.A(n_1400),
.Y(n_1695)
);

AO31x2_ASAP7_75t_L g1696 ( 
.A1(n_1426),
.A2(n_1444),
.A3(n_1456),
.B(n_1450),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1697)
);

AOI21xp5_ASAP7_75t_L g1698 ( 
.A1(n_1441),
.A2(n_1447),
.B(n_1417),
.Y(n_1698)
);

BUFx2_ASAP7_75t_L g1699 ( 
.A(n_1483),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1416),
.Y(n_1700)
);

BUFx2_ASAP7_75t_L g1701 ( 
.A(n_1483),
.Y(n_1701)
);

INVx5_ASAP7_75t_L g1702 ( 
.A(n_1483),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1483),
.Y(n_1703)
);

AO31x2_ASAP7_75t_L g1704 ( 
.A1(n_1426),
.A2(n_1444),
.A3(n_1450),
.B(n_1456),
.Y(n_1704)
);

AND2x4_ASAP7_75t_L g1705 ( 
.A(n_1513),
.B(n_1495),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1513),
.B(n_1514),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1513),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1513),
.B(n_1495),
.Y(n_1708)
);

OAI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1431),
.A2(n_1482),
.B1(n_1448),
.B2(n_1469),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1513),
.B(n_1514),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1473),
.A2(n_1481),
.B1(n_1490),
.B2(n_1425),
.C(n_1404),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1369),
.Y(n_1712)
);

OAI221xp5_ASAP7_75t_L g1713 ( 
.A1(n_1525),
.A2(n_1490),
.B1(n_1473),
.B2(n_1481),
.C(n_1425),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1640),
.A2(n_1649),
.B1(n_1550),
.B2(n_1648),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1671),
.Y(n_1715)
);

OAI33xp33_ASAP7_75t_L g1716 ( 
.A1(n_1650),
.A2(n_1545),
.A3(n_1622),
.B1(n_1625),
.B2(n_1639),
.B3(n_1631),
.Y(n_1716)
);

A2O1A1Ixp33_ASAP7_75t_L g1717 ( 
.A1(n_1646),
.A2(n_1522),
.B(n_1505),
.C(n_1496),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1634),
.A2(n_1518),
.B1(n_1524),
.B2(n_1429),
.C(n_1430),
.Y(n_1718)
);

OAI211xp5_ASAP7_75t_L g1719 ( 
.A1(n_1629),
.A2(n_1473),
.B(n_1481),
.C(n_1490),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1667),
.A2(n_1453),
.B(n_1354),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1536),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1668),
.B(n_1448),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1542),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1574),
.B(n_1369),
.Y(n_1724)
);

AOI211xp5_ASAP7_75t_L g1725 ( 
.A1(n_1545),
.A2(n_1522),
.B(n_1505),
.C(n_1496),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_R g1726 ( 
.A(n_1643),
.B(n_1569),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1584),
.B(n_1482),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1559),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1543),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1634),
.A2(n_1481),
.B1(n_1473),
.B2(n_1425),
.Y(n_1730)
);

BUFx12f_ASAP7_75t_L g1731 ( 
.A(n_1553),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1527),
.B(n_1514),
.Y(n_1732)
);

OR2x6_ASAP7_75t_L g1733 ( 
.A(n_1549),
.B(n_1348),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1659),
.A2(n_1645),
.B1(n_1663),
.B2(n_1665),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1587),
.B(n_1514),
.Y(n_1735)
);

AOI222xp33_ASAP7_75t_L g1736 ( 
.A1(n_1651),
.A2(n_1657),
.B1(n_1629),
.B2(n_1649),
.C1(n_1645),
.C2(n_1615),
.Y(n_1736)
);

AO21x2_ASAP7_75t_L g1737 ( 
.A1(n_1562),
.A2(n_1487),
.B(n_1429),
.Y(n_1737)
);

AOI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1651),
.A2(n_1524),
.B1(n_1430),
.B2(n_1457),
.C(n_1459),
.Y(n_1738)
);

HB1xp67_ASAP7_75t_L g1739 ( 
.A(n_1678),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1646),
.A2(n_1348),
.B(n_1511),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1541),
.B(n_1514),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_L g1742 ( 
.A(n_1660),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1608),
.A2(n_1482),
.B1(n_1425),
.B2(n_1404),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1553),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1604),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1661),
.A2(n_1490),
.B1(n_1404),
.B2(n_1441),
.C(n_1447),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1657),
.A2(n_1459),
.B1(n_1457),
.B2(n_1369),
.C(n_1404),
.Y(n_1747)
);

AOI21xp33_ASAP7_75t_L g1748 ( 
.A1(n_1526),
.A2(n_1441),
.B(n_1521),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1528),
.A2(n_1521),
.B1(n_1511),
.B2(n_1510),
.Y(n_1749)
);

AOI22xp33_ASAP7_75t_SL g1750 ( 
.A1(n_1663),
.A2(n_1521),
.B1(n_1510),
.B2(n_1467),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1568),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_SL g1752 ( 
.A1(n_1548),
.A2(n_1467),
.B1(n_1436),
.B2(n_1354),
.Y(n_1752)
);

OAI21xp33_ASAP7_75t_L g1753 ( 
.A1(n_1654),
.A2(n_1365),
.B(n_1374),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1647),
.B(n_1477),
.Y(n_1754)
);

BUFx6f_ASAP7_75t_L g1755 ( 
.A(n_1660),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1575),
.B(n_1477),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1598),
.A2(n_1380),
.B1(n_1381),
.B2(n_1479),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_L g1758 ( 
.A1(n_1551),
.A2(n_1541),
.B1(n_1564),
.B2(n_1533),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1584),
.A2(n_1380),
.B1(n_1381),
.B2(n_1394),
.C(n_1397),
.Y(n_1759)
);

AOI222xp33_ASAP7_75t_L g1760 ( 
.A1(n_1531),
.A2(n_1394),
.B1(n_1397),
.B2(n_1388),
.C1(n_1390),
.C2(n_1432),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1591),
.Y(n_1761)
);

AOI22xp5_ASAP7_75t_L g1762 ( 
.A1(n_1601),
.A2(n_1479),
.B1(n_1390),
.B2(n_1388),
.Y(n_1762)
);

A2O1A1Ixp33_ASAP7_75t_L g1763 ( 
.A1(n_1621),
.A2(n_1570),
.B(n_1641),
.C(n_1529),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1597),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_L g1765 ( 
.A1(n_1608),
.A2(n_1432),
.B1(n_1436),
.B2(n_1635),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1599),
.B(n_1539),
.Y(n_1766)
);

AOI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1635),
.A2(n_1653),
.B1(n_1601),
.B2(n_1556),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1560),
.A2(n_1600),
.B1(n_1532),
.B2(n_1547),
.Y(n_1768)
);

AOI21xp33_ASAP7_75t_L g1769 ( 
.A1(n_1612),
.A2(n_1588),
.B(n_1596),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1590),
.A2(n_1580),
.B1(n_1560),
.B2(n_1588),
.Y(n_1770)
);

CKINVDCx11_ASAP7_75t_R g1771 ( 
.A(n_1607),
.Y(n_1771)
);

CKINVDCx20_ASAP7_75t_R g1772 ( 
.A(n_1644),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1600),
.A2(n_1633),
.B1(n_1642),
.B2(n_1583),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1579),
.A2(n_1558),
.B(n_1698),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1605),
.B(n_1534),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1658),
.A2(n_1670),
.B1(n_1538),
.B2(n_1647),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1618),
.B(n_1672),
.Y(n_1777)
);

OAI211xp5_ASAP7_75t_L g1778 ( 
.A1(n_1544),
.A2(n_1555),
.B(n_1563),
.C(n_1637),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1607),
.B(n_1543),
.Y(n_1779)
);

INVx4_ASAP7_75t_L g1780 ( 
.A(n_1666),
.Y(n_1780)
);

AO31x2_ASAP7_75t_L g1781 ( 
.A1(n_1674),
.A2(n_1690),
.A3(n_1677),
.B(n_1712),
.Y(n_1781)
);

BUFx12f_ASAP7_75t_L g1782 ( 
.A(n_1602),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1595),
.B(n_1664),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1558),
.A2(n_1544),
.B(n_1606),
.C(n_1652),
.Y(n_1784)
);

OAI221xp5_ASAP7_75t_L g1785 ( 
.A1(n_1643),
.A2(n_1600),
.B1(n_1552),
.B2(n_1693),
.C(n_1610),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1670),
.A2(n_1616),
.B1(n_1613),
.B2(n_1585),
.Y(n_1786)
);

OAI211xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1693),
.A2(n_1552),
.B(n_1711),
.C(n_1617),
.Y(n_1787)
);

OAI22xp33_ASAP7_75t_L g1788 ( 
.A1(n_1637),
.A2(n_1656),
.B1(n_1603),
.B2(n_1623),
.Y(n_1788)
);

OA21x2_ASAP7_75t_L g1789 ( 
.A1(n_1546),
.A2(n_1571),
.B(n_1627),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1602),
.Y(n_1790)
);

HB1xp67_ASAP7_75t_L g1791 ( 
.A(n_1678),
.Y(n_1791)
);

OAI211xp5_ASAP7_75t_L g1792 ( 
.A1(n_1637),
.A2(n_1581),
.B(n_1585),
.C(n_1554),
.Y(n_1792)
);

INVx3_ASAP7_75t_L g1793 ( 
.A(n_1660),
.Y(n_1793)
);

AOI222xp33_ASAP7_75t_L g1794 ( 
.A1(n_1586),
.A2(n_1593),
.B1(n_1658),
.B2(n_1612),
.C1(n_1572),
.C2(n_1565),
.Y(n_1794)
);

OAI22xp33_ASAP7_75t_L g1795 ( 
.A1(n_1613),
.A2(n_1616),
.B1(n_1586),
.B2(n_1593),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1557),
.B(n_1577),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1658),
.A2(n_1581),
.B1(n_1652),
.B2(n_1638),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1624),
.A2(n_1578),
.B1(n_1582),
.B2(n_1557),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1594),
.A2(n_1577),
.B1(n_1578),
.B2(n_1582),
.Y(n_1799)
);

OAI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1619),
.A2(n_1694),
.B1(n_1673),
.B2(n_1702),
.Y(n_1800)
);

OAI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1619),
.A2(n_1694),
.B1(n_1673),
.B2(n_1702),
.Y(n_1801)
);

AOI22xp33_ASAP7_75t_L g1802 ( 
.A1(n_1602),
.A2(n_1535),
.B1(n_1537),
.B2(n_1606),
.Y(n_1802)
);

OAI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1554),
.A2(n_1690),
.B(n_1697),
.C(n_1679),
.Y(n_1803)
);

OA21x2_ASAP7_75t_L g1804 ( 
.A1(n_1684),
.A2(n_1685),
.B(n_1589),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1682),
.B(n_1687),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1688),
.B(n_1535),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1691),
.A2(n_1695),
.B1(n_1530),
.B2(n_1537),
.Y(n_1807)
);

BUFx8_ASAP7_75t_L g1808 ( 
.A(n_1699),
.Y(n_1808)
);

AOI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1535),
.A2(n_1537),
.B1(n_1662),
.B2(n_1636),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1573),
.A2(n_1630),
.B1(n_1662),
.B2(n_1636),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1576),
.B(n_1628),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1701),
.B(n_1695),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1709),
.A2(n_1689),
.B(n_1683),
.Y(n_1813)
);

CKINVDCx6p67_ASAP7_75t_R g1814 ( 
.A(n_1666),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1576),
.A2(n_1620),
.B1(n_1632),
.B2(n_1630),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1675),
.A2(n_1703),
.B(n_1655),
.Y(n_1816)
);

OAI211xp5_ASAP7_75t_SL g1817 ( 
.A1(n_1679),
.A2(n_1592),
.B(n_1626),
.C(n_1632),
.Y(n_1817)
);

INVxp33_ASAP7_75t_L g1818 ( 
.A(n_1660),
.Y(n_1818)
);

AOI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1706),
.A2(n_1710),
.B1(n_1681),
.B2(n_1628),
.C(n_1626),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1705),
.A2(n_1708),
.B1(n_1609),
.B2(n_1611),
.Y(n_1820)
);

OAI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1666),
.A2(n_1702),
.B1(n_1620),
.B2(n_1609),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1705),
.A2(n_1708),
.B1(n_1686),
.B2(n_1680),
.Y(n_1822)
);

OAI22xp5_ASAP7_75t_L g1823 ( 
.A1(n_1540),
.A2(n_1561),
.B1(n_1702),
.B2(n_1666),
.Y(n_1823)
);

BUFx12f_ASAP7_75t_L g1824 ( 
.A(n_1707),
.Y(n_1824)
);

AOI221xp5_ASAP7_75t_L g1825 ( 
.A1(n_1681),
.A2(n_1611),
.B1(n_1592),
.B2(n_1676),
.C(n_1708),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1669),
.B(n_1680),
.Y(n_1826)
);

AOI221xp5_ASAP7_75t_L g1827 ( 
.A1(n_1705),
.A2(n_1692),
.B1(n_1700),
.B2(n_1707),
.C(n_1561),
.Y(n_1827)
);

AOI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1692),
.A2(n_1700),
.B1(n_1707),
.B2(n_1540),
.C(n_1567),
.Y(n_1828)
);

OR2x2_ASAP7_75t_L g1829 ( 
.A(n_1696),
.B(n_1704),
.Y(n_1829)
);

CKINVDCx5p33_ASAP7_75t_R g1830 ( 
.A(n_1704),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1566),
.A2(n_1614),
.B1(n_1567),
.B2(n_1704),
.Y(n_1831)
);

AND2x4_ASAP7_75t_L g1832 ( 
.A(n_1704),
.B(n_1567),
.Y(n_1832)
);

AOI221xp5_ASAP7_75t_L g1833 ( 
.A1(n_1567),
.A2(n_884),
.B1(n_666),
.B2(n_668),
.C(n_1035),
.Y(n_1833)
);

INVx3_ASAP7_75t_L g1834 ( 
.A(n_1566),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1640),
.A2(n_1198),
.B1(n_1052),
.B2(n_1525),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1671),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1640),
.A2(n_1198),
.B1(n_1052),
.B2(n_1525),
.Y(n_1837)
);

AOI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1640),
.A2(n_1198),
.B1(n_1052),
.B2(n_1525),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1640),
.A2(n_1198),
.B1(n_1052),
.B2(n_1525),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1634),
.A2(n_884),
.B1(n_666),
.B2(n_668),
.C(n_1035),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1574),
.B(n_1587),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1525),
.A2(n_1035),
.B1(n_1018),
.B2(n_1205),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1640),
.A2(n_1198),
.B1(n_1052),
.B2(n_1525),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1640),
.A2(n_1198),
.B1(n_1052),
.B2(n_1525),
.Y(n_1844)
);

OAI22xp5_ASAP7_75t_L g1845 ( 
.A1(n_1525),
.A2(n_1035),
.B1(n_1018),
.B2(n_1205),
.Y(n_1845)
);

CKINVDCx6p67_ASAP7_75t_R g1846 ( 
.A(n_1553),
.Y(n_1846)
);

OA21x2_ASAP7_75t_L g1847 ( 
.A1(n_1667),
.A2(n_1562),
.B(n_1579),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1587),
.B(n_1351),
.Y(n_1848)
);

OAI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1643),
.A2(n_1351),
.B1(n_862),
.B2(n_1659),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1587),
.B(n_1351),
.Y(n_1850)
);

BUFx2_ASAP7_75t_L g1851 ( 
.A(n_1543),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1553),
.Y(n_1852)
);

OR2x6_ASAP7_75t_L g1853 ( 
.A(n_1549),
.B(n_1575),
.Y(n_1853)
);

AOI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1545),
.A2(n_1035),
.B(n_1018),
.C(n_884),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1536),
.Y(n_1855)
);

AOI222xp33_ASAP7_75t_L g1856 ( 
.A1(n_1650),
.A2(n_1198),
.B1(n_1052),
.B2(n_666),
.C1(n_668),
.C2(n_606),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1525),
.A2(n_1052),
.B1(n_1640),
.B2(n_1035),
.Y(n_1857)
);

INVx5_ASAP7_75t_L g1858 ( 
.A(n_1660),
.Y(n_1858)
);

AOI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1525),
.A2(n_1018),
.B(n_1035),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1525),
.A2(n_1052),
.B1(n_1640),
.B2(n_1035),
.Y(n_1860)
);

OAI221xp5_ASAP7_75t_SL g1861 ( 
.A1(n_1634),
.A2(n_1198),
.B1(n_826),
.B2(n_1018),
.C(n_586),
.Y(n_1861)
);

INVx6_ASAP7_75t_L g1862 ( 
.A(n_1613),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1634),
.A2(n_884),
.B1(n_666),
.B2(n_668),
.C(n_1035),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1574),
.B(n_1587),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1527),
.B(n_1528),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1525),
.A2(n_1052),
.B1(n_1640),
.B2(n_1035),
.Y(n_1866)
);

AOI22xp33_ASAP7_75t_L g1867 ( 
.A1(n_1525),
.A2(n_1052),
.B1(n_1640),
.B2(n_1035),
.Y(n_1867)
);

OAI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1525),
.A2(n_1035),
.B1(n_1018),
.B2(n_1205),
.Y(n_1868)
);

OAI211xp5_ASAP7_75t_SL g1869 ( 
.A1(n_1640),
.A2(n_1525),
.B(n_1353),
.C(n_1320),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1525),
.A2(n_1035),
.B1(n_1018),
.B2(n_1205),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1574),
.B(n_1587),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1671),
.Y(n_1872)
);

BUFx3_ASAP7_75t_L g1873 ( 
.A(n_1543),
.Y(n_1873)
);

OA21x2_ASAP7_75t_L g1874 ( 
.A1(n_1667),
.A2(n_1562),
.B(n_1579),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1830),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1832),
.B(n_1732),
.Y(n_1876)
);

NOR2x1_ASAP7_75t_L g1877 ( 
.A(n_1795),
.B(n_1785),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1832),
.B(n_1775),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1745),
.B(n_1848),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1829),
.Y(n_1880)
);

INVx4_ASAP7_75t_L g1881 ( 
.A(n_1858),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1834),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1834),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1781),
.B(n_1804),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1781),
.B(n_1804),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1735),
.B(n_1741),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1715),
.B(n_1836),
.Y(n_1887)
);

AOI22xp33_ASAP7_75t_L g1888 ( 
.A1(n_1869),
.A2(n_1837),
.B1(n_1844),
.B2(n_1835),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1739),
.Y(n_1889)
);

AO31x2_ASAP7_75t_L g1890 ( 
.A1(n_1717),
.A2(n_1743),
.A3(n_1774),
.B(n_1763),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1723),
.Y(n_1891)
);

OAI33xp33_ASAP7_75t_L g1892 ( 
.A1(n_1842),
.A2(n_1845),
.A3(n_1868),
.B1(n_1870),
.B2(n_1869),
.B3(n_1770),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1728),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1781),
.B(n_1865),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1751),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1761),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1872),
.B(n_1841),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1781),
.Y(n_1898)
);

OR2x2_ASAP7_75t_L g1899 ( 
.A(n_1724),
.B(n_1864),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1764),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1853),
.B(n_1831),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1853),
.B(n_1831),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_L g1903 ( 
.A1(n_1835),
.A2(n_1839),
.B1(n_1837),
.B2(n_1838),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1789),
.Y(n_1904)
);

AOI33xp33_ASAP7_75t_L g1905 ( 
.A1(n_1838),
.A2(n_1843),
.A3(n_1844),
.B1(n_1839),
.B2(n_1854),
.B3(n_1857),
.Y(n_1905)
);

INVx5_ASAP7_75t_L g1906 ( 
.A(n_1853),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1756),
.B(n_1847),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1847),
.B(n_1874),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1874),
.B(n_1737),
.Y(n_1909)
);

BUFx3_ASAP7_75t_L g1910 ( 
.A(n_1851),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1871),
.B(n_1739),
.Y(n_1911)
);

NOR2xp33_ASAP7_75t_L g1912 ( 
.A(n_1850),
.B(n_1859),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1737),
.B(n_1733),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1791),
.B(n_1805),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1733),
.B(n_1766),
.Y(n_1915)
);

AND2x4_ASAP7_75t_L g1916 ( 
.A(n_1733),
.B(n_1754),
.Y(n_1916)
);

OR2x2_ASAP7_75t_L g1917 ( 
.A(n_1791),
.B(n_1788),
.Y(n_1917)
);

INVx3_ASAP7_75t_L g1918 ( 
.A(n_1720),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1855),
.Y(n_1919)
);

INVxp67_ASAP7_75t_L g1920 ( 
.A(n_1721),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1752),
.B(n_1769),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1822),
.B(n_1740),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1752),
.B(n_1720),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1757),
.B(n_1813),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1777),
.B(n_1819),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1760),
.B(n_1820),
.Y(n_1926)
);

AND2x2_ASAP7_75t_L g1927 ( 
.A(n_1747),
.B(n_1762),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1758),
.B(n_1828),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1862),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1811),
.Y(n_1930)
);

AOI22xp33_ASAP7_75t_L g1931 ( 
.A1(n_1843),
.A2(n_1714),
.B1(n_1736),
.B2(n_1856),
.Y(n_1931)
);

INVxp67_ASAP7_75t_L g1932 ( 
.A(n_1727),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1788),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1794),
.B(n_1748),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1817),
.Y(n_1935)
);

BUFx2_ASAP7_75t_L g1936 ( 
.A(n_1795),
.Y(n_1936)
);

INVxp67_ASAP7_75t_SL g1937 ( 
.A(n_1825),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1730),
.B(n_1749),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1817),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1730),
.B(n_1806),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1810),
.Y(n_1941)
);

AND2x4_ASAP7_75t_L g1942 ( 
.A(n_1799),
.B(n_1722),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1759),
.B(n_1750),
.Y(n_1943)
);

AND2x2_ASAP7_75t_L g1944 ( 
.A(n_1750),
.B(n_1778),
.Y(n_1944)
);

AOI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1860),
.A2(n_1867),
.B1(n_1866),
.B2(n_1840),
.Y(n_1945)
);

AND2x2_ASAP7_75t_L g1946 ( 
.A(n_1809),
.B(n_1803),
.Y(n_1946)
);

INVxp67_ASAP7_75t_L g1947 ( 
.A(n_1816),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1746),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1833),
.B(n_1810),
.Y(n_1949)
);

NOR2xp67_ASAP7_75t_L g1950 ( 
.A(n_1792),
.B(n_1713),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1826),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1815),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1719),
.B(n_1797),
.Y(n_1953)
);

AOI22xp33_ASAP7_75t_L g1954 ( 
.A1(n_1863),
.A2(n_1734),
.B1(n_1716),
.B2(n_1849),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1783),
.B(n_1827),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1849),
.B(n_1798),
.Y(n_1956)
);

NOR2x1_ASAP7_75t_SL g1957 ( 
.A(n_1765),
.B(n_1786),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1797),
.B(n_1725),
.Y(n_1958)
);

INVxp67_ASAP7_75t_SL g1959 ( 
.A(n_1821),
.Y(n_1959)
);

BUFx8_ASAP7_75t_SL g1960 ( 
.A(n_1731),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1798),
.B(n_1768),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1753),
.B(n_1768),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1738),
.B(n_1773),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1773),
.B(n_1718),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1821),
.B(n_1784),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1793),
.B(n_1802),
.Y(n_1966)
);

AOI33xp33_ASAP7_75t_L g1967 ( 
.A1(n_1888),
.A2(n_1903),
.A3(n_1931),
.B1(n_1954),
.B2(n_1945),
.B3(n_1944),
.Y(n_1967)
);

OA21x2_ASAP7_75t_L g1968 ( 
.A1(n_1898),
.A2(n_1802),
.B(n_1776),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1919),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1891),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1919),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1919),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1894),
.B(n_1812),
.Y(n_1973)
);

OAI21x1_ASAP7_75t_L g1974 ( 
.A1(n_1918),
.A2(n_1823),
.B(n_1807),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1891),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1904),
.Y(n_1976)
);

NOR2xp33_ASAP7_75t_L g1977 ( 
.A(n_1932),
.B(n_1790),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1932),
.B(n_1729),
.Y(n_1978)
);

AOI22xp33_ASAP7_75t_L g1979 ( 
.A1(n_1892),
.A2(n_1734),
.B1(n_1716),
.B2(n_1767),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1912),
.B(n_1782),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1916),
.Y(n_1981)
);

AND2x4_ASAP7_75t_L g1982 ( 
.A(n_1916),
.B(n_1873),
.Y(n_1982)
);

OAI22xp5_ASAP7_75t_L g1983 ( 
.A1(n_1877),
.A2(n_1861),
.B1(n_1767),
.B2(n_1772),
.Y(n_1983)
);

OAI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1950),
.A2(n_1861),
.B1(n_1779),
.B2(n_1787),
.C(n_1852),
.Y(n_1984)
);

INVx2_ASAP7_75t_L g1985 ( 
.A(n_1904),
.Y(n_1985)
);

OAI31xp33_ASAP7_75t_L g1986 ( 
.A1(n_1958),
.A2(n_1787),
.A3(n_1801),
.B(n_1800),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1893),
.Y(n_1987)
);

AO21x2_ASAP7_75t_L g1988 ( 
.A1(n_1908),
.A2(n_1801),
.B(n_1800),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1956),
.A2(n_1846),
.B1(n_1814),
.B2(n_1862),
.Y(n_1989)
);

AOI221xp5_ASAP7_75t_L g1990 ( 
.A1(n_1892),
.A2(n_1726),
.B1(n_1796),
.B2(n_1818),
.C(n_1744),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_SL g1991 ( 
.A1(n_1877),
.A2(n_1862),
.B1(n_1771),
.B2(n_1780),
.Y(n_1991)
);

OR2x2_ASAP7_75t_L g1992 ( 
.A(n_1899),
.B(n_1911),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1895),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1950),
.A2(n_1780),
.B1(n_1858),
.B2(n_1824),
.Y(n_1994)
);

AOI211xp5_ASAP7_75t_SL g1995 ( 
.A1(n_1944),
.A2(n_1808),
.B(n_1858),
.C(n_1742),
.Y(n_1995)
);

AND2x4_ASAP7_75t_L g1996 ( 
.A(n_1916),
.B(n_1858),
.Y(n_1996)
);

NAND3xp33_ASAP7_75t_L g1997 ( 
.A(n_1905),
.B(n_1948),
.C(n_1934),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1895),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1894),
.B(n_1742),
.Y(n_1999)
);

AO21x2_ASAP7_75t_L g2000 ( 
.A1(n_1908),
.A2(n_1742),
.B(n_1755),
.Y(n_2000)
);

AOI211x1_ASAP7_75t_L g2001 ( 
.A1(n_1955),
.A2(n_1755),
.B(n_1808),
.C(n_1944),
.Y(n_2001)
);

OAI22xp5_ASAP7_75t_L g2002 ( 
.A1(n_1965),
.A2(n_1755),
.B1(n_1958),
.B2(n_1956),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1894),
.B(n_1755),
.Y(n_2003)
);

INVx3_ASAP7_75t_L g2004 ( 
.A(n_1882),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1896),
.Y(n_2005)
);

AOI21xp5_ASAP7_75t_L g2006 ( 
.A1(n_1906),
.A2(n_1937),
.B(n_1949),
.Y(n_2006)
);

AOI22xp5_ASAP7_75t_L g2007 ( 
.A1(n_1928),
.A2(n_1958),
.B1(n_1964),
.B2(n_1927),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_SL g2008 ( 
.A1(n_1934),
.A2(n_1964),
.B(n_1927),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1878),
.B(n_1876),
.Y(n_2009)
);

NAND3xp33_ASAP7_75t_L g2010 ( 
.A(n_1948),
.B(n_1934),
.C(n_1947),
.Y(n_2010)
);

OAI22xp33_ASAP7_75t_SL g2011 ( 
.A1(n_1947),
.A2(n_1937),
.B1(n_1965),
.B2(n_1963),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1928),
.A2(n_1964),
.B1(n_1927),
.B2(n_1921),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1897),
.B(n_1886),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1928),
.A2(n_1963),
.B1(n_1961),
.B2(n_1955),
.Y(n_2014)
);

AND2x2_ASAP7_75t_L g2015 ( 
.A(n_1878),
.B(n_1876),
.Y(n_2015)
);

INVxp67_ASAP7_75t_SL g2016 ( 
.A(n_1889),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_R g2017 ( 
.A(n_1929),
.B(n_1879),
.Y(n_2017)
);

NOR2x1p5_ASAP7_75t_L g2018 ( 
.A(n_1961),
.B(n_1897),
.Y(n_2018)
);

AOI33xp33_ASAP7_75t_L g2019 ( 
.A1(n_1943),
.A2(n_1921),
.A3(n_1933),
.B1(n_1948),
.B2(n_1953),
.B3(n_1962),
.Y(n_2019)
);

NAND3xp33_ASAP7_75t_L g2020 ( 
.A(n_1943),
.B(n_1949),
.C(n_1921),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_1878),
.B(n_1876),
.Y(n_2021)
);

BUFx3_ASAP7_75t_L g2022 ( 
.A(n_1929),
.Y(n_2022)
);

OAI211xp5_ASAP7_75t_L g2023 ( 
.A1(n_1943),
.A2(n_1933),
.B(n_1953),
.C(n_1962),
.Y(n_2023)
);

AOI221xp5_ASAP7_75t_L g2024 ( 
.A1(n_1924),
.A2(n_1953),
.B1(n_1962),
.B2(n_1926),
.C(n_1946),
.Y(n_2024)
);

CKINVDCx16_ASAP7_75t_R g2025 ( 
.A(n_1910),
.Y(n_2025)
);

AOI221xp5_ASAP7_75t_L g2026 ( 
.A1(n_1924),
.A2(n_1926),
.B1(n_1946),
.B2(n_1938),
.C(n_1939),
.Y(n_2026)
);

OR2x2_ASAP7_75t_L g2027 ( 
.A(n_1899),
.B(n_1911),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1882),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1889),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1900),
.Y(n_2030)
);

AOI221xp5_ASAP7_75t_L g2031 ( 
.A1(n_1924),
.A2(n_1926),
.B1(n_1946),
.B2(n_1938),
.C(n_1935),
.Y(n_2031)
);

OAI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1924),
.A2(n_1938),
.B(n_1939),
.Y(n_2032)
);

AOI221xp5_ASAP7_75t_L g2033 ( 
.A1(n_1924),
.A2(n_1935),
.B1(n_1922),
.B2(n_1936),
.C(n_1952),
.Y(n_2033)
);

NAND3xp33_ASAP7_75t_L g2034 ( 
.A(n_1941),
.B(n_1952),
.C(n_1909),
.Y(n_2034)
);

AOI221xp5_ASAP7_75t_L g2035 ( 
.A1(n_1922),
.A2(n_1936),
.B1(n_1941),
.B2(n_1886),
.C(n_1925),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1920),
.B(n_1887),
.Y(n_2036)
);

INVx2_ASAP7_75t_L g2037 ( 
.A(n_1883),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_2009),
.B(n_1923),
.Y(n_2038)
);

AND2x2_ASAP7_75t_L g2039 ( 
.A(n_2009),
.B(n_1923),
.Y(n_2039)
);

INVx2_ASAP7_75t_L g2040 ( 
.A(n_1976),
.Y(n_2040)
);

BUFx2_ASAP7_75t_L g2041 ( 
.A(n_1981),
.Y(n_2041)
);

HB1xp67_ASAP7_75t_L g2042 ( 
.A(n_2028),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2015),
.B(n_1923),
.Y(n_2043)
);

CKINVDCx16_ASAP7_75t_R g2044 ( 
.A(n_2025),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1976),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1969),
.Y(n_2046)
);

OR2x2_ASAP7_75t_L g2047 ( 
.A(n_1992),
.B(n_1899),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_1992),
.B(n_1911),
.Y(n_2048)
);

NOR2xp33_ASAP7_75t_L g2049 ( 
.A(n_1980),
.B(n_1960),
.Y(n_2049)
);

OR2x2_ASAP7_75t_L g2050 ( 
.A(n_2027),
.B(n_1917),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1969),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1971),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1971),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1972),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_2027),
.B(n_1917),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1972),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1987),
.Y(n_2057)
);

NOR2x1_ASAP7_75t_L g2058 ( 
.A(n_2034),
.B(n_2010),
.Y(n_2058)
);

OR2x2_ASAP7_75t_L g2059 ( 
.A(n_2029),
.B(n_1917),
.Y(n_2059)
);

INVx2_ASAP7_75t_SL g2060 ( 
.A(n_1985),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2016),
.B(n_1880),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_2013),
.B(n_1914),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1987),
.Y(n_2063)
);

BUFx3_ASAP7_75t_L g2064 ( 
.A(n_2022),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2015),
.B(n_1885),
.Y(n_2065)
);

AND2x4_ASAP7_75t_L g2066 ( 
.A(n_1981),
.B(n_1906),
.Y(n_2066)
);

NOR2x1_ASAP7_75t_L g2067 ( 
.A(n_2020),
.B(n_1910),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_1993),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2006),
.B(n_1880),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_2021),
.B(n_1999),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2021),
.B(n_1884),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1999),
.B(n_1884),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1993),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2003),
.B(n_1884),
.Y(n_2074)
);

INVx4_ASAP7_75t_L g2075 ( 
.A(n_2022),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1998),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2036),
.B(n_1920),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_1998),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_2003),
.B(n_1885),
.Y(n_2079)
);

AND2x2_ASAP7_75t_L g2080 ( 
.A(n_1973),
.B(n_1885),
.Y(n_2080)
);

AND2x2_ASAP7_75t_L g2081 ( 
.A(n_1973),
.B(n_1915),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1982),
.B(n_1915),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2004),
.B(n_1907),
.Y(n_2083)
);

AOI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_1997),
.A2(n_1922),
.B1(n_1942),
.B2(n_1940),
.Y(n_2084)
);

AND2x4_ASAP7_75t_L g2085 ( 
.A(n_1996),
.B(n_1906),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1996),
.B(n_1906),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_2004),
.B(n_1907),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2005),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_SL g2089 ( 
.A(n_2011),
.B(n_2019),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_1974),
.B(n_1907),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_2005),
.B(n_1930),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_2030),
.B(n_1930),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2030),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2018),
.B(n_1970),
.Y(n_2094)
);

OR2x2_ASAP7_75t_L g2095 ( 
.A(n_2028),
.B(n_1914),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1975),
.Y(n_2096)
);

AND2x4_ASAP7_75t_SL g2097 ( 
.A(n_2075),
.B(n_1982),
.Y(n_2097)
);

OAI21xp33_ASAP7_75t_L g2098 ( 
.A1(n_2058),
.A2(n_2089),
.B(n_2019),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2058),
.B(n_2035),
.Y(n_2099)
);

NOR2x1_ASAP7_75t_L g2100 ( 
.A(n_2067),
.B(n_2023),
.Y(n_2100)
);

AOI211x1_ASAP7_75t_L g2101 ( 
.A1(n_2094),
.A2(n_1984),
.B(n_2014),
.C(n_2032),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2057),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_2040),
.Y(n_2103)
);

OR2x2_ASAP7_75t_L g2104 ( 
.A(n_2050),
.B(n_2037),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2050),
.B(n_2037),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2094),
.B(n_2008),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2038),
.B(n_1982),
.Y(n_2107)
);

INVx2_ASAP7_75t_SL g2108 ( 
.A(n_2064),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2040),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2077),
.B(n_2033),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2057),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2038),
.B(n_1988),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2063),
.Y(n_2113)
);

NAND2x1p5_ASAP7_75t_L g2114 ( 
.A(n_2067),
.B(n_1906),
.Y(n_2114)
);

AND2x4_ASAP7_75t_L g2115 ( 
.A(n_2085),
.B(n_1974),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_L g2116 ( 
.A(n_2077),
.B(n_2007),
.Y(n_2116)
);

OAI32xp33_ASAP7_75t_L g2117 ( 
.A1(n_2069),
.A2(n_1983),
.A3(n_2012),
.B1(n_1979),
.B2(n_2044),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_2063),
.Y(n_2118)
);

INVx2_ASAP7_75t_SL g2119 ( 
.A(n_2064),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2040),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2038),
.B(n_1988),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_L g2122 ( 
.A(n_2049),
.B(n_2044),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_2045),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2068),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2039),
.B(n_2043),
.Y(n_2125)
);

AND2x2_ASAP7_75t_L g2126 ( 
.A(n_2039),
.B(n_1988),
.Y(n_2126)
);

OR2x2_ASAP7_75t_L g2127 ( 
.A(n_2055),
.B(n_1890),
.Y(n_2127)
);

NAND4xp25_ASAP7_75t_L g2128 ( 
.A(n_2084),
.B(n_1967),
.C(n_2024),
.D(n_2026),
.Y(n_2128)
);

INVx2_ASAP7_75t_SL g2129 ( 
.A(n_2064),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2068),
.Y(n_2130)
);

AND2x4_ASAP7_75t_L g2131 ( 
.A(n_2085),
.B(n_1996),
.Y(n_2131)
);

AND2x2_ASAP7_75t_L g2132 ( 
.A(n_2039),
.B(n_1916),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2043),
.B(n_1916),
.Y(n_2133)
);

NOR2xp33_ASAP7_75t_SL g2134 ( 
.A(n_2075),
.B(n_1986),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_2062),
.B(n_2031),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2073),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2062),
.B(n_1978),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2073),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_2076),
.Y(n_2139)
);

INVxp67_ASAP7_75t_L g2140 ( 
.A(n_2061),
.Y(n_2140)
);

INVxp67_ASAP7_75t_L g2141 ( 
.A(n_2061),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2076),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_2045),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2078),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2078),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2043),
.B(n_1957),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2080),
.B(n_1957),
.Y(n_2147)
);

AOI21xp33_ASAP7_75t_SL g2148 ( 
.A1(n_2069),
.A2(n_1991),
.B(n_1989),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2047),
.B(n_1951),
.Y(n_2149)
);

AOI21xp33_ASAP7_75t_L g2150 ( 
.A1(n_2117),
.A2(n_2090),
.B(n_2002),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2098),
.B(n_2047),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2111),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2110),
.B(n_2081),
.Y(n_2153)
);

NAND3xp33_ASAP7_75t_SL g2154 ( 
.A(n_2099),
.B(n_1967),
.C(n_2017),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2111),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_2116),
.B(n_2081),
.Y(n_2156)
);

AND2x4_ASAP7_75t_L g2157 ( 
.A(n_2131),
.B(n_2085),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2106),
.B(n_2048),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_L g2159 ( 
.A(n_2128),
.B(n_1977),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2135),
.B(n_2048),
.Y(n_2160)
);

AND2x4_ASAP7_75t_L g2161 ( 
.A(n_2131),
.B(n_2085),
.Y(n_2161)
);

NAND2xp33_ASAP7_75t_SL g2162 ( 
.A(n_2100),
.B(n_2075),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2113),
.Y(n_2163)
);

OAI33xp33_ASAP7_75t_L g2164 ( 
.A1(n_2140),
.A2(n_2096),
.A3(n_2059),
.B1(n_2093),
.B2(n_2088),
.B3(n_2092),
.Y(n_2164)
);

NOR3xp33_ASAP7_75t_L g2165 ( 
.A(n_2117),
.B(n_1990),
.C(n_1994),
.Y(n_2165)
);

OR2x2_ASAP7_75t_L g2166 ( 
.A(n_2127),
.B(n_2055),
.Y(n_2166)
);

OR2x2_ASAP7_75t_L g2167 ( 
.A(n_2137),
.B(n_2059),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2101),
.B(n_2070),
.Y(n_2168)
);

OR2x2_ASAP7_75t_L g2169 ( 
.A(n_2141),
.B(n_2095),
.Y(n_2169)
);

INVx2_ASAP7_75t_L g2170 ( 
.A(n_2125),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_2125),
.B(n_2080),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2149),
.B(n_2095),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_2097),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_2103),
.Y(n_2174)
);

OR2x2_ASAP7_75t_L g2175 ( 
.A(n_2127),
.B(n_2070),
.Y(n_2175)
);

BUFx2_ASAP7_75t_L g2176 ( 
.A(n_2108),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2113),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_2118),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2148),
.B(n_2070),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_2146),
.B(n_2080),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2118),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_L g2182 ( 
.A(n_2108),
.B(n_2065),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_2130),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2119),
.B(n_2065),
.Y(n_2184)
);

OR2x2_ASAP7_75t_L g2185 ( 
.A(n_2104),
.B(n_2105),
.Y(n_2185)
);

OAI33xp33_ASAP7_75t_L g2186 ( 
.A1(n_2130),
.A2(n_2142),
.A3(n_2138),
.B1(n_2139),
.B2(n_2145),
.B3(n_2144),
.Y(n_2186)
);

INVxp67_ASAP7_75t_L g2187 ( 
.A(n_2134),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2136),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2146),
.B(n_2147),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2147),
.B(n_2065),
.Y(n_2190)
);

OR2x2_ASAP7_75t_L g2191 ( 
.A(n_2104),
.B(n_1951),
.Y(n_2191)
);

AND2x2_ASAP7_75t_L g2192 ( 
.A(n_2132),
.B(n_2071),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2103),
.Y(n_2193)
);

OR2x2_ASAP7_75t_L g2194 ( 
.A(n_2105),
.B(n_2114),
.Y(n_2194)
);

NOR4xp25_ASAP7_75t_SL g2195 ( 
.A(n_2114),
.B(n_2041),
.C(n_1875),
.D(n_1959),
.Y(n_2195)
);

INVx1_ASAP7_75t_SL g2196 ( 
.A(n_2097),
.Y(n_2196)
);

AND2x2_ASAP7_75t_L g2197 ( 
.A(n_2132),
.B(n_2133),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2136),
.Y(n_2198)
);

OAI211xp5_ASAP7_75t_L g2199 ( 
.A1(n_2112),
.A2(n_2001),
.B(n_1875),
.C(n_1959),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2138),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2139),
.Y(n_2201)
);

AND2x4_ASAP7_75t_L g2202 ( 
.A(n_2131),
.B(n_2086),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2119),
.B(n_2071),
.Y(n_2203)
);

NAND2xp5_ASAP7_75t_L g2204 ( 
.A(n_2159),
.B(n_2129),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_2176),
.Y(n_2205)
);

OAI22xp5_ASAP7_75t_L g2206 ( 
.A1(n_2187),
.A2(n_2114),
.B1(n_2122),
.B2(n_2129),
.Y(n_2206)
);

A2O1A1Ixp33_ASAP7_75t_L g2207 ( 
.A1(n_2165),
.A2(n_1995),
.B(n_2112),
.C(n_2121),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_L g2208 ( 
.A(n_2159),
.B(n_2107),
.Y(n_2208)
);

INVx2_ASAP7_75t_L g2209 ( 
.A(n_2170),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_2178),
.Y(n_2210)
);

AND2x4_ASAP7_75t_L g2211 ( 
.A(n_2157),
.B(n_2107),
.Y(n_2211)
);

INVxp67_ASAP7_75t_L g2212 ( 
.A(n_2154),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2178),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2152),
.Y(n_2214)
);

XNOR2x1_ASAP7_75t_SL g2215 ( 
.A(n_2162),
.B(n_2121),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2157),
.B(n_2133),
.Y(n_2216)
);

AND2x2_ASAP7_75t_L g2217 ( 
.A(n_2157),
.B(n_2082),
.Y(n_2217)
);

NAND4xp25_ASAP7_75t_L g2218 ( 
.A(n_2150),
.B(n_2126),
.C(n_2115),
.D(n_1922),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2155),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2163),
.Y(n_2220)
);

AOI221xp5_ASAP7_75t_L g2221 ( 
.A1(n_2162),
.A2(n_2126),
.B1(n_2115),
.B2(n_2124),
.C(n_2102),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_2168),
.B(n_2072),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2177),
.Y(n_2223)
);

INVx1_ASAP7_75t_SL g2224 ( 
.A(n_2173),
.Y(n_2224)
);

AOI22xp5_ASAP7_75t_L g2225 ( 
.A1(n_2199),
.A2(n_2115),
.B1(n_2086),
.B2(n_2090),
.Y(n_2225)
);

INVxp67_ASAP7_75t_L g2226 ( 
.A(n_2179),
.Y(n_2226)
);

INVx1_ASAP7_75t_L g2227 ( 
.A(n_2181),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_2161),
.B(n_2086),
.Y(n_2228)
);

OAI322xp33_ASAP7_75t_L g2229 ( 
.A1(n_2151),
.A2(n_2145),
.A3(n_2144),
.B1(n_2142),
.B2(n_2143),
.C1(n_2109),
.C2(n_2123),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2183),
.Y(n_2230)
);

OR2x2_ASAP7_75t_L g2231 ( 
.A(n_2158),
.B(n_2090),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2153),
.B(n_2082),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2170),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_2160),
.B(n_2072),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2161),
.B(n_2086),
.Y(n_2235)
);

AOI322xp5_ASAP7_75t_L g2236 ( 
.A1(n_2171),
.A2(n_2071),
.A3(n_2079),
.B1(n_2074),
.B2(n_2072),
.C1(n_1922),
.C2(n_1925),
.Y(n_2236)
);

OAI21xp33_ASAP7_75t_L g2237 ( 
.A1(n_2156),
.A2(n_2090),
.B(n_1925),
.Y(n_2237)
);

OAI21xp5_ASAP7_75t_L g2238 ( 
.A1(n_2196),
.A2(n_2090),
.B(n_2066),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_2164),
.A2(n_1968),
.B1(n_1901),
.B2(n_1902),
.Y(n_2239)
);

OR2x2_ASAP7_75t_L g2240 ( 
.A(n_2167),
.B(n_2090),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_L g2241 ( 
.A(n_2182),
.B(n_2074),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_2161),
.B(n_2074),
.Y(n_2242)
);

NAND2xp5_ASAP7_75t_L g2243 ( 
.A(n_2184),
.B(n_2079),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2211),
.Y(n_2244)
);

OAI32xp33_ASAP7_75t_L g2245 ( 
.A1(n_2212),
.A2(n_2218),
.A3(n_2215),
.B1(n_2226),
.B2(n_2204),
.Y(n_2245)
);

INVx2_ASAP7_75t_SL g2246 ( 
.A(n_2205),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2210),
.Y(n_2247)
);

OAI21xp33_ASAP7_75t_SL g2248 ( 
.A1(n_2215),
.A2(n_2212),
.B(n_2221),
.Y(n_2248)
);

NOR2xp33_ASAP7_75t_L g2249 ( 
.A(n_2224),
.B(n_2202),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2211),
.B(n_2202),
.Y(n_2250)
);

INVx1_ASAP7_75t_L g2251 ( 
.A(n_2213),
.Y(n_2251)
);

OAI22xp5_ASAP7_75t_L g2252 ( 
.A1(n_2207),
.A2(n_2195),
.B1(n_2202),
.B2(n_2203),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_2207),
.A2(n_2194),
.B(n_2200),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_2205),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2226),
.B(n_2186),
.Y(n_2255)
);

AOI222xp33_ASAP7_75t_L g2256 ( 
.A1(n_2237),
.A2(n_2171),
.B1(n_2198),
.B2(n_2201),
.C1(n_2188),
.C2(n_2192),
.Y(n_2256)
);

OAI22xp5_ASAP7_75t_L g2257 ( 
.A1(n_2239),
.A2(n_2175),
.B1(n_2189),
.B2(n_2169),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_2242),
.Y(n_2258)
);

AND2x2_ASAP7_75t_L g2259 ( 
.A(n_2217),
.B(n_2189),
.Y(n_2259)
);

CKINVDCx14_ASAP7_75t_R g2260 ( 
.A(n_2206),
.Y(n_2260)
);

OAI21xp33_ASAP7_75t_L g2261 ( 
.A1(n_2208),
.A2(n_2194),
.B(n_2166),
.Y(n_2261)
);

OAI31xp33_ASAP7_75t_L g2262 ( 
.A1(n_2208),
.A2(n_2066),
.A3(n_2197),
.B(n_2166),
.Y(n_2262)
);

INVx1_ASAP7_75t_L g2263 ( 
.A(n_2214),
.Y(n_2263)
);

INVx3_ASAP7_75t_L g2264 ( 
.A(n_2216),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2222),
.B(n_2192),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2219),
.Y(n_2266)
);

AOI22xp5_ASAP7_75t_SL g2267 ( 
.A1(n_2228),
.A2(n_2075),
.B1(n_2066),
.B2(n_2041),
.Y(n_2267)
);

AOI221xp5_ASAP7_75t_L g2268 ( 
.A1(n_2229),
.A2(n_2193),
.B1(n_2174),
.B2(n_2185),
.C(n_2180),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_SL g2269 ( 
.A(n_2225),
.B(n_2066),
.Y(n_2269)
);

NOR2x1_ASAP7_75t_L g2270 ( 
.A(n_2220),
.B(n_2174),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2228),
.A2(n_1942),
.B1(n_2197),
.B2(n_1913),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_L g2272 ( 
.A(n_2232),
.B(n_2180),
.Y(n_2272)
);

AND2x2_ASAP7_75t_SL g2273 ( 
.A(n_2255),
.B(n_2249),
.Y(n_2273)
);

OAI31xp33_ASAP7_75t_SL g2274 ( 
.A1(n_2252),
.A2(n_2238),
.A3(n_2235),
.B(n_2216),
.Y(n_2274)
);

AOI211xp5_ASAP7_75t_L g2275 ( 
.A1(n_2248),
.A2(n_2227),
.B(n_2223),
.C(n_2230),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_L g2276 ( 
.A(n_2249),
.B(n_2232),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2254),
.Y(n_2277)
);

AND2x2_ASAP7_75t_L g2278 ( 
.A(n_2244),
.B(n_2209),
.Y(n_2278)
);

INVx1_ASAP7_75t_L g2279 ( 
.A(n_2254),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2246),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_L g2281 ( 
.A(n_2246),
.B(n_2209),
.Y(n_2281)
);

OR2x2_ASAP7_75t_L g2282 ( 
.A(n_2265),
.B(n_2234),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2270),
.Y(n_2283)
);

INVx1_ASAP7_75t_L g2284 ( 
.A(n_2263),
.Y(n_2284)
);

OAI211xp5_ASAP7_75t_SL g2285 ( 
.A1(n_2253),
.A2(n_2236),
.B(n_2239),
.C(n_2231),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2266),
.Y(n_2286)
);

OAI22xp5_ASAP7_75t_L g2287 ( 
.A1(n_2260),
.A2(n_2243),
.B1(n_2241),
.B2(n_2240),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2255),
.B(n_2233),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2247),
.Y(n_2289)
);

AOI21x1_ASAP7_75t_L g2290 ( 
.A1(n_2251),
.A2(n_2233),
.B(n_2193),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_2244),
.B(n_2190),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2244),
.Y(n_2292)
);

INVx2_ASAP7_75t_L g2293 ( 
.A(n_2264),
.Y(n_2293)
);

INVx1_ASAP7_75t_L g2294 ( 
.A(n_2264),
.Y(n_2294)
);

CKINVDCx20_ASAP7_75t_R g2295 ( 
.A(n_2260),
.Y(n_2295)
);

AND2x2_ASAP7_75t_L g2296 ( 
.A(n_2273),
.B(n_2250),
.Y(n_2296)
);

NAND4xp25_ASAP7_75t_L g2297 ( 
.A(n_2275),
.B(n_2245),
.C(n_2262),
.D(n_2261),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2278),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2273),
.B(n_2258),
.Y(n_2299)
);

AND3x1_ASAP7_75t_L g2300 ( 
.A(n_2274),
.B(n_2264),
.C(n_2258),
.Y(n_2300)
);

NOR2xp33_ASAP7_75t_L g2301 ( 
.A(n_2295),
.B(n_2269),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_2293),
.Y(n_2302)
);

O2A1O1Ixp33_ASAP7_75t_L g2303 ( 
.A1(n_2288),
.A2(n_2269),
.B(n_2257),
.C(n_2256),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2293),
.B(n_2259),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2295),
.B(n_2272),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2278),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2280),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_L g2308 ( 
.A(n_2288),
.B(n_2268),
.Y(n_2308)
);

NOR3xp33_ASAP7_75t_L g2309 ( 
.A(n_2287),
.B(n_2271),
.C(n_2267),
.Y(n_2309)
);

AOI222xp33_ASAP7_75t_L g2310 ( 
.A1(n_2308),
.A2(n_2285),
.B1(n_2276),
.B2(n_2283),
.C1(n_2289),
.C2(n_2284),
.Y(n_2310)
);

OAI221xp5_ASAP7_75t_L g2311 ( 
.A1(n_2297),
.A2(n_2276),
.B1(n_2294),
.B2(n_2292),
.C(n_2291),
.Y(n_2311)
);

AND2x2_ASAP7_75t_L g2312 ( 
.A(n_2296),
.B(n_2277),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2302),
.Y(n_2313)
);

NOR2xp33_ASAP7_75t_R g2314 ( 
.A(n_2299),
.B(n_2279),
.Y(n_2314)
);

O2A1O1Ixp33_ASAP7_75t_L g2315 ( 
.A1(n_2303),
.A2(n_2305),
.B(n_2301),
.C(n_2307),
.Y(n_2315)
);

HB1xp67_ASAP7_75t_L g2316 ( 
.A(n_2302),
.Y(n_2316)
);

AOI22xp33_ASAP7_75t_L g2317 ( 
.A1(n_2309),
.A2(n_2282),
.B1(n_2286),
.B2(n_2281),
.Y(n_2317)
);

OAI22x1_ASAP7_75t_L g2318 ( 
.A1(n_2301),
.A2(n_2290),
.B1(n_2190),
.B2(n_2120),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2305),
.B(n_2304),
.Y(n_2319)
);

OAI211xp5_ASAP7_75t_SL g2320 ( 
.A1(n_2298),
.A2(n_2172),
.B(n_2109),
.C(n_2143),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2316),
.Y(n_2321)
);

AND2x2_ASAP7_75t_L g2322 ( 
.A(n_2312),
.B(n_2306),
.Y(n_2322)
);

INVx2_ASAP7_75t_L g2323 ( 
.A(n_2313),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_2310),
.B(n_2300),
.Y(n_2324)
);

AOI211xp5_ASAP7_75t_L g2325 ( 
.A1(n_2315),
.A2(n_1908),
.B(n_1913),
.C(n_1929),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2319),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2317),
.B(n_2120),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_2311),
.A2(n_1906),
.B1(n_1968),
.B2(n_1901),
.Y(n_2328)
);

OR2x2_ASAP7_75t_L g2329 ( 
.A(n_2321),
.B(n_2318),
.Y(n_2329)
);

NAND5xp2_ASAP7_75t_L g2330 ( 
.A(n_2324),
.B(n_2315),
.C(n_2314),
.D(n_2320),
.E(n_1966),
.Y(n_2330)
);

AOI21xp5_ASAP7_75t_L g2331 ( 
.A1(n_2324),
.A2(n_2123),
.B(n_2191),
.Y(n_2331)
);

OAI211xp5_ASAP7_75t_L g2332 ( 
.A1(n_2326),
.A2(n_1881),
.B(n_1906),
.C(n_1910),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2322),
.Y(n_2333)
);

AO22x1_ASAP7_75t_L g2334 ( 
.A1(n_2323),
.A2(n_2079),
.B1(n_1881),
.B2(n_2087),
.Y(n_2334)
);

INVx2_ASAP7_75t_L g2335 ( 
.A(n_2327),
.Y(n_2335)
);

XNOR2x2_ASAP7_75t_L g2336 ( 
.A(n_2325),
.B(n_2083),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2329),
.Y(n_2337)
);

NOR3xp33_ASAP7_75t_L g2338 ( 
.A(n_2333),
.B(n_2328),
.C(n_1881),
.Y(n_2338)
);

AOI22xp5_ASAP7_75t_L g2339 ( 
.A1(n_2335),
.A2(n_2083),
.B1(n_2087),
.B2(n_2096),
.Y(n_2339)
);

OAI322xp33_ASAP7_75t_L g2340 ( 
.A1(n_2331),
.A2(n_2060),
.A3(n_2088),
.B1(n_2093),
.B2(n_2052),
.C1(n_2053),
.C2(n_2046),
.Y(n_2340)
);

NOR3xp33_ASAP7_75t_L g2341 ( 
.A(n_2330),
.B(n_1881),
.C(n_1887),
.Y(n_2341)
);

NOR4xp25_ASAP7_75t_L g2342 ( 
.A(n_2332),
.B(n_2330),
.C(n_2336),
.D(n_2334),
.Y(n_2342)
);

AOI211xp5_ASAP7_75t_L g2343 ( 
.A1(n_2342),
.A2(n_2087),
.B(n_2083),
.C(n_1913),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2337),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2341),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2339),
.Y(n_2346)
);

OAI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_2344),
.A2(n_2343),
.B1(n_2345),
.B2(n_2346),
.Y(n_2347)
);

INVx2_ASAP7_75t_L g2348 ( 
.A(n_2344),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2348),
.Y(n_2349)
);

AND2x4_ASAP7_75t_L g2350 ( 
.A(n_2349),
.B(n_2338),
.Y(n_2350)
);

NAND3xp33_ASAP7_75t_L g2351 ( 
.A(n_2349),
.B(n_2347),
.C(n_2340),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2351),
.Y(n_2352)
);

OR2x6_ASAP7_75t_L g2353 ( 
.A(n_2350),
.B(n_1881),
.Y(n_2353)
);

AOI22xp33_ASAP7_75t_L g2354 ( 
.A1(n_2352),
.A2(n_2000),
.B1(n_2060),
.B2(n_2052),
.Y(n_2354)
);

AOI322xp5_ASAP7_75t_L g2355 ( 
.A1(n_2354),
.A2(n_2353),
.A3(n_2060),
.B1(n_2042),
.B2(n_2051),
.C1(n_2046),
.C2(n_2053),
.Y(n_2355)
);

AOI221xp5_ASAP7_75t_L g2356 ( 
.A1(n_2355),
.A2(n_2051),
.B1(n_2042),
.B2(n_2056),
.C(n_2054),
.Y(n_2356)
);

AOI211xp5_ASAP7_75t_L g2357 ( 
.A1(n_2356),
.A2(n_2092),
.B(n_2091),
.C(n_2054),
.Y(n_2357)
);


endmodule