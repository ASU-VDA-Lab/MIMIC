module real_jpeg_30684_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_47;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_0),
.B(n_1),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx2_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

AOI222xp33_ASAP7_75t_SL g36 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_43),
.C1(n_44),
.C2(n_47),
.Y(n_36)
);

AND2x4_ASAP7_75t_SL g11 ( 
.A(n_4),
.B(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_4),
.B(n_16),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_4),
.B(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g15 ( 
.A1(n_6),
.A2(n_7),
.B1(n_16),
.B2(n_17),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

OAI221xp5_ASAP7_75t_L g8 ( 
.A1(n_9),
.A2(n_21),
.B1(n_26),
.B2(n_32),
.C(n_36),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_10),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_20),
.Y(n_10)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OA22x2_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_15),
.B1(n_18),
.B2(n_19),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_31),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_31),
.Y(n_46)
);

OR2x2_ASAP7_75t_L g40 ( 
.A(n_18),
.B(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_19),
.B(n_31),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_25),
.Y(n_22)
);

AND2x4_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_35),
.Y(n_37)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_30),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

AND2x4_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);


endmodule