module fake_jpeg_22534_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_37),
.B(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

CKINVDCx11_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_40),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_30),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_46),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_17),
.B(n_9),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_21),
.A2(n_31),
.B1(n_25),
.B2(n_24),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_31),
.B1(n_21),
.B2(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_25),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_59),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_62),
.A2(n_45),
.B1(n_18),
.B2(n_28),
.Y(n_106)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_70),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_31),
.B1(n_25),
.B2(n_21),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_36),
.B1(n_28),
.B2(n_18),
.Y(n_83)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

AO22x1_ASAP7_75t_SL g71 ( 
.A1(n_47),
.A2(n_24),
.B1(n_23),
.B2(n_29),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_71),
.A2(n_37),
.B1(n_45),
.B2(n_24),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_53),
.A2(n_43),
.B(n_47),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_89),
.B(n_30),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_77),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_47),
.C(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_80),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_79),
.B(n_50),
.Y(n_114)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_81),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_96),
.B1(n_100),
.B2(n_106),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_84),
.B(n_85),
.Y(n_127)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_53),
.B(n_46),
.Y(n_86)
);

BUFx24_ASAP7_75t_SL g124 ( 
.A(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_55),
.B(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_87),
.B(n_42),
.Y(n_125)
);

AND2x4_ASAP7_75t_SL g89 ( 
.A(n_64),
.B(n_24),
.Y(n_89)
);

INVx4_ASAP7_75t_SL g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_97),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_58),
.B(n_43),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_98),
.Y(n_134)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_93),
.B(n_94),
.Y(n_130)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_51),
.A2(n_27),
.B1(n_18),
.B2(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_101),
.Y(n_116)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_42),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_132),
.Y(n_159)
);

OA22x2_ASAP7_75t_SL g109 ( 
.A1(n_81),
.A2(n_38),
.B1(n_41),
.B2(n_48),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_135),
.B1(n_93),
.B2(n_100),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_112),
.A2(n_123),
.B(n_17),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_122),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_72),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_119),
.B(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_69),
.B(n_30),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_129),
.Y(n_167)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_48),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_78),
.A2(n_37),
.B1(n_45),
.B2(n_59),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_118),
.B(n_77),
.C(n_88),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_151),
.C(n_155),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_149),
.B1(n_150),
.B2(n_156),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_114),
.B(n_44),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_139),
.B(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_142),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_131),
.A2(n_84),
.B1(n_89),
.B2(n_76),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_141),
.A2(n_148),
.B1(n_161),
.B2(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

AND2x4_ASAP7_75t_SL g146 ( 
.A(n_112),
.B(n_76),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_146),
.A2(n_121),
.B(n_115),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_131),
.A2(n_45),
.B1(n_105),
.B2(n_70),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_95),
.B1(n_68),
.B2(n_97),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_111),
.A2(n_95),
.B1(n_102),
.B2(n_99),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_99),
.C(n_75),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_116),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_162),
.Y(n_187)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_154),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_48),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_44),
.B1(n_36),
.B2(n_28),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_116),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_158),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_125),
.B(n_122),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_109),
.A2(n_90),
.B1(n_91),
.B2(n_17),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_166),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_85),
.B1(n_80),
.B2(n_26),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_48),
.C(n_41),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_109),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_41),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_168),
.B(n_169),
.Y(n_223)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_163),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_108),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_170),
.B(n_184),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_171),
.B(n_172),
.Y(n_232)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

INVxp67_ASAP7_75t_SL g211 ( 
.A(n_174),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_183),
.C(n_155),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_189),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_170),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_108),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_124),
.B1(n_119),
.B2(n_128),
.C(n_121),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_198),
.B(n_160),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_141),
.A2(n_115),
.B1(n_132),
.B2(n_107),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_196),
.B1(n_200),
.B2(n_126),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_138),
.A2(n_110),
.B1(n_107),
.B2(n_120),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_192),
.A2(n_144),
.B1(n_142),
.B2(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_23),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_154),
.Y(n_195)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_195),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_153),
.A2(n_110),
.B1(n_26),
.B2(n_19),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_197),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_159),
.A2(n_120),
.B(n_26),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_162),
.A2(n_110),
.B1(n_38),
.B2(n_41),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_201),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_203),
.A2(n_209),
.B1(n_215),
.B2(n_228),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_219),
.C(n_220),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_207),
.A2(n_217),
.B(n_231),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_222),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_172),
.A2(n_151),
.B1(n_143),
.B2(n_147),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_181),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_221),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_192),
.A2(n_158),
.B1(n_145),
.B2(n_126),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_185),
.A2(n_126),
.B(n_34),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_174),
.B1(n_178),
.B2(n_194),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_183),
.C(n_189),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_103),
.C(n_29),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_35),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_35),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_198),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_227),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_180),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_226),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_179),
.A2(n_34),
.B1(n_27),
.B2(n_23),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_187),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_229),
.B(n_230),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

OA21x2_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_29),
.B(n_20),
.Y(n_231)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_223),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_236),
.Y(n_265)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_249),
.B1(n_227),
.B2(n_212),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_210),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_247),
.B(n_251),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_171),
.B1(n_193),
.B2(n_169),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_241),
.A2(n_243),
.B1(n_224),
.B2(n_202),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_188),
.B1(n_200),
.B2(n_187),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_245),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_182),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_211),
.A2(n_178),
.B1(n_168),
.B2(n_191),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_215),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_208),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_250),
.C(n_256),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_207),
.A2(n_195),
.B1(n_2),
.B2(n_3),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_29),
.C(n_20),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_218),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_20),
.C(n_35),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_206),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_258),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_259),
.B(n_260),
.Y(n_286)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_252),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_214),
.B(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_SL g294 ( 
.A(n_262),
.B(n_10),
.C(n_16),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_270),
.B1(n_273),
.B2(n_234),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_231),
.Y(n_269)
);

OAI22x1_ASAP7_75t_L g290 ( 
.A1(n_269),
.A2(n_279),
.B1(n_259),
.B2(n_273),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_205),
.B1(n_231),
.B2(n_216),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_237),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_272),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_249),
.A2(n_216),
.B1(n_2),
.B2(n_3),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_20),
.C(n_35),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_277),
.C(n_256),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_243),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_245),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_20),
.C(n_35),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_278),
.A2(n_255),
.B(n_250),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_244),
.B(n_1),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_280),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_265),
.B(n_238),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_281),
.B(n_284),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_291),
.C(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_290),
.B(n_278),
.Y(n_300)
);

BUFx12_ASAP7_75t_L g284 ( 
.A(n_262),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_248),
.C(n_234),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_295),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_255),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_288),
.A2(n_268),
.B1(n_266),
.B2(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_33),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_267),
.B(n_10),
.Y(n_293)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_294),
.A2(n_290),
.B(n_292),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_263),
.B(n_279),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_261),
.B(n_33),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_10),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_298),
.B(n_13),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_300),
.A2(n_305),
.B(n_310),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_261),
.C(n_277),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_301),
.C(n_300),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_304),
.B(n_308),
.Y(n_320)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_284),
.B(n_286),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_309),
.B(n_312),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_284),
.A2(n_269),
.B(n_279),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_291),
.B(n_269),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_305),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_314),
.B(n_322),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_307),
.A2(n_302),
.B(n_306),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_315),
.A2(n_324),
.B(n_311),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_299),
.A2(n_295),
.B1(n_285),
.B2(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_8),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_310),
.B(n_11),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_318),
.C(n_321),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_11),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_303),
.B(n_1),
.C(n_3),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_326),
.B(n_328),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_313),
.B(n_4),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_327),
.A2(n_330),
.B(n_9),
.Y(n_335)
);

AOI221xp5_ASAP7_75t_L g328 ( 
.A1(n_323),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.C(n_7),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g329 ( 
.A1(n_317),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_329),
.B(n_324),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_7),
.B(n_8),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_334),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_320),
.B(n_33),
.Y(n_334)
);

NAND3xp33_ASAP7_75t_L g343 ( 
.A(n_335),
.B(n_337),
.C(n_341),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_333),
.A2(n_321),
.B(n_325),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_336),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_318),
.Y(n_340)
);

A2O1A1O1Ixp25_ASAP7_75t_L g344 ( 
.A1(n_340),
.A2(n_12),
.B(n_13),
.C(n_14),
.D(n_15),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_333),
.B(n_12),
.Y(n_341)
);

OAI21xp33_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_339),
.B(n_16),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_345),
.Y(n_346)
);

AOI321xp33_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_342),
.A3(n_343),
.B1(n_338),
.B2(n_12),
.C(n_33),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_33),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_33),
.Y(n_349)
);


endmodule