module fake_jpeg_15342_n_156 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_156);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_156;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_25),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_14),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_25),
.B1(n_15),
.B2(n_28),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_15),
.B1(n_26),
.B2(n_21),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_0),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_26),
.B(n_21),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_25),
.B1(n_15),
.B2(n_28),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_48),
.A2(n_32),
.B1(n_24),
.B2(n_18),
.Y(n_64)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_18),
.C(n_20),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_59),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_51),
.A2(n_64),
.B1(n_65),
.B2(n_17),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_56),
.Y(n_75)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_20),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_43),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_67),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_61),
.B(n_14),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_16),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_63),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_27),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_43),
.A2(n_24),
.B1(n_27),
.B2(n_22),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_37),
.C(n_31),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_31),
.C(n_29),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_22),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_17),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_74),
.Y(n_91)
);

XNOR2x2_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_17),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_83),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_80),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_60),
.Y(n_81)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_58),
.B1(n_51),
.B2(n_53),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_97),
.Y(n_106)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_95),
.Y(n_110)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_57),
.B1(n_68),
.B2(n_67),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_98),
.B(n_100),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_43),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_79),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_72),
.A2(n_29),
.B1(n_6),
.B2(n_7),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_76),
.A3(n_75),
.B1(n_87),
.B2(n_83),
.C1(n_86),
.C2(n_78),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_72),
.C(n_70),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_113),
.C(n_114),
.Y(n_124)
);

AO21x1_ASAP7_75t_L g125 ( 
.A1(n_107),
.A2(n_99),
.B(n_95),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_80),
.C(n_73),
.Y(n_108)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_115),
.C(n_3),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_117),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_91),
.A2(n_86),
.B(n_84),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_111),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_93),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_85),
.C(n_6),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_85),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g115 ( 
.A(n_103),
.B(n_0),
.C(n_2),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_2),
.B(n_3),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_101),
.Y(n_121)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_125),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_123),
.B(n_127),
.Y(n_134)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_126),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_116),
.B(n_92),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_128),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_120),
.A2(n_106),
.B1(n_110),
.B2(n_113),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_119),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_124),
.A2(n_111),
.B1(n_117),
.B2(n_97),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_124),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_138),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_125),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_135),
.A2(n_128),
.B(n_115),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_141),
.A2(n_136),
.B(n_130),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_9),
.C(n_10),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_142),
.B(n_129),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_4),
.Y(n_151)
);

AOI322xp5_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_131),
.A3(n_134),
.B1(n_10),
.B2(n_11),
.C1(n_5),
.C2(n_3),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_142),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_150),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_137),
.B(n_11),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_148),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_145),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_152),
.C(n_147),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_5),
.Y(n_156)
);


endmodule