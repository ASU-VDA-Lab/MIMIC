module fake_ariane_2658_n_1802 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1802);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1802;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_784;
wire n_648;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_51),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_10),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_115),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_152),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_39),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_48),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_24),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_44),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_106),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_84),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_5),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_42),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_130),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_113),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_134),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_149),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_36),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_52),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_47),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_119),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_8),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g188 ( 
.A(n_11),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_101),
.Y(n_189)
);

BUFx8_ASAP7_75t_SL g190 ( 
.A(n_28),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_158),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_99),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_60),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_151),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_124),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_62),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_36),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_57),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_20),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g202 ( 
.A(n_74),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_51),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_137),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_45),
.Y(n_208)
);

INVxp67_ASAP7_75t_SL g209 ( 
.A(n_29),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_121),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_107),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_148),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_79),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_13),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_90),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_114),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_17),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_66),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_45),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_159),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_52),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_132),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_26),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_59),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_93),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_72),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_92),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_73),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_2),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_41),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_87),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_75),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_164),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_68),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_70),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g236 ( 
.A(n_50),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_129),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_15),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_54),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_146),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_82),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_7),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_31),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_85),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_42),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_156),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_120),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_102),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_150),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_29),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_13),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

BUFx10_ASAP7_75t_L g253 ( 
.A(n_49),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_53),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_19),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_91),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_154),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_143),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_20),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_21),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_77),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_104),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_83),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_117),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_103),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_131),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_96),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_100),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_4),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_88),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_55),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_98),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_37),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_71),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_53),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_118),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_140),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_89),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_19),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_21),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_163),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_126),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_24),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_26),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_65),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_2),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_76),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_9),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_105),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_8),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_23),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_54),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_139),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_50),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g297 ( 
.A(n_80),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_16),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_9),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_44),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_128),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_6),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_17),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_28),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_123),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_48),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_142),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_147),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_95),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_4),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_27),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_34),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_81),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_144),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_27),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_136),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_0),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_31),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_40),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_46),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_46),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_125),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_78),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_64),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_162),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_38),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_245),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_190),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_229),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_1),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_192),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_165),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_320),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_250),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_245),
.B(n_1),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_220),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_225),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_228),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_231),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_245),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_257),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_261),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_245),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_326),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_203),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_252),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_219),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_240),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_320),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_245),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_167),
.B(n_3),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_171),
.B(n_3),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_173),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_184),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_221),
.Y(n_359)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_184),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_223),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_184),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_184),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_168),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_184),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_185),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_201),
.Y(n_367)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_238),
.B(n_5),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_239),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_207),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_242),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_189),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_243),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_254),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_185),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_185),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_236),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_259),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_185),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_269),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_169),
.B(n_193),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_271),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_230),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_273),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_185),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_312),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_255),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_236),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_312),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

NAND2xp33_ASAP7_75t_R g391 ( 
.A(n_170),
.B(n_176),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_189),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_276),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_236),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_281),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_200),
.B(n_7),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_172),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_285),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_168),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_172),
.B(n_11),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_208),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_287),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_R g405 ( 
.A(n_179),
.B(n_56),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_401),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_335),
.B(n_208),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_342),
.Y(n_408)
);

OAI21x1_ASAP7_75t_L g409 ( 
.A1(n_339),
.A2(n_182),
.B(n_218),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_206),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_401),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_342),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_381),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_372),
.B(n_251),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_342),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_331),
.B(n_251),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_334),
.A2(n_289),
.B1(n_322),
.B2(n_321),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_328),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_249),
.Y(n_420)
);

AND2x4_ASAP7_75t_L g421 ( 
.A(n_360),
.B(n_260),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_342),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_332),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_342),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_224),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_332),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_336),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_336),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_338),
.Y(n_429)
);

BUFx8_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_338),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_344),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_347),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_347),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_354),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_354),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_358),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_358),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_362),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_399),
.B(n_260),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_L g443 ( 
.A(n_355),
.B(n_202),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_399),
.B(n_280),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_363),
.Y(n_445)
);

INVx5_ASAP7_75t_L g446 ( 
.A(n_405),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_363),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_365),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_365),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_403),
.B(n_280),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_350),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_366),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_366),
.B(n_232),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_403),
.B(n_352),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_404),
.B(n_249),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_352),
.B(n_293),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_398),
.B(n_182),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_376),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_376),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_379),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_379),
.B(n_241),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_385),
.B(n_389),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_385),
.A2(n_258),
.B(n_256),
.Y(n_465)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_389),
.A2(n_264),
.B(n_263),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_357),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_390),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_392),
.B(n_293),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_393),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_393),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_377),
.B(n_298),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_349),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_402),
.B(n_266),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_402),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_368),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_368),
.Y(n_479)
);

NOR2x1p5_ASAP7_75t_L g480 ( 
.A(n_475),
.B(n_330),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_475),
.B(n_351),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_432),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_429),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_359),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_L g485 ( 
.A(n_418),
.B(n_209),
.C(n_188),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_432),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_475),
.B(n_361),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_415),
.B(n_364),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_429),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_429),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_415),
.B(n_388),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_432),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_456),
.B(n_414),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_427),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_475),
.B(n_369),
.Y(n_495)
);

BUFx6f_ASAP7_75t_SL g496 ( 
.A(n_475),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_429),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_435),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

NOR2x1p5_ASAP7_75t_L g500 ( 
.A(n_454),
.B(n_337),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_435),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_435),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_454),
.B(n_371),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_427),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_454),
.B(n_373),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_457),
.Y(n_506)
);

INVx3_ASAP7_75t_L g507 ( 
.A(n_432),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_414),
.B(n_374),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_430),
.Y(n_509)
);

BUFx10_ASAP7_75t_L g510 ( 
.A(n_411),
.Y(n_510)
);

BUFx6f_ASAP7_75t_SL g511 ( 
.A(n_417),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_411),
.B(n_378),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_457),
.B(n_380),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

OAI22xp33_ASAP7_75t_L g515 ( 
.A1(n_418),
.A2(n_391),
.B1(n_396),
.B2(n_166),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_478),
.B(n_382),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_438),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_459),
.A2(n_298),
.B1(n_356),
.B2(n_284),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_459),
.A2(n_214),
.B1(n_217),
.B2(n_316),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_469),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_478),
.B(n_479),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_415),
.B(n_384),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_430),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_457),
.B(n_395),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_478),
.B(n_397),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_407),
.B(n_400),
.Y(n_526)
);

BUFx4f_ASAP7_75t_L g527 ( 
.A(n_427),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_438),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_407),
.B(n_253),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_417),
.A2(n_303),
.B1(n_294),
.B2(n_199),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_425),
.B(n_345),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_469),
.Y(n_532)
);

AND2x6_ASAP7_75t_L g533 ( 
.A(n_417),
.B(n_262),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_410),
.B(n_268),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_469),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_410),
.B(n_319),
.C(n_275),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_438),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_474),
.B(n_170),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_479),
.B(n_175),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_407),
.B(n_186),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_419),
.B(n_233),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_438),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_410),
.Y(n_543)
);

NAND3xp33_ASAP7_75t_L g544 ( 
.A(n_431),
.B(n_278),
.C(n_270),
.Y(n_544)
);

AOI22xp33_ASAP7_75t_L g545 ( 
.A1(n_417),
.A2(n_253),
.B1(n_204),
.B2(n_248),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_417),
.A2(n_253),
.B1(n_204),
.B2(n_292),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_452),
.Y(n_547)
);

BUFx4f_ASAP7_75t_L g548 ( 
.A(n_427),
.Y(n_548)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_446),
.B(n_176),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_451),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_432),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_474),
.B(n_446),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_417),
.A2(n_204),
.B1(n_327),
.B2(n_296),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_474),
.B(n_383),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_425),
.B(n_333),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_419),
.B(n_423),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_431),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_451),
.B(n_174),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_431),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_476),
.A2(n_299),
.B1(n_291),
.B2(n_178),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_446),
.B(n_180),
.Y(n_561)
);

AOI22xp33_ASAP7_75t_L g562 ( 
.A1(n_476),
.A2(n_302),
.B1(n_304),
.B2(n_174),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_427),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_467),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_433),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_427),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_433),
.B(n_290),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_452),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_433),
.Y(n_570)
);

BUFx3_ASAP7_75t_L g571 ( 
.A(n_434),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_477),
.A2(n_310),
.B1(n_177),
.B2(n_178),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_477),
.B(n_262),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_406),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_423),
.B(n_180),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_452),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_434),
.Y(n_577)
);

OR2x6_ASAP7_75t_L g578 ( 
.A(n_442),
.B(n_274),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_413),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_434),
.B(n_295),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_426),
.B(n_314),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_452),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_462),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_427),
.Y(n_584)
);

CKINVDCx16_ASAP7_75t_R g585 ( 
.A(n_467),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_426),
.B(n_181),
.Y(n_586)
);

INVx5_ASAP7_75t_L g587 ( 
.A(n_413),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_439),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_406),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_462),
.Y(n_590)
);

NOR2x1p5_ASAP7_75t_L g591 ( 
.A(n_412),
.B(n_177),
.Y(n_591)
);

BUFx10_ASAP7_75t_L g592 ( 
.A(n_421),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_439),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_421),
.B(n_274),
.Y(n_594)
);

INVx6_ASAP7_75t_L g595 ( 
.A(n_430),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_446),
.B(n_181),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_421),
.A2(n_315),
.B1(n_302),
.B2(n_187),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_462),
.Y(n_598)
);

INVxp33_ASAP7_75t_L g599 ( 
.A(n_412),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_455),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_462),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_441),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_441),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_421),
.A2(n_300),
.B1(n_304),
.B2(n_187),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_428),
.B(n_317),
.C(n_325),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_446),
.B(n_191),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_442),
.B(n_444),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_445),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_446),
.B(n_191),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_446),
.B(n_246),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_421),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_455),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_473),
.Y(n_613)
);

BUFx3_ASAP7_75t_L g614 ( 
.A(n_428),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_473),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_473),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_473),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_413),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_436),
.B(n_246),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_436),
.B(n_340),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_430),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_442),
.B(n_183),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_430),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_437),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_437),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_430),
.A2(n_183),
.B1(n_306),
.B2(n_310),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_445),
.Y(n_627)
);

BUFx8_ASAP7_75t_SL g628 ( 
.A(n_444),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_444),
.B(n_300),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_455),
.Y(n_630)
);

BUFx6f_ASAP7_75t_SL g631 ( 
.A(n_550),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_588),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_L g633 ( 
.A(n_494),
.B(n_446),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_493),
.B(n_420),
.Y(n_634)
);

INVx4_ASAP7_75t_L g635 ( 
.A(n_511),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_588),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_512),
.B(n_446),
.Y(n_637)
);

NAND2x1_ASAP7_75t_L g638 ( 
.A(n_595),
.B(n_424),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_508),
.B(n_420),
.Y(n_639)
);

NAND2xp33_ASAP7_75t_L g640 ( 
.A(n_494),
.B(n_301),
.Y(n_640)
);

AOI22xp5_ASAP7_75t_L g641 ( 
.A1(n_524),
.A2(n_531),
.B1(n_526),
.B2(n_506),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_484),
.B(n_540),
.Y(n_642)
);

O2A1O1Ixp5_ASAP7_75t_L g643 ( 
.A1(n_527),
.A2(n_453),
.B(n_463),
.C(n_447),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_510),
.B(n_443),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_529),
.B(n_470),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_529),
.B(n_470),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_510),
.B(n_443),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_510),
.B(n_301),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_483),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_510),
.B(n_305),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_550),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_526),
.B(n_470),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_506),
.B(n_450),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_483),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_497),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_541),
.B(n_521),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_607),
.B(n_450),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_607),
.B(n_450),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g659 ( 
.A(n_516),
.B(n_453),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_497),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_554),
.B(n_341),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_515),
.B(n_305),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_626),
.B(n_323),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_624),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_555),
.A2(n_308),
.B1(n_307),
.B2(n_309),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_525),
.B(n_463),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_514),
.B(n_307),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_513),
.B(n_306),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_514),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_611),
.B(n_455),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_611),
.B(n_409),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_554),
.Y(n_672)
);

NAND2xp33_ASAP7_75t_L g673 ( 
.A(n_494),
.B(n_308),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_482),
.B(n_409),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_624),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_574),
.B(n_343),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_625),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_539),
.B(n_409),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_625),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_482),
.B(n_486),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_522),
.B(n_447),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_574),
.B(n_346),
.Y(n_682)
);

OR2x6_ASAP7_75t_L g683 ( 
.A(n_578),
.B(n_348),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_517),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_600),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_517),
.Y(n_686)
);

AND2x4_ASAP7_75t_SL g687 ( 
.A(n_514),
.B(n_592),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_496),
.B(n_311),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_522),
.B(n_449),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_593),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_600),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_528),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_528),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_514),
.B(n_309),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_482),
.B(n_449),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_537),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_486),
.B(n_460),
.Y(n_697)
);

OAI21xp5_ASAP7_75t_L g698 ( 
.A1(n_543),
.A2(n_466),
.B(n_465),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_486),
.B(n_460),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_492),
.B(n_461),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_592),
.B(n_313),
.Y(n_701)
);

OAI21xp5_ASAP7_75t_L g702 ( 
.A1(n_543),
.A2(n_559),
.B(n_557),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_557),
.A2(n_461),
.B(n_464),
.C(n_324),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_593),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_589),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_492),
.B(n_313),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_494),
.B(n_311),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_492),
.B(n_465),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_507),
.B(n_465),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_600),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_589),
.B(n_367),
.Y(n_711)
);

OR2x6_ASAP7_75t_L g712 ( 
.A(n_578),
.B(n_466),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_507),
.B(n_464),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_L g714 ( 
.A(n_494),
.B(n_315),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_507),
.B(n_318),
.Y(n_715)
);

INVx8_ASAP7_75t_L g716 ( 
.A(n_594),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_551),
.B(n_318),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_551),
.B(n_491),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_L g719 ( 
.A1(n_599),
.A2(n_321),
.B1(n_322),
.B2(n_329),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_500),
.Y(n_720)
);

NOR2xp67_ASAP7_75t_L g721 ( 
.A(n_620),
.B(n_472),
.Y(n_721)
);

INVx3_ASAP7_75t_L g722 ( 
.A(n_592),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_551),
.B(n_491),
.Y(n_723)
);

BUFx6f_ASAP7_75t_L g724 ( 
.A(n_600),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_571),
.B(n_194),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_592),
.B(n_195),
.Y(n_726)
);

OAI22xp5_ASAP7_75t_L g727 ( 
.A1(n_571),
.A2(n_197),
.B1(n_196),
.B2(n_198),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_602),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_537),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_503),
.B(n_12),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_500),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_480),
.B(n_370),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_542),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_542),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_571),
.B(n_205),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_481),
.B(n_487),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_603),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_594),
.B(n_210),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_547),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_495),
.B(n_211),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_505),
.B(n_14),
.Y(n_741)
);

NOR2x1p5_ASAP7_75t_L g742 ( 
.A(n_558),
.B(n_387),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_565),
.B(n_14),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_594),
.B(n_212),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_594),
.A2(n_297),
.B1(n_466),
.B2(n_468),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_547),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_569),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_556),
.A2(n_408),
.B(n_422),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_L g749 ( 
.A1(n_527),
.A2(n_424),
.B(n_408),
.C(n_422),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_553),
.B(n_213),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_629),
.B(n_215),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_538),
.B(n_15),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_569),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_594),
.B(n_216),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_603),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_608),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_504),
.B(n_440),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_511),
.B(n_18),
.Y(n_758)
);

INVx8_ASAP7_75t_L g759 ( 
.A(n_594),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_629),
.B(n_222),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_488),
.B(n_18),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_608),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_594),
.B(n_226),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_558),
.B(n_597),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_485),
.A2(n_297),
.B1(n_23),
.B2(n_25),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_614),
.B(n_227),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_614),
.B(n_244),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_614),
.B(n_237),
.Y(n_768)
);

INVx8_ASAP7_75t_L g769 ( 
.A(n_533),
.Y(n_769)
);

OAI22xp33_ASAP7_75t_L g770 ( 
.A1(n_578),
.A2(n_283),
.B1(n_267),
.B2(n_272),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_600),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_604),
.B(n_288),
.Y(n_772)
);

A2O1A1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_559),
.A2(n_424),
.B(n_422),
.C(n_408),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_511),
.B(n_552),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_576),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_SL g776 ( 
.A(n_565),
.B(n_234),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_573),
.B(n_286),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_575),
.B(n_22),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_627),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_585),
.Y(n_780)
);

INVx2_ASAP7_75t_SL g781 ( 
.A(n_488),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_SL g782 ( 
.A(n_496),
.B(n_480),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_627),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_622),
.B(n_22),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_520),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_586),
.B(n_25),
.Y(n_786)
);

INVx2_ASAP7_75t_SL g787 ( 
.A(n_591),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_573),
.B(n_235),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_576),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_573),
.B(n_247),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_573),
.B(n_265),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_504),
.B(n_440),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_533),
.B(n_619),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_533),
.B(n_277),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_520),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_612),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_622),
.B(n_30),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_578),
.B(n_30),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_533),
.B(n_279),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_582),
.Y(n_800)
);

BUFx3_ASAP7_75t_L g801 ( 
.A(n_612),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_634),
.B(n_533),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_641),
.B(n_612),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_643),
.A2(n_577),
.B(n_570),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_642),
.B(n_585),
.Y(n_805)
);

AOI22xp33_ASAP7_75t_L g806 ( 
.A1(n_663),
.A2(n_533),
.B1(n_578),
.B2(n_591),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_674),
.A2(n_548),
.B(n_527),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_632),
.Y(n_808)
);

AOI21x1_ASAP7_75t_L g809 ( 
.A1(n_708),
.A2(n_566),
.B(n_570),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_634),
.A2(n_577),
.B1(n_566),
.B2(n_496),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_711),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_663),
.A2(n_764),
.B1(n_672),
.B2(n_797),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_661),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_639),
.B(n_659),
.Y(n_814)
);

BUFx6f_ASAP7_75t_L g815 ( 
.A(n_685),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_674),
.A2(n_501),
.B(n_490),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_716),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_639),
.B(n_533),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_659),
.B(n_545),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_708),
.A2(n_709),
.B(n_680),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_SL g821 ( 
.A(n_780),
.B(n_628),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_636),
.Y(n_822)
);

A2O1A1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_797),
.A2(n_581),
.B(n_568),
.C(n_534),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_666),
.B(n_546),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_666),
.A2(n_581),
.B(n_568),
.C(n_534),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_676),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_SL g827 ( 
.A(n_665),
.B(n_562),
.C(n_560),
.Y(n_827)
);

OAI22xp5_ASAP7_75t_L g828 ( 
.A1(n_785),
.A2(n_535),
.B1(n_532),
.B2(n_580),
.Y(n_828)
);

OR2x6_ASAP7_75t_L g829 ( 
.A(n_683),
.B(n_623),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_656),
.B(n_518),
.Y(n_830)
);

AOI21x1_ASAP7_75t_L g831 ( 
.A1(n_709),
.A2(n_535),
.B(n_532),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_651),
.B(n_572),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_718),
.B(n_530),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_702),
.A2(n_548),
.B(n_567),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_649),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_778),
.A2(n_580),
.B(n_489),
.C(n_490),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_798),
.A2(n_519),
.B1(n_612),
.B2(n_630),
.Y(n_837)
);

BUFx2_ASAP7_75t_L g838 ( 
.A(n_682),
.Y(n_838)
);

OAI22xp5_ASAP7_75t_L g839 ( 
.A1(n_795),
.A2(n_501),
.B1(n_489),
.B2(n_498),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_631),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_649),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_781),
.Y(n_842)
);

NAND2x1p5_ASAP7_75t_L g843 ( 
.A(n_635),
.B(n_612),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_723),
.B(n_498),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_645),
.B(n_499),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_690),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_646),
.B(n_499),
.Y(n_847)
);

NAND2x1_ASAP7_75t_L g848 ( 
.A(n_654),
.B(n_502),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_704),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_705),
.B(n_623),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_631),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_637),
.A2(n_548),
.B(n_567),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_654),
.Y(n_853)
);

INVx4_ASAP7_75t_L g854 ( 
.A(n_716),
.Y(n_854)
);

AOI22xp5_ASAP7_75t_L g855 ( 
.A1(n_798),
.A2(n_630),
.B1(n_536),
.B2(n_605),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_680),
.A2(n_502),
.B(n_584),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_761),
.B(n_536),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_757),
.A2(n_609),
.B(n_561),
.Y(n_858)
);

BUFx4f_ASAP7_75t_L g859 ( 
.A(n_683),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_655),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_678),
.A2(n_584),
.B(n_564),
.Y(n_861)
);

AOI21xp5_ASAP7_75t_L g862 ( 
.A1(n_713),
.A2(n_584),
.B(n_564),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_757),
.A2(n_792),
.B(n_697),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_635),
.B(n_509),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_657),
.B(n_658),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_728),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_792),
.A2(n_567),
.B(n_564),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_685),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_695),
.A2(n_606),
.B(n_596),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_655),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_749),
.A2(n_583),
.B(n_590),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_699),
.A2(n_610),
.B(n_549),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_700),
.A2(n_563),
.B(n_504),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_652),
.B(n_582),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_683),
.B(n_583),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_751),
.B(n_760),
.Y(n_876)
);

INVx11_ASAP7_75t_L g877 ( 
.A(n_776),
.Y(n_877)
);

AOI21xp33_ASAP7_75t_L g878 ( 
.A1(n_668),
.A2(n_621),
.B(n_523),
.Y(n_878)
);

A2O1A1Ixp33_ASAP7_75t_L g879 ( 
.A1(n_778),
.A2(n_786),
.B(n_752),
.C(n_730),
.Y(n_879)
);

AOI33xp33_ASAP7_75t_L g880 ( 
.A1(n_784),
.A2(n_590),
.A3(n_598),
.B1(n_601),
.B2(n_613),
.B3(n_615),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_660),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_687),
.B(n_563),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_698),
.A2(n_598),
.B(n_617),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_668),
.B(n_504),
.Y(n_884)
);

OAI21xp33_ASAP7_75t_L g885 ( 
.A1(n_786),
.A2(n_605),
.B(n_544),
.Y(n_885)
);

INVx3_ASAP7_75t_L g886 ( 
.A(n_687),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_685),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_720),
.B(n_601),
.Y(n_888)
);

BUFx10_ASAP7_75t_L g889 ( 
.A(n_732),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_681),
.B(n_613),
.Y(n_890)
);

NOR2x1p5_ASAP7_75t_L g891 ( 
.A(n_732),
.B(n_544),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_743),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_689),
.B(n_617),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_653),
.B(n_616),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_662),
.B(n_504),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_737),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_755),
.B(n_616),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_787),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_748),
.A2(n_563),
.B(n_615),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_660),
.Y(n_900)
);

OR2x2_ASAP7_75t_L g901 ( 
.A(n_742),
.B(n_32),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_756),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_762),
.B(n_563),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_779),
.B(n_563),
.Y(n_904)
);

NOR2xp67_ASAP7_75t_SL g905 ( 
.A(n_669),
.B(n_595),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_716),
.Y(n_906)
);

OAI21xp5_ASAP7_75t_L g907 ( 
.A1(n_671),
.A2(n_579),
.B(n_587),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_731),
.B(n_587),
.Y(n_908)
);

AOI33xp33_ASAP7_75t_L g909 ( 
.A1(n_719),
.A2(n_32),
.A3(n_33),
.B1(n_34),
.B2(n_35),
.B3(n_37),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_752),
.A2(n_424),
.B(n_440),
.C(n_448),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_644),
.A2(n_618),
.B(n_587),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_644),
.A2(n_618),
.B(n_587),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_783),
.B(n_595),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_664),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_647),
.A2(n_618),
.B(n_587),
.Y(n_915)
);

NAND2x1p5_ASAP7_75t_L g916 ( 
.A(n_669),
.B(n_618),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_730),
.A2(n_424),
.B(n_440),
.C(n_448),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_793),
.A2(n_579),
.B(n_587),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_670),
.B(n_595),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_647),
.A2(n_618),
.B(n_579),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_741),
.B(n_648),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_736),
.A2(n_618),
.B(n_579),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_664),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_725),
.A2(n_579),
.B(n_422),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_722),
.B(n_579),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_741),
.A2(n_282),
.B1(n_471),
.B2(n_468),
.Y(n_926)
);

BUFx4f_ASAP7_75t_L g927 ( 
.A(n_759),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_SL g928 ( 
.A(n_759),
.B(n_440),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_722),
.B(n_33),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_735),
.A2(n_408),
.B(n_413),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_766),
.A2(n_413),
.B(n_416),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_767),
.A2(n_413),
.B(n_416),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_715),
.B(n_35),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_758),
.Y(n_934)
);

AOI22xp33_ASAP7_75t_L g935 ( 
.A1(n_765),
.A2(n_440),
.B1(n_471),
.B2(n_468),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_770),
.B(n_440),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_773),
.A2(n_472),
.B(n_471),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_768),
.A2(n_413),
.B(n_416),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_675),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_759),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_717),
.B(n_38),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_675),
.B(n_39),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_706),
.A2(n_413),
.B(n_416),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_677),
.B(n_40),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_650),
.B(n_41),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_758),
.B(n_448),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_782),
.B(n_448),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_684),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_688),
.B(n_448),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_677),
.A2(n_679),
.B(n_800),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_684),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_679),
.A2(n_416),
.B(n_471),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_765),
.A2(n_448),
.B1(n_471),
.B2(n_468),
.Y(n_953)
);

INVx6_ASAP7_75t_L g954 ( 
.A(n_685),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_777),
.B(n_43),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_788),
.B(n_448),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_686),
.A2(n_416),
.B(n_471),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_790),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_692),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_692),
.A2(n_416),
.B(n_471),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_693),
.A2(n_416),
.B(n_471),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_791),
.B(n_43),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_772),
.B(n_47),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_693),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_712),
.A2(n_468),
.B(n_458),
.Y(n_965)
);

INVx3_ASAP7_75t_L g966 ( 
.A(n_769),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_750),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_696),
.B(n_49),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_696),
.B(n_55),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_769),
.B(n_468),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_769),
.A2(n_468),
.B1(n_458),
.B2(n_448),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_729),
.A2(n_468),
.B(n_458),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_729),
.B(n_733),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_724),
.B(n_796),
.Y(n_974)
);

INVx4_ASAP7_75t_L g975 ( 
.A(n_724),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_733),
.A2(n_746),
.B(n_800),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_734),
.A2(n_458),
.B(n_440),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_734),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_703),
.A2(n_458),
.B(n_228),
.C(n_472),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_739),
.A2(n_228),
.B(n_458),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_746),
.A2(n_228),
.B(n_458),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_747),
.A2(n_228),
.B(n_472),
.C(n_202),
.Y(n_982)
);

AND2x2_ASAP7_75t_SL g983 ( 
.A(n_745),
.B(n_202),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_747),
.B(n_202),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_765),
.B(n_472),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_753),
.B(n_202),
.Y(n_986)
);

BUFx12f_ASAP7_75t_L g987 ( 
.A(n_712),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_753),
.B(n_202),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_667),
.B(n_472),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_775),
.A2(n_472),
.B(n_202),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_827),
.A2(n_774),
.B1(n_701),
.B2(n_694),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_814),
.B(n_789),
.Y(n_992)
);

INVx3_ASAP7_75t_L g993 ( 
.A(n_817),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_879),
.A2(n_745),
.B1(n_712),
.B2(n_726),
.Y(n_994)
);

AOI22xp5_ASAP7_75t_L g995 ( 
.A1(n_805),
.A2(n_921),
.B1(n_824),
.B2(n_832),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_865),
.B(n_775),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_808),
.Y(n_997)
);

AND2x2_ASAP7_75t_SL g998 ( 
.A(n_859),
.B(n_774),
.Y(n_998)
);

INVx2_ASAP7_75t_SL g999 ( 
.A(n_877),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_825),
.B(n_819),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_874),
.B(n_789),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_934),
.B(n_721),
.Y(n_1002)
);

CKINVDCx6p67_ASAP7_75t_R g1003 ( 
.A(n_889),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_815),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_845),
.B(n_724),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_847),
.B(n_796),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_830),
.B(n_796),
.Y(n_1007)
);

AO22x1_ASAP7_75t_L g1008 ( 
.A1(n_840),
.A2(n_738),
.B1(n_744),
.B2(n_763),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_822),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_846),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_802),
.B(n_796),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_R g1012 ( 
.A(n_821),
.B(n_710),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_849),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_806),
.B(n_801),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_SL g1015 ( 
.A(n_859),
.B(n_889),
.Y(n_1015)
);

A2O1A1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_945),
.A2(n_740),
.B(n_691),
.C(n_710),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_958),
.B(n_727),
.Y(n_1017)
);

A2O1A1Ixp33_ASAP7_75t_L g1018 ( 
.A1(n_885),
.A2(n_801),
.B(n_691),
.C(n_771),
.Y(n_1018)
);

OAI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_909),
.A2(n_707),
.B(n_714),
.Y(n_1019)
);

OAI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_818),
.A2(n_754),
.B(n_794),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_810),
.A2(n_673),
.B(n_640),
.Y(n_1021)
);

BUFx2_ASAP7_75t_L g1022 ( 
.A(n_811),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_807),
.A2(n_633),
.B(n_771),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_SL g1024 ( 
.A1(n_804),
.A2(n_799),
.B(n_638),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_838),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_813),
.A2(n_202),
.B1(n_472),
.B2(n_63),
.Y(n_1026)
);

INVx4_ASAP7_75t_L g1027 ( 
.A(n_886),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_823),
.A2(n_58),
.B1(n_61),
.B2(n_67),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_812),
.B(n_69),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_866),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_820),
.A2(n_86),
.B(n_94),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_826),
.B(n_967),
.Y(n_1032)
);

INVx4_ASAP7_75t_L g1033 ( 
.A(n_886),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_983),
.A2(n_97),
.B1(n_109),
.B2(n_110),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_892),
.B(n_111),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_890),
.B(n_112),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_807),
.A2(n_116),
.B(n_122),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_820),
.A2(n_127),
.B(n_133),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_891),
.B(n_138),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_852),
.A2(n_141),
.B(n_145),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_955),
.A2(n_160),
.B(n_962),
.C(n_941),
.Y(n_1041)
);

INVx2_ASAP7_75t_SL g1042 ( 
.A(n_851),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_896),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_911),
.A2(n_912),
.B(n_834),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_857),
.B(n_902),
.Y(n_1045)
);

OAI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_863),
.A2(n_861),
.B(n_862),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_875),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_911),
.A2(n_912),
.B(n_828),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_L g1049 ( 
.A(n_876),
.B(n_842),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_933),
.A2(n_963),
.B(n_836),
.C(n_803),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_835),
.Y(n_1051)
);

CKINVDCx11_ASAP7_75t_R g1052 ( 
.A(n_898),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_893),
.B(n_844),
.Y(n_1053)
);

AO32x1_ASAP7_75t_L g1054 ( 
.A1(n_985),
.A2(n_839),
.A3(n_914),
.B1(n_939),
.B2(n_923),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_L g1055 ( 
.A(n_815),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_841),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_829),
.B(n_901),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_853),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_888),
.B(n_829),
.Y(n_1059)
);

INVx5_ASAP7_75t_L g1060 ( 
.A(n_970),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_SL g1061 ( 
.A(n_864),
.B(n_878),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_833),
.B(n_894),
.Y(n_1062)
);

AOI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_864),
.A2(n_884),
.B1(n_953),
.B2(n_888),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_861),
.A2(n_907),
.B(n_920),
.Y(n_1064)
);

CKINVDCx6p67_ASAP7_75t_R g1065 ( 
.A(n_829),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_915),
.A2(n_873),
.B(n_883),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_860),
.Y(n_1067)
);

CKINVDCx11_ASAP7_75t_R g1068 ( 
.A(n_987),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_873),
.A2(n_862),
.B(n_863),
.Y(n_1069)
);

NAND3xp33_ASAP7_75t_SL g1070 ( 
.A(n_935),
.B(n_855),
.C(n_929),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_908),
.B(n_959),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_978),
.B(n_870),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_942),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_895),
.A2(n_880),
.B(n_913),
.C(n_837),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_944),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_908),
.B(n_817),
.Y(n_1076)
);

HB1xp67_ASAP7_75t_L g1077 ( 
.A(n_968),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_881),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_927),
.B(n_815),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_900),
.B(n_948),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_951),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_897),
.B(n_964),
.Y(n_1082)
);

INVx4_ASAP7_75t_L g1083 ( 
.A(n_927),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_854),
.B(n_940),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_868),
.B(n_887),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_973),
.B(n_850),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_969),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_954),
.Y(n_1088)
);

BUFx4f_ASAP7_75t_L g1089 ( 
.A(n_868),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_899),
.A2(n_816),
.B(n_872),
.Y(n_1090)
);

OAI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_856),
.A2(n_903),
.B(n_904),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_848),
.Y(n_1092)
);

O2A1O1Ixp5_ASAP7_75t_L g1093 ( 
.A1(n_949),
.A2(n_956),
.B(n_882),
.C(n_943),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_899),
.A2(n_872),
.B(n_943),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_946),
.B(n_917),
.C(n_910),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_868),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_887),
.B(n_954),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_970),
.A2(n_954),
.B1(n_919),
.B2(n_940),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_871),
.A2(n_867),
.B(n_869),
.Y(n_1099)
);

BUFx4f_ASAP7_75t_L g1100 ( 
.A(n_887),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_843),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_975),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_950),
.B(n_975),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_950),
.B(n_976),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_843),
.Y(n_1105)
);

NOR3xp33_ASAP7_75t_SL g1106 ( 
.A(n_856),
.B(n_867),
.C(n_947),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_854),
.Y(n_1107)
);

INVx1_ASAP7_75t_SL g1108 ( 
.A(n_974),
.Y(n_1108)
);

A2O1A1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_869),
.A2(n_989),
.B(n_979),
.C(n_922),
.Y(n_1109)
);

NOR2xp67_ASAP7_75t_L g1110 ( 
.A(n_926),
.B(n_906),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_809),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_906),
.B(n_966),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_966),
.B(n_916),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_990),
.A2(n_972),
.B(n_977),
.C(n_936),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_916),
.B(n_905),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_R g1116 ( 
.A(n_928),
.B(n_965),
.Y(n_1116)
);

O2A1O1Ixp5_ASAP7_75t_L g1117 ( 
.A1(n_931),
.A2(n_938),
.B(n_932),
.C(n_924),
.Y(n_1117)
);

CKINVDCx20_ASAP7_75t_R g1118 ( 
.A(n_970),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_925),
.B(n_918),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_984),
.B(n_988),
.Y(n_1120)
);

INVxp67_ASAP7_75t_SL g1121 ( 
.A(n_971),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_986),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_858),
.Y(n_1123)
);

CKINVDCx20_ASAP7_75t_R g1124 ( 
.A(n_937),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_952),
.A2(n_957),
.B(n_960),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_990),
.B(n_977),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_L g1127 ( 
.A1(n_952),
.A2(n_980),
.B1(n_981),
.B2(n_960),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_SL g1128 ( 
.A(n_957),
.B(n_961),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_982),
.A2(n_814),
.B1(n_879),
.B2(n_865),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_930),
.B(n_814),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_814),
.A2(n_802),
.B(n_825),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_814),
.A2(n_802),
.B(n_825),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_808),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_817),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_808),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_809),
.A2(n_831),
.B(n_883),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_808),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_835),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_814),
.B(n_634),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_814),
.B(n_345),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_814),
.A2(n_802),
.B(n_825),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_814),
.B(n_634),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_814),
.B(n_634),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1044),
.A2(n_1136),
.B(n_1094),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1089),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1139),
.B(n_1143),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1140),
.A2(n_1143),
.B(n_1129),
.C(n_1050),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1048),
.A2(n_1132),
.B(n_1131),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_997),
.Y(n_1149)
);

AOI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_995),
.A2(n_1049),
.B1(n_1124),
.B2(n_1032),
.Y(n_1150)
);

OAI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_1141),
.A2(n_1121),
.B(n_1000),
.Y(n_1151)
);

AO32x2_ASAP7_75t_L g1152 ( 
.A1(n_1129),
.A2(n_994),
.A3(n_1028),
.B1(n_1034),
.B2(n_1098),
.Y(n_1152)
);

OAI22xp33_ASAP7_75t_L g1153 ( 
.A1(n_1017),
.A2(n_1045),
.B1(n_994),
.B2(n_1022),
.Y(n_1153)
);

BUFx3_ASAP7_75t_L g1154 ( 
.A(n_1052),
.Y(n_1154)
);

AND2x4_ASAP7_75t_L g1155 ( 
.A(n_1083),
.B(n_1076),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1047),
.B(n_1025),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_999),
.B(n_1027),
.Y(n_1157)
);

NAND2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1012),
.B(n_1083),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1125),
.A2(n_1111),
.A3(n_1064),
.B(n_1126),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_1000),
.A2(n_1041),
.B(n_991),
.C(n_1070),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1074),
.A2(n_1011),
.B(n_992),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1011),
.A2(n_992),
.B(n_1053),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_998),
.B(n_1009),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1028),
.A2(n_1029),
.B(n_1019),
.C(n_1034),
.Y(n_1164)
);

AND2x2_ASAP7_75t_SL g1165 ( 
.A(n_1015),
.B(n_1039),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1010),
.B(n_1013),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_1089),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_1031),
.A2(n_1038),
.B(n_1109),
.C(n_1053),
.Y(n_1168)
);

AO21x2_ASAP7_75t_L g1169 ( 
.A1(n_1066),
.A2(n_1046),
.B(n_1069),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1003),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1076),
.B(n_1084),
.Y(n_1171)
);

OAI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1063),
.A2(n_1026),
.B1(n_1118),
.B2(n_1030),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1114),
.A2(n_1090),
.A3(n_1099),
.B(n_1104),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1005),
.A2(n_1006),
.B(n_1095),
.Y(n_1174)
);

OR2x2_ASAP7_75t_L g1175 ( 
.A(n_1043),
.B(n_1133),
.Y(n_1175)
);

AO22x1_ASAP7_75t_L g1176 ( 
.A1(n_1059),
.A2(n_1057),
.B1(n_1035),
.B2(n_1033),
.Y(n_1176)
);

AOI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1128),
.A2(n_1008),
.B(n_1021),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1027),
.B(n_1033),
.Y(n_1178)
);

BUFx10_ASAP7_75t_L g1179 ( 
.A(n_1042),
.Y(n_1179)
);

BUFx10_ASAP7_75t_L g1180 ( 
.A(n_1004),
.Y(n_1180)
);

OR2x6_ASAP7_75t_L g1181 ( 
.A(n_1061),
.B(n_1071),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1135),
.B(n_1137),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_1072),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_SL g1184 ( 
.A1(n_1062),
.A2(n_996),
.B(n_1098),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1130),
.A2(n_1119),
.B(n_1036),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1130),
.A2(n_1036),
.B(n_1006),
.Y(n_1186)
);

OA22x2_ASAP7_75t_L g1187 ( 
.A1(n_1077),
.A2(n_1075),
.B1(n_1087),
.B2(n_1073),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1051),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_996),
.A2(n_1062),
.B1(n_1005),
.B2(n_1016),
.C(n_1007),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_1068),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_1007),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1080),
.B(n_1065),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1023),
.A2(n_1091),
.B(n_1117),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1056),
.Y(n_1194)
);

AO21x2_ASAP7_75t_L g1195 ( 
.A1(n_1020),
.A2(n_1024),
.B(n_1116),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1018),
.A2(n_1093),
.B(n_1106),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1088),
.B(n_1102),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1110),
.A2(n_1086),
.B(n_1002),
.C(n_1122),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1103),
.A2(n_1115),
.B(n_1120),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1001),
.B(n_1138),
.Y(n_1200)
);

NOR2x1_ASAP7_75t_R g1201 ( 
.A(n_1060),
.B(n_1096),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1127),
.A2(n_1040),
.B(n_1037),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_SL g1203 ( 
.A1(n_1115),
.A2(n_1113),
.B(n_1112),
.C(n_1079),
.Y(n_1203)
);

BUFx6f_ASAP7_75t_L g1204 ( 
.A(n_1100),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1001),
.B(n_1067),
.Y(n_1205)
);

AOI221xp5_ASAP7_75t_L g1206 ( 
.A1(n_1014),
.A2(n_1082),
.B1(n_1108),
.B2(n_1120),
.C(n_1072),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1058),
.B(n_1078),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1054),
.A2(n_1081),
.A3(n_1092),
.B(n_1123),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1112),
.A2(n_1113),
.B(n_1100),
.Y(n_1209)
);

BUFx12f_ASAP7_75t_L g1210 ( 
.A(n_1004),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_993),
.A2(n_1107),
.B(n_1134),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1060),
.A2(n_1123),
.B(n_1054),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_993),
.A2(n_1107),
.B(n_1134),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1123),
.A2(n_1054),
.B(n_1060),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1097),
.B(n_1004),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1101),
.A2(n_1084),
.B(n_1060),
.C(n_1105),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_1105),
.A2(n_1055),
.B(n_1096),
.C(n_1085),
.Y(n_1217)
);

AOI221x1_ASAP7_75t_L g1218 ( 
.A1(n_1105),
.A2(n_879),
.B1(n_1028),
.B2(n_1034),
.C(n_994),
.Y(n_1218)
);

INVx1_ASAP7_75t_SL g1219 ( 
.A(n_1055),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1055),
.B(n_1096),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1044),
.A2(n_1136),
.B(n_1094),
.Y(n_1221)
);

INVx2_ASAP7_75t_SL g1222 ( 
.A(n_999),
.Y(n_1222)
);

NAND3xp33_ASAP7_75t_L g1223 ( 
.A(n_1140),
.B(n_879),
.C(n_814),
.Y(n_1223)
);

CKINVDCx8_ASAP7_75t_R g1224 ( 
.A(n_1025),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1048),
.A2(n_814),
.B(n_879),
.Y(n_1225)
);

AO21x2_ASAP7_75t_L g1226 ( 
.A1(n_1064),
.A2(n_1094),
.B(n_1044),
.Y(n_1226)
);

INVx5_ASAP7_75t_L g1227 ( 
.A(n_1060),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1140),
.A2(n_661),
.B1(n_565),
.B2(n_663),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1052),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1044),
.A2(n_1136),
.B(n_1094),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1140),
.B(n_661),
.Y(n_1231)
);

INVx1_ASAP7_75t_SL g1232 ( 
.A(n_1052),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1044),
.A2(n_1136),
.B(n_1094),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_997),
.Y(n_1234)
);

AOI211x1_ASAP7_75t_L g1235 ( 
.A1(n_1139),
.A2(n_827),
.B(n_1143),
.C(n_1142),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_995),
.A2(n_879),
.B(n_814),
.Y(n_1236)
);

INVxp67_ASAP7_75t_SL g1237 ( 
.A(n_1118),
.Y(n_1237)
);

AO31x2_ASAP7_75t_L g1238 ( 
.A1(n_1125),
.A2(n_1111),
.A3(n_1064),
.B(n_1126),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1125),
.A2(n_1111),
.A3(n_1064),
.B(n_1126),
.Y(n_1239)
);

O2A1O1Ixp33_ASAP7_75t_L g1240 ( 
.A1(n_1140),
.A2(n_814),
.B(n_879),
.C(n_512),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1125),
.A2(n_1111),
.A3(n_1064),
.B(n_1126),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_1052),
.Y(n_1242)
);

AO31x2_ASAP7_75t_L g1243 ( 
.A1(n_1125),
.A2(n_1111),
.A3(n_1064),
.B(n_1126),
.Y(n_1243)
);

AOI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1128),
.A2(n_1044),
.B(n_1066),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1048),
.A2(n_814),
.B(n_879),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1089),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1142),
.B(n_814),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_995),
.A2(n_814),
.B1(n_879),
.B2(n_1139),
.Y(n_1248)
);

AOI221x1_ASAP7_75t_L g1249 ( 
.A1(n_1028),
.A2(n_879),
.B1(n_1034),
.B2(n_994),
.C(n_765),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1142),
.B(n_814),
.Y(n_1250)
);

OAI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_995),
.A2(n_814),
.B1(n_879),
.B2(n_1139),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1048),
.A2(n_814),
.B(n_879),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1089),
.Y(n_1253)
);

BUFx3_ASAP7_75t_L g1254 ( 
.A(n_1052),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_997),
.Y(n_1255)
);

AO21x1_ASAP7_75t_L g1256 ( 
.A1(n_1034),
.A2(n_994),
.B(n_1050),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_SL g1257 ( 
.A1(n_1139),
.A2(n_879),
.B(n_814),
.C(n_1143),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_997),
.Y(n_1258)
);

AOI221x1_ASAP7_75t_L g1259 ( 
.A1(n_1028),
.A2(n_879),
.B1(n_1034),
.B2(n_994),
.C(n_765),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_997),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_997),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_SL g1262 ( 
.A(n_995),
.B(n_814),
.Y(n_1262)
);

INVx4_ASAP7_75t_SL g1263 ( 
.A(n_999),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_995),
.A2(n_814),
.B1(n_879),
.B2(n_1139),
.Y(n_1264)
);

INVx3_ASAP7_75t_L g1265 ( 
.A(n_1083),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1044),
.A2(n_1136),
.B(n_1094),
.Y(n_1266)
);

OAI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_995),
.A2(n_879),
.B(n_814),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1142),
.B(n_814),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1048),
.A2(n_814),
.B(n_879),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_SL g1270 ( 
.A1(n_1139),
.A2(n_879),
.B(n_814),
.C(n_1143),
.Y(n_1270)
);

BUFx4f_ASAP7_75t_SL g1271 ( 
.A(n_1003),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1048),
.A2(n_814),
.B(n_879),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1140),
.B(n_879),
.C(n_814),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1140),
.B(n_585),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1052),
.Y(n_1275)
);

AOI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_1048),
.A2(n_814),
.B(n_879),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1125),
.A2(n_1111),
.A3(n_1064),
.B(n_1126),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1140),
.B(n_585),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1048),
.A2(n_814),
.B(n_879),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_L g1280 ( 
.A1(n_995),
.A2(n_879),
.B(n_814),
.C(n_921),
.Y(n_1280)
);

INVx3_ASAP7_75t_SL g1281 ( 
.A(n_1003),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1083),
.B(n_1076),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_995),
.A2(n_879),
.B(n_814),
.C(n_921),
.Y(n_1283)
);

NAND3x1_ASAP7_75t_L g1284 ( 
.A(n_995),
.B(n_1140),
.C(n_909),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1052),
.Y(n_1285)
);

BUFx6f_ASAP7_75t_L g1286 ( 
.A(n_1089),
.Y(n_1286)
);

INVxp67_ASAP7_75t_L g1287 ( 
.A(n_1025),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_L g1288 ( 
.A(n_1140),
.B(n_585),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1044),
.A2(n_1136),
.B(n_1094),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1142),
.B(n_814),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_995),
.A2(n_879),
.B(n_814),
.C(n_921),
.Y(n_1291)
);

AOI21x1_ASAP7_75t_SL g1292 ( 
.A1(n_1139),
.A2(n_814),
.B(n_933),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_995),
.A2(n_879),
.B(n_814),
.C(n_921),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_997),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1025),
.Y(n_1295)
);

AO22x2_ASAP7_75t_L g1296 ( 
.A1(n_994),
.A2(n_1034),
.B1(n_1070),
.B2(n_565),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1275),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1231),
.A2(n_1228),
.B1(n_1256),
.B2(n_1296),
.Y(n_1298)
);

BUFx12f_ASAP7_75t_L g1299 ( 
.A(n_1190),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1224),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_SL g1301 ( 
.A1(n_1296),
.A2(n_1165),
.B1(n_1267),
.B2(n_1236),
.Y(n_1301)
);

BUFx8_ASAP7_75t_L g1302 ( 
.A(n_1154),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1175),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1150),
.B(n_1237),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1166),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1249),
.A2(n_1259),
.B1(n_1273),
.B2(n_1223),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1182),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1271),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1172),
.A2(n_1153),
.B1(n_1187),
.B2(n_1274),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1149),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_1229),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1145),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1264),
.A2(n_1278),
.B1(n_1288),
.B2(n_1152),
.Y(n_1314)
);

OAI21xp33_ASAP7_75t_L g1315 ( 
.A1(n_1280),
.A2(n_1283),
.B(n_1293),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1262),
.A2(n_1181),
.B1(n_1206),
.B2(n_1188),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1145),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1234),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_SL g1319 ( 
.A1(n_1152),
.A2(n_1163),
.B1(n_1284),
.B2(n_1151),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1254),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1255),
.Y(n_1321)
);

CKINVDCx6p67_ASAP7_75t_R g1322 ( 
.A(n_1281),
.Y(n_1322)
);

BUFx6f_ASAP7_75t_SL g1323 ( 
.A(n_1167),
.Y(n_1323)
);

CKINVDCx11_ASAP7_75t_R g1324 ( 
.A(n_1232),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1291),
.A2(n_1240),
.B1(n_1147),
.B2(n_1146),
.Y(n_1325)
);

INVx3_ASAP7_75t_L g1326 ( 
.A(n_1167),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_L g1327 ( 
.A1(n_1181),
.A2(n_1247),
.B1(n_1290),
.B2(n_1268),
.Y(n_1327)
);

CKINVDCx11_ASAP7_75t_R g1328 ( 
.A(n_1242),
.Y(n_1328)
);

CKINVDCx20_ASAP7_75t_R g1329 ( 
.A(n_1285),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1258),
.Y(n_1330)
);

BUFx8_ASAP7_75t_SL g1331 ( 
.A(n_1210),
.Y(n_1331)
);

CKINVDCx16_ASAP7_75t_R g1332 ( 
.A(n_1158),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1260),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1183),
.B(n_1162),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1204),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1225),
.A2(n_1252),
.B1(n_1272),
.B2(n_1245),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1261),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1152),
.A2(n_1161),
.B1(n_1250),
.B2(n_1218),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1171),
.B(n_1155),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1156),
.A2(n_1287),
.B1(n_1192),
.B2(n_1222),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1294),
.Y(n_1341)
);

CKINVDCx11_ASAP7_75t_R g1342 ( 
.A(n_1179),
.Y(n_1342)
);

BUFx4_ASAP7_75t_SL g1343 ( 
.A(n_1263),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1207),
.Y(n_1344)
);

NAND2x1p5_ASAP7_75t_L g1345 ( 
.A(n_1171),
.B(n_1155),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_SL g1346 ( 
.A1(n_1183),
.A2(n_1196),
.B1(n_1276),
.B2(n_1279),
.Y(n_1346)
);

OAI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1204),
.A2(n_1246),
.B1(n_1286),
.B2(n_1253),
.Y(n_1347)
);

OAI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1246),
.A2(n_1253),
.B1(n_1286),
.B2(n_1170),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1200),
.A2(n_1205),
.B1(n_1189),
.B2(n_1191),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1246),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1174),
.A2(n_1199),
.B1(n_1269),
.B2(n_1282),
.Y(n_1351)
);

BUFx10_ASAP7_75t_L g1352 ( 
.A(n_1197),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_L g1353 ( 
.A1(n_1195),
.A2(n_1212),
.B1(n_1186),
.B2(n_1286),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_1201),
.Y(n_1354)
);

BUFx8_ASAP7_75t_SL g1355 ( 
.A(n_1253),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1195),
.A2(n_1215),
.B1(n_1209),
.B2(n_1214),
.Y(n_1356)
);

CKINVDCx11_ASAP7_75t_R g1357 ( 
.A(n_1179),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1184),
.B(n_1270),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1185),
.A2(n_1157),
.B1(n_1219),
.B2(n_1263),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1235),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1265),
.A2(n_1178),
.B1(n_1220),
.B2(n_1164),
.Y(n_1361)
);

BUFx2_ASAP7_75t_SL g1362 ( 
.A(n_1265),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1176),
.A2(n_1169),
.B1(n_1148),
.B2(n_1180),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_SL g1364 ( 
.A1(n_1168),
.A2(n_1160),
.B(n_1177),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1169),
.A2(n_1180),
.B1(n_1202),
.B2(n_1198),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1208),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1226),
.A2(n_1257),
.B1(n_1193),
.B2(n_1213),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1226),
.A2(n_1211),
.B1(n_1292),
.B2(n_1144),
.Y(n_1368)
);

OAI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1203),
.A2(n_1244),
.B1(n_1216),
.B2(n_1217),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1221),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1173),
.A2(n_1159),
.B1(n_1277),
.B2(n_1243),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1173),
.A2(n_1159),
.B1(n_1277),
.B2(n_1243),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1230),
.A2(n_1289),
.B1(n_1266),
.B2(n_1233),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1238),
.A2(n_1239),
.B1(n_1241),
.B2(n_1243),
.Y(n_1374)
);

INVx8_ASAP7_75t_L g1375 ( 
.A(n_1239),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1173),
.A2(n_1239),
.B1(n_1241),
.B2(n_1277),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1175),
.Y(n_1377)
);

INVx8_ASAP7_75t_L g1378 ( 
.A(n_1210),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1231),
.B(n_1150),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1275),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1175),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1280),
.A2(n_814),
.B1(n_1291),
.B2(n_1283),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1145),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1385)
);

BUFx2_ASAP7_75t_SL g1386 ( 
.A(n_1224),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1175),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_1145),
.Y(n_1388)
);

NAND2x1p5_ASAP7_75t_L g1389 ( 
.A(n_1227),
.B(n_1060),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1179),
.Y(n_1390)
);

INVx4_ASAP7_75t_L g1391 ( 
.A(n_1145),
.Y(n_1391)
);

INVx8_ASAP7_75t_L g1392 ( 
.A(n_1210),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1296),
.A2(n_1165),
.B1(n_765),
.B2(n_340),
.Y(n_1393)
);

BUFx12f_ASAP7_75t_L g1394 ( 
.A(n_1275),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1275),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1295),
.Y(n_1396)
);

AOI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1284),
.A2(n_1140),
.B1(n_805),
.B2(n_1150),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1175),
.Y(n_1398)
);

BUFx12f_ASAP7_75t_L g1399 ( 
.A(n_1275),
.Y(n_1399)
);

INVx3_ASAP7_75t_L g1400 ( 
.A(n_1145),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1280),
.A2(n_814),
.B1(n_1291),
.B2(n_1283),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1175),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1194),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1275),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1231),
.A2(n_663),
.B1(n_467),
.B2(n_1228),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_SL g1406 ( 
.A1(n_1165),
.A2(n_333),
.B1(n_341),
.B2(n_340),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1231),
.A2(n_663),
.B1(n_467),
.B2(n_1228),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1274),
.A2(n_1278),
.B1(n_1288),
.B2(n_1150),
.Y(n_1408)
);

AOI22xp33_ASAP7_75t_SL g1409 ( 
.A1(n_1296),
.A2(n_1165),
.B1(n_765),
.B2(n_340),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_L g1410 ( 
.A1(n_1231),
.A2(n_663),
.B1(n_467),
.B2(n_1228),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1248),
.B(n_1251),
.Y(n_1411)
);

CKINVDCx11_ASAP7_75t_R g1412 ( 
.A(n_1275),
.Y(n_1412)
);

CKINVDCx11_ASAP7_75t_R g1413 ( 
.A(n_1275),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1150),
.A2(n_1249),
.B1(n_1259),
.B2(n_995),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1231),
.A2(n_663),
.B1(n_467),
.B2(n_1228),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1295),
.Y(n_1416)
);

INVx4_ASAP7_75t_L g1417 ( 
.A(n_1145),
.Y(n_1417)
);

CKINVDCx20_ASAP7_75t_R g1418 ( 
.A(n_1275),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1374),
.B(n_1311),
.Y(n_1419)
);

AOI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1336),
.A2(n_1383),
.B(n_1305),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1366),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_L g1422 ( 
.A(n_1408),
.B(n_1352),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1303),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1334),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1397),
.A2(n_1401),
.B(n_1382),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1378),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1334),
.Y(n_1427)
);

INVx11_ASAP7_75t_L g1428 ( 
.A(n_1302),
.Y(n_1428)
);

OA21x2_ASAP7_75t_L g1429 ( 
.A1(n_1364),
.A2(n_1367),
.B(n_1358),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1371),
.B(n_1372),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1318),
.Y(n_1431)
);

AOI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1336),
.A2(n_1372),
.B(n_1371),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_SL g1433 ( 
.A1(n_1382),
.A2(n_1401),
.B1(n_1325),
.B2(n_1379),
.Y(n_1433)
);

CKINVDCx6p67_ASAP7_75t_R g1434 ( 
.A(n_1300),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1321),
.B(n_1330),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1333),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1377),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1306),
.B(n_1308),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1337),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1341),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1376),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1376),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1338),
.B(n_1319),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1305),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1375),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1383),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1385),
.Y(n_1447)
);

OA21x2_ASAP7_75t_L g1448 ( 
.A1(n_1373),
.A2(n_1368),
.B(n_1385),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1375),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1411),
.A2(n_1315),
.B(n_1325),
.Y(n_1450)
);

BUFx2_ASAP7_75t_L g1451 ( 
.A(n_1375),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1338),
.B(n_1319),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1370),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1411),
.A2(n_1365),
.B(n_1353),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1378),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1363),
.A2(n_1351),
.B(n_1356),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1360),
.A2(n_1389),
.B(n_1361),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1346),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1346),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1389),
.A2(n_1349),
.B(n_1359),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1344),
.Y(n_1461)
);

AO31x2_ASAP7_75t_L g1462 ( 
.A1(n_1403),
.A2(n_1398),
.A3(n_1381),
.B(n_1402),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1307),
.A2(n_1414),
.B(n_1314),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1314),
.B(n_1304),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1387),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1309),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1378),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1369),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1301),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1327),
.B(n_1396),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1301),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1298),
.B(n_1416),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1393),
.B(n_1409),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1352),
.B(n_1310),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1339),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1362),
.Y(n_1476)
);

INVx4_ASAP7_75t_L g1477 ( 
.A(n_1332),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1316),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1354),
.B(n_1384),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1340),
.A2(n_1347),
.B(n_1348),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1386),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1390),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_1392),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1405),
.B(n_1407),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1339),
.B(n_1345),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1345),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1313),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1317),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1406),
.A2(n_1410),
.B1(n_1415),
.B2(n_1323),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1326),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1350),
.B(n_1400),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1343),
.A2(n_1323),
.B(n_1335),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1388),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1335),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1391),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1417),
.Y(n_1496)
);

OR2x6_ASAP7_75t_L g1497 ( 
.A(n_1392),
.B(n_1399),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1342),
.B(n_1357),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1392),
.A2(n_1355),
.B(n_1331),
.Y(n_1499)
);

INVxp67_ASAP7_75t_R g1500 ( 
.A(n_1322),
.Y(n_1500)
);

CKINVDCx20_ASAP7_75t_R g1501 ( 
.A(n_1434),
.Y(n_1501)
);

INVxp67_ASAP7_75t_L g1502 ( 
.A(n_1424),
.Y(n_1502)
);

OR2x2_ASAP7_75t_L g1503 ( 
.A(n_1423),
.B(n_1297),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1441),
.Y(n_1504)
);

OAI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1425),
.A2(n_1394),
.B1(n_1418),
.B2(n_1404),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1437),
.B(n_1328),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1465),
.B(n_1324),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1473),
.A2(n_1302),
.B1(n_1329),
.B2(n_1413),
.Y(n_1508)
);

NOR2x1_ASAP7_75t_SL g1509 ( 
.A(n_1480),
.B(n_1477),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1473),
.A2(n_1312),
.B1(n_1320),
.B2(n_1299),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1465),
.B(n_1380),
.Y(n_1511)
);

NOR2xp33_ASAP7_75t_L g1512 ( 
.A(n_1450),
.B(n_1433),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1435),
.B(n_1395),
.Y(n_1513)
);

OA21x2_ASAP7_75t_L g1514 ( 
.A1(n_1420),
.A2(n_1412),
.B(n_1458),
.Y(n_1514)
);

OA21x2_ASAP7_75t_L g1515 ( 
.A1(n_1458),
.A2(n_1459),
.B(n_1456),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1451),
.B(n_1445),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1481),
.B(n_1422),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1444),
.B(n_1446),
.Y(n_1518)
);

NAND2x1_ASAP7_75t_L g1519 ( 
.A(n_1477),
.B(n_1476),
.Y(n_1519)
);

A2O1A1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1463),
.A2(n_1443),
.B(n_1452),
.C(n_1464),
.Y(n_1520)
);

OAI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1459),
.A2(n_1468),
.B(n_1456),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1444),
.B(n_1446),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1447),
.B(n_1424),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1468),
.A2(n_1443),
.B(n_1452),
.Y(n_1524)
);

OAI211xp5_ASAP7_75t_L g1525 ( 
.A1(n_1447),
.A2(n_1464),
.B(n_1471),
.C(n_1469),
.Y(n_1525)
);

A2O1A1Ixp33_ASAP7_75t_L g1526 ( 
.A1(n_1469),
.A2(n_1471),
.B(n_1484),
.C(n_1474),
.Y(n_1526)
);

BUFx2_ASAP7_75t_L g1527 ( 
.A(n_1476),
.Y(n_1527)
);

NOR4xp25_ASAP7_75t_SL g1528 ( 
.A(n_1495),
.B(n_1494),
.C(n_1493),
.D(n_1487),
.Y(n_1528)
);

AOI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1474),
.A2(n_1478),
.B1(n_1472),
.B2(n_1480),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1427),
.B(n_1482),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1427),
.B(n_1441),
.Y(n_1531)
);

CKINVDCx20_ASAP7_75t_R g1532 ( 
.A(n_1434),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1442),
.B(n_1431),
.Y(n_1533)
);

AOI221xp5_ASAP7_75t_L g1534 ( 
.A1(n_1442),
.A2(n_1484),
.B1(n_1489),
.B2(n_1478),
.C(n_1430),
.Y(n_1534)
);

INVxp67_ASAP7_75t_L g1535 ( 
.A(n_1429),
.Y(n_1535)
);

OAI211xp5_ASAP7_75t_SL g1536 ( 
.A1(n_1470),
.A2(n_1483),
.B(n_1487),
.C(n_1490),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1436),
.B(n_1439),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1472),
.A2(n_1480),
.B1(n_1486),
.B2(n_1419),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1440),
.B(n_1461),
.Y(n_1539)
);

NOR2xp33_ASAP7_75t_L g1540 ( 
.A(n_1429),
.B(n_1495),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_SL g1541 ( 
.A1(n_1483),
.A2(n_1428),
.B(n_1496),
.C(n_1500),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1429),
.B(n_1488),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1419),
.B(n_1491),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1454),
.B(n_1438),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1462),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1485),
.B(n_1493),
.Y(n_1546)
);

NAND4xp25_ASAP7_75t_L g1547 ( 
.A(n_1498),
.B(n_1455),
.C(n_1467),
.D(n_1426),
.Y(n_1547)
);

OA21x2_ASAP7_75t_L g1548 ( 
.A1(n_1457),
.A2(n_1460),
.B(n_1432),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1504),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1502),
.B(n_1454),
.Y(n_1551)
);

INVxp67_ASAP7_75t_L g1552 ( 
.A(n_1540),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1543),
.B(n_1448),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1502),
.B(n_1454),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1512),
.A2(n_1454),
.B1(n_1486),
.B2(n_1497),
.C(n_1448),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1522),
.B(n_1448),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1519),
.Y(n_1557)
);

NOR2x1_ASAP7_75t_L g1558 ( 
.A(n_1536),
.B(n_1497),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1542),
.B(n_1448),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1523),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1540),
.B(n_1453),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1539),
.Y(n_1562)
);

AOI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1512),
.A2(n_1460),
.B1(n_1475),
.B2(n_1479),
.Y(n_1563)
);

INVxp67_ASAP7_75t_SL g1564 ( 
.A(n_1535),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1527),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1545),
.Y(n_1566)
);

AND2x4_ASAP7_75t_L g1567 ( 
.A(n_1516),
.B(n_1449),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1531),
.Y(n_1568)
);

INVx2_ASAP7_75t_SL g1569 ( 
.A(n_1537),
.Y(n_1569)
);

INVxp67_ASAP7_75t_L g1570 ( 
.A(n_1509),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1533),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1544),
.B(n_1421),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1553),
.B(n_1530),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1568),
.B(n_1560),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1556),
.B(n_1544),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1549),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1553),
.B(n_1530),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1549),
.Y(n_1578)
);

INVx4_ASAP7_75t_L g1579 ( 
.A(n_1557),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1550),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1557),
.Y(n_1581)
);

INVx5_ASAP7_75t_SL g1582 ( 
.A(n_1567),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1556),
.B(n_1518),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1550),
.Y(n_1584)
);

AND2x2_ASAP7_75t_SL g1585 ( 
.A(n_1559),
.B(n_1514),
.Y(n_1585)
);

INVx2_ASAP7_75t_L g1586 ( 
.A(n_1566),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1551),
.B(n_1520),
.C(n_1514),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1572),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1565),
.B(n_1505),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1553),
.B(n_1515),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_R g1591 ( 
.A(n_1559),
.B(n_1528),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1572),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1552),
.B(n_1515),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1555),
.A2(n_1534),
.B1(n_1524),
.B2(n_1529),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1552),
.B(n_1533),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1559),
.B(n_1546),
.Y(n_1596)
);

AOI222xp33_ASAP7_75t_L g1597 ( 
.A1(n_1555),
.A2(n_1534),
.B1(n_1525),
.B2(n_1505),
.C1(n_1508),
.C2(n_1526),
.Y(n_1597)
);

OR2x6_ASAP7_75t_L g1598 ( 
.A(n_1570),
.B(n_1525),
.Y(n_1598)
);

AOI221xp5_ASAP7_75t_L g1599 ( 
.A1(n_1551),
.A2(n_1508),
.B1(n_1521),
.B2(n_1538),
.C(n_1510),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1561),
.B(n_1548),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1586),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1576),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1583),
.B(n_1571),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1576),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1583),
.B(n_1571),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1586),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1593),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1583),
.B(n_1562),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_SL g1609 ( 
.A(n_1585),
.B(n_1558),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1576),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1581),
.Y(n_1611)
);

NAND4xp25_ASAP7_75t_L g1612 ( 
.A(n_1589),
.B(n_1517),
.C(n_1503),
.D(n_1513),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1600),
.B(n_1564),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1589),
.B(n_1565),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1582),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1573),
.B(n_1577),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1575),
.B(n_1554),
.Y(n_1617)
);

INVx3_ASAP7_75t_L g1618 ( 
.A(n_1582),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1573),
.B(n_1577),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1573),
.B(n_1569),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_1581),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1578),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1578),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1575),
.B(n_1554),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1597),
.A2(n_1594),
.B1(n_1587),
.B2(n_1599),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1588),
.B(n_1562),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1596),
.B(n_1569),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1615),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1622),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1616),
.B(n_1585),
.Y(n_1630)
);

HB1xp67_ASAP7_75t_L g1631 ( 
.A(n_1622),
.Y(n_1631)
);

NOR2x1_ASAP7_75t_L g1632 ( 
.A(n_1615),
.B(n_1501),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1615),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1616),
.B(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1623),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1623),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1625),
.B(n_1588),
.Y(n_1637)
);

OAI21xp33_ASAP7_75t_L g1638 ( 
.A1(n_1625),
.A2(n_1597),
.B(n_1587),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1603),
.B(n_1588),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1602),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1616),
.B(n_1585),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1601),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1616),
.B(n_1581),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1602),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1619),
.B(n_1581),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1604),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1604),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1619),
.B(n_1615),
.Y(n_1648)
);

CKINVDCx20_ASAP7_75t_R g1649 ( 
.A(n_1614),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1601),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1603),
.B(n_1592),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1601),
.Y(n_1652)
);

INVx2_ASAP7_75t_SL g1653 ( 
.A(n_1615),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1604),
.Y(n_1654)
);

INVx2_ASAP7_75t_SL g1655 ( 
.A(n_1615),
.Y(n_1655)
);

CKINVDCx16_ASAP7_75t_R g1656 ( 
.A(n_1614),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1610),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1610),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1618),
.B(n_1579),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1617),
.B(n_1595),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1610),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1618),
.B(n_1607),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1605),
.B(n_1592),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1601),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1606),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1606),
.Y(n_1666)
);

OAI33xp33_ASAP7_75t_L g1667 ( 
.A1(n_1612),
.A2(n_1595),
.A3(n_1574),
.B1(n_1584),
.B2(n_1580),
.B3(n_1592),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1631),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1638),
.B(n_1607),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1618),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1605),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1642),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1630),
.B(n_1618),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1660),
.B(n_1608),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1642),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1630),
.B(n_1618),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1656),
.B(n_1608),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1631),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1656),
.B(n_1617),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1660),
.B(n_1617),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1648),
.B(n_1618),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1634),
.B(n_1611),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1634),
.B(n_1611),
.Y(n_1683)
);

NAND4xp25_ASAP7_75t_L g1684 ( 
.A(n_1662),
.B(n_1612),
.C(n_1621),
.D(n_1613),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1649),
.B(n_1620),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1634),
.B(n_1627),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1647),
.Y(n_1687)
);

OR2x6_ASAP7_75t_L g1688 ( 
.A(n_1632),
.B(n_1558),
.Y(n_1688)
);

HB1xp67_ASAP7_75t_L g1689 ( 
.A(n_1629),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1660),
.B(n_1639),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1637),
.B(n_1624),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1642),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1641),
.B(n_1627),
.Y(n_1694)
);

NAND3xp33_ASAP7_75t_L g1695 ( 
.A(n_1649),
.B(n_1635),
.C(n_1629),
.Y(n_1695)
);

INVxp67_ASAP7_75t_SL g1696 ( 
.A(n_1662),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1641),
.B(n_1627),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1641),
.B(n_1627),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1635),
.B(n_1624),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1647),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1648),
.B(n_1621),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1636),
.B(n_1626),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1648),
.B(n_1621),
.Y(n_1703)
);

INVx1_ASAP7_75t_SL g1704 ( 
.A(n_1679),
.Y(n_1704)
);

AOI222xp33_ASAP7_75t_L g1705 ( 
.A1(n_1669),
.A2(n_1667),
.B1(n_1599),
.B2(n_1594),
.C1(n_1593),
.C2(n_1609),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1679),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1687),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1687),
.Y(n_1708)
);

AOI21xp5_ASAP7_75t_L g1709 ( 
.A1(n_1669),
.A2(n_1667),
.B(n_1609),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1684),
.A2(n_1632),
.B(n_1662),
.Y(n_1710)
);

NAND2x1_ASAP7_75t_SL g1711 ( 
.A(n_1670),
.B(n_1659),
.Y(n_1711)
);

A2O1A1Ixp33_ASAP7_75t_L g1712 ( 
.A1(n_1671),
.A2(n_1684),
.B(n_1692),
.C(n_1690),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1670),
.B(n_1643),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1671),
.A2(n_1612),
.B(n_1628),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1700),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1700),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1690),
.A2(n_1692),
.B1(n_1591),
.B2(n_1695),
.Y(n_1717)
);

OAI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1695),
.A2(n_1696),
.B(n_1633),
.Y(n_1718)
);

OAI322xp33_ASAP7_75t_L g1719 ( 
.A1(n_1677),
.A2(n_1636),
.A3(n_1591),
.B1(n_1655),
.B2(n_1653),
.C1(n_1651),
.C2(n_1639),
.Y(n_1719)
);

OAI21xp33_ASAP7_75t_L g1720 ( 
.A1(n_1677),
.A2(n_1645),
.B(n_1643),
.Y(n_1720)
);

OAI322xp33_ASAP7_75t_L g1721 ( 
.A1(n_1691),
.A2(n_1653),
.A3(n_1655),
.B1(n_1651),
.B2(n_1663),
.C1(n_1661),
.C2(n_1644),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1673),
.B(n_1643),
.Y(n_1722)
);

AOI22xp33_ASAP7_75t_L g1723 ( 
.A1(n_1672),
.A2(n_1598),
.B1(n_1590),
.B2(n_1593),
.Y(n_1723)
);

OAI21xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1673),
.A2(n_1655),
.B(n_1653),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1676),
.A2(n_1598),
.B1(n_1682),
.B2(n_1683),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1680),
.B(n_1663),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1672),
.Y(n_1727)
);

NOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1668),
.B(n_1532),
.Y(n_1728)
);

OAI22xp33_ASAP7_75t_L g1729 ( 
.A1(n_1688),
.A2(n_1598),
.B1(n_1563),
.B2(n_1628),
.Y(n_1729)
);

AOI21xp33_ASAP7_75t_SL g1730 ( 
.A1(n_1705),
.A2(n_1685),
.B(n_1688),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1704),
.B(n_1691),
.Y(n_1731)
);

AOI221xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1712),
.A2(n_1668),
.B1(n_1678),
.B2(n_1683),
.C(n_1682),
.Y(n_1732)
);

AND2x4_ASAP7_75t_L g1733 ( 
.A(n_1728),
.B(n_1681),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1717),
.A2(n_1676),
.B(n_1680),
.C(n_1590),
.Y(n_1734)
);

INVx1_ASAP7_75t_SL g1735 ( 
.A(n_1706),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1714),
.B(n_1686),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1711),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1713),
.B(n_1686),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1727),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1722),
.B(n_1694),
.Y(n_1740)
);

AOI31xp33_ASAP7_75t_L g1741 ( 
.A1(n_1718),
.A2(n_1678),
.A3(n_1701),
.B(n_1703),
.Y(n_1741)
);

NOR3xp33_ASAP7_75t_L g1742 ( 
.A(n_1719),
.B(n_1710),
.C(n_1729),
.Y(n_1742)
);

AOI33xp33_ASAP7_75t_L g1743 ( 
.A1(n_1723),
.A2(n_1703),
.A3(n_1701),
.B1(n_1681),
.B2(n_1694),
.B3(n_1697),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1726),
.B(n_1697),
.Y(n_1744)
);

O2A1O1Ixp5_ASAP7_75t_L g1745 ( 
.A1(n_1709),
.A2(n_1681),
.B(n_1699),
.C(n_1702),
.Y(n_1745)
);

AOI221xp5_ASAP7_75t_L g1746 ( 
.A1(n_1721),
.A2(n_1699),
.B1(n_1672),
.B2(n_1693),
.C(n_1675),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1707),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1727),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1720),
.B(n_1698),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1723),
.B(n_1689),
.C(n_1633),
.Y(n_1750)
);

XNOR2xp5_ASAP7_75t_L g1751 ( 
.A(n_1735),
.B(n_1725),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1739),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1748),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1731),
.B(n_1698),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1744),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1747),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_SL g1757 ( 
.A1(n_1741),
.A2(n_1715),
.B(n_1708),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1738),
.Y(n_1758)
);

NOR4xp25_ASAP7_75t_L g1759 ( 
.A(n_1743),
.B(n_1716),
.C(n_1724),
.D(n_1729),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1740),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1749),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1756),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1754),
.B(n_1732),
.Y(n_1763)
);

NOR5xp2_ASAP7_75t_L g1764 ( 
.A(n_1757),
.B(n_1750),
.C(n_1734),
.D(n_1753),
.E(n_1752),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1751),
.Y(n_1765)
);

NAND3xp33_ASAP7_75t_L g1766 ( 
.A(n_1757),
.B(n_1732),
.C(n_1742),
.Y(n_1766)
);

NAND4xp25_ASAP7_75t_L g1767 ( 
.A(n_1761),
.B(n_1745),
.C(n_1736),
.D(n_1733),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1755),
.Y(n_1768)
);

NOR3xp33_ASAP7_75t_L g1769 ( 
.A(n_1760),
.B(n_1730),
.C(n_1746),
.Y(n_1769)
);

NAND4xp25_ASAP7_75t_L g1770 ( 
.A(n_1758),
.B(n_1733),
.C(n_1681),
.D(n_1628),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_SL g1771 ( 
.A(n_1766),
.B(n_1759),
.Y(n_1771)
);

NAND3xp33_ASAP7_75t_SL g1772 ( 
.A(n_1764),
.B(n_1633),
.C(n_1466),
.Y(n_1772)
);

CKINVDCx20_ASAP7_75t_R g1773 ( 
.A(n_1765),
.Y(n_1773)
);

XNOR2xp5_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1499),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1762),
.B(n_1737),
.Y(n_1775)
);

OAI211xp5_ASAP7_75t_SL g1776 ( 
.A1(n_1771),
.A2(n_1763),
.B(n_1769),
.C(n_1768),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1773),
.Y(n_1777)
);

OAI221xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1774),
.A2(n_1770),
.B1(n_1688),
.B2(n_1693),
.C(n_1675),
.Y(n_1778)
);

AND4x1_ASAP7_75t_L g1779 ( 
.A(n_1775),
.B(n_1498),
.C(n_1428),
.D(n_1500),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_SL g1780 ( 
.A(n_1772),
.B(n_1466),
.Y(n_1780)
);

NAND4xp25_ASAP7_75t_L g1781 ( 
.A(n_1772),
.B(n_1467),
.C(n_1455),
.D(n_1426),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1777),
.B(n_1674),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1779),
.B(n_1645),
.Y(n_1783)
);

NAND4xp75_ASAP7_75t_L g1784 ( 
.A(n_1780),
.B(n_1693),
.C(n_1675),
.D(n_1702),
.Y(n_1784)
);

NOR3xp33_ASAP7_75t_L g1785 ( 
.A(n_1776),
.B(n_1499),
.C(n_1674),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1781),
.Y(n_1786)
);

NOR3xp33_ASAP7_75t_L g1787 ( 
.A(n_1785),
.B(n_1778),
.C(n_1652),
.Y(n_1787)
);

OAI221xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1782),
.A2(n_1688),
.B1(n_1511),
.B2(n_1665),
.C(n_1664),
.Y(n_1788)
);

OR2x2_ASAP7_75t_L g1789 ( 
.A(n_1784),
.B(n_1645),
.Y(n_1789)
);

OAI22xp33_ASAP7_75t_L g1790 ( 
.A1(n_1789),
.A2(n_1786),
.B1(n_1783),
.B2(n_1688),
.Y(n_1790)
);

AOI22xp5_ASAP7_75t_L g1791 ( 
.A1(n_1790),
.A2(n_1787),
.B1(n_1788),
.B2(n_1666),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1791),
.A2(n_1506),
.B1(n_1507),
.B2(n_1644),
.Y(n_1792)
);

XNOR2xp5_ASAP7_75t_L g1793 ( 
.A(n_1791),
.B(n_1492),
.Y(n_1793)
);

XNOR2xp5_ASAP7_75t_L g1794 ( 
.A(n_1793),
.B(n_1492),
.Y(n_1794)
);

OAI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1792),
.A2(n_1666),
.B1(n_1665),
.B2(n_1664),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1794),
.A2(n_1652),
.B(n_1650),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1795),
.A2(n_1666),
.B1(n_1665),
.B2(n_1664),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_R g1798 ( 
.A1(n_1797),
.A2(n_1650),
.B1(n_1652),
.B2(n_1658),
.Y(n_1798)
);

AOI21xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1798),
.A2(n_1796),
.B(n_1659),
.Y(n_1799)
);

OAI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1650),
.B1(n_1640),
.B2(n_1658),
.Y(n_1800)
);

AOI221xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1661),
.B1(n_1646),
.B2(n_1657),
.C(n_1654),
.Y(n_1801)
);

AOI211xp5_ASAP7_75t_L g1802 ( 
.A1(n_1801),
.A2(n_1541),
.B(n_1659),
.C(n_1547),
.Y(n_1802)
);


endmodule