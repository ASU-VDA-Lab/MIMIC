module real_jpeg_25370_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_355, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_355;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_1),
.A2(n_30),
.B1(n_33),
.B2(n_49),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_1),
.A2(n_49),
.B1(n_66),
.B2(n_69),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_1),
.A2(n_49),
.B1(n_90),
.B2(n_305),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_2),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_32)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_2),
.A2(n_34),
.B1(n_47),
.B2(n_48),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g295 ( 
.A1(n_2),
.A2(n_34),
.B1(n_66),
.B2(n_69),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_2),
.A2(n_34),
.B1(n_96),
.B2(n_97),
.Y(n_324)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_30),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_5),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_5),
.A2(n_40),
.B1(n_66),
.B2(n_69),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_L g287 ( 
.A1(n_5),
.A2(n_40),
.B1(n_80),
.B2(n_88),
.Y(n_287)
);

INVx8_ASAP7_75t_SL g86 ( 
.A(n_6),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_7),
.A2(n_61),
.B1(n_66),
.B2(n_69),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_7),
.A2(n_30),
.B1(n_33),
.B2(n_61),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_7),
.A2(n_61),
.B1(n_81),
.B2(n_90),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_8),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_68),
.B1(n_81),
.B2(n_90),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_8),
.A2(n_30),
.B1(n_33),
.B2(n_68),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_9),
.A2(n_66),
.B1(n_69),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_9),
.A2(n_30),
.B1(n_33),
.B2(n_77),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_77),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_9),
.A2(n_77),
.B1(n_81),
.B2(n_90),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_10),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_10),
.B(n_91),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_10),
.B(n_30),
.C(n_44),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_82),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_10),
.B(n_75),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_10),
.A2(n_29),
.B1(n_173),
.B2(n_174),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_11),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_12),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_12),
.A2(n_66),
.B1(n_69),
.B2(n_95),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_12),
.A2(n_47),
.B1(n_48),
.B2(n_95),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_12),
.A2(n_30),
.B1(n_33),
.B2(n_95),
.Y(n_173)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_13),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_15),
.Y(n_176)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_348),
.C(n_353),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_346),
.B(n_351),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_333),
.B(n_345),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_299),
.A3(n_326),
.B1(n_331),
.B2(n_332),
.C(n_355),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_274),
.B(n_298),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_250),
.B(n_273),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_135),
.B(n_224),
.C(n_249),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_119),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_24),
.B(n_119),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_99),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_55),
.B2(n_56),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_26),
.B(n_56),
.C(n_99),
.Y(n_225)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_41),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_28),
.B(n_41),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_32),
.B(n_35),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_29),
.A2(n_32),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_29),
.B(n_39),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_29),
.A2(n_156),
.B(n_157),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_29),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_29),
.A2(n_115),
.B1(n_164),
.B2(n_173),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_29),
.A2(n_31),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_30),
.A2(n_33),
.B1(n_43),
.B2(n_44),
.Y(n_42)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx5_ASAP7_75t_L g180 ( 
.A(n_31),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_33),
.B(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_36),
.A2(n_158),
.B(n_162),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_37),
.Y(n_133)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_46),
.B(n_50),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_42),
.A2(n_53),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_42),
.A2(n_53),
.B1(n_147),
.B2(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_42),
.B(n_82),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_42),
.A2(n_46),
.B1(n_53),
.B2(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_42),
.A2(n_53),
.B(n_59),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_43),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_54)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx24_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_48),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_47),
.B(n_66),
.C(n_73),
.Y(n_192)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_48),
.B(n_143),
.Y(n_142)
);

A2O1A1Ixp33_ASAP7_75t_L g190 ( 
.A1(n_48),
.A2(n_72),
.B(n_191),
.C(n_192),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_50),
.B(n_214),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_52),
.A2(n_63),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_53),
.A2(n_59),
.B(n_62),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_53),
.A2(n_213),
.B(n_214),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_53),
.A2(n_62),
.B(n_245),
.Y(n_258)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_64),
.C(n_78),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_57),
.A2(n_58),
.B1(n_64),
.B2(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_60),
.B(n_63),
.Y(n_214)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_75),
.B2(n_76),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_65),
.Y(n_128)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_69),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_66),
.A2(n_79),
.B(n_85),
.C(n_117),
.Y(n_116)
);

HAxp5_ASAP7_75t_SL g191 ( 
.A(n_66),
.B(n_82),
.CON(n_191),
.SN(n_191)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_80),
.C(n_86),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_70),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_70),
.A2(n_75),
.B1(n_127),
.B2(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_70),
.B(n_238),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_70),
.A2(n_75),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_70),
.A2(n_75),
.B(n_110),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_74),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_71),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_108),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_71),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_75),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_75),
.B(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g120 ( 
.A(n_78),
.B(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_83),
.B1(n_91),
.B2(n_92),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_82),
.CON(n_79),
.SN(n_79)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_80),
.Y(n_305)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_82),
.B(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_83),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_83),
.A2(n_91),
.B1(n_105),
.B2(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_83),
.B(n_287),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_83),
.A2(n_91),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_83),
.A2(n_324),
.B(n_340),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_83),
.A2(n_91),
.B(n_266),
.Y(n_353)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_87),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_84),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_93),
.B1(n_103),
.B2(n_104),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_84),
.A2(n_304),
.B(n_306),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_L g87 ( 
.A1(n_85),
.A2(n_86),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_91),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_91),
.B(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_111),
.B2(n_118),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_106),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_102),
.B(n_106),
.C(n_118),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_103),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_103),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B(n_109),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g235 ( 
.A1(n_108),
.A2(n_236),
.B(n_237),
.Y(n_235)
);

OAI21xp33_ASAP7_75t_L g309 ( 
.A1(n_108),
.A2(n_237),
.B(n_295),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_109),
.B(n_269),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_110),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_111),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_112),
.B(n_116),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_114),
.A2(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_123),
.C(n_124),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_120),
.B(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_123),
.B(n_124),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.C(n_131),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_125),
.B(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_134),
.B(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_223),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_218),
.B(n_222),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_203),
.B(n_217),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_187),
.B(n_202),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_159),
.B(n_186),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_148),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_148),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_144),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_142),
.Y(n_169)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_155),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_153),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_154),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_156),
.Y(n_167)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_157),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_158),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_170),
.B(n_185),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_165),
.B2(n_167),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_181),
.B(n_184),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_182),
.B(n_183),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_188),
.B(n_201),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_201),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_196),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_189),
.B(n_197),
.C(n_200),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_190),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_195),
.Y(n_211)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_193),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_204),
.B(n_205),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_212),
.C(n_215),
.Y(n_221)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_215),
.B2(n_216),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_221),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_225),
.B(n_226),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_248),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_239),
.B1(n_246),
.B2(n_247),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_232),
.C(n_234),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_234),
.B2(n_235),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_239),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_246),
.C(n_248),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_244),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_240),
.B(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_252),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_251),
.B(n_252),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_272),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_260),
.C(n_272),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_255),
.A2(n_256),
.B1(n_283),
.B2(n_284),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_255),
.A2(n_280),
.B(n_284),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_256),
.B(n_258),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_258),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_261),
.A2(n_262),
.B1(n_270),
.B2(n_271),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_263),
.B(n_267),
.C(n_271),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_265),
.B(n_306),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_266),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_270),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_275),
.B(n_276),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_297),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_289),
.B2(n_290),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_289),
.C(n_297),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_288),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_282),
.Y(n_288)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_286),
.Y(n_340)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B(n_296),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_292),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_296),
.A2(n_301),
.B1(n_313),
.B2(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_315),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_315),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_313),
.C(n_314),
.Y(n_300)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_301),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_307),
.B2(n_312),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_302),
.A2(n_303),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_303),
.B(n_308),
.C(n_311),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_303),
.B(n_318),
.C(n_325),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_304),
.Y(n_323)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_310),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_310),
.A2(n_311),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_310),
.B(n_320),
.C(n_322),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_329),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_325),
.Y(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_335),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_336),
.A2(n_337),
.B1(n_343),
.B2(n_344),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_338),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_339),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_339),
.B(n_341),
.C(n_343),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g343 ( 
.A(n_344),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_349),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_348),
.Y(n_352)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_350),
.B(n_352),
.Y(n_351)
);


endmodule