module real_aes_6399_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g171 ( .A1(n_0), .A2(n_172), .B(n_175), .C(n_179), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_1), .B(n_163), .Y(n_182) );
INVx1_ASAP7_75t_L g105 ( .A(n_2), .Y(n_105) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_3), .B(n_173), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g520 ( .A1(n_4), .A2(n_136), .B(n_139), .C(n_521), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_5), .A2(n_131), .B(n_546), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_6), .A2(n_131), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_7), .B(n_163), .Y(n_552) );
AO21x2_ASAP7_75t_L g236 ( .A1(n_8), .A2(n_165), .B(n_237), .Y(n_236) );
AND2x6_ASAP7_75t_L g136 ( .A(n_9), .B(n_137), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_10), .A2(n_136), .B(n_139), .C(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g512 ( .A(n_11), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_12), .B(n_111), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g448 ( .A(n_12), .B(n_39), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g523 ( .A(n_13), .B(n_178), .Y(n_523) );
INVx1_ASAP7_75t_L g157 ( .A(n_14), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_15), .B(n_173), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_16), .A2(n_174), .B(n_532), .C(n_534), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_17), .B(n_163), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_18), .B(n_151), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g138 ( .A1(n_19), .A2(n_139), .B(n_142), .C(n_150), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_L g561 ( .A1(n_20), .A2(n_177), .B(n_245), .C(n_562), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_21), .B(n_178), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_22), .A2(n_74), .B1(n_454), .B2(n_743), .C1(n_746), .C2(n_747), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_23), .B(n_178), .Y(n_474) );
CKINVDCx16_ASAP7_75t_R g493 ( .A(n_24), .Y(n_493) );
INVx1_ASAP7_75t_L g473 ( .A(n_25), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_26), .A2(n_139), .B(n_150), .C(n_240), .Y(n_239) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_27), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g519 ( .A(n_28), .Y(n_519) );
INVx1_ASAP7_75t_L g487 ( .A(n_29), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_30), .A2(n_131), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g134 ( .A(n_31), .Y(n_134) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_32), .A2(n_189), .B(n_190), .C(n_194), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_33), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_34), .A2(n_177), .B(n_549), .C(n_551), .Y(n_548) );
INVxp67_ASAP7_75t_L g488 ( .A(n_35), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_36), .B(n_242), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g471 ( .A1(n_37), .A2(n_139), .B(n_150), .C(n_472), .Y(n_471) );
CKINVDCx14_ASAP7_75t_R g547 ( .A(n_38), .Y(n_547) );
INVx1_ASAP7_75t_L g111 ( .A(n_39), .Y(n_111) );
A2O1A1Ixp33_ASAP7_75t_L g509 ( .A1(n_40), .A2(n_179), .B(n_510), .C(n_511), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g129 ( .A(n_41), .B(n_130), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g258 ( .A(n_42), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_43), .B(n_173), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_44), .B(n_131), .Y(n_238) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_45), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_46), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_47), .B(n_450), .Y(n_449) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_48), .A2(n_189), .B(n_194), .C(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g176 ( .A(n_49), .Y(n_176) );
INVx1_ASAP7_75t_L g220 ( .A(n_50), .Y(n_220) );
INVx1_ASAP7_75t_L g560 ( .A(n_51), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_52), .B(n_131), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_53), .Y(n_159) );
CKINVDCx14_ASAP7_75t_R g508 ( .A(n_54), .Y(n_508) );
INVx1_ASAP7_75t_L g137 ( .A(n_55), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_56), .B(n_131), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_57), .B(n_163), .Y(n_233) );
A2O1A1Ixp33_ASAP7_75t_L g230 ( .A1(n_58), .A2(n_149), .B(n_205), .C(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g156 ( .A(n_59), .Y(n_156) );
INVx1_ASAP7_75t_SL g550 ( .A(n_60), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_61), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_62), .B(n_173), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_63), .B(n_163), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_64), .B(n_174), .Y(n_255) );
INVx1_ASAP7_75t_L g496 ( .A(n_65), .Y(n_496) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_66), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_67), .B(n_144), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_68), .A2(n_139), .B(n_194), .C(n_203), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g229 ( .A(n_69), .Y(n_229) );
INVx1_ASAP7_75t_L g108 ( .A(n_70), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_71), .A2(n_131), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_72), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_73), .A2(n_131), .B(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_74), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_75), .A2(n_130), .B(n_483), .Y(n_482) );
CKINVDCx16_ASAP7_75t_R g470 ( .A(n_76), .Y(n_470) );
INVx1_ASAP7_75t_L g530 ( .A(n_77), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_78), .B(n_147), .Y(n_146) );
AOI22xp5_ASAP7_75t_L g99 ( .A1(n_79), .A2(n_100), .B1(n_112), .B2(n_751), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_80), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_81), .A2(n_131), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g533 ( .A(n_82), .Y(n_533) );
INVx2_ASAP7_75t_L g154 ( .A(n_83), .Y(n_154) );
INVx1_ASAP7_75t_L g522 ( .A(n_84), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_85), .Y(n_212) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_86), .B(n_178), .Y(n_256) );
NAND3xp33_ASAP7_75t_SL g104 ( .A(n_87), .B(n_105), .C(n_106), .Y(n_104) );
OR2x2_ASAP7_75t_L g445 ( .A(n_87), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g457 ( .A(n_87), .B(n_447), .Y(n_457) );
INVx2_ASAP7_75t_L g462 ( .A(n_87), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_88), .A2(n_139), .B(n_194), .C(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_89), .B(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g191 ( .A(n_90), .Y(n_191) );
INVxp67_ASAP7_75t_L g232 ( .A(n_91), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_92), .A2(n_119), .B1(n_441), .B2(n_442), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_92), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_93), .B(n_165), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_94), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g204 ( .A(n_95), .Y(n_204) );
INVx1_ASAP7_75t_L g251 ( .A(n_96), .Y(n_251) );
INVx2_ASAP7_75t_L g563 ( .A(n_97), .Y(n_563) );
AND2x2_ASAP7_75t_L g222 ( .A(n_98), .B(n_153), .Y(n_222) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
BUFx4f_ASAP7_75t_SL g751 ( .A(n_101), .Y(n_751) );
INVx2_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_109), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
AND2x2_ASAP7_75t_L g447 ( .A(n_105), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
AO21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_452), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g750 ( .A(n_114), .Y(n_750) );
INVx2_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI21xp5_ASAP7_75t_SL g117 ( .A1(n_118), .A2(n_443), .B(n_449), .Y(n_117) );
INVx1_ASAP7_75t_L g442 ( .A(n_119), .Y(n_442) );
INVx2_ASAP7_75t_L g458 ( .A(n_119), .Y(n_458) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_119), .A2(n_455), .B1(n_744), .B2(n_745), .Y(n_743) );
AND2x2_ASAP7_75t_SL g119 ( .A(n_120), .B(n_396), .Y(n_119) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_121), .B(n_331), .Y(n_120) );
NAND4xp25_ASAP7_75t_SL g121 ( .A(n_122), .B(n_276), .C(n_300), .D(n_323), .Y(n_121) );
AOI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_213), .B1(n_247), .B2(n_260), .C(n_263), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_183), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g266 ( .A1(n_125), .A2(n_161), .B1(n_214), .B2(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_125), .B(n_184), .Y(n_334) );
AND2x2_ASAP7_75t_L g353 ( .A(n_125), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_125), .B(n_337), .Y(n_423) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_161), .Y(n_125) );
AND2x2_ASAP7_75t_L g291 ( .A(n_126), .B(n_184), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_126), .B(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g314 ( .A(n_126), .B(n_315), .Y(n_314) );
AND2x2_ASAP7_75t_L g319 ( .A(n_126), .B(n_162), .Y(n_319) );
INVx2_ASAP7_75t_L g351 ( .A(n_126), .Y(n_351) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_126), .Y(n_395) );
AND2x2_ASAP7_75t_L g412 ( .A(n_126), .B(n_289), .Y(n_412) );
INVx5_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g330 ( .A(n_127), .B(n_289), .Y(n_330) );
AND2x4_ASAP7_75t_L g344 ( .A(n_127), .B(n_161), .Y(n_344) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_127), .Y(n_348) );
AND2x2_ASAP7_75t_L g368 ( .A(n_127), .B(n_283), .Y(n_368) );
AND2x2_ASAP7_75t_L g418 ( .A(n_127), .B(n_185), .Y(n_418) );
AND2x2_ASAP7_75t_L g428 ( .A(n_127), .B(n_162), .Y(n_428) );
OR2x6_ASAP7_75t_L g127 ( .A(n_128), .B(n_158), .Y(n_127) );
AOI21xp5_ASAP7_75t_SL g128 ( .A1(n_129), .A2(n_138), .B(n_151), .Y(n_128) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_136), .Y(n_131) );
NAND2x1p5_ASAP7_75t_L g252 ( .A(n_132), .B(n_136), .Y(n_252) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx1_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_L g140 ( .A(n_134), .Y(n_140) );
INVx1_ASAP7_75t_L g246 ( .A(n_134), .Y(n_246) );
INVx1_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_135), .Y(n_145) );
INVx3_ASAP7_75t_L g174 ( .A(n_135), .Y(n_174) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_135), .Y(n_178) );
INVx1_ASAP7_75t_L g242 ( .A(n_135), .Y(n_242) );
BUFx3_ASAP7_75t_L g150 ( .A(n_136), .Y(n_150) );
INVx4_ASAP7_75t_SL g181 ( .A(n_136), .Y(n_181) );
INVx5_ASAP7_75t_L g170 ( .A(n_139), .Y(n_170) );
AND2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
BUFx3_ASAP7_75t_L g180 ( .A(n_140), .Y(n_180) );
BUFx6f_ASAP7_75t_L g209 ( .A(n_140), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B(n_148), .Y(n_142) );
INVx2_ASAP7_75t_L g147 ( .A(n_144), .Y(n_147) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g206 ( .A(n_145), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g190 ( .A1(n_147), .A2(n_191), .B(n_192), .C(n_193), .Y(n_190) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_147), .A2(n_193), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_147), .A2(n_496), .B(n_497), .C(n_498), .Y(n_495) );
O2A1O1Ixp5_ASAP7_75t_L g521 ( .A1(n_147), .A2(n_498), .B(n_522), .C(n_523), .Y(n_521) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_148), .A2(n_173), .B(n_473), .C(n_474), .Y(n_472) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_149), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g499 ( .A(n_152), .B(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx1_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_153), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_153), .A2(n_217), .B(n_218), .Y(n_216) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_153), .A2(n_252), .B(n_470), .C(n_471), .Y(n_469) );
OA21x2_ASAP7_75t_L g505 ( .A1(n_153), .A2(n_506), .B(n_513), .Y(n_505) );
AND2x2_ASAP7_75t_SL g153 ( .A(n_154), .B(n_155), .Y(n_153) );
AND2x2_ASAP7_75t_L g166 ( .A(n_154), .B(n_155), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AO21x2_ASAP7_75t_L g517 ( .A1(n_160), .A2(n_518), .B(n_524), .Y(n_517) );
AND2x2_ASAP7_75t_L g284 ( .A(n_161), .B(n_184), .Y(n_284) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_161), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_161), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g374 ( .A(n_161), .Y(n_374) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g262 ( .A(n_162), .B(n_199), .Y(n_262) );
AND2x2_ASAP7_75t_L g289 ( .A(n_162), .B(n_200), .Y(n_289) );
OA21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_167), .B(n_182), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_164), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g200 ( .A1(n_164), .A2(n_201), .B(n_211), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_164), .B(n_212), .Y(n_211) );
AO21x2_ASAP7_75t_L g249 ( .A1(n_164), .A2(n_250), .B(n_257), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_164), .B(n_476), .Y(n_475) );
AO21x2_ASAP7_75t_L g491 ( .A1(n_164), .A2(n_492), .B(n_499), .Y(n_491) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_164), .B(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_165), .A2(n_238), .B(n_239), .Y(n_237) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx1_ASAP7_75t_L g259 ( .A(n_166), .Y(n_259) );
O2A1O1Ixp33_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B(n_171), .C(n_181), .Y(n_168) );
INVx2_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_170), .A2(n_181), .B(n_229), .C(n_230), .Y(n_228) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_170), .A2(n_181), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_170), .A2(n_181), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_SL g529 ( .A1(n_170), .A2(n_181), .B(n_530), .C(n_531), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_170), .A2(n_181), .B(n_547), .C(n_548), .Y(n_546) );
O2A1O1Ixp33_ASAP7_75t_SL g559 ( .A1(n_170), .A2(n_181), .B(n_560), .C(n_561), .Y(n_559) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_173), .B(n_232), .Y(n_231) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_173), .A2(n_206), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx5_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_174), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_176), .B(n_177), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_177), .B(n_550), .Y(n_549) );
INVx4_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx2_ASAP7_75t_L g510 ( .A(n_178), .Y(n_510) );
INVx2_ASAP7_75t_L g498 ( .A(n_179), .Y(n_498) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_180), .Y(n_193) );
INVx1_ASAP7_75t_L g534 ( .A(n_180), .Y(n_534) );
INVx1_ASAP7_75t_L g194 ( .A(n_181), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_183), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_197), .Y(n_183) );
OR2x2_ASAP7_75t_L g315 ( .A(n_184), .B(n_198), .Y(n_315) );
AND2x2_ASAP7_75t_L g352 ( .A(n_184), .B(n_262), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_184), .B(n_283), .Y(n_363) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_184), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_184), .B(n_319), .Y(n_436) );
INVx5_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g261 ( .A(n_185), .Y(n_261) );
AND2x2_ASAP7_75t_L g270 ( .A(n_185), .B(n_198), .Y(n_270) );
AND2x2_ASAP7_75t_L g386 ( .A(n_185), .B(n_281), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_185), .B(n_319), .Y(n_408) );
OR2x6_ASAP7_75t_L g185 ( .A(n_186), .B(n_195), .Y(n_185) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
HB1xp67_ASAP7_75t_L g354 ( .A(n_198), .Y(n_354) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_199), .Y(n_306) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx2_ASAP7_75t_L g283 ( .A(n_200), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_207), .C(n_208), .Y(n_203) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_206), .B(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_206), .B(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx3_ASAP7_75t_L g551 ( .A(n_209), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_223), .Y(n_213) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_214), .B(n_296), .Y(n_415) );
HB1xp67_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_215), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g267 ( .A(n_215), .B(n_268), .Y(n_267) );
INVx5_ASAP7_75t_SL g275 ( .A(n_215), .Y(n_275) );
OR2x2_ASAP7_75t_L g298 ( .A(n_215), .B(n_268), .Y(n_298) );
OR2x2_ASAP7_75t_L g308 ( .A(n_215), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g371 ( .A(n_215), .B(n_225), .Y(n_371) );
AND2x2_ASAP7_75t_SL g409 ( .A(n_215), .B(n_224), .Y(n_409) );
NOR4xp25_ASAP7_75t_L g430 ( .A(n_215), .B(n_351), .C(n_431), .D(n_432), .Y(n_430) );
AND2x2_ASAP7_75t_L g440 ( .A(n_215), .B(n_272), .Y(n_440) );
OR2x6_ASAP7_75t_L g215 ( .A(n_216), .B(n_222), .Y(n_215) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g265 ( .A(n_224), .B(n_261), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_224), .B(n_267), .Y(n_434) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_234), .Y(n_224) );
OR2x2_ASAP7_75t_L g274 ( .A(n_225), .B(n_275), .Y(n_274) );
INVx3_ASAP7_75t_L g281 ( .A(n_225), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_225), .B(n_249), .Y(n_293) );
INVxp67_ASAP7_75t_L g296 ( .A(n_225), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_225), .B(n_268), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_225), .B(n_235), .Y(n_362) );
AND2x2_ASAP7_75t_L g377 ( .A(n_225), .B(n_272), .Y(n_377) );
OR2x2_ASAP7_75t_L g406 ( .A(n_225), .B(n_235), .Y(n_406) );
OA21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_233), .Y(n_225) );
OA21x2_ASAP7_75t_L g527 ( .A1(n_226), .A2(n_528), .B(n_535), .Y(n_527) );
OA21x2_ASAP7_75t_L g544 ( .A1(n_226), .A2(n_545), .B(n_552), .Y(n_544) );
OA21x2_ASAP7_75t_L g557 ( .A1(n_226), .A2(n_558), .B(n_564), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_234), .B(n_311), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_234), .B(n_275), .Y(n_414) );
OR2x2_ASAP7_75t_L g435 ( .A(n_234), .B(n_312), .Y(n_435) );
INVx1_ASAP7_75t_SL g234 ( .A(n_235), .Y(n_234) );
OR2x2_ASAP7_75t_L g248 ( .A(n_235), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g272 ( .A(n_235), .B(n_268), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_235), .B(n_249), .Y(n_287) );
AND2x2_ASAP7_75t_L g357 ( .A(n_235), .B(n_281), .Y(n_357) );
AND2x2_ASAP7_75t_L g391 ( .A(n_235), .B(n_275), .Y(n_391) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_236), .B(n_275), .Y(n_294) );
AND2x2_ASAP7_75t_L g322 ( .A(n_236), .B(n_249), .Y(n_322) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_243), .B(n_244), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_244), .A2(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx3_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_247), .B(n_330), .Y(n_329) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_248), .A2(n_337), .B1(n_373), .B2(n_390), .C(n_392), .Y(n_389) );
INVx5_ASAP7_75t_SL g268 ( .A(n_249), .Y(n_268) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_252), .B(n_253), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g492 ( .A1(n_252), .A2(n_493), .B(n_494), .Y(n_492) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_252), .A2(n_519), .B(n_520), .Y(n_518) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g481 ( .A(n_259), .Y(n_481) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OAI33xp33_ASAP7_75t_L g288 ( .A1(n_261), .A2(n_289), .A3(n_290), .B1(n_292), .B2(n_295), .B3(n_299), .Y(n_288) );
OR2x2_ASAP7_75t_L g304 ( .A(n_261), .B(n_305), .Y(n_304) );
AOI322xp5_ASAP7_75t_L g413 ( .A1(n_261), .A2(n_330), .A3(n_337), .B1(n_414), .B2(n_415), .C1(n_416), .C2(n_419), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_261), .B(n_289), .Y(n_431) );
A2O1A1Ixp33_ASAP7_75t_SL g437 ( .A1(n_261), .A2(n_289), .B(n_438), .C(n_440), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g276 ( .A1(n_262), .A2(n_277), .B1(n_282), .B2(n_285), .C(n_288), .Y(n_276) );
INVx1_ASAP7_75t_L g369 ( .A(n_262), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_262), .B(n_418), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_266), .B1(n_269), .B2(n_271), .Y(n_263) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g346 ( .A(n_267), .B(n_281), .Y(n_346) );
AND2x2_ASAP7_75t_L g404 ( .A(n_267), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_275), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_268), .B(n_281), .Y(n_340) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_270), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_270), .B(n_348), .Y(n_402) );
OAI321xp33_ASAP7_75t_L g421 ( .A1(n_270), .A2(n_343), .A3(n_422), .B1(n_423), .B2(n_424), .C(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g388 ( .A(n_271), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_272), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g327 ( .A(n_272), .B(n_275), .Y(n_327) );
AOI321xp33_ASAP7_75t_L g385 ( .A1(n_272), .A2(n_289), .A3(n_386), .B1(n_387), .B2(n_388), .C(n_389), .Y(n_385) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g302 ( .A(n_274), .B(n_287), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_275), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_275), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_275), .B(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g321 ( .A(n_279), .B(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g286 ( .A(n_280), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g394 ( .A(n_281), .Y(n_394) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_284), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g317 ( .A(n_289), .Y(n_317) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_291), .B(n_326), .Y(n_375) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OR2x2_ASAP7_75t_L g339 ( .A(n_294), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_SL g384 ( .A(n_294), .Y(n_384) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_295), .A2(n_342), .B1(n_345), .B2(n_347), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g439 ( .A(n_298), .B(n_362), .Y(n_439) );
AOI221xp5_ASAP7_75t_L g300 ( .A1(n_301), .A2(n_303), .B1(n_307), .B2(n_313), .C(n_316), .Y(n_300) );
INVx1_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g337 ( .A(n_306), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_SL g383 ( .A(n_309), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_311), .B(n_361), .Y(n_360) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_311), .A2(n_379), .B(n_381), .Y(n_378) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g424 ( .A(n_312), .B(n_406), .Y(n_424) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_SL g326 ( .A(n_315), .Y(n_326) );
AOI21xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B(n_320), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_SL g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g370 ( .A(n_322), .B(n_371), .Y(n_370) );
INVxp67_ASAP7_75t_L g432 ( .A(n_322), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B(n_328), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_326), .B(n_344), .Y(n_380) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g401 ( .A(n_330), .Y(n_401) );
NAND5xp2_ASAP7_75t_L g331 ( .A(n_332), .B(n_349), .C(n_358), .D(n_378), .E(n_385), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B(n_338), .C(n_341), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g373 ( .A(n_337), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
NOR2xp33_ASAP7_75t_L g410 ( .A(n_345), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
OAI21xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_353), .B(n_355), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_350), .A2(n_404), .B1(n_407), .B2(n_409), .C(n_410), .Y(n_403) );
AND2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
AOI321xp33_ASAP7_75t_L g358 ( .A1(n_351), .A2(n_359), .A3(n_363), .B1(n_364), .B2(n_370), .C(n_372), .Y(n_358) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g429 ( .A(n_363), .Y(n_429) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_369), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g381 ( .A(n_366), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
NOR2xp67_ASAP7_75t_SL g393 ( .A(n_367), .B(n_374), .Y(n_393) );
AOI321xp33_ASAP7_75t_SL g425 ( .A1(n_370), .A2(n_426), .A3(n_427), .B1(n_428), .B2(n_429), .C(n_430), .Y(n_425) );
O2A1O1Ixp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_374), .B(n_375), .C(n_376), .Y(n_372) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_383), .B(n_391), .Y(n_420) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND3xp33_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .C(n_395), .Y(n_392) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_421), .C(n_433), .Y(n_396) );
OAI211xp5_ASAP7_75t_SL g397 ( .A1(n_398), .A2(n_399), .B(n_403), .C(n_413), .Y(n_397) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_SL g400 ( .A(n_401), .B(n_402), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_402), .A2(n_434), .B1(n_435), .B2(n_436), .C(n_437), .Y(n_433) );
INVx1_ASAP7_75t_L g422 ( .A(n_404), .Y(n_422) );
INVx1_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_SL g426 ( .A(n_424), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
CKINVDCx14_ASAP7_75t_R g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_445), .Y(n_451) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_446), .B(n_462), .Y(n_749) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g461 ( .A(n_447), .B(n_462), .Y(n_461) );
AOI21xp33_ASAP7_75t_L g452 ( .A1(n_449), .A2(n_453), .B(n_750), .Y(n_452) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_455), .A2(n_458), .B1(n_459), .B2(n_463), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx2_ASAP7_75t_L g745 ( .A(n_460), .Y(n_745) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g744 ( .A(n_463), .Y(n_744) );
OR4x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_633), .C(n_680), .D(n_720), .Y(n_463) );
NAND3xp33_ASAP7_75t_SL g464 ( .A(n_465), .B(n_579), .C(n_608), .Y(n_464) );
AOI211xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_501), .B(n_536), .C(n_572), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_L g608 ( .A1(n_466), .A2(n_592), .B(n_609), .C(n_613), .Y(n_608) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_468), .B(n_477), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_468), .B(n_571), .Y(n_570) );
INVx3_ASAP7_75t_SL g575 ( .A(n_468), .Y(n_575) );
HB1xp67_ASAP7_75t_L g587 ( .A(n_468), .Y(n_587) );
AND2x4_ASAP7_75t_L g591 ( .A(n_468), .B(n_543), .Y(n_591) );
AND2x2_ASAP7_75t_L g602 ( .A(n_468), .B(n_491), .Y(n_602) );
OR2x2_ASAP7_75t_L g626 ( .A(n_468), .B(n_539), .Y(n_626) );
AND2x2_ASAP7_75t_L g639 ( .A(n_468), .B(n_544), .Y(n_639) );
AND2x2_ASAP7_75t_L g679 ( .A(n_468), .B(n_665), .Y(n_679) );
AND2x2_ASAP7_75t_L g686 ( .A(n_468), .B(n_649), .Y(n_686) );
AND2x2_ASAP7_75t_L g716 ( .A(n_468), .B(n_478), .Y(n_716) );
OR2x6_ASAP7_75t_L g468 ( .A(n_469), .B(n_475), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_477), .B(n_643), .Y(n_655) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_490), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_478), .B(n_586), .Y(n_585) );
OR2x2_ASAP7_75t_L g593 ( .A(n_478), .B(n_490), .Y(n_593) );
BUFx3_ASAP7_75t_L g601 ( .A(n_478), .Y(n_601) );
OR2x2_ASAP7_75t_L g622 ( .A(n_478), .B(n_504), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_478), .B(n_643), .Y(n_733) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_482), .B(n_489), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_480), .A2(n_540), .B(n_541), .Y(n_539) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g540 ( .A(n_482), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_489), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_490), .B(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g586 ( .A(n_490), .Y(n_586) );
AND2x2_ASAP7_75t_L g649 ( .A(n_490), .B(n_544), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_490), .A2(n_652), .B1(n_654), .B2(n_656), .C(n_657), .Y(n_651) );
AND2x2_ASAP7_75t_L g665 ( .A(n_490), .B(n_539), .Y(n_665) );
AND2x2_ASAP7_75t_L g691 ( .A(n_490), .B(n_575), .Y(n_691) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g571 ( .A(n_491), .B(n_544), .Y(n_571) );
BUFx2_ASAP7_75t_L g705 ( .A(n_491), .Y(n_705) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI32xp33_ASAP7_75t_L g671 ( .A1(n_502), .A2(n_632), .A3(n_646), .B1(n_672), .B2(n_673), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_514), .Y(n_502) );
AND2x2_ASAP7_75t_L g612 ( .A(n_503), .B(n_556), .Y(n_612) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
OR2x2_ASAP7_75t_L g594 ( .A(n_504), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_504), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g666 ( .A(n_504), .B(n_556), .Y(n_666) );
AND2x2_ASAP7_75t_L g677 ( .A(n_504), .B(n_569), .Y(n_677) );
BUFx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g578 ( .A(n_505), .B(n_557), .Y(n_578) );
AND2x2_ASAP7_75t_L g582 ( .A(n_505), .B(n_557), .Y(n_582) );
AND2x2_ASAP7_75t_L g617 ( .A(n_505), .B(n_568), .Y(n_617) );
AND2x2_ASAP7_75t_L g624 ( .A(n_505), .B(n_526), .Y(n_624) );
OAI211xp5_ASAP7_75t_L g629 ( .A1(n_505), .A2(n_575), .B(n_586), .C(n_630), .Y(n_629) );
INVx2_ASAP7_75t_L g683 ( .A(n_505), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_505), .B(n_516), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_514), .B(n_566), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_514), .B(n_582), .Y(n_672) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g577 ( .A(n_515), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .Y(n_515) );
AND2x2_ASAP7_75t_L g569 ( .A(n_516), .B(n_527), .Y(n_569) );
OR2x2_ASAP7_75t_L g584 ( .A(n_516), .B(n_527), .Y(n_584) );
AND2x2_ASAP7_75t_L g607 ( .A(n_516), .B(n_568), .Y(n_607) );
INVx1_ASAP7_75t_L g611 ( .A(n_516), .Y(n_611) );
AND2x2_ASAP7_75t_L g630 ( .A(n_516), .B(n_567), .Y(n_630) );
OAI22xp33_ASAP7_75t_L g640 ( .A1(n_516), .A2(n_595), .B1(n_641), .B2(n_642), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_516), .B(n_683), .Y(n_707) );
AND2x2_ASAP7_75t_L g722 ( .A(n_516), .B(n_582), .Y(n_722) );
INVx4_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx3_ASAP7_75t_L g554 ( .A(n_517), .Y(n_554) );
AND2x2_ASAP7_75t_L g596 ( .A(n_517), .B(n_527), .Y(n_596) );
AND2x2_ASAP7_75t_L g598 ( .A(n_517), .B(n_556), .Y(n_598) );
AND3x2_ASAP7_75t_L g660 ( .A(n_517), .B(n_624), .C(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g695 ( .A(n_526), .B(n_567), .Y(n_695) );
INVx1_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g556 ( .A(n_527), .B(n_557), .Y(n_556) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_527), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_527), .B(n_566), .Y(n_628) );
NAND3xp33_ASAP7_75t_L g735 ( .A(n_527), .B(n_607), .C(n_683), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_553), .B1(n_565), .B2(n_570), .Y(n_536) );
INVx1_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_542), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_539), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_SL g647 ( .A(n_539), .Y(n_647) );
OAI31xp33_ASAP7_75t_L g663 ( .A1(n_542), .A2(n_664), .A3(n_665), .B(n_666), .Y(n_663) );
AND2x2_ASAP7_75t_L g688 ( .A(n_542), .B(n_575), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_542), .B(n_601), .Y(n_734) );
AND2x2_ASAP7_75t_L g643 ( .A(n_543), .B(n_575), .Y(n_643) );
AND2x2_ASAP7_75t_L g704 ( .A(n_543), .B(n_705), .Y(n_704) );
INVx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g574 ( .A(n_544), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g632 ( .A(n_544), .Y(n_632) );
OR2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
CKINVDCx16_ASAP7_75t_R g653 ( .A(n_554), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_555), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
AOI221x1_ASAP7_75t_SL g620 ( .A1(n_556), .A2(n_621), .B1(n_623), .B2(n_625), .C(n_627), .Y(n_620) );
INVx2_ASAP7_75t_L g568 ( .A(n_557), .Y(n_568) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_557), .Y(n_662) );
INVx1_ASAP7_75t_L g650 ( .A(n_565), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_569), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_566), .B(n_583), .Y(n_675) );
INVx1_ASAP7_75t_SL g738 ( .A(n_566), .Y(n_738) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g656 ( .A(n_569), .B(n_582), .Y(n_656) );
INVx1_ASAP7_75t_L g724 ( .A(n_570), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_570), .B(n_653), .Y(n_737) );
INVx2_ASAP7_75t_SL g576 ( .A(n_571), .Y(n_576) );
AND2x2_ASAP7_75t_L g619 ( .A(n_571), .B(n_575), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_571), .B(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_571), .B(n_646), .Y(n_673) );
AOI21xp33_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_576), .B(n_577), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_574), .B(n_646), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_574), .B(n_601), .Y(n_742) );
OR2x2_ASAP7_75t_L g614 ( .A(n_575), .B(n_593), .Y(n_614) );
AND2x2_ASAP7_75t_L g713 ( .A(n_575), .B(n_704), .Y(n_713) );
OAI22xp5_ASAP7_75t_SL g588 ( .A1(n_576), .A2(n_589), .B1(n_594), .B2(n_597), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_576), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g636 ( .A(n_578), .B(n_584), .Y(n_636) );
INVx1_ASAP7_75t_L g700 ( .A(n_578), .Y(n_700) );
AOI311xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_585), .A3(n_587), .B(n_588), .C(n_599), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_583), .A2(n_715), .B1(n_727), .B2(n_730), .C(n_732), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_583), .B(n_738), .Y(n_740) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g637 ( .A(n_585), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g627 ( .A1(n_586), .A2(n_628), .B(n_629), .C(n_631), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_592), .Y(n_589) );
O2A1O1Ixp33_ASAP7_75t_SL g696 ( .A1(n_590), .A2(n_592), .B(n_697), .C(n_698), .Y(n_696) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_591), .B(n_665), .Y(n_731) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g613 ( .A1(n_594), .A2(n_614), .B1(n_615), .B2(n_618), .C(n_620), .Y(n_613) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g616 ( .A(n_596), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g699 ( .A(n_596), .B(n_700), .Y(n_699) );
INVx1_ASAP7_75t_SL g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_600), .B(n_603), .Y(n_599) );
A2O1A1Ixp33_ASAP7_75t_L g657 ( .A1(n_600), .A2(n_658), .B(n_659), .C(n_663), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_601), .B(n_602), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_601), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_601), .B(n_704), .Y(n_703) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AND2x2_ASAP7_75t_L g623 ( .A(n_607), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_611), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g725 ( .A(n_614), .Y(n_725) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_617), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g652 ( .A(n_617), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g729 ( .A(n_617), .Y(n_729) );
INVx1_ASAP7_75t_SL g618 ( .A(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g670 ( .A(n_619), .B(n_646), .Y(n_670) );
INVx1_ASAP7_75t_SL g664 ( .A(n_626), .Y(n_664) );
INVx1_ASAP7_75t_L g641 ( .A(n_632), .Y(n_641) );
NAND3xp33_ASAP7_75t_SL g633 ( .A(n_634), .B(n_651), .C(n_667), .Y(n_633) );
AOI322xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_637), .A3(n_638), .B1(n_640), .B2(n_644), .C1(n_648), .C2(n_650), .Y(n_634) );
AOI211xp5_ASAP7_75t_L g687 ( .A1(n_635), .A2(n_688), .B(n_689), .C(n_696), .Y(n_687) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g689 ( .A1(n_638), .A2(n_659), .B1(n_690), .B2(n_692), .Y(n_689) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
AND2x2_ASAP7_75t_L g648 ( .A(n_646), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g685 ( .A(n_646), .B(n_686), .Y(n_685) );
AOI32xp33_ASAP7_75t_L g736 ( .A1(n_646), .A2(n_737), .A3(n_738), .B1(n_739), .B2(n_741), .Y(n_736) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g658 ( .A(n_649), .Y(n_658) );
AOI221xp5_ASAP7_75t_L g701 ( .A1(n_649), .A2(n_702), .B1(n_706), .B2(n_708), .C(n_711), .Y(n_701) );
AND2x2_ASAP7_75t_L g715 ( .A(n_649), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_L g718 ( .A(n_653), .B(n_719), .Y(n_718) );
OR2x2_ASAP7_75t_L g728 ( .A(n_653), .B(n_729), .Y(n_728) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AND2x2_ASAP7_75t_L g719 ( .A(n_662), .B(n_683), .Y(n_719) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B(n_671), .C(n_674), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI211xp5_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_684), .B(n_687), .C(n_701), .Y(n_680) );
INVxp67_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_695), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g710 ( .A(n_707), .Y(n_710) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B(n_717), .Y(n_711) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
OAI211xp5_ASAP7_75t_SL g720 ( .A1(n_721), .A2(n_723), .B(n_726), .C(n_736), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AOI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_735), .Y(n_732) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
endmodule