module fake_jpeg_3622_n_68 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_68);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_68;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_5),
.B(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_24),
.B(n_0),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_24),
.B(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_23),
.Y(n_29)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_29),
.A2(n_33),
.B(n_28),
.Y(n_37)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_22),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_26),
.B1(n_27),
.B2(n_33),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_30),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_31),
.A2(n_22),
.B1(n_20),
.B2(n_19),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_42),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_3),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_40),
.B1(n_7),
.B2(n_8),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_40),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_6),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_18),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_13),
.B1(n_17),
.B2(n_16),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_51),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_41),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_54),
.C(n_58),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_11),
.C(n_15),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_8),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_6),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_47),
.C(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_62),
.Y(n_64)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_63),
.A2(n_59),
.B(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_66),
.A2(n_64),
.B(n_63),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_9),
.Y(n_68)
);


endmodule