module fake_jpeg_3089_n_231 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_231);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_231;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_16),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_16),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_23),
.B(n_50),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_3),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_19),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_34),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_0),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_72),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_55),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_84),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_1),
.Y(n_84)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_77),
.B1(n_60),
.B2(n_56),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_SL g110 ( 
.A1(n_91),
.A2(n_99),
.B(n_93),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_85),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_79),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_83),
.A2(n_77),
.B1(n_56),
.B2(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_105),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_117),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_82),
.B1(n_63),
.B2(n_75),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_108),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_81),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_107),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_52),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_93),
.A2(n_82),
.B1(n_63),
.B2(n_75),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_110),
.A2(n_114),
.B1(n_119),
.B2(n_78),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_111),
.B(n_115),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_54),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_112),
.B(n_113),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_82),
.C(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_114),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_97),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_87),
.B(n_57),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_65),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_119),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_96),
.B1(n_95),
.B2(n_86),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_128),
.B1(n_61),
.B2(n_53),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_114),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_79),
.Y(n_146)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_125),
.A2(n_141),
.B(n_127),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_35),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_130),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_113),
.B1(n_103),
.B2(n_109),
.Y(n_128)
);

AND2x6_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_36),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_109),
.B(n_73),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_131),
.B(n_139),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_33),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_51),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_96),
.B1(n_70),
.B2(n_76),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_133),
.A2(n_74),
.B1(n_64),
.B2(n_59),
.Y(n_151)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

INVx13_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_116),
.Y(n_139)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_136),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_156),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_146),
.A2(n_147),
.B(n_150),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_73),
.B(n_69),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g148 ( 
.A1(n_123),
.A2(n_96),
.B1(n_76),
.B2(n_57),
.Y(n_148)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_66),
.B(n_68),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_153),
.B1(n_160),
.B2(n_164),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_129),
.A2(n_71),
.B(n_78),
.C(n_67),
.Y(n_152)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_26),
.B(n_14),
.C(n_15),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_129),
.A2(n_74),
.B1(n_64),
.B2(n_67),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_154),
.B(n_158),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_61),
.B(n_53),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_155),
.A2(n_162),
.B(n_166),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_62),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_1),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_159),
.B(n_2),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_128),
.B1(n_141),
.B2(n_140),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_42),
.B(n_49),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_166),
.B1(n_138),
.B2(n_3),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_71),
.B1(n_47),
.B2(n_45),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_39),
.B1(n_38),
.B2(n_37),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_181),
.B(n_183),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_172),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_2),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_173),
.B(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_142),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_27),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_165),
.A2(n_4),
.B(n_5),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_155),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_152),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_27),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_25),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_149),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_164),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_186)
);

AOI221xp5_ASAP7_75t_L g190 ( 
.A1(n_187),
.A2(n_162),
.B1(n_152),
.B2(n_148),
.C(n_151),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_13),
.B1(n_15),
.B2(n_17),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_18),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_191),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g191 ( 
.A1(n_167),
.A2(n_152),
.B(n_148),
.C(n_143),
.D(n_20),
.Y(n_191)
);

AO22x1_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_178),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_198),
.B(n_199),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_170),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_201),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_196),
.A2(n_178),
.B1(n_188),
.B2(n_183),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_202),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_167),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_204),
.C(n_209),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_173),
.C(n_184),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_20),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_197),
.B(n_176),
.C(n_169),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_203),
.B(n_189),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_213),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_195),
.A3(n_191),
.B1(n_192),
.B2(n_190),
.C1(n_194),
.C2(n_187),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_206),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_215),
.A2(n_211),
.B1(n_205),
.B2(n_23),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_209),
.B(n_202),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_217),
.C(n_216),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_221),
.A2(n_217),
.B1(n_212),
.B2(n_204),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_224),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_222),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_220),
.C(n_221),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_227),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_219),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_21),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_230),
.A2(n_21),
.B(n_22),
.Y(n_231)
);


endmodule