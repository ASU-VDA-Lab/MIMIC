module fake_jpeg_595_n_373 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_373);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_373;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_44),
.Y(n_113)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_SL g115 ( 
.A(n_46),
.Y(n_115)
);

INVx11_ASAP7_75t_SL g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_47),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_21),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_49),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_50),
.Y(n_140)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_51),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_34),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_52),
.B(n_53),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_54),
.Y(n_102)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_59),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_17),
.B(n_6),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_74),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_20),
.B(n_6),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_60),
.B(n_65),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_21),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_67),
.B(n_80),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_69),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_24),
.B(n_7),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_15),
.Y(n_77)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_78),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_24),
.B(n_12),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_86),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_22),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_81),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_82),
.Y(n_128)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_85),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_26),
.B(n_11),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_8),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_88),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_30),
.B(n_9),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_90),
.B(n_92),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_30),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_37),
.B(n_0),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_37),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_94),
.Y(n_148)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_95),
.B(n_23),
.Y(n_106)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_96),
.B(n_97),
.Y(n_129)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_38),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_87),
.A2(n_43),
.B1(n_32),
.B2(n_28),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_105),
.A2(n_108),
.B1(n_139),
.B2(n_151),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_106),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_46),
.A2(n_43),
.B1(n_19),
.B2(n_28),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_45),
.B(n_32),
.C(n_19),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_120),
.B(n_121),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_60),
.B(n_78),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_56),
.A2(n_77),
.B1(n_89),
.B2(n_73),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_135),
.B1(n_51),
.B2(n_95),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_54),
.B(n_0),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_131),
.B(n_136),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_63),
.A2(n_35),
.B1(n_42),
.B2(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_47),
.B(n_66),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_64),
.A2(n_35),
.B1(n_42),
.B2(n_2),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_55),
.B(n_0),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_152),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_50),
.A2(n_75),
.B1(n_62),
.B2(n_61),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_61),
.B(n_1),
.Y(n_152)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_154),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_44),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_166),
.Y(n_209)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_157),
.Y(n_212)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_158),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_159),
.Y(n_203)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_164),
.Y(n_206)
);

INVx11_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_161),
.Y(n_213)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_163),
.Y(n_218)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_149),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_106),
.A2(n_130),
.B1(n_124),
.B2(n_110),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_165),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_112),
.B(n_94),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_167),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_168),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_170),
.B(n_175),
.Y(n_207)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_171),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_103),
.Y(n_173)
);

INVx11_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_85),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_176),
.B(n_179),
.Y(n_210)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_109),
.Y(n_179)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_100),
.B(n_82),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_186),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_183),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_122),
.A2(n_71),
.B1(n_68),
.B2(n_76),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_184),
.A2(n_193),
.B1(n_151),
.B2(n_140),
.Y(n_223)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_1),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_189),
.C(n_190),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_111),
.B(n_72),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_3),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_145),
.B(n_3),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_115),
.B(n_81),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_191),
.Y(n_211)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_128),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_122),
.A2(n_70),
.B1(n_83),
.B2(n_88),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_162),
.A2(n_132),
.B1(n_138),
.B2(n_113),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_194),
.A2(n_200),
.B1(n_156),
.B2(n_140),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_178),
.A2(n_108),
.B1(n_132),
.B2(n_113),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_199),
.A2(n_204),
.B1(n_172),
.B2(n_115),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_155),
.A2(n_116),
.B1(n_126),
.B2(n_146),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_193),
.B1(n_153),
.B2(n_176),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_126),
.B1(n_104),
.B2(n_150),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_202),
.B(n_153),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_237),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_156),
.C(n_167),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_230),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_227),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_187),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_235),
.Y(n_263)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_222),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_229),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_185),
.C(n_157),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_190),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_234),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_232),
.A2(n_203),
.B1(n_223),
.B2(n_194),
.Y(n_247)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_195),
.Y(n_233)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_211),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_204),
.B(n_192),
.Y(n_235)
);

NOR2x1_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_163),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_240),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_211),
.B(n_183),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_171),
.C(n_123),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_242),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_199),
.A2(n_177),
.B1(n_182),
.B2(n_168),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_239),
.A2(n_197),
.B1(n_215),
.B2(n_196),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_180),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_245),
.B1(n_213),
.B2(n_197),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_158),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_114),
.C(n_144),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_164),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_246),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_248),
.B1(n_228),
.B2(n_230),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_235),
.B1(n_240),
.B2(n_239),
.Y(n_248)
);

OAI22x1_ASAP7_75t_L g252 ( 
.A1(n_245),
.A2(n_206),
.B1(n_221),
.B2(n_101),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_252),
.Y(n_280)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_255),
.Y(n_274)
);

AO22x1_ASAP7_75t_L g258 ( 
.A1(n_226),
.A2(n_195),
.B1(n_219),
.B2(n_206),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_259),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_261),
.B(n_264),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_SL g265 ( 
.A1(n_236),
.A2(n_213),
.B(n_196),
.C(n_215),
.Y(n_265)
);

AO21x1_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_218),
.B(n_246),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_233),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_219),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_286),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_267),
.C(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_277),
.C(n_259),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_225),
.B(n_238),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_282),
.B(n_258),
.Y(n_294)
);

NAND3xp33_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_207),
.C(n_227),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_272),
.B(n_285),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_207),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_250),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_254),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_278),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_256),
.C(n_262),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_254),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_249),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_249),
.Y(n_283)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_283),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_250),
.B(n_217),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_248),
.A2(n_229),
.B1(n_243),
.B2(n_205),
.Y(n_286)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_256),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_288),
.A2(n_281),
.B1(n_274),
.B2(n_273),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_291),
.B(n_292),
.C(n_300),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_263),
.C(n_247),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_294),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_280),
.A2(n_255),
.B1(n_253),
.B2(n_266),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_297),
.A2(n_276),
.B1(n_278),
.B2(n_282),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_301),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_205),
.C(n_252),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_258),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_304),
.B(n_279),
.C(n_283),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_275),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_306),
.C(n_307),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_273),
.B(n_198),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_274),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_290),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_310),
.B(n_315),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_208),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_312),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_286),
.B1(n_282),
.B2(n_287),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_313),
.A2(n_309),
.B1(n_319),
.B2(n_293),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_291),
.B(n_257),
.C(n_253),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_292),
.C(n_300),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_265),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_319),
.Y(n_329)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_295),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_321),
.Y(n_325)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_298),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_309),
.A2(n_296),
.B(n_307),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_315),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_322),
.C(n_314),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_328),
.A2(n_305),
.B1(n_322),
.B2(n_314),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_308),
.Y(n_330)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_330),
.Y(n_335)
);

A2O1A1Ixp33_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_293),
.B(n_304),
.C(n_265),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_313),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_317),
.Y(n_334)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_334),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_336),
.B(n_340),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_339),
.Y(n_348)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_332),
.B(n_316),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_342),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_333),
.B(n_299),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_344),
.A2(n_323),
.B1(n_328),
.B2(n_331),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_338),
.A2(n_334),
.B(n_330),
.Y(n_345)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_345),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_336),
.A2(n_326),
.B(n_327),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_208),
.C(n_265),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_344),
.A2(n_323),
.B(n_329),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_351),
.A2(n_217),
.B(n_219),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_335),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_346),
.B(n_343),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_354),
.B(n_357),
.Y(n_364)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_356),
.A2(n_359),
.B(n_349),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_347),
.B(n_221),
.C(n_198),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_349),
.A2(n_265),
.B1(n_161),
.B2(n_174),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_358),
.B(n_353),
.Y(n_361)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_360),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_212),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_358),
.B(n_348),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_363),
.A2(n_212),
.B(n_154),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_365),
.B(n_125),
.Y(n_369)
);

OAI321xp33_ASAP7_75t_L g368 ( 
.A1(n_366),
.A2(n_364),
.A3(n_362),
.B1(n_101),
.B2(n_102),
.C(n_125),
.Y(n_368)
);

OA21x2_ASAP7_75t_SL g370 ( 
.A1(n_368),
.A2(n_369),
.B(n_367),
.Y(n_370)
);

AOI321xp33_ASAP7_75t_L g371 ( 
.A1(n_370),
.A2(n_88),
.A3(n_146),
.B1(n_70),
.B2(n_142),
.C(n_3),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g372 ( 
.A1(n_371),
.A2(n_3),
.B(n_4),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_372),
.B(n_4),
.Y(n_373)
);


endmodule