module fake_jpeg_328_n_168 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_168);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_168;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx2_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx14_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_31),
.B(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_33),
.Y(n_86)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_37),
.Y(n_80)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_45),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_44),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_0),
.C(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_1),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_53),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_15),
.B(n_2),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_30),
.Y(n_59)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_13),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_10),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_29),
.C(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_57),
.B(n_59),
.Y(n_101)
);

AO22x2_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_29),
.B1(n_28),
.B2(n_23),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_64),
.B1(n_86),
.B2(n_81),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_20),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_61),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_20),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_62),
.B(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_38),
.A2(n_26),
.B1(n_21),
.B2(n_30),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_87),
.B1(n_67),
.B2(n_81),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_40),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_41),
.A2(n_16),
.B1(n_23),
.B2(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_73),
.A2(n_74),
.B1(n_85),
.B2(n_86),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_43),
.A2(n_21),
.B1(n_27),
.B2(n_7),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_78),
.B(n_79),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_10),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_43),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_4),
.B1(n_5),
.B2(n_44),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_75),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_90),
.Y(n_118)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_91),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_33),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_105),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_60),
.A2(n_44),
.B1(n_33),
.B2(n_5),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_96),
.B1(n_107),
.B2(n_64),
.Y(n_109)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_61),
.A2(n_70),
.B1(n_80),
.B2(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_102),
.Y(n_124)
);

OAI21x1_ASAP7_75t_R g111 ( 
.A1(n_98),
.A2(n_75),
.B(n_58),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_69),
.B1(n_80),
.B2(n_83),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_108),
.B1(n_95),
.B2(n_102),
.Y(n_122)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_103),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_57),
.B(n_77),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_106),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_58),
.B(n_76),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_65),
.A2(n_76),
.B1(n_66),
.B2(n_58),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_122),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_75),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_123),
.C(n_97),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_104),
.B(n_68),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_97),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_106),
.A2(n_65),
.B(n_66),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_91),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_88),
.A2(n_90),
.B(n_97),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_101),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_125),
.B(n_101),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_126),
.A2(n_128),
.B(n_130),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_96),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_129),
.B(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_123),
.C(n_124),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_120),
.B(n_103),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_134),
.B(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_112),
.B(n_107),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_135),
.A2(n_109),
.B1(n_119),
.B2(n_110),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_142),
.C(n_146),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_141),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g141 ( 
.A1(n_131),
.A2(n_111),
.B(n_118),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_116),
.C(n_117),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_130),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_114),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_117),
.C(n_115),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_131),
.B(n_136),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_149),
.A2(n_151),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_150),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_144),
.A2(n_111),
.B(n_136),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_128),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_139),
.C(n_141),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_156),
.C(n_121),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_155),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_127),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_157),
.A2(n_150),
.B(n_121),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_159),
.B(n_161),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_156),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_99),
.B(n_113),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_153),
.Y(n_162)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_162),
.B(n_164),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_165),
.A2(n_100),
.B(n_113),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_167),
.B(n_166),
.Y(n_168)
);


endmodule