module real_jpeg_24110_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_1),
.A2(n_35),
.B1(n_64),
.B2(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_1),
.A2(n_35),
.B1(n_59),
.B2(n_170),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_3),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_3),
.B(n_63),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g230 ( 
.A1(n_3),
.A2(n_67),
.B(n_83),
.C(n_231),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_3),
.A2(n_64),
.B1(n_67),
.B2(n_171),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_3),
.B(n_28),
.C(n_45),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_3),
.A2(n_40),
.B1(n_42),
.B2(n_171),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_3),
.A2(n_25),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_3),
.B(n_125),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_61),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_61),
.Y(n_191)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_60),
.B1(n_72),
.B2(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_7),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_7),
.A2(n_64),
.B1(n_67),
.B2(n_110),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_110),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_110),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_10),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_40),
.B1(n_42),
.B2(n_74),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_10),
.A2(n_64),
.B1(n_67),
.B2(n_74),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_74),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_11),
.A2(n_50),
.B1(n_64),
.B2(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_11),
.A2(n_50),
.B1(n_57),
.B2(n_60),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_12),
.A2(n_64),
.B1(n_67),
.B2(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_12),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_40),
.B1(n_42),
.B2(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_12),
.A2(n_60),
.B1(n_87),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_87),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_13),
.A2(n_64),
.B1(n_67),
.B2(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_13),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_161),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_13),
.A2(n_40),
.B1(n_42),
.B2(n_161),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_161),
.Y(n_258)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_39),
.B1(n_64),
.B2(n_67),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_15),
.A2(n_39),
.B1(n_72),
.B2(n_73),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_179)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_16),
.A2(n_26),
.B1(n_177),
.B2(n_179),
.Y(n_176)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_16),
.Y(n_194)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_16),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_16),
.A2(n_26),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_347),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_334),
.B(n_346),
.Y(n_18)
);

OAI31xp33_ASAP7_75t_SL g19 ( 
.A1(n_20),
.A2(n_136),
.A3(n_150),
.B(n_331),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_21),
.B(n_114),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.C(n_94),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_22),
.A2(n_78),
.B1(n_79),
.B2(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_22),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_24),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_25),
.A2(n_34),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_25),
.A2(n_178),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_25),
.A2(n_31),
.B1(n_99),
.B2(n_208),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_25),
.A2(n_260),
.B(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_26),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_27),
.B(n_264),
.Y(n_263)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_32),
.B(n_171),
.Y(n_264)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_38),
.A2(n_43),
.B1(n_51),
.B2(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_42),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_40),
.B(n_252),
.Y(n_251)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_42),
.A2(n_84),
.B(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_43),
.A2(n_51),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_43),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_43),
.A2(n_51),
.B1(n_226),
.B2(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_48),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_48),
.A2(n_90),
.B1(n_104),
.B2(n_165),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_48),
.B(n_171),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_48),
.A2(n_166),
.B(n_241),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_51),
.B(n_167),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_69),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_56),
.A2(n_62),
.B1(n_111),
.B2(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_57),
.Y(n_170)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_SL g182 ( 
.A(n_58),
.B(n_66),
.C(n_67),
.Y(n_182)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_71),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_62),
.A2(n_111),
.B1(n_133),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_62),
.A2(n_69),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_63),
.A2(n_76),
.B1(n_109),
.B2(n_203),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_63),
.A2(n_76),
.B1(n_341),
.B2(n_342),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_63),
.A2(n_76),
.B1(n_342),
.B2(n_351),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_67),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_64),
.A2(n_68),
.B(n_172),
.C(n_182),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_68),
.B1(n_72),
.B2(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_73),
.B(n_171),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_76),
.A2(n_113),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_89),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_88),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_81),
.A2(n_82),
.B1(n_127),
.B2(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_81),
.A2(n_199),
.B(n_200),
.Y(n_198)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_81),
.A2(n_200),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_82),
.A2(n_185),
.B(n_186),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_82),
.A2(n_106),
.B(n_186),
.Y(n_310)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_90),
.A2(n_225),
.B(n_227),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_90),
.A2(n_227),
.B(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_94),
.A2(n_95),
.B1(n_326),
.B2(n_328),
.Y(n_325)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.C(n_107),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_96),
.A2(n_97),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_98),
.Y(n_303)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_100),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_100),
.A2(n_234),
.B(n_258),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_105),
.B(n_107),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_112),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_117),
.C(n_119),
.Y(n_149)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_135),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_122),
.B(n_129),
.C(n_132),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_125),
.B1(n_160),
.B2(n_162),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_124),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_124),
.A2(n_125),
.B(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_125),
.B(n_187),
.Y(n_200)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_129),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_129),
.B(n_143),
.C(n_147),
.Y(n_345)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_132),
.A2(n_135),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_132),
.B(n_139),
.C(n_142),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_137),
.A2(n_332),
.B(n_333),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_149),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_138),
.B(n_149),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_144),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_148),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_324),
.B(n_330),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_314),
.B(n_323),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_212),
.B(n_297),
.C(n_313),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_195),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_154),
.B(n_195),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_173),
.C(n_183),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_155),
.A2(n_156),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_168),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_163),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_163),
.C(n_168),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_171),
.B(n_172),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_173),
.A2(n_174),
.B1(n_183),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_180),
.B2(n_181),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_180),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_183),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_188),
.C(n_190),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_220),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_221),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_191),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_204),
.B1(n_205),
.B2(n_211),
.Y(n_195)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_196),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.CI(n_201),
.CON(n_196),
.SN(n_196)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_197),
.B(n_198),
.C(n_201),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_210),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_207),
.B(n_209),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_290),
.B(n_296),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_245),
.B(n_289),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_237),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_217),
.B(n_237),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_236),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_218),
.B(n_224),
.C(n_228),
.Y(n_295)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_230),
.B(n_232),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_267),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.C(n_242),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_285),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_239),
.A2(n_242),
.B1(n_243),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_283),
.B(n_288),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_273),
.B(n_282),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_261),
.B(n_272),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_256),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_268),
.B(n_271),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_265),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_269),
.B(n_270),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_281),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_274),
.B(n_281),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_280),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_278),
.B2(n_279),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_279),
.C(n_280),
.Y(n_287)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_287),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_295),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_312),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_312),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_302),
.C(n_304),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_309),
.C(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_316),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_318),
.B(n_319),
.C(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_329),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_329),
.Y(n_330)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_326),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_335),
.B(n_336),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_345),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_340),
.B1(n_343),
.B2(n_344),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_338),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_340),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_343),
.C(n_345),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_352),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_350),
.B(n_352),
.Y(n_353)
);


endmodule