module fake_jpeg_19102_n_86 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_86);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_86;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx11_ASAP7_75t_SL g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx14_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

BUFx10_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_18),
.B(n_0),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_15),
.B(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_25),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_10),
.Y(n_36)
);

OAI32xp33_ASAP7_75t_L g35 ( 
.A1(n_28),
.A2(n_23),
.A3(n_9),
.B1(n_17),
.B2(n_10),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_11),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_11),
.B(n_12),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_25),
.C(n_20),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_39),
.C(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_17),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_27),
.B(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_16),
.Y(n_46)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_30),
.B1(n_13),
.B2(n_20),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_47),
.A2(n_56),
.B1(n_39),
.B2(n_42),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_37),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_59),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_60),
.B(n_61),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_52),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_65),
.C(n_53),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_1),
.B(n_2),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_40),
.C(n_11),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_55),
.C(n_53),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_71),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_65),
.C(n_62),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_61),
.A2(n_48),
.B(n_47),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_75),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_74),
.C(n_64),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_57),
.C(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_77),
.B(n_78),
.Y(n_80)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_79),
.B(n_76),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_82),
.A2(n_83),
.B(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_78),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_3),
.B(n_7),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_85),
.B(n_11),
.Y(n_86)
);


endmodule