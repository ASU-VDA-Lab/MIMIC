module fake_jpeg_11860_n_579 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_579);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_579;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_12),
.B(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx3_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_33),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_55),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_57),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_58),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_59),
.Y(n_168)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_63),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_35),
.B(n_17),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_64),
.B(n_87),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_65),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_71),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_67),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_68),
.Y(n_111)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_53),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_89),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_78),
.Y(n_164)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_80),
.Y(n_169)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_53),
.Y(n_82)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_84),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_30),
.B1(n_39),
.B2(n_37),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_86),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_0),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_34),
.B(n_44),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_103),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_53),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_26),
.B(n_0),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_27),
.B(n_0),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_107),
.Y(n_150)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_27),
.Y(n_93)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx11_ASAP7_75t_L g132 ( 
.A(n_95),
.Y(n_132)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_27),
.Y(n_96)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_96),
.Y(n_158)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_44),
.Y(n_97)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_97),
.Y(n_170)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_32),
.Y(n_99)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_52),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_46),
.B(n_1),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_46),
.Y(n_104)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_105),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

INVx4_ASAP7_75t_SL g151 ( 
.A(n_106),
.Y(n_151)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_108),
.Y(n_156)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_109),
.Y(n_176)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_27),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_123),
.A2(n_50),
.B1(n_37),
.B2(n_36),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_26),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_131),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_82),
.A2(n_30),
.B1(n_43),
.B2(n_27),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_129),
.A2(n_79),
.B1(n_84),
.B2(n_60),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_92),
.B(n_48),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_130),
.B(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_48),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_98),
.B(n_25),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_147),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_57),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_92),
.B(n_48),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_162),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_103),
.B(n_25),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_88),
.B(n_40),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_152),
.B(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_63),
.B(n_40),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_61),
.B(n_41),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_161),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_72),
.B(n_97),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_63),
.B(n_42),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_68),
.B(n_41),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_167),
.B(n_172),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_68),
.B(n_19),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_175),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_76),
.B(n_19),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_110),
.B(n_42),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_105),
.B1(n_57),
.B2(n_95),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_177),
.B(n_227),
.Y(n_246)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_179),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_137),
.A2(n_109),
.B1(n_78),
.B2(n_80),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_180),
.A2(n_199),
.B1(n_222),
.B2(n_233),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_107),
.B1(n_56),
.B2(n_106),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_181),
.A2(n_133),
.B1(n_146),
.B2(n_115),
.Y(n_250)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_163),
.Y(n_183)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_2),
.B(n_3),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_184),
.B(n_197),
.Y(n_282)
);

OAI22x1_ASAP7_75t_L g272 ( 
.A1(n_185),
.A2(n_196),
.B1(n_206),
.B2(n_217),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_186),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_114),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_214),
.Y(n_245)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_151),
.Y(n_188)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_188),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_189),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_113),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_191),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_112),
.B(n_96),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_192),
.Y(n_276)
);

INVx11_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_193),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_127),
.A2(n_55),
.B1(n_43),
.B2(n_104),
.Y(n_196)
);

AND2x4_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_69),
.Y(n_197)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_166),
.Y(n_198)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_198),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_138),
.A2(n_67),
.B1(n_100),
.B2(n_99),
.Y(n_199)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_200),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_149),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_SL g253 ( 
.A(n_203),
.B(n_226),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_154),
.Y(n_204)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_204),
.Y(n_294)
);

OR2x2_ASAP7_75t_SL g205 ( 
.A(n_121),
.B(n_70),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_205),
.A2(n_168),
.B(n_158),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_127),
.A2(n_93),
.B1(n_22),
.B2(n_47),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_145),
.Y(n_207)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_207),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_149),
.Y(n_208)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_209),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_142),
.Y(n_211)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_211),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_124),
.B(n_73),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_212),
.B(n_234),
.Y(n_271)
);

BUFx2_ASAP7_75t_L g213 ( 
.A(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

CKINVDCx9p33_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_134),
.B(n_65),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_215),
.B(n_218),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_216),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_118),
.B(n_62),
.Y(n_218)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_224),
.Y(n_249)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_122),
.A2(n_31),
.B(n_28),
.C(n_36),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_221),
.B(n_120),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_125),
.A2(n_94),
.B1(n_86),
.B2(n_83),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_145),
.A2(n_22),
.B1(n_28),
.B2(n_47),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_223),
.A2(n_146),
.B1(n_133),
.B2(n_136),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_148),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_228),
.Y(n_260)
);

BUFx2_ASAP7_75t_R g226 ( 
.A(n_174),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g227 ( 
.A(n_118),
.B(n_59),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_176),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_230),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_231),
.B(n_232),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_165),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_125),
.A2(n_77),
.B1(n_75),
.B2(n_58),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_119),
.B(n_45),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_119),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_237),
.Y(n_275)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_153),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_140),
.B(n_45),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_238),
.B(n_2),
.Y(n_290)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_140),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_239),
.B(n_3),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_123),
.A2(n_50),
.B1(n_39),
.B2(n_31),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_240),
.A2(n_160),
.B1(n_132),
.B2(n_108),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_241),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_129),
.B1(n_173),
.B2(n_170),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_243),
.A2(n_250),
.B1(n_262),
.B2(n_256),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_215),
.A2(n_165),
.B(n_135),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_247),
.A2(n_248),
.B(n_295),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_178),
.A2(n_135),
.B(n_126),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_197),
.B(n_236),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_252),
.B(n_268),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_227),
.A2(n_136),
.B1(n_111),
.B2(n_126),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_257),
.A2(n_265),
.B(n_286),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_181),
.A2(n_115),
.B1(n_173),
.B2(n_169),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_227),
.A2(n_111),
.B1(n_116),
.B2(n_120),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_197),
.B(n_170),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_197),
.B(n_158),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_270),
.B(n_280),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_218),
.A2(n_169),
.B1(n_153),
.B2(n_164),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g318 ( 
.A1(n_273),
.A2(n_287),
.B1(n_188),
.B2(n_182),
.Y(n_318)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_177),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_166),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_281),
.B(n_284),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_202),
.B(n_164),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_289),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_194),
.B(n_2),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_185),
.A2(n_223),
.B(n_196),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_210),
.B(n_160),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_290),
.B(n_293),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_217),
.A2(n_52),
.B1(n_4),
.B2(n_5),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_245),
.B(n_195),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_296),
.B(n_299),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_SL g386 ( 
.A1(n_297),
.A2(n_320),
.B(n_337),
.Y(n_386)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_275),
.Y(n_298)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_298),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_284),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_260),
.Y(n_300)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_300),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_201),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_301),
.B(n_313),
.Y(n_374)
);

INVx13_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

BUFx4f_ASAP7_75t_SL g387 ( 
.A(n_303),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_272),
.A2(n_186),
.B1(n_190),
.B2(n_224),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_246),
.A2(n_206),
.B1(n_177),
.B2(n_217),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_305),
.A2(n_323),
.B1(n_328),
.B2(n_329),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_279),
.Y(n_306)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_306),
.Y(n_357)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_308),
.Y(n_364)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_205),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_309),
.B(n_314),
.Y(n_360)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_242),
.Y(n_310)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_310),
.Y(n_367)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_242),
.Y(n_311)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_311),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_312),
.A2(n_342),
.B1(n_259),
.B2(n_258),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_192),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_261),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_251),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_266),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_317),
.B(n_321),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_232),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_319),
.B(n_326),
.Y(n_378)
);

INVx5_ASAP7_75t_L g321 ( 
.A(n_255),
.Y(n_321)
);

AOI21xp33_ASAP7_75t_L g322 ( 
.A1(n_248),
.A2(n_184),
.B(n_226),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_324),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_246),
.A2(n_237),
.B1(n_231),
.B2(n_225),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_249),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_292),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_325),
.B(n_339),
.Y(n_368)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_282),
.B(n_203),
.C(n_208),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_288),
.C(n_277),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_280),
.A2(n_200),
.B1(n_198),
.B2(n_191),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_268),
.A2(n_216),
.B1(n_211),
.B2(n_219),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_254),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_331),
.Y(n_358)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_282),
.A2(n_207),
.B(n_204),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_338),
.B(n_285),
.Y(n_366)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_253),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_336),
.B(n_341),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_270),
.B(n_179),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_337),
.B(n_286),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_282),
.A2(n_189),
.B(n_209),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_269),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_264),
.B(n_213),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_340),
.B(n_267),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_243),
.A2(n_193),
.B1(n_52),
.B2(n_5),
.Y(n_342)
);

INVx4_ASAP7_75t_SL g343 ( 
.A(n_285),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g385 ( 
.A(n_343),
.Y(n_385)
);

INVx13_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_344),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_274),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_346),
.A2(n_386),
.B(n_366),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_333),
.B(n_345),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_350),
.B(n_375),
.C(n_376),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_305),
.A2(n_250),
.B1(n_272),
.B2(n_262),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_353),
.A2(n_373),
.B1(n_377),
.B2(n_382),
.Y(n_412)
);

OAI32xp33_ASAP7_75t_L g354 ( 
.A1(n_341),
.A2(n_264),
.A3(n_276),
.B1(n_295),
.B2(n_247),
.Y(n_354)
);

AOI221xp5_ASAP7_75t_L g405 ( 
.A1(n_354),
.A2(n_388),
.B1(n_340),
.B2(n_335),
.C(n_329),
.Y(n_405)
);

OAI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_297),
.A2(n_287),
.B1(n_257),
.B2(n_265),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_355),
.A2(n_379),
.B1(n_383),
.B2(n_339),
.Y(n_424)
);

OR2x2_ASAP7_75t_SL g393 ( 
.A(n_359),
.B(n_302),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_366),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_369),
.A2(n_337),
.B(n_309),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_372),
.B(n_384),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_323),
.A2(n_263),
.B1(n_291),
.B2(n_279),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_244),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_244),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_328),
.A2(n_263),
.B1(n_291),
.B2(n_259),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_380),
.B(n_381),
.C(n_338),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_327),
.B(n_336),
.C(n_334),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_312),
.A2(n_292),
.B1(n_288),
.B2(n_277),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_320),
.A2(n_292),
.B1(n_258),
.B2(n_267),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_314),
.B(n_294),
.Y(n_384)
);

OAI32xp33_ASAP7_75t_L g388 ( 
.A1(n_335),
.A2(n_294),
.A3(n_255),
.B1(n_5),
.B2(n_6),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_353),
.A2(n_332),
.B1(n_342),
.B2(n_324),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_389),
.A2(n_398),
.B1(n_420),
.B2(n_421),
.Y(n_427)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_367),
.Y(n_390)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_390),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_362),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_391),
.B(n_392),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_SL g456 ( 
.A1(n_393),
.A2(n_413),
.B(n_423),
.Y(n_456)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_367),
.Y(n_394)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_394),
.Y(n_434)
);

INVx13_ASAP7_75t_L g395 ( 
.A(n_387),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_395),
.Y(n_458)
);

O2A1O1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_396),
.A2(n_346),
.B(n_351),
.C(n_385),
.Y(n_448)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_397),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_352),
.A2(n_332),
.B1(n_302),
.B2(n_317),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_298),
.Y(n_401)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_401),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_380),
.C(n_376),
.Y(n_440)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_370),
.Y(n_403)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_403),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_405),
.B(n_414),
.Y(n_433)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_361),
.Y(n_406)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_406),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_374),
.B(n_365),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_407),
.B(n_409),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_378),
.B(n_300),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_410),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_347),
.B(n_315),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_358),
.Y(n_410)
);

INVx5_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_411),
.Y(n_436)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_360),
.B(n_318),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_321),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_358),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_415),
.B(n_416),
.Y(n_439)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_356),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_417),
.Y(n_426)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_357),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_418),
.A2(n_424),
.B1(n_377),
.B2(n_351),
.Y(n_437)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_419),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_371),
.A2(n_318),
.B1(n_306),
.B2(n_330),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_371),
.A2(n_318),
.B1(n_306),
.B2(n_326),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_308),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_422),
.Y(n_451)
);

AND2x6_ASAP7_75t_L g423 ( 
.A(n_359),
.B(n_343),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_425),
.A2(n_349),
.B1(n_364),
.B2(n_316),
.Y(n_452)
);

OA22x2_ASAP7_75t_L g428 ( 
.A1(n_424),
.A2(n_352),
.B1(n_382),
.B2(n_373),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g484 ( 
.A(n_428),
.Y(n_484)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_437),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_389),
.A2(n_379),
.B1(n_383),
.B2(n_348),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_438),
.A2(n_445),
.B1(n_449),
.B2(n_404),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_440),
.B(n_454),
.C(n_399),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_386),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_441),
.B(n_442),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_400),
.B(n_402),
.Y(n_442)
);

OAI22x1_ASAP7_75t_L g444 ( 
.A1(n_413),
.A2(n_348),
.B1(n_346),
.B2(n_388),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g462 ( 
.A1(n_444),
.A2(n_457),
.B(n_439),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_398),
.A2(n_369),
.B1(n_375),
.B2(n_354),
.Y(n_445)
);

XOR2x1_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_452),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_412),
.A2(n_421),
.B1(n_420),
.B2(n_410),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_392),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_453),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_396),
.B(n_425),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_399),
.B(n_364),
.C(n_310),
.Y(n_454)
);

OAI21xp33_ASAP7_75t_L g457 ( 
.A1(n_393),
.A2(n_349),
.B(n_343),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_408),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_459),
.B(n_440),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_429),
.B(n_419),
.Y(n_460)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_460),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_461),
.A2(n_471),
.B1(n_486),
.B2(n_448),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_462),
.A2(n_472),
.B(n_485),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_451),
.B(n_407),
.Y(n_463)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_463),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_454),
.C(n_452),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_430),
.B(n_404),
.Y(n_465)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_465),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_429),
.B(n_417),
.Y(n_467)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_467),
.Y(n_503)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_468),
.B(n_476),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_311),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_470),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_449),
.A2(n_423),
.B1(n_394),
.B2(n_403),
.Y(n_471)
);

NOR2xp67_ASAP7_75t_SL g472 ( 
.A(n_453),
.B(n_418),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_SL g473 ( 
.A1(n_458),
.A2(n_397),
.B1(n_390),
.B2(n_411),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_479),
.B1(n_481),
.B2(n_482),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_307),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_474),
.Y(n_495)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_434),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_416),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_477),
.B(n_478),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_436),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_458),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_427),
.A2(n_406),
.B1(n_368),
.B2(n_395),
.Y(n_481)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_436),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_450),
.B(n_387),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_483),
.A2(n_487),
.B1(n_445),
.B2(n_435),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_457),
.A2(n_387),
.B(n_344),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_427),
.A2(n_325),
.B1(n_387),
.B2(n_303),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_426),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_500),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_441),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_SL g522 ( 
.A(n_492),
.B(n_499),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_493),
.B(n_496),
.Y(n_513)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_494),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_464),
.B(n_456),
.C(n_428),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_498),
.A2(n_501),
.B1(n_460),
.B2(n_479),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_456),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_480),
.B(n_444),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_484),
.A2(n_428),
.B1(n_438),
.B2(n_432),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_469),
.B(n_428),
.C(n_455),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_511),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_462),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_504),
.B(n_505),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_471),
.B(n_447),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_484),
.A2(n_325),
.B1(n_4),
.B2(n_6),
.Y(n_507)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_507),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_466),
.B(n_3),
.C(n_7),
.Y(n_511)
);

INVx1_ASAP7_75t_SL g512 ( 
.A(n_510),
.Y(n_512)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_512),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g514 ( 
.A(n_491),
.B(n_477),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_514),
.A2(n_520),
.B1(n_526),
.B2(n_529),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_510),
.B(n_467),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_517),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_503),
.B(n_485),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g545 ( 
.A(n_518),
.B(n_528),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_489),
.A2(n_484),
.B1(n_466),
.B2(n_487),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_504),
.B(n_472),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_523),
.B(n_497),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g525 ( 
.A(n_509),
.B(n_476),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_525),
.B(n_530),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_498),
.A2(n_475),
.B1(n_468),
.B2(n_486),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_527),
.A2(n_503),
.B1(n_475),
.B2(n_501),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_506),
.B(n_482),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_506),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_490),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_515),
.B(n_495),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_532),
.B(n_533),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_516),
.B(n_488),
.C(n_493),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_522),
.B(n_499),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_535),
.B(n_537),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_502),
.C(n_496),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_536),
.B(n_538),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_522),
.B(n_492),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_513),
.B(n_505),
.C(n_500),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_541),
.B(n_542),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_521),
.B(n_508),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_511),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_543),
.B(n_546),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_544),
.A2(n_512),
.B1(n_526),
.B2(n_517),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_497),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_531),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_547),
.B(n_558),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_545),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_540),
.A2(n_518),
.B(n_545),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g563 ( 
.A1(n_549),
.A2(n_550),
.B(n_537),
.Y(n_563)
);

AOI21x1_ASAP7_75t_L g550 ( 
.A1(n_539),
.A2(n_518),
.B(n_528),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_519),
.C(n_523),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_551),
.A2(n_557),
.B(n_8),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_536),
.B(n_524),
.C(n_9),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_534),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_559),
.B(n_564),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_552),
.A2(n_538),
.B1(n_546),
.B2(n_535),
.Y(n_560)
);

AOI322xp5_ASAP7_75t_L g569 ( 
.A1(n_560),
.A2(n_553),
.A3(n_551),
.B1(n_554),
.B2(n_557),
.C1(n_15),
.C2(n_14),
.Y(n_569)
);

CKINVDCx16_ASAP7_75t_R g562 ( 
.A(n_555),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_562),
.A2(n_565),
.B(n_549),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g568 ( 
.A1(n_563),
.A2(n_550),
.B(n_548),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_556),
.B(n_8),
.C(n_10),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_567),
.B(n_569),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_568),
.A2(n_563),
.B(n_561),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_SL g574 ( 
.A(n_571),
.B(n_572),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g572 ( 
.A1(n_566),
.A2(n_565),
.B(n_559),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_570),
.B(n_554),
.Y(n_573)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_573),
.A2(n_574),
.B(n_13),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_L g576 ( 
.A1(n_575),
.A2(n_8),
.B(n_13),
.Y(n_576)
);

AOI21x1_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_8),
.B(n_13),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_14),
.C(n_15),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_15),
.Y(n_579)
);


endmodule