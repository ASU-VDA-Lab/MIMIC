module fake_jpeg_7961_n_98 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx11_ASAP7_75t_SL g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

OR2x2_ASAP7_75t_SL g32 ( 
.A(n_23),
.B(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_36),
.Y(n_47)
);

NOR2x1_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_20),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_41),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_44),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_45),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_27),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_50),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_38),
.A2(n_24),
.B1(n_25),
.B2(n_14),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_51),
.A2(n_35),
.B1(n_34),
.B2(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_28),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_36),
.C(n_32),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_55),
.B(n_56),
.Y(n_68)
);

NOR2xp67_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_26),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_35),
.B(n_24),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_16),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_48),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_0),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_34),
.B1(n_51),
.B2(n_49),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_53),
.C(n_43),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_69),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_58),
.B1(n_54),
.B2(n_49),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_61),
.Y(n_69)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_71),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_74),
.B1(n_45),
.B2(n_52),
.Y(n_84)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_67),
.A2(n_62),
.B(n_39),
.C(n_20),
.Y(n_74)
);

AOI322xp5_ASAP7_75t_SL g75 ( 
.A1(n_68),
.A2(n_16),
.A3(n_22),
.B1(n_19),
.B2(n_12),
.C1(n_4),
.C2(n_5),
.Y(n_75)
);

AOI322xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_77),
.A3(n_22),
.B1(n_19),
.B2(n_9),
.C1(n_5),
.C2(n_8),
.Y(n_83)
);

A2O1A1O1Ixp25_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_65),
.B(n_58),
.C(n_17),
.D(n_13),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_72),
.B(n_70),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_80),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_71),
.C(n_46),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_46),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_74),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_82),
.A2(n_83),
.B(n_84),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_87),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_81),
.B(n_74),
.Y(n_87)
);

AOI321xp33_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C(n_28),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_93),
.B(n_92),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_82),
.B(n_3),
.C(n_2),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_94),
.Y(n_98)
);


endmodule