module fake_ariane_2179_n_2110 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_2110);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_2110;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_279;
wire n_958;
wire n_813;
wire n_419;
wire n_1985;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_851;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2072;
wire n_306;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_2100;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_1802;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_1906;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1966;
wire n_1243;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1429;
wire n_1324;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_914;
wire n_330;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1955;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_1986;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_1956;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1967;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_67),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_52),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_33),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_138),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_192),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_96),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_106),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_60),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_187),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_72),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_142),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_201),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_171),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_131),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_126),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_47),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_48),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_105),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_39),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_151),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_140),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_102),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_159),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_1),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_209),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_32),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_34),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_76),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_191),
.Y(n_248)
);

INVx2_ASAP7_75t_SL g249 ( 
.A(n_82),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_134),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_89),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_135),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_95),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_84),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_3),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_52),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_197),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_45),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_139),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_9),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_154),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_180),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_30),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_136),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_32),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_120),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_77),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_48),
.Y(n_269)
);

BUFx10_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_157),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_18),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_161),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_34),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_38),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_155),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_39),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_144),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_110),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_17),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_94),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_196),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_66),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_189),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_86),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_121),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_30),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_193),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_90),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_38),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_125),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_141),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_214),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_88),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_9),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_116),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_107),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_20),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_33),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_25),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_68),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_49),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_62),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_19),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_55),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_170),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_25),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_2),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_113),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_68),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_11),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_74),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_14),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_182),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_16),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_167),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_43),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_112),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_117),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_183),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_53),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_75),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_63),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_203),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_130),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_11),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_145),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_168),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_53),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_123),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_69),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_59),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_104),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_56),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_91),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_19),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_166),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_100),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_103),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_76),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_18),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_164),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_128),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_163),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_185),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_208),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_99),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_174),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_122),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_186),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_14),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_43),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_160),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_172),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_70),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_8),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_50),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_108),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_21),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_195),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_206),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_69),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_67),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_65),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_66),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_188),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_13),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_85),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_109),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_204),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_26),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_26),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_8),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_5),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_44),
.Y(n_377)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_71),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_200),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_36),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_56),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_82),
.Y(n_382)
);

BUFx10_ASAP7_75t_L g383 ( 
.A(n_59),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_118),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_212),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_150),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_3),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_194),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_176),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_181),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_31),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_98),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_173),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_190),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_42),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_10),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_156),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g398 ( 
.A(n_78),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_23),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_84),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_57),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_54),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_213),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_198),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_93),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_210),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_71),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_80),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_28),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_41),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_137),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_80),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_72),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_73),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_51),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_179),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_70),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_44),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_24),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_47),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_0),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_101),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_50),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_177),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_232),
.Y(n_425)
);

BUFx2_ASAP7_75t_SL g426 ( 
.A(n_243),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_240),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_251),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_219),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_287),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_350),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_371),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_250),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g434 ( 
.A(n_269),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_404),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_215),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_219),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_268),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_220),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_220),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_223),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_R g442 ( 
.A(n_337),
.B(n_87),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g443 ( 
.A(n_249),
.B(n_0),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_380),
.Y(n_444)
);

INVxp33_ASAP7_75t_L g445 ( 
.A(n_247),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_328),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_380),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_229),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_229),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_315),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_239),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_239),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_331),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_245),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_245),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_258),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_398),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_216),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_223),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_258),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_269),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_249),
.B(n_1),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_315),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_359),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_275),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_217),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_273),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_273),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_225),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_235),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_278),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_278),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_237),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_244),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_282),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_255),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_231),
.B(n_2),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_275),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_414),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_282),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_292),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_231),
.B(n_4),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_292),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_256),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_308),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_259),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_308),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_262),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_264),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_262),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_315),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_272),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_353),
.B(n_4),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_316),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_243),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_316),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_277),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_233),
.Y(n_499)
);

CKINVDCx16_ASAP7_75t_R g500 ( 
.A(n_242),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_320),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_320),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_321),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_243),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_243),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_222),
.B(n_5),
.Y(n_506)
);

NOR2xp67_ASAP7_75t_L g507 ( 
.A(n_374),
.B(n_6),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_270),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_321),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_288),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_326),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_326),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_291),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_296),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_270),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_309),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_300),
.B(n_6),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_315),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_299),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_301),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_270),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_233),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_349),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_349),
.B(n_7),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_351),
.Y(n_525)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_378),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_270),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_351),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g529 ( 
.A(n_374),
.B(n_7),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_356),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_356),
.Y(n_531)
);

CKINVDCx16_ASAP7_75t_R g532 ( 
.A(n_242),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_302),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_363),
.B(n_10),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_492),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_492),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_429),
.B(n_363),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_492),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_429),
.B(n_378),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_437),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_437),
.B(n_370),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_450),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_439),
.B(n_370),
.Y(n_543)
);

INVx5_ASAP7_75t_L g544 ( 
.A(n_433),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_450),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_439),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_440),
.B(n_300),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_440),
.B(n_325),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_433),
.Y(n_549)
);

BUFx8_ASAP7_75t_L g550 ( 
.A(n_462),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_478),
.B(n_315),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_448),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_448),
.Y(n_553)
);

BUFx8_ASAP7_75t_L g554 ( 
.A(n_462),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_449),
.B(n_379),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_449),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_451),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_451),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_453),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_455),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_464),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_433),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_433),
.Y(n_564)
);

CKINVDCx8_ASAP7_75t_R g565 ( 
.A(n_426),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_433),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_455),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_518),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_518),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g572 ( 
.A(n_436),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_456),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_457),
.B(n_379),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_444),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_457),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_461),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_447),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_461),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_468),
.B(n_469),
.Y(n_580)
);

BUFx2_ASAP7_75t_L g581 ( 
.A(n_458),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_469),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_452),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_472),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_472),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_473),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_473),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_476),
.B(n_388),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_466),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_476),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_500),
.B(n_311),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_481),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_481),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_482),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_484),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_484),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g599 ( 
.A(n_516),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_486),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_486),
.B(n_388),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_488),
.B(n_394),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_434),
.B(n_483),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g604 ( 
.A1(n_488),
.A2(n_397),
.B(n_394),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_495),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_495),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_497),
.Y(n_607)
);

CKINVDCx8_ASAP7_75t_R g608 ( 
.A(n_426),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_497),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_501),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_489),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_501),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_442),
.B(n_315),
.Y(n_613)
);

BUFx2_ASAP7_75t_L g614 ( 
.A(n_491),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_502),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_502),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_503),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_503),
.B(n_325),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_509),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_509),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_511),
.Y(n_621)
);

BUFx3_ASAP7_75t_L g622 ( 
.A(n_479),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_585),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_585),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_603),
.B(n_441),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_565),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_585),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_565),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_584),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_542),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_565),
.B(n_459),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_585),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_547),
.B(n_441),
.Y(n_633)
);

INVx5_ASAP7_75t_L g634 ( 
.A(n_549),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_608),
.B(n_467),
.Y(n_635)
);

BUFx10_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_585),
.B(n_534),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_585),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_542),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_585),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_591),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_613),
.A2(n_460),
.B1(n_524),
.B2(n_494),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_608),
.B(n_470),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_591),
.B(n_460),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_613),
.A2(n_445),
.B1(n_517),
.B2(n_463),
.Y(n_645)
);

INVx4_ASAP7_75t_SL g646 ( 
.A(n_586),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_586),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_572),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_584),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_547),
.B(n_548),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_586),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_591),
.B(n_600),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_L g653 ( 
.A1(n_608),
.A2(n_507),
.B1(n_529),
.B2(n_443),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_604),
.A2(n_517),
.B1(n_512),
.B2(n_511),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

BUFx6f_ASAP7_75t_L g656 ( 
.A(n_586),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_562),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_591),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_600),
.B(n_512),
.Y(n_659)
);

INVx4_ASAP7_75t_L g660 ( 
.A(n_600),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_592),
.B(n_532),
.Y(n_661)
);

NAND3xp33_ASAP7_75t_L g662 ( 
.A(n_586),
.B(n_525),
.C(n_523),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_586),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_R g664 ( 
.A(n_578),
.B(n_425),
.Y(n_664)
);

AND2x2_ASAP7_75t_SL g665 ( 
.A(n_604),
.B(n_389),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_539),
.Y(n_666)
);

OAI22x1_ASAP7_75t_L g667 ( 
.A1(n_599),
.A2(n_506),
.B1(n_430),
.B2(n_432),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_562),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_600),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_586),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_609),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_609),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_562),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_540),
.B(n_471),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_599),
.B(n_427),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_604),
.A2(n_525),
.B1(n_528),
.B2(n_523),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_609),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_540),
.B(n_474),
.Y(n_678)
);

BUFx8_ASAP7_75t_SL g679 ( 
.A(n_611),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_578),
.B(n_475),
.Y(n_680)
);

BUFx4f_ASAP7_75t_L g681 ( 
.A(n_587),
.Y(n_681)
);

NAND3xp33_ASAP7_75t_L g682 ( 
.A(n_587),
.B(n_530),
.C(n_528),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_570),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_581),
.B(n_477),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_587),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_609),
.B(n_530),
.Y(n_687)
);

INVx1_ASAP7_75t_SL g688 ( 
.A(n_581),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_604),
.A2(n_531),
.B1(n_504),
.B2(n_505),
.Y(n_689)
);

NAND2xp33_ASAP7_75t_L g690 ( 
.A(n_587),
.B(n_419),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_547),
.B(n_531),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_587),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_546),
.B(n_485),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_570),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_571),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_546),
.B(n_487),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_552),
.B(n_490),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_552),
.B(n_493),
.Y(n_698)
);

BUFx4f_ASAP7_75t_L g699 ( 
.A(n_587),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_575),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_553),
.B(n_498),
.Y(n_701)
);

AND2x6_ASAP7_75t_L g702 ( 
.A(n_573),
.B(n_397),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_553),
.B(n_510),
.Y(n_703)
);

NOR2x1p5_ASAP7_75t_L g704 ( 
.A(n_580),
.B(n_513),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_580),
.B(n_514),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_587),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_588),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_588),
.Y(n_708)
);

NAND3xp33_ASAP7_75t_L g709 ( 
.A(n_588),
.B(n_419),
.C(n_405),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_556),
.B(n_519),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_588),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_588),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_571),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_604),
.A2(n_618),
.B1(n_622),
.B2(n_590),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_588),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_588),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_548),
.B(n_539),
.Y(n_717)
);

BUFx4f_ASAP7_75t_L g718 ( 
.A(n_606),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_556),
.B(n_520),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_606),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_571),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_539),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_557),
.B(n_533),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_557),
.B(n_496),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_606),
.Y(n_725)
);

OR2x6_ASAP7_75t_L g726 ( 
.A(n_548),
.B(n_499),
.Y(n_726)
);

BUFx6f_ASAP7_75t_L g727 ( 
.A(n_606),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_618),
.A2(n_515),
.B1(n_521),
.B2(n_508),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_606),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_535),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_558),
.B(n_522),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_618),
.B(n_526),
.Y(n_732)
);

AND2x6_ASAP7_75t_L g733 ( 
.A(n_573),
.B(n_582),
.Y(n_733)
);

INVx4_ASAP7_75t_L g734 ( 
.A(n_606),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_558),
.B(n_435),
.Y(n_735)
);

INVx4_ASAP7_75t_SL g736 ( 
.A(n_606),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_536),
.Y(n_737)
);

INVx8_ASAP7_75t_L g738 ( 
.A(n_619),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_559),
.B(n_238),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_619),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_618),
.A2(n_527),
.B1(n_400),
.B2(n_423),
.Y(n_741)
);

BUFx10_ASAP7_75t_L g742 ( 
.A(n_618),
.Y(n_742)
);

BUFx10_ASAP7_75t_L g743 ( 
.A(n_559),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_536),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_619),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_619),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_560),
.B(n_406),
.Y(n_747)
);

INVx1_ASAP7_75t_SL g748 ( 
.A(n_611),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_614),
.B(n_506),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_619),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_619),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_619),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_550),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_560),
.B(n_406),
.Y(n_754)
);

OAI22xp33_ASAP7_75t_SL g755 ( 
.A1(n_537),
.A2(n_246),
.B1(n_254),
.B2(n_234),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_573),
.A2(n_373),
.B1(n_381),
.B2(n_319),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_561),
.B(n_295),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_538),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_614),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_590),
.A2(n_400),
.B1(n_423),
.B2(n_391),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_561),
.B(n_295),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_567),
.B(n_242),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_538),
.Y(n_763)
);

INVx3_ASAP7_75t_L g764 ( 
.A(n_582),
.Y(n_764)
);

NOR3xp33_ASAP7_75t_L g765 ( 
.A(n_537),
.B(n_412),
.C(n_246),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_545),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_582),
.B(n_389),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_590),
.A2(n_391),
.B1(n_254),
.B2(n_261),
.Y(n_768)
);

BUFx6f_ASAP7_75t_L g769 ( 
.A(n_569),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_593),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_545),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_593),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_567),
.B(n_428),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_568),
.B(n_431),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_568),
.B(n_242),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_636),
.B(n_622),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_743),
.B(n_576),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_630),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_674),
.B(n_576),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_656),
.B(n_577),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_678),
.B(n_577),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_693),
.B(n_579),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_630),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_626),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_698),
.B(n_579),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_636),
.B(n_705),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_730),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_626),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_701),
.B(n_583),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_743),
.B(n_583),
.Y(n_790)
);

NOR2xp67_ASAP7_75t_L g791 ( 
.A(n_675),
.B(n_593),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_703),
.B(n_594),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_625),
.B(n_594),
.Y(n_793)
);

BUFx8_ASAP7_75t_L g794 ( 
.A(n_629),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_691),
.B(n_595),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_737),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_737),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_743),
.B(n_595),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_744),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_744),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_639),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_691),
.B(n_596),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_636),
.B(n_641),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_675),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_666),
.B(n_596),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_666),
.B(n_597),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_628),
.B(n_622),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_641),
.B(n_597),
.Y(n_808)
);

NOR2xp67_ASAP7_75t_L g809 ( 
.A(n_629),
.B(n_607),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_628),
.B(n_598),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_688),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_641),
.B(n_598),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_L g813 ( 
.A1(n_714),
.A2(n_554),
.B1(n_550),
.B2(n_605),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_722),
.B(n_605),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_722),
.B(n_610),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_731),
.A2(n_755),
.B(n_644),
.C(n_687),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_655),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_696),
.B(n_610),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_700),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_717),
.B(n_612),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_758),
.Y(n_821)
);

NOR2xp67_ASAP7_75t_L g822 ( 
.A(n_649),
.B(n_607),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_697),
.B(n_612),
.Y(n_823)
);

INVx8_ASAP7_75t_L g824 ( 
.A(n_726),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_615),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_719),
.B(n_615),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_652),
.A2(n_551),
.B(n_543),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_739),
.B(n_717),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_649),
.B(n_700),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_655),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_650),
.B(n_621),
.Y(n_831)
);

BUFx8_ASAP7_75t_L g832 ( 
.A(n_749),
.Y(n_832)
);

BUFx6f_ASAP7_75t_SL g833 ( 
.A(n_700),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_650),
.B(n_658),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_748),
.B(n_541),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_658),
.B(n_607),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_660),
.B(n_616),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_657),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_657),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_665),
.A2(n_554),
.B1(n_550),
.B2(n_616),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_758),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_660),
.B(n_616),
.Y(n_842)
);

AND2x6_ASAP7_75t_L g843 ( 
.A(n_669),
.B(n_617),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_660),
.B(n_617),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_763),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_763),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_677),
.B(n_617),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_677),
.B(n_665),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_770),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_656),
.B(n_620),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_677),
.B(n_620),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_SL g852 ( 
.A(n_753),
.B(n_550),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_723),
.B(n_550),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_665),
.A2(n_554),
.B1(n_620),
.B2(n_286),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_654),
.B(n_669),
.Y(n_855)
);

AOI22xp33_ASAP7_75t_L g856 ( 
.A1(n_689),
.A2(n_554),
.B1(n_286),
.B2(n_384),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_724),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_671),
.B(n_541),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_671),
.B(n_543),
.Y(n_859)
);

INVx3_ASAP7_75t_L g860 ( 
.A(n_672),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_653),
.A2(n_554),
.B1(n_574),
.B2(n_555),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_672),
.B(n_555),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_668),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_656),
.B(n_574),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_656),
.B(n_589),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_772),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_659),
.B(n_589),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_656),
.B(n_601),
.Y(n_868)
);

INVx8_ASAP7_75t_L g869 ( 
.A(n_726),
.Y(n_869)
);

O2A1O1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_755),
.A2(n_602),
.B(n_601),
.C(n_261),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_668),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_773),
.B(n_438),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_741),
.A2(n_286),
.B1(n_384),
.B2(n_285),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_759),
.B(n_602),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_631),
.B(n_304),
.Y(n_875)
);

OR2x2_ASAP7_75t_SL g876 ( 
.A(n_749),
.B(n_446),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_673),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_670),
.B(n_392),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_772),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_635),
.B(n_305),
.Y(n_880)
);

NOR3xp33_ASAP7_75t_L g881 ( 
.A(n_680),
.B(n_266),
.C(n_234),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_664),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_764),
.Y(n_883)
);

AOI221xp5_ASAP7_75t_L g884 ( 
.A1(n_765),
.A2(n_324),
.B1(n_317),
.B2(n_306),
.C(n_303),
.Y(n_884)
);

INVx3_ASAP7_75t_L g885 ( 
.A(n_742),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_764),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_670),
.B(n_392),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_645),
.B(n_545),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_673),
.Y(n_889)
);

NOR2xp67_ASAP7_75t_L g890 ( 
.A(n_661),
.B(n_753),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_764),
.B(n_545),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_733),
.Y(n_892)
);

BUFx2_ASAP7_75t_L g893 ( 
.A(n_648),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_766),
.Y(n_894)
);

AND2x4_ASAP7_75t_L g895 ( 
.A(n_726),
.B(n_266),
.Y(n_895)
);

BUFx8_ASAP7_75t_L g896 ( 
.A(n_732),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_643),
.B(n_307),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_683),
.Y(n_898)
);

BUFx2_ASAP7_75t_L g899 ( 
.A(n_648),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_742),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_683),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_670),
.B(n_252),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_642),
.B(n_274),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_685),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_679),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_766),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_633),
.B(n_274),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_670),
.B(n_711),
.Y(n_908)
);

AND2x2_ASAP7_75t_SL g909 ( 
.A(n_676),
.B(n_252),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_637),
.A2(n_563),
.B(n_549),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_771),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_771),
.Y(n_912)
);

BUFx6f_ASAP7_75t_L g913 ( 
.A(n_670),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_742),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_726),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_685),
.Y(n_916)
);

OAI22xp33_ASAP7_75t_L g917 ( 
.A1(n_756),
.A2(n_324),
.B1(n_342),
.B2(n_281),
.Y(n_917)
);

AOI22xp5_ASAP7_75t_L g918 ( 
.A1(n_704),
.A2(n_290),
.B1(n_424),
.B2(n_422),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_694),
.Y(n_919)
);

NAND2x1_ASAP7_75t_L g920 ( 
.A(n_733),
.B(n_389),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_694),
.Y(n_921)
);

AND2x6_ASAP7_75t_L g922 ( 
.A(n_711),
.B(n_389),
.Y(n_922)
);

INVx2_ASAP7_75t_SL g923 ( 
.A(n_633),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_732),
.B(n_281),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_747),
.A2(n_303),
.B(n_408),
.C(n_306),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_757),
.B(n_284),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_735),
.B(n_310),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_695),
.Y(n_928)
);

INVxp67_ASAP7_75t_SL g929 ( 
.A(n_711),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_774),
.B(n_313),
.C(n_312),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_711),
.B(n_265),
.Y(n_931)
);

INVxp67_ASAP7_75t_L g932 ( 
.A(n_684),
.Y(n_932)
);

BUFx6f_ASAP7_75t_SL g933 ( 
.A(n_702),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_695),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_711),
.B(n_265),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_761),
.B(n_284),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_754),
.B(n_317),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_727),
.B(n_332),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_762),
.B(n_314),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_760),
.B(n_342),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_778),
.Y(n_941)
);

AOI22xp33_ASAP7_75t_L g942 ( 
.A1(n_909),
.A2(n_756),
.B1(n_702),
.B2(n_768),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_779),
.B(n_781),
.Y(n_943)
);

AO21x1_ASAP7_75t_L g944 ( 
.A1(n_848),
.A2(n_637),
.B(n_624),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_778),
.Y(n_945)
);

AOI22xp5_ASAP7_75t_L g946 ( 
.A1(n_857),
.A2(n_704),
.B1(n_775),
.B2(n_733),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_836),
.A2(n_699),
.B(n_681),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_782),
.B(n_632),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_786),
.A2(n_638),
.B(n_712),
.C(n_632),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_837),
.A2(n_699),
.B(n_681),
.Y(n_950)
);

INVx2_ASAP7_75t_L g951 ( 
.A(n_783),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_835),
.B(n_728),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_804),
.B(n_725),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_917),
.A2(n_413),
.A3(n_408),
.B1(n_407),
.B2(n_387),
.C(n_375),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_L g955 ( 
.A1(n_786),
.A2(n_638),
.B(n_712),
.C(n_632),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_828),
.B(n_785),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_874),
.B(n_667),
.Y(n_957)
);

NAND2xp33_ASAP7_75t_L g958 ( 
.A(n_843),
.B(n_733),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_847),
.A2(n_699),
.B(n_681),
.Y(n_959)
);

BUFx6f_ASAP7_75t_L g960 ( 
.A(n_913),
.Y(n_960)
);

AOI21x1_ASAP7_75t_L g961 ( 
.A1(n_908),
.A2(n_624),
.B(n_623),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_789),
.B(n_792),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_784),
.B(n_646),
.Y(n_963)
);

AOI22xp5_ASAP7_75t_L g964 ( 
.A1(n_791),
.A2(n_733),
.B1(n_667),
.B2(n_725),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_867),
.A2(n_718),
.B(n_738),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_811),
.Y(n_966)
);

HB1xp67_ASAP7_75t_L g967 ( 
.A(n_915),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_932),
.B(n_725),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_820),
.B(n_638),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_820),
.B(n_712),
.Y(n_970)
);

OAI21xp5_ASAP7_75t_L g971 ( 
.A1(n_827),
.A2(n_627),
.B(n_623),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_872),
.B(n_454),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_820),
.B(n_720),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_849),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_834),
.A2(n_823),
.B(n_825),
.C(n_818),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_826),
.B(n_882),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_776),
.B(n_720),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_824),
.B(n_738),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_853),
.A2(n_733),
.B1(n_746),
.B2(n_734),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_831),
.A2(n_367),
.B(n_375),
.C(n_365),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_776),
.B(n_720),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_923),
.B(n_734),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_892),
.B(n_727),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_810),
.B(n_750),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_L g985 ( 
.A(n_819),
.B(n_662),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_816),
.A2(n_751),
.B(n_750),
.C(n_640),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_864),
.A2(n_640),
.B(n_627),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_908),
.A2(n_738),
.B(n_651),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_892),
.B(n_727),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_864),
.A2(n_651),
.B(n_647),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_808),
.A2(n_663),
.B(n_647),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_885),
.B(n_727),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_808),
.A2(n_686),
.B(n_663),
.Y(n_993)
);

O2A1O1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_858),
.A2(n_367),
.B(n_387),
.C(n_365),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_801),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_810),
.B(n_750),
.Y(n_996)
);

AOI21x1_ASAP7_75t_L g997 ( 
.A1(n_842),
.A2(n_692),
.B(n_686),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_810),
.B(n_751),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_843),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_793),
.B(n_751),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_812),
.A2(n_706),
.B(n_692),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_829),
.B(n_465),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_859),
.A2(n_413),
.B(n_407),
.C(n_745),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_812),
.A2(n_707),
.B(n_706),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_853),
.A2(n_733),
.B1(n_734),
.B2(n_746),
.Y(n_1005)
);

NOR2x1_ASAP7_75t_L g1006 ( 
.A(n_784),
.B(n_662),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_842),
.A2(n_851),
.B(n_844),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_895),
.B(n_480),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_795),
.B(n_746),
.Y(n_1009)
);

INVxp67_ASAP7_75t_L g1010 ( 
.A(n_893),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_913),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_802),
.B(n_713),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_809),
.B(n_713),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_822),
.B(n_721),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_844),
.A2(n_851),
.B(n_790),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_777),
.A2(n_708),
.B(n_707),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_788),
.B(n_927),
.Y(n_1017)
);

NAND2x1_ASAP7_75t_L g1018 ( 
.A(n_843),
.B(n_913),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_865),
.A2(n_715),
.B(n_708),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_862),
.A2(n_745),
.B(n_740),
.C(n_715),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_895),
.B(n_383),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_895),
.B(n_383),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_905),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_899),
.B(n_383),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_807),
.B(n_721),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_L g1026 ( 
.A(n_788),
.B(n_927),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_890),
.B(n_383),
.Y(n_1027)
);

NOR2xp67_ASAP7_75t_L g1028 ( 
.A(n_930),
.B(n_918),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_924),
.B(n_682),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_777),
.A2(n_740),
.B(n_716),
.Y(n_1030)
);

NOR2x1_ASAP7_75t_L g1031 ( 
.A(n_807),
.B(n_682),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_807),
.B(n_716),
.Y(n_1032)
);

INVxp67_ASAP7_75t_L g1033 ( 
.A(n_896),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_885),
.B(n_727),
.Y(n_1034)
);

INVx6_ASAP7_75t_L g1035 ( 
.A(n_794),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_866),
.Y(n_1036)
);

O2A1O1Ixp33_ASAP7_75t_SL g1037 ( 
.A1(n_803),
.A2(n_332),
.B(n_345),
.C(n_709),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_817),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_870),
.A2(n_709),
.B(n_752),
.C(n_729),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_790),
.A2(n_752),
.B(n_729),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_879),
.Y(n_1041)
);

INVx3_ASAP7_75t_L g1042 ( 
.A(n_843),
.Y(n_1042)
);

OAI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_865),
.A2(n_702),
.B(n_690),
.Y(n_1043)
);

BUFx5_ASAP7_75t_L g1044 ( 
.A(n_843),
.Y(n_1044)
);

NOR2xp67_ASAP7_75t_L g1045 ( 
.A(n_875),
.B(n_634),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_900),
.B(n_729),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_798),
.A2(n_752),
.B(n_729),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_913),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_798),
.A2(n_752),
.B(n_729),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_868),
.A2(n_769),
.B(n_690),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_914),
.B(n_769),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_900),
.B(n_769),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_868),
.A2(n_345),
.B(n_702),
.C(n_646),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_794),
.Y(n_1054)
);

NOR2xp67_ASAP7_75t_L g1055 ( 
.A(n_875),
.B(n_634),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_824),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_805),
.B(n_702),
.Y(n_1057)
);

AOI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_861),
.A2(n_702),
.B1(n_767),
.B2(n_736),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_880),
.B(n_769),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_929),
.A2(n_634),
.B(n_221),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_794),
.Y(n_1061)
);

NAND2xp33_ASAP7_75t_L g1062 ( 
.A(n_860),
.B(n_702),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_860),
.Y(n_1063)
);

OAI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_910),
.A2(n_767),
.B(n_634),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_855),
.A2(n_409),
.B1(n_366),
.B2(n_376),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_880),
.B(n_323),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_897),
.A2(n_840),
.B1(n_869),
.B2(n_824),
.Y(n_1067)
);

AOI22xp33_ASAP7_75t_L g1068 ( 
.A1(n_909),
.A2(n_767),
.B1(n_285),
.B2(n_286),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_806),
.B(n_646),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_814),
.B(n_646),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_883),
.A2(n_634),
.B(n_224),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_787),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_854),
.A2(n_815),
.B1(n_813),
.B2(n_886),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_876),
.B(n_333),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_830),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_897),
.B(n_334),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_869),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_891),
.A2(n_906),
.B(n_894),
.Y(n_1078)
);

AO21x1_ASAP7_75t_L g1079 ( 
.A1(n_902),
.A2(n_736),
.B(n_767),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_830),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_911),
.A2(n_634),
.B(n_226),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_933),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_852),
.B(n_336),
.Y(n_1083)
);

INVx6_ASAP7_75t_L g1084 ( 
.A(n_896),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_937),
.B(n_903),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_796),
.B(n_736),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_933),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_912),
.A2(n_227),
.B(n_218),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_838),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_797),
.B(n_736),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_926),
.B(n_767),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_799),
.A2(n_767),
.B(n_544),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_850),
.A2(n_230),
.B(n_228),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_SL g1094 ( 
.A(n_800),
.B(n_419),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_838),
.Y(n_1095)
);

NOR2xp67_ASAP7_75t_L g1096 ( 
.A(n_936),
.B(n_236),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_821),
.A2(n_767),
.B(n_544),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_907),
.B(n_338),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_873),
.B(n_343),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_841),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_839),
.Y(n_1101)
);

BUFx4f_ASAP7_75t_L g1102 ( 
.A(n_869),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_939),
.B(n_354),
.Y(n_1103)
);

OAI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_939),
.A2(n_358),
.B(n_357),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_845),
.A2(n_248),
.B(n_241),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_881),
.B(n_294),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_846),
.Y(n_1107)
);

AOI21x1_ASAP7_75t_L g1108 ( 
.A1(n_902),
.A2(n_544),
.B(n_549),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_940),
.B(n_361),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_896),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_780),
.A2(n_257),
.B(n_253),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_839),
.A2(n_263),
.B(n_260),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_884),
.A2(n_364),
.B(n_401),
.C(n_402),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_888),
.B(n_369),
.Y(n_1114)
);

AOI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_856),
.A2(n_285),
.B1(n_384),
.B2(n_294),
.Y(n_1115)
);

INVx1_ASAP7_75t_SL g1116 ( 
.A(n_922),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_925),
.A2(n_322),
.B(n_417),
.C(n_377),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_863),
.A2(n_360),
.B(n_335),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_863),
.A2(n_362),
.B(n_339),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_871),
.A2(n_368),
.B(n_340),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_833),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_943),
.A2(n_887),
.B(n_878),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_966),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_956),
.B(n_832),
.Y(n_1124)
);

AOI22xp33_ASAP7_75t_L g1125 ( 
.A1(n_952),
.A2(n_832),
.B1(n_833),
.B2(n_916),
.Y(n_1125)
);

BUFx6f_ASAP7_75t_L g1126 ( 
.A(n_1056),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_1066),
.A2(n_920),
.B(n_878),
.C(n_887),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_957),
.A2(n_832),
.B1(n_871),
.B2(n_934),
.Y(n_1128)
);

NOR3xp33_ASAP7_75t_L g1129 ( 
.A(n_1066),
.B(n_396),
.C(n_399),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_956),
.B(n_877),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_SL g1131 ( 
.A1(n_962),
.A2(n_938),
.B(n_935),
.C(n_931),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_1017),
.B(n_877),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1076),
.A2(n_922),
.B1(n_420),
.B2(n_418),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1056),
.Y(n_1134)
);

AND2x4_ASAP7_75t_L g1135 ( 
.A(n_1056),
.B(n_889),
.Y(n_1135)
);

OAI22xp5_ASAP7_75t_L g1136 ( 
.A1(n_1076),
.A2(n_919),
.B1(n_889),
.B2(n_934),
.Y(n_1136)
);

AO21x1_ASAP7_75t_L g1137 ( 
.A1(n_1059),
.A2(n_938),
.B(n_935),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_966),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_975),
.A2(n_928),
.B(n_898),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_1084),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_1017),
.B(n_898),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_R g1142 ( 
.A(n_1023),
.B(n_922),
.Y(n_1142)
);

AOI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_1002),
.A2(n_922),
.B1(n_395),
.B2(n_382),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_965),
.A2(n_928),
.B(n_901),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_948),
.A2(n_901),
.B(n_921),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_976),
.B(n_904),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1026),
.A2(n_922),
.B1(n_421),
.B2(n_415),
.Y(n_1147)
);

INVx3_ASAP7_75t_L g1148 ( 
.A(n_978),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_SL g1149 ( 
.A1(n_1103),
.A2(n_285),
.B1(n_384),
.B2(n_410),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1056),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_976),
.B(n_904),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_1026),
.B(n_919),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_1084),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1008),
.B(n_921),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_SL g1155 ( 
.A(n_1054),
.B(n_419),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1061),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1062),
.A2(n_346),
.B(n_267),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1021),
.B(n_419),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_947),
.A2(n_347),
.B(n_271),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_941),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1010),
.A2(n_348),
.B1(n_280),
.B2(n_283),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_974),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_972),
.B(n_289),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_1010),
.B(n_293),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_950),
.A2(n_372),
.B(n_297),
.Y(n_1165)
);

OAI21xp33_ASAP7_75t_L g1166 ( 
.A1(n_1104),
.A2(n_419),
.B(n_322),
.Y(n_1166)
);

AOI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1083),
.A2(n_385),
.B1(n_298),
.B2(n_318),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_953),
.B(n_327),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_942),
.A2(n_352),
.B1(n_416),
.B2(n_411),
.Y(n_1169)
);

OAI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_986),
.A2(n_544),
.B(n_329),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_945),
.Y(n_1171)
);

OAI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_942),
.A2(n_344),
.B1(n_403),
.B2(n_393),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_978),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1068),
.A2(n_341),
.B1(n_390),
.B2(n_386),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_959),
.A2(n_330),
.B(n_355),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_967),
.B(n_12),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1022),
.B(n_569),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_967),
.B(n_12),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1098),
.B(n_13),
.Y(n_1179)
);

BUFx4f_ASAP7_75t_L g1180 ( 
.A(n_1084),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_SL g1181 ( 
.A1(n_953),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_968),
.B(n_569),
.Y(n_1182)
);

NAND2xp33_ASAP7_75t_R g1183 ( 
.A(n_963),
.B(n_1082),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_969),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_L g1185 ( 
.A(n_1113),
.B(n_1083),
.C(n_1028),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_1074),
.B(n_15),
.Y(n_1186)
);

INVxp67_ASAP7_75t_L g1187 ( 
.A(n_1024),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1085),
.B(n_20),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_L g1189 ( 
.A(n_1035),
.B(n_21),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1029),
.B(n_22),
.Y(n_1190)
);

INVx5_ASAP7_75t_L g1191 ( 
.A(n_978),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_968),
.B(n_22),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1035),
.B(n_23),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1036),
.B(n_1041),
.Y(n_1194)
);

BUFx8_ASAP7_75t_L g1195 ( 
.A(n_1027),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_1033),
.A2(n_1035),
.B1(n_1067),
.B2(n_1110),
.Y(n_1196)
);

NOR3xp33_ASAP7_75t_SL g1197 ( 
.A(n_1065),
.B(n_24),
.C(n_27),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_L g1198 ( 
.A(n_1059),
.B(n_27),
.Y(n_1198)
);

O2A1O1Ixp5_ASAP7_75t_L g1199 ( 
.A1(n_944),
.A2(n_29),
.B(n_31),
.C(n_35),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_980),
.A2(n_29),
.B(n_35),
.C(n_37),
.Y(n_1200)
);

INVxp67_ASAP7_75t_L g1201 ( 
.A(n_1110),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1102),
.B(n_569),
.Y(n_1202)
);

INVx3_ASAP7_75t_L g1203 ( 
.A(n_1077),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1033),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_SL g1205 ( 
.A(n_1099),
.B(n_37),
.C(n_40),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_985),
.A2(n_569),
.B1(n_250),
.B2(n_279),
.Y(n_1206)
);

NOR3xp33_ASAP7_75t_SL g1207 ( 
.A(n_954),
.B(n_40),
.C(n_41),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1015),
.A2(n_569),
.B(n_250),
.C(n_279),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1077),
.Y(n_1209)
);

INVx3_ASAP7_75t_L g1210 ( 
.A(n_1077),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1072),
.B(n_42),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1068),
.A2(n_279),
.B1(n_276),
.B2(n_250),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1102),
.B(n_569),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_946),
.A2(n_250),
.B(n_276),
.C(n_279),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_971),
.A2(n_279),
.B(n_276),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_994),
.A2(n_250),
.B(n_276),
.C(n_279),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1063),
.B(n_45),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_960),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_977),
.A2(n_544),
.B(n_276),
.Y(n_1219)
);

NAND2x1p5_ASAP7_75t_L g1220 ( 
.A(n_1082),
.B(n_544),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_SL g1221 ( 
.A(n_1116),
.B(n_46),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1063),
.B(n_46),
.Y(n_1222)
);

OAI21xp33_ASAP7_75t_SL g1223 ( 
.A1(n_970),
.A2(n_49),
.B(n_51),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_973),
.B(n_54),
.Y(n_1224)
);

NAND2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1018),
.B(n_55),
.Y(n_1225)
);

INVxp67_ASAP7_75t_L g1226 ( 
.A(n_1121),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_951),
.Y(n_1227)
);

BUFx6f_ASAP7_75t_L g1228 ( 
.A(n_960),
.Y(n_1228)
);

HB1xp67_ASAP7_75t_L g1229 ( 
.A(n_984),
.Y(n_1229)
);

O2A1O1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1117),
.A2(n_57),
.B(n_58),
.C(n_60),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1012),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.Y(n_1231)
);

OR2x2_ASAP7_75t_L g1232 ( 
.A(n_1109),
.B(n_61),
.Y(n_1232)
);

OA22x2_ASAP7_75t_L g1233 ( 
.A1(n_964),
.A2(n_64),
.B1(n_65),
.B2(n_73),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_981),
.A2(n_566),
.B(n_564),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1020),
.A2(n_566),
.B(n_564),
.C(n_563),
.Y(n_1235)
);

NOR2xp33_ASAP7_75t_L g1236 ( 
.A(n_1114),
.B(n_64),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1106),
.B(n_74),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1106),
.B(n_75),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1100),
.B(n_77),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1009),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_960),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1007),
.A2(n_566),
.B(n_564),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_999),
.Y(n_1243)
);

BUFx6f_ASAP7_75t_L g1244 ( 
.A(n_960),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_R g1245 ( 
.A(n_1087),
.B(n_143),
.Y(n_1245)
);

INVxp67_ASAP7_75t_L g1246 ( 
.A(n_1107),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_996),
.B(n_79),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1000),
.A2(n_566),
.B(n_564),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1003),
.A2(n_566),
.B(n_564),
.C(n_563),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_998),
.B(n_81),
.Y(n_1250)
);

AOI21x1_ASAP7_75t_L g1251 ( 
.A1(n_961),
.A2(n_566),
.B(n_564),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_995),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_988),
.A2(n_564),
.B(n_563),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_982),
.B(n_83),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_982),
.B(n_83),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1096),
.B(n_563),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1087),
.B(n_92),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_1011),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1011),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1091),
.A2(n_563),
.B(n_549),
.C(n_111),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1038),
.Y(n_1261)
);

AO21x1_ASAP7_75t_L g1262 ( 
.A1(n_1073),
.A2(n_1086),
.B(n_1090),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_SL g1263 ( 
.A(n_1044),
.B(n_549),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_SL g1264 ( 
.A(n_1044),
.B(n_549),
.Y(n_1264)
);

NOR2x1p5_ASAP7_75t_SL g1265 ( 
.A(n_1044),
.B(n_97),
.Y(n_1265)
);

AO32x1_ASAP7_75t_L g1266 ( 
.A1(n_1075),
.A2(n_114),
.A3(n_115),
.B1(n_119),
.B2(n_124),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_958),
.A2(n_127),
.B(n_129),
.Y(n_1267)
);

BUFx10_ASAP7_75t_L g1268 ( 
.A(n_1051),
.Y(n_1268)
);

AO32x1_ASAP7_75t_L g1269 ( 
.A1(n_1080),
.A2(n_132),
.A3(n_133),
.B1(n_146),
.B2(n_147),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1040),
.A2(n_148),
.B(n_152),
.Y(n_1270)
);

A2O1A1Ixp33_ASAP7_75t_L g1271 ( 
.A1(n_1057),
.A2(n_153),
.B(n_158),
.C(n_162),
.Y(n_1271)
);

O2A1O1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_949),
.A2(n_169),
.B(n_199),
.C(n_202),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1047),
.A2(n_211),
.B(n_1049),
.Y(n_1273)
);

OAI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1122),
.A2(n_1039),
.B(n_955),
.Y(n_1274)
);

AOI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1251),
.A2(n_1055),
.B(n_1045),
.Y(n_1275)
);

O2A1O1Ixp33_ASAP7_75t_L g1276 ( 
.A1(n_1129),
.A2(n_1046),
.B(n_992),
.C(n_1034),
.Y(n_1276)
);

O2A1O1Ixp33_ASAP7_75t_SL g1277 ( 
.A1(n_1168),
.A2(n_1034),
.B(n_1046),
.C(n_992),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1215),
.A2(n_997),
.B(n_1108),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1138),
.Y(n_1279)
);

O2A1O1Ixp33_ASAP7_75t_SL g1280 ( 
.A1(n_1192),
.A2(n_1052),
.B(n_983),
.C(n_989),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1146),
.B(n_1101),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1139),
.A2(n_1078),
.B(n_1050),
.Y(n_1282)
);

INVxp67_ASAP7_75t_SL g1283 ( 
.A(n_1123),
.Y(n_1283)
);

AO31x2_ASAP7_75t_L g1284 ( 
.A1(n_1262),
.A2(n_1079),
.A3(n_1070),
.B(n_1069),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1130),
.B(n_1095),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1236),
.A2(n_1115),
.B(n_1058),
.C(n_1051),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1137),
.A2(n_1089),
.A3(n_1081),
.B(n_1071),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1151),
.B(n_1011),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_L g1289 ( 
.A1(n_1185),
.A2(n_1186),
.B(n_1207),
.C(n_1188),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1198),
.A2(n_1043),
.B(n_979),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_SL g1291 ( 
.A1(n_1254),
.A2(n_1052),
.B(n_983),
.C(n_989),
.Y(n_1291)
);

OAI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1190),
.A2(n_1005),
.B(n_990),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1162),
.Y(n_1293)
);

AO31x2_ASAP7_75t_L g1294 ( 
.A1(n_1235),
.A2(n_1208),
.A3(n_1212),
.B(n_1214),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1212),
.A2(n_1014),
.A3(n_1013),
.B(n_1016),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1124),
.A2(n_1115),
.B1(n_1031),
.B2(n_1006),
.Y(n_1296)
);

OA21x2_ASAP7_75t_L g1297 ( 
.A1(n_1242),
.A2(n_987),
.B(n_1019),
.Y(n_1297)
);

NOR2xp67_ASAP7_75t_SL g1298 ( 
.A(n_1156),
.B(n_1048),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1179),
.A2(n_1105),
.B(n_1032),
.C(n_1088),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1273),
.A2(n_1064),
.B(n_1030),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1263),
.A2(n_991),
.B(n_993),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1180),
.Y(n_1302)
);

AOI22xp5_ASAP7_75t_L g1303 ( 
.A1(n_1163),
.A2(n_1187),
.B1(n_1237),
.B2(n_1221),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1233),
.A2(n_1025),
.B1(n_1086),
.B2(n_1090),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1263),
.A2(n_1001),
.B(n_1004),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1242),
.A2(n_1048),
.B(n_1092),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1184),
.B(n_1048),
.Y(n_1307)
);

O2A1O1Ixp33_ASAP7_75t_SL g1308 ( 
.A1(n_1255),
.A2(n_1127),
.B(n_1181),
.C(n_1182),
.Y(n_1308)
);

A2O1A1Ixp33_ASAP7_75t_L g1309 ( 
.A1(n_1230),
.A2(n_1042),
.B(n_1097),
.C(n_1119),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1234),
.A2(n_1248),
.B(n_1144),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1154),
.B(n_1042),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1184),
.B(n_1044),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1194),
.B(n_1044),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1160),
.Y(n_1314)
);

AO31x2_ASAP7_75t_L g1315 ( 
.A1(n_1136),
.A2(n_1060),
.A3(n_1118),
.B(n_1120),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1204),
.Y(n_1316)
);

BUFx3_ASAP7_75t_L g1317 ( 
.A(n_1180),
.Y(n_1317)
);

O2A1O1Ixp5_ASAP7_75t_SL g1318 ( 
.A1(n_1231),
.A2(n_1094),
.B(n_1037),
.C(n_1053),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1264),
.A2(n_1145),
.B(n_1170),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1229),
.B(n_1044),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_1246),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1170),
.A2(n_1053),
.B(n_1037),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1232),
.A2(n_1112),
.B(n_1094),
.C(n_1111),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1267),
.A2(n_1093),
.B(n_1253),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1171),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1140),
.Y(n_1326)
);

BUFx10_ASAP7_75t_L g1327 ( 
.A(n_1189),
.Y(n_1327)
);

BUFx2_ASAP7_75t_L g1328 ( 
.A(n_1195),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1195),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1227),
.Y(n_1330)
);

AO31x2_ASAP7_75t_L g1331 ( 
.A1(n_1249),
.A2(n_1260),
.A3(n_1219),
.B(n_1216),
.Y(n_1331)
);

NOR2xp33_ASAP7_75t_L g1332 ( 
.A(n_1201),
.B(n_1196),
.Y(n_1332)
);

OAI21xp33_ASAP7_75t_L g1333 ( 
.A1(n_1197),
.A2(n_1205),
.B(n_1133),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1132),
.B(n_1141),
.Y(n_1334)
);

AOI221xp5_ASAP7_75t_SL g1335 ( 
.A1(n_1231),
.A2(n_1240),
.B1(n_1200),
.B2(n_1223),
.C(n_1224),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1252),
.Y(n_1336)
);

OAI22x1_ASAP7_75t_L g1337 ( 
.A1(n_1143),
.A2(n_1238),
.B1(n_1193),
.B2(n_1176),
.Y(n_1337)
);

AO21x2_ASAP7_75t_L g1338 ( 
.A1(n_1131),
.A2(n_1166),
.B(n_1152),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1261),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1270),
.A2(n_1272),
.B(n_1173),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1240),
.A2(n_1149),
.B(n_1178),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1125),
.B(n_1158),
.Y(n_1342)
);

A2O1A1Ixp33_ASAP7_75t_L g1343 ( 
.A1(n_1247),
.A2(n_1250),
.B(n_1222),
.C(n_1217),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1211),
.Y(n_1344)
);

CKINVDCx20_ASAP7_75t_R g1345 ( 
.A(n_1142),
.Y(n_1345)
);

OA21x2_ASAP7_75t_L g1346 ( 
.A1(n_1199),
.A2(n_1206),
.B(n_1271),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1239),
.Y(n_1347)
);

INVx2_ASAP7_75t_L g1348 ( 
.A(n_1135),
.Y(n_1348)
);

BUFx8_ASAP7_75t_L g1349 ( 
.A(n_1153),
.Y(n_1349)
);

INVxp67_ASAP7_75t_SL g1350 ( 
.A(n_1218),
.Y(n_1350)
);

AOI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1221),
.A2(n_1167),
.B1(n_1155),
.B2(n_1174),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1233),
.A2(n_1147),
.B1(n_1128),
.B2(n_1169),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1257),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1225),
.A2(n_1269),
.B(n_1266),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1257),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1148),
.A2(n_1173),
.B(n_1243),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1177),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1148),
.A2(n_1243),
.B(n_1256),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1191),
.Y(n_1359)
);

A2O1A1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1265),
.A2(n_1174),
.B(n_1169),
.C(n_1172),
.Y(n_1360)
);

AOI221x1_ASAP7_75t_L g1361 ( 
.A1(n_1172),
.A2(n_1159),
.B1(n_1175),
.B2(n_1165),
.C(n_1157),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1220),
.A2(n_1213),
.B(n_1202),
.Y(n_1362)
);

AOI221x1_ASAP7_75t_L g1363 ( 
.A1(n_1241),
.A2(n_1218),
.B1(n_1244),
.B2(n_1228),
.C(n_1210),
.Y(n_1363)
);

AO32x2_ASAP7_75t_L g1364 ( 
.A1(n_1241),
.A2(n_1258),
.A3(n_1259),
.B1(n_1268),
.B2(n_1266),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1126),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1266),
.A2(n_1269),
.B(n_1244),
.Y(n_1366)
);

A2O1A1Ixp33_ASAP7_75t_L g1367 ( 
.A1(n_1161),
.A2(n_1164),
.B(n_1209),
.C(n_1210),
.Y(n_1367)
);

AO31x2_ASAP7_75t_L g1368 ( 
.A1(n_1269),
.A2(n_1268),
.A3(n_1183),
.B(n_1191),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1191),
.A2(n_1226),
.B1(n_1203),
.B2(n_1209),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1126),
.B(n_1134),
.Y(n_1370)
);

NAND3x1_ASAP7_75t_L g1371 ( 
.A(n_1203),
.B(n_1245),
.C(n_1150),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1244),
.B(n_1218),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1228),
.A2(n_1134),
.B(n_1150),
.Y(n_1373)
);

A2O1A1Ixp33_ASAP7_75t_L g1374 ( 
.A1(n_1134),
.A2(n_1076),
.B(n_1066),
.C(n_1236),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1150),
.B(n_1228),
.Y(n_1375)
);

O2A1O1Ixp33_ASAP7_75t_L g1376 ( 
.A1(n_1129),
.A2(n_857),
.B(n_1076),
.C(n_1066),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1124),
.B(n_857),
.Y(n_1377)
);

AOI21xp5_ASAP7_75t_L g1378 ( 
.A1(n_1263),
.A2(n_962),
.B(n_943),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1160),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1129),
.A2(n_857),
.B(n_1076),
.C(n_1066),
.Y(n_1380)
);

O2A1O1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1129),
.A2(n_857),
.B(n_1076),
.C(n_1066),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1156),
.Y(n_1382)
);

INVxp67_ASAP7_75t_SL g1383 ( 
.A(n_1123),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1146),
.B(n_956),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1146),
.B(n_956),
.Y(n_1385)
);

BUFx2_ASAP7_75t_L g1386 ( 
.A(n_1138),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1146),
.B(n_956),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1263),
.A2(n_962),
.B(n_943),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1122),
.A2(n_956),
.B(n_986),
.Y(n_1389)
);

AOI221xp5_ASAP7_75t_SL g1390 ( 
.A1(n_1231),
.A2(n_1240),
.B1(n_1200),
.B2(n_1230),
.C(n_1066),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1160),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1273),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1138),
.Y(n_1393)
);

OAI21xp5_ASAP7_75t_L g1394 ( 
.A1(n_1122),
.A2(n_956),
.B(n_986),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1154),
.B(n_952),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1162),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1162),
.Y(n_1397)
);

OAI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1122),
.A2(n_956),
.B(n_986),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1191),
.B(n_1056),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1263),
.A2(n_962),
.B(n_943),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1162),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1263),
.A2(n_962),
.B(n_943),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1146),
.B(n_956),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_SL g1404 ( 
.A(n_1124),
.B(n_1017),
.Y(n_1404)
);

AOI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1129),
.A2(n_1076),
.B1(n_1066),
.B2(n_872),
.Y(n_1405)
);

A2O1A1Ixp33_ASAP7_75t_L g1406 ( 
.A1(n_1236),
.A2(n_1076),
.B(n_1066),
.C(n_956),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1236),
.A2(n_1076),
.B(n_1066),
.C(n_956),
.Y(n_1407)
);

AO21x2_ASAP7_75t_L g1408 ( 
.A1(n_1242),
.A2(n_1262),
.B(n_1251),
.Y(n_1408)
);

NAND2x1p5_ASAP7_75t_L g1409 ( 
.A(n_1191),
.B(n_1056),
.Y(n_1409)
);

BUFx12f_ASAP7_75t_L g1410 ( 
.A(n_1156),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1251),
.A2(n_1234),
.B(n_1273),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1273),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1273),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_SL g1414 ( 
.A(n_1124),
.B(n_1017),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1160),
.Y(n_1415)
);

NOR2x1_ASAP7_75t_SL g1416 ( 
.A(n_1191),
.B(n_978),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1263),
.A2(n_962),
.B(n_943),
.Y(n_1417)
);

NOR4xp25_ASAP7_75t_L g1418 ( 
.A(n_1231),
.B(n_1200),
.C(n_1240),
.D(n_1230),
.Y(n_1418)
);

INVx4_ASAP7_75t_L g1419 ( 
.A(n_1180),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1162),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1273),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1263),
.A2(n_962),
.B(n_943),
.Y(n_1422)
);

AO31x2_ASAP7_75t_L g1423 ( 
.A1(n_1262),
.A2(n_1137),
.A3(n_944),
.B(n_1235),
.Y(n_1423)
);

AO31x2_ASAP7_75t_L g1424 ( 
.A1(n_1262),
.A2(n_1137),
.A3(n_944),
.B(n_1235),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1273),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1273),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1122),
.A2(n_956),
.B(n_986),
.Y(n_1427)
);

A2O1A1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1236),
.A2(n_1076),
.B(n_1066),
.C(n_956),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1236),
.A2(n_1076),
.B(n_1066),
.C(n_956),
.Y(n_1429)
);

O2A1O1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1129),
.A2(n_857),
.B(n_1076),
.C(n_1066),
.Y(n_1430)
);

NOR2xp33_ASAP7_75t_L g1431 ( 
.A(n_1124),
.B(n_857),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1180),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1215),
.A2(n_1251),
.B(n_1273),
.Y(n_1433)
);

INVx3_ASAP7_75t_L g1434 ( 
.A(n_1191),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1191),
.B(n_1056),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1263),
.A2(n_962),
.B(n_943),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1162),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_SL g1438 ( 
.A1(n_1405),
.A2(n_1303),
.B1(n_1377),
.B2(n_1431),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1293),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1410),
.Y(n_1440)
);

CKINVDCx11_ASAP7_75t_R g1441 ( 
.A(n_1345),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1352),
.A2(n_1342),
.B1(n_1337),
.B2(n_1395),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1328),
.Y(n_1443)
);

CKINVDCx20_ASAP7_75t_R g1444 ( 
.A(n_1382),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1329),
.Y(n_1445)
);

AOI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1341),
.A2(n_1406),
.B1(n_1407),
.B2(n_1428),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_SL g1447 ( 
.A1(n_1352),
.A2(n_1387),
.B1(n_1385),
.B2(n_1384),
.Y(n_1447)
);

CKINVDCx11_ASAP7_75t_R g1448 ( 
.A(n_1365),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1384),
.B(n_1385),
.Y(n_1449)
);

BUFx4_ASAP7_75t_SL g1450 ( 
.A(n_1317),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1387),
.A2(n_1403),
.B1(n_1333),
.B2(n_1351),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1403),
.A2(n_1332),
.B1(n_1347),
.B2(n_1344),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1396),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1316),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1397),
.Y(n_1455)
);

BUFx12f_ASAP7_75t_L g1456 ( 
.A(n_1302),
.Y(n_1456)
);

BUFx8_ASAP7_75t_SL g1457 ( 
.A(n_1302),
.Y(n_1457)
);

INVx1_ASAP7_75t_SL g1458 ( 
.A(n_1316),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1341),
.A2(n_1429),
.B1(n_1343),
.B2(n_1374),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1404),
.A2(n_1414),
.B1(n_1390),
.B2(n_1289),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_SL g1461 ( 
.A1(n_1327),
.A2(n_1321),
.B1(n_1292),
.B2(n_1290),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1432),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1327),
.A2(n_1292),
.B1(n_1357),
.B2(n_1290),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1376),
.A2(n_1430),
.B1(n_1381),
.B2(n_1380),
.Y(n_1464)
);

INVx1_ASAP7_75t_SL g1465 ( 
.A(n_1386),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1281),
.A2(n_1437),
.B1(n_1401),
.B2(n_1420),
.Y(n_1466)
);

INVx4_ASAP7_75t_L g1467 ( 
.A(n_1432),
.Y(n_1467)
);

AOI22x1_ASAP7_75t_SL g1468 ( 
.A1(n_1419),
.A2(n_1353),
.B1(n_1355),
.B2(n_1283),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1326),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1314),
.A2(n_1330),
.B1(n_1325),
.B2(n_1379),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1339),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1279),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1391),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1415),
.A2(n_1281),
.B1(n_1296),
.B2(n_1348),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1346),
.A2(n_1418),
.B1(n_1388),
.B2(n_1422),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1383),
.B(n_1393),
.Y(n_1476)
);

INVx2_ASAP7_75t_SL g1477 ( 
.A(n_1349),
.Y(n_1477)
);

CKINVDCx11_ASAP7_75t_R g1478 ( 
.A(n_1419),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1312),
.A2(n_1311),
.B1(n_1285),
.B2(n_1304),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1307),
.B(n_1378),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1360),
.A2(n_1286),
.B1(n_1436),
.B2(n_1400),
.Y(n_1481)
);

AOI22xp33_ASAP7_75t_L g1482 ( 
.A1(n_1312),
.A2(n_1285),
.B1(n_1320),
.B2(n_1307),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_1349),
.Y(n_1483)
);

CKINVDCx11_ASAP7_75t_R g1484 ( 
.A(n_1375),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1402),
.A2(n_1417),
.B1(n_1398),
.B2(n_1427),
.Y(n_1485)
);

AOI22xp33_ASAP7_75t_L g1486 ( 
.A1(n_1389),
.A2(n_1394),
.B1(n_1427),
.B2(n_1398),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1288),
.Y(n_1487)
);

OAI21xp5_ASAP7_75t_SL g1488 ( 
.A1(n_1354),
.A2(n_1389),
.B(n_1394),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1334),
.Y(n_1489)
);

OAI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1313),
.A2(n_1320),
.B1(n_1390),
.B2(n_1322),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1372),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1370),
.Y(n_1492)
);

OAI21xp33_ASAP7_75t_L g1493 ( 
.A1(n_1418),
.A2(n_1367),
.B(n_1299),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1372),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_SL g1495 ( 
.A1(n_1346),
.A2(n_1335),
.B1(n_1274),
.B2(n_1313),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_SL g1496 ( 
.A1(n_1335),
.A2(n_1274),
.B1(n_1369),
.B2(n_1338),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1369),
.A2(n_1338),
.B1(n_1399),
.B2(n_1359),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1356),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1350),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1358),
.Y(n_1500)
);

INVxp67_ASAP7_75t_SL g1501 ( 
.A(n_1297),
.Y(n_1501)
);

OAI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1361),
.A2(n_1297),
.B1(n_1366),
.B2(n_1363),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1359),
.Y(n_1503)
);

INVx6_ASAP7_75t_L g1504 ( 
.A(n_1371),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1434),
.A2(n_1408),
.B1(n_1319),
.B2(n_1435),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1434),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1409),
.B(n_1373),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1277),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_SL g1509 ( 
.A1(n_1416),
.A2(n_1364),
.B1(n_1408),
.B2(n_1340),
.Y(n_1509)
);

CKINVDCx6p67_ASAP7_75t_R g1510 ( 
.A(n_1308),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1276),
.Y(n_1511)
);

AOI22xp33_ASAP7_75t_SL g1512 ( 
.A1(n_1364),
.A2(n_1306),
.B1(n_1282),
.B2(n_1368),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1282),
.A2(n_1305),
.B1(n_1301),
.B2(n_1362),
.Y(n_1513)
);

INVx6_ASAP7_75t_L g1514 ( 
.A(n_1280),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1324),
.A2(n_1300),
.B1(n_1278),
.B2(n_1310),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1423),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1364),
.A2(n_1295),
.B1(n_1318),
.B2(n_1294),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1291),
.Y(n_1518)
);

INVx6_ASAP7_75t_L g1519 ( 
.A(n_1323),
.Y(n_1519)
);

BUFx6f_ASAP7_75t_L g1520 ( 
.A(n_1275),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1309),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1295),
.A2(n_1294),
.B1(n_1423),
.B2(n_1424),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1411),
.A2(n_1294),
.B1(n_1424),
.B2(n_1331),
.Y(n_1523)
);

BUFx8_ASAP7_75t_L g1524 ( 
.A(n_1424),
.Y(n_1524)
);

BUFx12f_ASAP7_75t_L g1525 ( 
.A(n_1287),
.Y(n_1525)
);

AOI22xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1295),
.A2(n_1413),
.B1(n_1426),
.B2(n_1425),
.Y(n_1526)
);

BUFx2_ASAP7_75t_SL g1527 ( 
.A(n_1284),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1315),
.Y(n_1528)
);

BUFx3_ASAP7_75t_L g1529 ( 
.A(n_1315),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1392),
.Y(n_1530)
);

BUFx3_ASAP7_75t_L g1531 ( 
.A(n_1412),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1421),
.A2(n_1433),
.B1(n_872),
.B2(n_856),
.Y(n_1532)
);

BUFx8_ASAP7_75t_L g1533 ( 
.A(n_1328),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1352),
.A2(n_1212),
.B1(n_554),
.B2(n_550),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1382),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1352),
.A2(n_872),
.B1(n_856),
.B2(n_1066),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1293),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1406),
.A2(n_1407),
.B1(n_1429),
.B2(n_1428),
.Y(n_1539)
);

INVxp67_ASAP7_75t_SL g1540 ( 
.A(n_1288),
.Y(n_1540)
);

OAI21xp33_ASAP7_75t_L g1541 ( 
.A1(n_1406),
.A2(n_1428),
.B(n_1407),
.Y(n_1541)
);

BUFx12f_ASAP7_75t_L g1542 ( 
.A(n_1365),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1352),
.A2(n_1212),
.B1(n_554),
.B2(n_550),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1352),
.A2(n_872),
.B1(n_856),
.B2(n_1066),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1352),
.A2(n_872),
.B1(n_856),
.B2(n_1066),
.Y(n_1545)
);

BUFx8_ASAP7_75t_L g1546 ( 
.A(n_1328),
.Y(n_1546)
);

INVx6_ASAP7_75t_L g1547 ( 
.A(n_1302),
.Y(n_1547)
);

CKINVDCx6p67_ASAP7_75t_R g1548 ( 
.A(n_1317),
.Y(n_1548)
);

OAI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1406),
.A2(n_1428),
.B(n_1407),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1293),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1293),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1336),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1406),
.A2(n_1407),
.B1(n_1429),
.B2(n_1428),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_L g1554 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1555)
);

BUFx3_ASAP7_75t_L g1556 ( 
.A(n_1410),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1406),
.A2(n_1407),
.B1(n_1429),
.B2(n_1428),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1293),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_L g1560 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1293),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_SL g1562 ( 
.A1(n_1352),
.A2(n_1212),
.B1(n_554),
.B2(n_550),
.Y(n_1562)
);

BUFx10_ASAP7_75t_L g1563 ( 
.A(n_1382),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_SL g1564 ( 
.A1(n_1405),
.A2(n_1341),
.B(n_1406),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1384),
.B(n_1385),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1566)
);

BUFx6f_ASAP7_75t_L g1567 ( 
.A(n_1365),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1384),
.B(n_1385),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1298),
.B(n_1191),
.Y(n_1569)
);

INVx5_ASAP7_75t_L g1570 ( 
.A(n_1359),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1293),
.Y(n_1573)
);

INVx6_ASAP7_75t_L g1574 ( 
.A(n_1302),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1293),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1382),
.Y(n_1576)
);

NAND2x1p5_ASAP7_75t_L g1577 ( 
.A(n_1298),
.B(n_1191),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1293),
.Y(n_1578)
);

INVx6_ASAP7_75t_L g1579 ( 
.A(n_1302),
.Y(n_1579)
);

CKINVDCx11_ASAP7_75t_R g1580 ( 
.A(n_1410),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1395),
.B(n_957),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1423),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1405),
.A2(n_1352),
.B1(n_952),
.B2(n_872),
.Y(n_1583)
);

CKINVDCx11_ASAP7_75t_R g1584 ( 
.A(n_1410),
.Y(n_1584)
);

INVxp67_ASAP7_75t_L g1585 ( 
.A(n_1476),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1540),
.Y(n_1586)
);

INVx6_ASAP7_75t_L g1587 ( 
.A(n_1456),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1472),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1540),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1499),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1454),
.Y(n_1591)
);

AO21x2_ASAP7_75t_L g1592 ( 
.A1(n_1502),
.A2(n_1528),
.B(n_1481),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1487),
.Y(n_1593)
);

NOR2xp33_ASAP7_75t_SL g1594 ( 
.A(n_1542),
.B(n_1457),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1452),
.B(n_1449),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1480),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1458),
.Y(n_1597)
);

OAI21x1_ASAP7_75t_L g1598 ( 
.A1(n_1515),
.A2(n_1513),
.B(n_1523),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1452),
.B(n_1565),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1498),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1504),
.B(n_1527),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1530),
.Y(n_1602)
);

INVx3_ASAP7_75t_L g1603 ( 
.A(n_1531),
.Y(n_1603)
);

CKINVDCx5p33_ASAP7_75t_R g1604 ( 
.A(n_1441),
.Y(n_1604)
);

INVx5_ASAP7_75t_L g1605 ( 
.A(n_1514),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1500),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1486),
.B(n_1439),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1516),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1564),
.A2(n_1554),
.B1(n_1583),
.B2(n_1536),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1582),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1568),
.B(n_1489),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1582),
.Y(n_1612)
);

OAI21x1_ASAP7_75t_L g1613 ( 
.A1(n_1485),
.A2(n_1505),
.B(n_1517),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1465),
.B(n_1451),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1518),
.Y(n_1615)
);

INVx2_ASAP7_75t_SL g1616 ( 
.A(n_1570),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1486),
.A2(n_1553),
.B(n_1539),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1525),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1511),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1453),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1455),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1529),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1505),
.A2(n_1517),
.B(n_1508),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1538),
.Y(n_1624)
);

INVx4_ASAP7_75t_L g1625 ( 
.A(n_1504),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1550),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1501),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1551),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1501),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1524),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1520),
.Y(n_1631)
);

INVxp33_ASAP7_75t_L g1632 ( 
.A(n_1469),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1488),
.A2(n_1493),
.B(n_1549),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_L g1634 ( 
.A1(n_1532),
.A2(n_1507),
.B(n_1557),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1558),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1561),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1471),
.Y(n_1637)
);

AO21x2_ASAP7_75t_L g1638 ( 
.A1(n_1502),
.A2(n_1490),
.B(n_1446),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1573),
.Y(n_1639)
);

NAND2x1p5_ASAP7_75t_L g1640 ( 
.A(n_1570),
.B(n_1518),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1575),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1491),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1524),
.Y(n_1643)
);

AOI22xp33_ASAP7_75t_L g1644 ( 
.A1(n_1534),
.A2(n_1562),
.B1(n_1543),
.B2(n_1566),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1578),
.Y(n_1645)
);

OA21x2_ASAP7_75t_L g1646 ( 
.A1(n_1541),
.A2(n_1463),
.B(n_1459),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1451),
.B(n_1447),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1519),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1490),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1495),
.B(n_1496),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1494),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1522),
.Y(n_1652)
);

OAI21x1_ASAP7_75t_L g1653 ( 
.A1(n_1497),
.A2(n_1463),
.B(n_1482),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1519),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1522),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1466),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1447),
.B(n_1466),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1495),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1460),
.B(n_1581),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1519),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1442),
.B(n_1536),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1438),
.Y(n_1662)
);

CKINVDCx8_ASAP7_75t_R g1663 ( 
.A(n_1483),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1552),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1473),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1461),
.B(n_1554),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_L g1667 ( 
.A1(n_1534),
.A2(n_1562),
.B1(n_1543),
.B2(n_1583),
.Y(n_1667)
);

OA21x2_ASAP7_75t_L g1668 ( 
.A1(n_1479),
.A2(n_1506),
.B(n_1503),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1496),
.B(n_1512),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1521),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1512),
.Y(n_1671)
);

HB1xp67_ASAP7_75t_L g1672 ( 
.A(n_1464),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1461),
.B(n_1559),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1475),
.B(n_1509),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1509),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1475),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1555),
.B(n_1571),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1510),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1570),
.Y(n_1679)
);

OAI21x1_ASAP7_75t_L g1680 ( 
.A1(n_1569),
.A2(n_1577),
.B(n_1474),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1492),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1555),
.B(n_1560),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1559),
.B(n_1572),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1560),
.A2(n_1572),
.B1(n_1571),
.B2(n_1566),
.Y(n_1684)
);

AOI22xp33_ASAP7_75t_L g1685 ( 
.A1(n_1537),
.A2(n_1545),
.B1(n_1544),
.B2(n_1470),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1526),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1468),
.Y(n_1687)
);

CKINVDCx9p33_ASAP7_75t_R g1688 ( 
.A(n_1450),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1567),
.B(n_1484),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1567),
.B(n_1462),
.Y(n_1690)
);

INVx3_ASAP7_75t_L g1691 ( 
.A(n_1467),
.Y(n_1691)
);

CKINVDCx12_ASAP7_75t_R g1692 ( 
.A(n_1450),
.Y(n_1692)
);

AOI22xp33_ASAP7_75t_L g1693 ( 
.A1(n_1478),
.A2(n_1574),
.B1(n_1579),
.B2(n_1547),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1547),
.Y(n_1694)
);

HB1xp67_ASAP7_75t_L g1695 ( 
.A(n_1574),
.Y(n_1695)
);

AND2x6_ASAP7_75t_L g1696 ( 
.A(n_1440),
.B(n_1556),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1467),
.Y(n_1697)
);

AOI21x1_ASAP7_75t_L g1698 ( 
.A1(n_1477),
.A2(n_1548),
.B(n_1546),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1533),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1533),
.Y(n_1700)
);

INVx3_ASAP7_75t_L g1701 ( 
.A(n_1563),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1546),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1563),
.Y(n_1703)
);

AOI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1662),
.A2(n_1535),
.B(n_1576),
.C(n_1448),
.Y(n_1704)
);

A2O1A1Ixp33_ASAP7_75t_L g1705 ( 
.A1(n_1609),
.A2(n_1444),
.B(n_1580),
.C(n_1584),
.Y(n_1705)
);

OR2x6_ASAP7_75t_L g1706 ( 
.A(n_1601),
.B(n_1443),
.Y(n_1706)
);

NOR2x1_ASAP7_75t_SL g1707 ( 
.A(n_1605),
.B(n_1445),
.Y(n_1707)
);

INVx4_ASAP7_75t_L g1708 ( 
.A(n_1678),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1585),
.B(n_1642),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1609),
.A2(n_1617),
.B(n_1647),
.C(n_1673),
.Y(n_1710)
);

INVx3_ASAP7_75t_L g1711 ( 
.A(n_1679),
.Y(n_1711)
);

OA21x2_ASAP7_75t_L g1712 ( 
.A1(n_1598),
.A2(n_1613),
.B(n_1623),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1672),
.A2(n_1644),
.B1(n_1667),
.B2(n_1684),
.Y(n_1713)
);

O2A1O1Ixp33_ASAP7_75t_SL g1714 ( 
.A1(n_1678),
.A2(n_1657),
.B(n_1666),
.C(n_1700),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1637),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1690),
.B(n_1607),
.Y(n_1716)
);

OAI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1646),
.A2(n_1633),
.B(n_1650),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1627),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1611),
.B(n_1595),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1637),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1607),
.B(n_1591),
.Y(n_1721)
);

OAI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1633),
.A2(n_1650),
.B(n_1646),
.C(n_1686),
.Y(n_1722)
);

AO32x2_ASAP7_75t_L g1723 ( 
.A1(n_1590),
.A2(n_1625),
.A3(n_1616),
.B1(n_1655),
.B2(n_1652),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1597),
.B(n_1588),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1646),
.A2(n_1633),
.B(n_1669),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1689),
.B(n_1669),
.Y(n_1726)
);

OA21x2_ASAP7_75t_L g1727 ( 
.A1(n_1613),
.A2(n_1623),
.B(n_1634),
.Y(n_1727)
);

AO32x1_ASAP7_75t_L g1728 ( 
.A1(n_1674),
.A2(n_1590),
.A3(n_1671),
.B1(n_1675),
.B2(n_1676),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1689),
.B(n_1674),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1646),
.A2(n_1633),
.B(n_1638),
.Y(n_1730)
);

O2A1O1Ixp33_ASAP7_75t_L g1731 ( 
.A1(n_1599),
.A2(n_1614),
.B(n_1676),
.C(n_1658),
.Y(n_1731)
);

OAI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1658),
.A2(n_1653),
.B(n_1649),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1645),
.Y(n_1733)
);

A2O1A1Ixp33_ASAP7_75t_L g1734 ( 
.A1(n_1677),
.A2(n_1683),
.B(n_1653),
.C(n_1682),
.Y(n_1734)
);

OAI22xp33_ASAP7_75t_SL g1735 ( 
.A1(n_1670),
.A2(n_1661),
.B1(n_1671),
.B2(n_1675),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1670),
.B(n_1702),
.Y(n_1736)
);

CKINVDCx5p33_ASAP7_75t_R g1737 ( 
.A(n_1688),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1596),
.B(n_1651),
.Y(n_1738)
);

CKINVDCx11_ASAP7_75t_R g1739 ( 
.A(n_1663),
.Y(n_1739)
);

A2O1A1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1677),
.A2(n_1683),
.B(n_1685),
.C(n_1661),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1627),
.Y(n_1741)
);

INVxp67_ASAP7_75t_L g1742 ( 
.A(n_1586),
.Y(n_1742)
);

CKINVDCx20_ASAP7_75t_R g1743 ( 
.A(n_1692),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1702),
.B(n_1681),
.Y(n_1744)
);

CKINVDCx5p33_ASAP7_75t_R g1745 ( 
.A(n_1692),
.Y(n_1745)
);

O2A1O1Ixp33_ASAP7_75t_SL g1746 ( 
.A1(n_1678),
.A2(n_1700),
.B(n_1699),
.C(n_1615),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1596),
.B(n_1651),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1620),
.B(n_1621),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1593),
.B(n_1624),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1626),
.B(n_1628),
.Y(n_1750)
);

OAI22xp5_ASAP7_75t_L g1751 ( 
.A1(n_1678),
.A2(n_1654),
.B1(n_1659),
.B2(n_1693),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1628),
.B(n_1635),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_L g1753 ( 
.A1(n_1640),
.A2(n_1680),
.B(n_1619),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1618),
.B(n_1630),
.Y(n_1754)
);

O2A1O1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1649),
.A2(n_1638),
.B(n_1686),
.C(n_1654),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1593),
.B(n_1635),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1636),
.B(n_1639),
.Y(n_1757)
);

A2O1A1Ixp33_ASAP7_75t_L g1758 ( 
.A1(n_1654),
.A2(n_1687),
.B(n_1660),
.C(n_1652),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1641),
.B(n_1586),
.Y(n_1759)
);

O2A1O1Ixp33_ASAP7_75t_SL g1760 ( 
.A1(n_1615),
.A2(n_1632),
.B(n_1701),
.C(n_1703),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1589),
.B(n_1648),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1695),
.B(n_1703),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1604),
.Y(n_1763)
);

AND2x6_ASAP7_75t_L g1764 ( 
.A(n_1643),
.B(n_1679),
.Y(n_1764)
);

NOR2xp33_ASAP7_75t_L g1765 ( 
.A(n_1701),
.B(n_1619),
.Y(n_1765)
);

O2A1O1Ixp33_ASAP7_75t_SL g1766 ( 
.A1(n_1701),
.A2(n_1616),
.B(n_1691),
.C(n_1697),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1715),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1720),
.Y(n_1768)
);

AND2x4_ASAP7_75t_L g1769 ( 
.A(n_1764),
.B(n_1627),
.Y(n_1769)
);

AOI22xp33_ASAP7_75t_L g1770 ( 
.A1(n_1725),
.A2(n_1655),
.B1(n_1656),
.B2(n_1592),
.Y(n_1770)
);

AOI22xp33_ASAP7_75t_L g1771 ( 
.A1(n_1717),
.A2(n_1592),
.B1(n_1643),
.B2(n_1622),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1733),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1742),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1742),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1629),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1716),
.B(n_1629),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1718),
.Y(n_1777)
);

OR2x2_ASAP7_75t_L g1778 ( 
.A(n_1721),
.B(n_1610),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1712),
.B(n_1629),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1712),
.B(n_1606),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1718),
.Y(n_1781)
);

AND2x2_ASAP7_75t_L g1782 ( 
.A(n_1712),
.B(n_1606),
.Y(n_1782)
);

AND2x4_ASAP7_75t_L g1783 ( 
.A(n_1764),
.B(n_1603),
.Y(n_1783)
);

INVx1_ASAP7_75t_SL g1784 ( 
.A(n_1762),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1748),
.B(n_1600),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1741),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1741),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1747),
.B(n_1610),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1713),
.A2(n_1643),
.B1(n_1668),
.B2(n_1625),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1759),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1719),
.B(n_1612),
.Y(n_1791)
);

OR2x2_ASAP7_75t_L g1792 ( 
.A(n_1709),
.B(n_1612),
.Y(n_1792)
);

OAI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1710),
.A2(n_1640),
.B1(n_1625),
.B2(n_1619),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1750),
.B(n_1631),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_1631),
.Y(n_1795)
);

INVxp67_ASAP7_75t_SL g1796 ( 
.A(n_1761),
.Y(n_1796)
);

NOR2xp33_ASAP7_75t_L g1797 ( 
.A(n_1737),
.B(n_1698),
.Y(n_1797)
);

OAI21xp33_ASAP7_75t_L g1798 ( 
.A1(n_1710),
.A2(n_1594),
.B(n_1694),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1706),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1757),
.B(n_1668),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1749),
.Y(n_1801)
);

NAND2x1_ASAP7_75t_L g1802 ( 
.A(n_1706),
.B(n_1602),
.Y(n_1802)
);

INVxp67_ASAP7_75t_SL g1803 ( 
.A(n_1730),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1756),
.Y(n_1804)
);

BUFx3_ASAP7_75t_L g1805 ( 
.A(n_1764),
.Y(n_1805)
);

AOI222xp33_ASAP7_75t_L g1806 ( 
.A1(n_1740),
.A2(n_1696),
.B1(n_1665),
.B2(n_1608),
.C1(n_1664),
.C2(n_1587),
.Y(n_1806)
);

INVxp67_ASAP7_75t_L g1807 ( 
.A(n_1724),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1805),
.B(n_1706),
.Y(n_1808)
);

INVx1_ASAP7_75t_SL g1809 ( 
.A(n_1792),
.Y(n_1809)
);

OR2x2_ASAP7_75t_L g1810 ( 
.A(n_1778),
.B(n_1732),
.Y(n_1810)
);

AOI31xp33_ASAP7_75t_L g1811 ( 
.A1(n_1789),
.A2(n_1705),
.A3(n_1745),
.B(n_1714),
.Y(n_1811)
);

BUFx2_ASAP7_75t_L g1812 ( 
.A(n_1805),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1767),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1779),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1770),
.A2(n_1735),
.B1(n_1729),
.B2(n_1726),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1779),
.Y(n_1816)
);

AND2x4_ASAP7_75t_L g1817 ( 
.A(n_1805),
.B(n_1783),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1796),
.B(n_1773),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1780),
.Y(n_1819)
);

NOR2xp67_ASAP7_75t_L g1820 ( 
.A(n_1800),
.B(n_1708),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1767),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1768),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1777),
.Y(n_1823)
);

INVx4_ASAP7_75t_L g1824 ( 
.A(n_1799),
.Y(n_1824)
);

BUFx2_ASAP7_75t_L g1825 ( 
.A(n_1799),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1776),
.B(n_1723),
.Y(n_1826)
);

CKINVDCx20_ASAP7_75t_R g1827 ( 
.A(n_1784),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1776),
.B(n_1723),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1796),
.B(n_1734),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1768),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1797),
.B(n_1739),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1773),
.B(n_1734),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1783),
.B(n_1753),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1774),
.B(n_1722),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1777),
.Y(n_1835)
);

AOI211xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1798),
.A2(n_1705),
.B(n_1714),
.C(n_1746),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1772),
.Y(n_1837)
);

AOI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1803),
.A2(n_1728),
.B(n_1755),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_SL g1839 ( 
.A1(n_1803),
.A2(n_1751),
.B1(n_1728),
.B2(n_1727),
.Y(n_1839)
);

AOI221xp5_ASAP7_75t_L g1840 ( 
.A1(n_1798),
.A2(n_1740),
.B1(n_1731),
.B2(n_1758),
.C(n_1760),
.Y(n_1840)
);

OR2x2_ASAP7_75t_SL g1841 ( 
.A(n_1792),
.B(n_1587),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1778),
.B(n_1744),
.Y(n_1842)
);

OAI221xp5_ASAP7_75t_SL g1843 ( 
.A1(n_1789),
.A2(n_1806),
.B1(n_1771),
.B2(n_1758),
.C(n_1807),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1807),
.B(n_1723),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1776),
.B(n_1723),
.Y(n_1845)
);

INVxp67_ASAP7_75t_SL g1846 ( 
.A(n_1781),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1775),
.Y(n_1847)
);

AND2x2_ASAP7_75t_L g1848 ( 
.A(n_1794),
.B(n_1795),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1801),
.B(n_1804),
.Y(n_1849)
);

BUFx6f_ASAP7_75t_L g1850 ( 
.A(n_1802),
.Y(n_1850)
);

OAI21x1_ASAP7_75t_SL g1851 ( 
.A1(n_1793),
.A2(n_1707),
.B(n_1708),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1801),
.B(n_1711),
.Y(n_1852)
);

INVxp67_ASAP7_75t_SL g1853 ( 
.A(n_1781),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1813),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1844),
.B(n_1786),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1844),
.B(n_1786),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1813),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1826),
.B(n_1787),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1847),
.B(n_1849),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1821),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1819),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1821),
.Y(n_1862)
);

INVx3_ASAP7_75t_L g1863 ( 
.A(n_1850),
.Y(n_1863)
);

INVx2_ASAP7_75t_L g1864 ( 
.A(n_1819),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1826),
.B(n_1787),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1826),
.B(n_1828),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1828),
.B(n_1780),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1847),
.B(n_1804),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1849),
.B(n_1780),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1819),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1834),
.B(n_1782),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1828),
.B(n_1782),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_L g1873 ( 
.A(n_1831),
.B(n_1743),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1845),
.B(n_1782),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1818),
.B(n_1800),
.Y(n_1875)
);

OR2x2_ASAP7_75t_L g1876 ( 
.A(n_1818),
.B(n_1775),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1845),
.B(n_1848),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1814),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1834),
.B(n_1791),
.Y(n_1879)
);

OR2x2_ASAP7_75t_L g1880 ( 
.A(n_1832),
.B(n_1791),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1832),
.B(n_1788),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1845),
.B(n_1785),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1814),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1848),
.B(n_1785),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1809),
.B(n_1788),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1848),
.B(n_1785),
.Y(n_1886)
);

AND2x4_ASAP7_75t_L g1887 ( 
.A(n_1817),
.B(n_1769),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1822),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1814),
.Y(n_1889)
);

BUFx2_ASAP7_75t_L g1890 ( 
.A(n_1850),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1822),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1816),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1830),
.Y(n_1893)
);

INVxp67_ASAP7_75t_SL g1894 ( 
.A(n_1829),
.Y(n_1894)
);

NOR2xp33_ASAP7_75t_L g1895 ( 
.A(n_1824),
.B(n_1743),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1809),
.B(n_1830),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1837),
.B(n_1790),
.Y(n_1897)
);

INVx3_ASAP7_75t_L g1898 ( 
.A(n_1850),
.Y(n_1898)
);

BUFx2_ASAP7_75t_L g1899 ( 
.A(n_1854),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1854),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1894),
.B(n_1810),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1894),
.B(n_1880),
.Y(n_1902)
);

AOI32xp33_ASAP7_75t_L g1903 ( 
.A1(n_1866),
.A2(n_1836),
.A3(n_1840),
.B1(n_1839),
.B2(n_1829),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1895),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1861),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1877),
.B(n_1817),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1879),
.A2(n_1811),
.B1(n_1843),
.B2(n_1840),
.Y(n_1907)
);

OR2x2_ASAP7_75t_L g1908 ( 
.A(n_1881),
.B(n_1810),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1861),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1881),
.B(n_1852),
.Y(n_1910)
);

AND2x4_ASAP7_75t_L g1911 ( 
.A(n_1887),
.B(n_1833),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1877),
.B(n_1817),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1854),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1877),
.B(n_1817),
.Y(n_1914)
);

INVx2_ASAP7_75t_L g1915 ( 
.A(n_1861),
.Y(n_1915)
);

OR2x2_ASAP7_75t_L g1916 ( 
.A(n_1881),
.B(n_1852),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1857),
.Y(n_1917)
);

NOR2xp67_ASAP7_75t_L g1918 ( 
.A(n_1887),
.B(n_1863),
.Y(n_1918)
);

AND2x2_ASAP7_75t_L g1919 ( 
.A(n_1866),
.B(n_1825),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1879),
.Y(n_1920)
);

HB1xp67_ASAP7_75t_L g1921 ( 
.A(n_1879),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1861),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1880),
.B(n_1823),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_SL g1924 ( 
.A(n_1895),
.B(n_1808),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1880),
.B(n_1884),
.Y(n_1925)
);

NOR2x1_ASAP7_75t_L g1926 ( 
.A(n_1863),
.B(n_1824),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1857),
.Y(n_1927)
);

INVx2_ASAP7_75t_SL g1928 ( 
.A(n_1887),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1857),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1859),
.B(n_1823),
.Y(n_1930)
);

AOI21xp33_ASAP7_75t_SL g1931 ( 
.A1(n_1873),
.A2(n_1811),
.B(n_1737),
.Y(n_1931)
);

OAI211xp5_ASAP7_75t_L g1932 ( 
.A1(n_1871),
.A2(n_1836),
.B(n_1839),
.C(n_1824),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1884),
.B(n_1825),
.Y(n_1933)
);

OR2x2_ASAP7_75t_L g1934 ( 
.A(n_1871),
.B(n_1842),
.Y(n_1934)
);

AND2x2_ASAP7_75t_L g1935 ( 
.A(n_1866),
.B(n_1824),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1896),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1896),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1884),
.B(n_1812),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1859),
.B(n_1835),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1860),
.Y(n_1940)
);

NOR2xp33_ASAP7_75t_L g1941 ( 
.A(n_1873),
.B(n_1739),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_L g1942 ( 
.A(n_1868),
.B(n_1835),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1864),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1860),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1864),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1941),
.B(n_1763),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1899),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1899),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1900),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1908),
.B(n_1902),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1907),
.A2(n_1838),
.B(n_1843),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1906),
.B(n_1886),
.Y(n_1952)
);

NOR2x1_ASAP7_75t_L g1953 ( 
.A(n_1932),
.B(n_1890),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_L g1954 ( 
.A(n_1920),
.B(n_1886),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1900),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1921),
.B(n_1886),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1913),
.Y(n_1957)
);

NOR2x1_ASAP7_75t_L g1958 ( 
.A(n_1907),
.B(n_1890),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1906),
.B(n_1882),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1908),
.B(n_1876),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1903),
.B(n_1882),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1912),
.B(n_1882),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1913),
.Y(n_1963)
);

OR2x2_ASAP7_75t_L g1964 ( 
.A(n_1902),
.B(n_1876),
.Y(n_1964)
);

HB1xp67_ASAP7_75t_L g1965 ( 
.A(n_1904),
.Y(n_1965)
);

AOI211x1_ASAP7_75t_SL g1966 ( 
.A1(n_1918),
.A2(n_1870),
.B(n_1864),
.C(n_1869),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1917),
.Y(n_1967)
);

NOR2xp33_ASAP7_75t_L g1968 ( 
.A(n_1931),
.B(n_1763),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1917),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1912),
.B(n_1887),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1919),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1931),
.B(n_1903),
.Y(n_1972)
);

AOI221xp5_ASAP7_75t_L g1973 ( 
.A1(n_1901),
.A2(n_1838),
.B1(n_1874),
.B2(n_1867),
.C(n_1872),
.Y(n_1973)
);

NOR3xp33_ASAP7_75t_L g1974 ( 
.A(n_1923),
.B(n_1890),
.C(n_1863),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1927),
.Y(n_1975)
);

HB1xp67_ASAP7_75t_L g1976 ( 
.A(n_1936),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1927),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1929),
.Y(n_1978)
);

INVx4_ASAP7_75t_L g1979 ( 
.A(n_1919),
.Y(n_1979)
);

OAI21x1_ASAP7_75t_SL g1980 ( 
.A1(n_1926),
.A2(n_1851),
.B(n_1698),
.Y(n_1980)
);

OAI211xp5_ASAP7_75t_SL g1981 ( 
.A1(n_1923),
.A2(n_1926),
.B(n_1939),
.C(n_1930),
.Y(n_1981)
);

AND2x2_ASAP7_75t_L g1982 ( 
.A(n_1914),
.B(n_1887),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1929),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1914),
.B(n_1887),
.Y(n_1984)
);

AOI22xp33_ASAP7_75t_L g1985 ( 
.A1(n_1951),
.A2(n_1937),
.B1(n_1815),
.B2(n_1874),
.Y(n_1985)
);

OAI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1961),
.A2(n_1924),
.B1(n_1928),
.B2(n_1841),
.Y(n_1986)
);

OR2x2_ASAP7_75t_L g1987 ( 
.A(n_1960),
.B(n_1925),
.Y(n_1987)
);

AO221x1_ASAP7_75t_L g1988 ( 
.A1(n_1980),
.A2(n_1863),
.B1(n_1898),
.B2(n_1850),
.C(n_1851),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1947),
.Y(n_1989)
);

OAI22xp33_ASAP7_75t_SL g1990 ( 
.A1(n_1972),
.A2(n_1928),
.B1(n_1934),
.B2(n_1910),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1947),
.Y(n_1991)
);

NOR2xp33_ASAP7_75t_SL g1992 ( 
.A(n_1946),
.B(n_1745),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1955),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_L g1994 ( 
.A1(n_1958),
.A2(n_1841),
.B1(n_1933),
.B2(n_1938),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1965),
.B(n_1938),
.Y(n_1995)
);

OR2x2_ASAP7_75t_L g1996 ( 
.A(n_1960),
.B(n_1910),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1955),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1976),
.B(n_1950),
.Y(n_1998)
);

NOR2xp33_ASAP7_75t_L g1999 ( 
.A(n_1979),
.B(n_1663),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1950),
.B(n_1971),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1957),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1971),
.B(n_1935),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1957),
.Y(n_2003)
);

CKINVDCx14_ASAP7_75t_R g2004 ( 
.A(n_1968),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1963),
.Y(n_2005)
);

OAI322xp33_ASAP7_75t_L g2006 ( 
.A1(n_1964),
.A2(n_1948),
.A3(n_1954),
.B1(n_1956),
.B2(n_1979),
.C1(n_1939),
.C2(n_1930),
.Y(n_2006)
);

INVx2_ASAP7_75t_SL g2007 ( 
.A(n_1979),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1964),
.B(n_1935),
.Y(n_2008)
);

INVx1_ASAP7_75t_SL g2009 ( 
.A(n_1953),
.Y(n_2009)
);

NOR2x1_ASAP7_75t_L g2010 ( 
.A(n_1981),
.B(n_1918),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1973),
.A2(n_1874),
.B1(n_1872),
.B2(n_1867),
.Y(n_2011)
);

OAI22xp5_ASAP7_75t_L g2012 ( 
.A1(n_1959),
.A2(n_1827),
.B1(n_1911),
.B2(n_1934),
.Y(n_2012)
);

CKINVDCx14_ASAP7_75t_R g2013 ( 
.A(n_1970),
.Y(n_2013)
);

INVxp67_ASAP7_75t_L g2014 ( 
.A(n_2007),
.Y(n_2014)
);

OAI221xp5_ASAP7_75t_L g2015 ( 
.A1(n_1985),
.A2(n_1966),
.B1(n_1974),
.B2(n_1975),
.C(n_1978),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1995),
.B(n_1959),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1993),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1997),
.Y(n_2018)
);

AOI322xp5_ASAP7_75t_L g2019 ( 
.A1(n_1985),
.A2(n_1874),
.A3(n_1867),
.B1(n_1872),
.B2(n_1865),
.C1(n_1858),
.C2(n_1855),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_2013),
.B(n_1962),
.Y(n_2020)
);

AND2x2_ASAP7_75t_L g2021 ( 
.A(n_2013),
.B(n_1962),
.Y(n_2021)
);

OAI322xp33_ASAP7_75t_L g2022 ( 
.A1(n_2009),
.A2(n_1977),
.A3(n_1963),
.B1(n_1975),
.B2(n_1978),
.C1(n_1967),
.C2(n_1949),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_L g2023 ( 
.A1(n_2011),
.A2(n_1984),
.B1(n_1970),
.B2(n_1982),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_2000),
.B(n_1952),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_2001),
.Y(n_2025)
);

NOR2xp33_ASAP7_75t_L g2026 ( 
.A(n_1992),
.B(n_1916),
.Y(n_2026)
);

NOR2xp33_ASAP7_75t_L g2027 ( 
.A(n_2004),
.B(n_1916),
.Y(n_2027)
);

AOI221xp5_ASAP7_75t_L g2028 ( 
.A1(n_1990),
.A2(n_1977),
.B1(n_1969),
.B2(n_1983),
.C(n_1905),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_2003),
.Y(n_2029)
);

AOI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1994),
.A2(n_1806),
.B1(n_1984),
.B2(n_1982),
.Y(n_2030)
);

OAI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1998),
.A2(n_1875),
.B1(n_1922),
.B2(n_1905),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1999),
.B(n_1952),
.Y(n_2032)
);

OAI21xp33_ASAP7_75t_SL g2033 ( 
.A1(n_2010),
.A2(n_1942),
.B(n_1909),
.Y(n_2033)
);

AOI222xp33_ASAP7_75t_L g2034 ( 
.A1(n_2011),
.A2(n_1942),
.B1(n_1856),
.B2(n_1855),
.C1(n_1943),
.C2(n_1909),
.Y(n_2034)
);

OR2x2_ASAP7_75t_L g2035 ( 
.A(n_1996),
.B(n_1987),
.Y(n_2035)
);

AOI21xp33_ASAP7_75t_SL g2036 ( 
.A1(n_1999),
.A2(n_1980),
.B(n_1898),
.Y(n_2036)
);

AOI32xp33_ASAP7_75t_L g2037 ( 
.A1(n_2033),
.A2(n_1986),
.A3(n_2012),
.B1(n_2005),
.B2(n_1991),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_2027),
.B(n_2008),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_2035),
.Y(n_2039)
);

OAI21xp5_ASAP7_75t_SL g2040 ( 
.A1(n_2020),
.A2(n_2002),
.B(n_1989),
.Y(n_2040)
);

AOI321xp33_ASAP7_75t_SL g2041 ( 
.A1(n_2027),
.A2(n_2006),
.A3(n_1988),
.B1(n_1911),
.B2(n_1905),
.C(n_1943),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_2021),
.B(n_1858),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2017),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2024),
.B(n_1858),
.Y(n_2044)
);

NAND3xp33_ASAP7_75t_L g2045 ( 
.A(n_2028),
.B(n_1915),
.C(n_1909),
.Y(n_2045)
);

XOR2x2_ASAP7_75t_L g2046 ( 
.A(n_2026),
.B(n_1704),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_2014),
.B(n_1865),
.Y(n_2047)
);

OR2x2_ASAP7_75t_L g2048 ( 
.A(n_2016),
.B(n_1875),
.Y(n_2048)
);

XNOR2xp5_ASAP7_75t_L g2049 ( 
.A(n_2032),
.B(n_1754),
.Y(n_2049)
);

XNOR2x1_ASAP7_75t_L g2050 ( 
.A(n_2030),
.B(n_1808),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_2018),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_2014),
.Y(n_2052)
);

AOI211xp5_ASAP7_75t_SL g2053 ( 
.A1(n_2039),
.A2(n_2022),
.B(n_2015),
.C(n_2031),
.Y(n_2053)
);

NAND5xp2_ASAP7_75t_L g2054 ( 
.A(n_2041),
.B(n_2019),
.C(n_2034),
.D(n_2029),
.E(n_2025),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_2052),
.B(n_2031),
.Y(n_2055)
);

NAND4xp25_ASAP7_75t_L g2056 ( 
.A(n_2037),
.B(n_2023),
.C(n_2036),
.D(n_1911),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_2040),
.B(n_2038),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_2047),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_2042),
.B(n_1915),
.Y(n_2059)
);

NOR4xp25_ASAP7_75t_L g2060 ( 
.A(n_2043),
.B(n_1945),
.C(n_1943),
.D(n_1915),
.Y(n_2060)
);

NAND4xp25_ASAP7_75t_L g2061 ( 
.A(n_2044),
.B(n_1911),
.C(n_1945),
.D(n_1922),
.Y(n_2061)
);

AND2x2_ASAP7_75t_SL g2062 ( 
.A(n_2051),
.B(n_2048),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_2045),
.B(n_1875),
.Y(n_2063)
);

AOI21xp5_ASAP7_75t_L g2064 ( 
.A1(n_2045),
.A2(n_2046),
.B(n_2049),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_2050),
.B(n_1865),
.Y(n_2065)
);

NOR3xp33_ASAP7_75t_L g2066 ( 
.A(n_2052),
.B(n_1945),
.C(n_1922),
.Y(n_2066)
);

NOR3xp33_ASAP7_75t_L g2067 ( 
.A(n_2052),
.B(n_1944),
.C(n_1940),
.Y(n_2067)
);

NAND3xp33_ASAP7_75t_L g2068 ( 
.A(n_2052),
.B(n_1944),
.C(n_1940),
.Y(n_2068)
);

OAI211xp5_ASAP7_75t_L g2069 ( 
.A1(n_2053),
.A2(n_1898),
.B(n_1863),
.C(n_1864),
.Y(n_2069)
);

O2A1O1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_2055),
.A2(n_1870),
.B(n_1863),
.C(n_1898),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_2062),
.Y(n_2071)
);

OAI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2057),
.A2(n_1898),
.B(n_1870),
.C(n_1746),
.Y(n_2072)
);

NAND4xp25_ASAP7_75t_L g2073 ( 
.A(n_2054),
.B(n_1898),
.C(n_1870),
.D(n_1760),
.Y(n_2073)
);

AOI211x1_ASAP7_75t_SL g2074 ( 
.A1(n_2056),
.A2(n_1869),
.B(n_1897),
.C(n_1820),
.Y(n_2074)
);

NAND2x1_ASAP7_75t_SL g2075 ( 
.A(n_2065),
.B(n_1808),
.Y(n_2075)
);

AO22x1_ASAP7_75t_L g2076 ( 
.A1(n_2066),
.A2(n_1696),
.B1(n_1808),
.B2(n_1853),
.Y(n_2076)
);

NAND3xp33_ASAP7_75t_L g2077 ( 
.A(n_2064),
.B(n_1862),
.C(n_1860),
.Y(n_2077)
);

OAI22xp33_ASAP7_75t_L g2078 ( 
.A1(n_2063),
.A2(n_1892),
.B1(n_1883),
.B2(n_1889),
.Y(n_2078)
);

AOI222xp33_ASAP7_75t_L g2079 ( 
.A1(n_2069),
.A2(n_2068),
.B1(n_2059),
.B2(n_2058),
.C1(n_2060),
.C2(n_2067),
.Y(n_2079)
);

CKINVDCx16_ASAP7_75t_R g2080 ( 
.A(n_2071),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_2077),
.A2(n_2068),
.B1(n_1855),
.B2(n_1856),
.Y(n_2081)
);

OAI211xp5_ASAP7_75t_L g2082 ( 
.A1(n_2073),
.A2(n_2061),
.B(n_1820),
.C(n_1812),
.Y(n_2082)
);

OAI222xp33_ASAP7_75t_L g2083 ( 
.A1(n_2070),
.A2(n_1889),
.B1(n_1878),
.B2(n_1892),
.C1(n_1883),
.C2(n_1876),
.Y(n_2083)
);

NAND5xp2_ASAP7_75t_L g2084 ( 
.A(n_2072),
.B(n_1696),
.C(n_1856),
.D(n_1765),
.E(n_1766),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2075),
.Y(n_2085)
);

AOI221xp5_ASAP7_75t_L g2086 ( 
.A1(n_2078),
.A2(n_1878),
.B1(n_1889),
.B2(n_1883),
.C(n_1892),
.Y(n_2086)
);

AOI211xp5_ASAP7_75t_L g2087 ( 
.A1(n_2076),
.A2(n_1850),
.B(n_1696),
.C(n_1833),
.Y(n_2087)
);

NAND3xp33_ASAP7_75t_L g2088 ( 
.A(n_2079),
.B(n_2074),
.C(n_1888),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2080),
.Y(n_2089)
);

NAND4xp75_ASAP7_75t_L g2090 ( 
.A(n_2085),
.B(n_1696),
.C(n_1736),
.D(n_1878),
.Y(n_2090)
);

INVx1_ASAP7_75t_SL g2091 ( 
.A(n_2081),
.Y(n_2091)
);

INVxp33_ASAP7_75t_L g2092 ( 
.A(n_2086),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_2082),
.B(n_1862),
.Y(n_2093)
);

INVx2_ASAP7_75t_SL g2094 ( 
.A(n_2083),
.Y(n_2094)
);

CKINVDCx16_ASAP7_75t_R g2095 ( 
.A(n_2089),
.Y(n_2095)
);

AND2x2_ASAP7_75t_L g2096 ( 
.A(n_2091),
.B(n_2087),
.Y(n_2096)
);

NOR2x1p5_ASAP7_75t_L g2097 ( 
.A(n_2088),
.B(n_2084),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_2096),
.Y(n_2098)
);

AO22x1_ASAP7_75t_L g2099 ( 
.A1(n_2098),
.A2(n_2094),
.B1(n_2092),
.B2(n_2095),
.Y(n_2099)
);

AOI22xp5_ASAP7_75t_L g2100 ( 
.A1(n_2099),
.A2(n_2097),
.B1(n_2093),
.B2(n_2090),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2099),
.Y(n_2101)
);

CKINVDCx20_ASAP7_75t_R g2102 ( 
.A(n_2101),
.Y(n_2102)
);

OAI22xp5_ASAP7_75t_L g2103 ( 
.A1(n_2100),
.A2(n_1883),
.B1(n_1889),
.B2(n_1892),
.Y(n_2103)
);

AOI22xp33_ASAP7_75t_L g2104 ( 
.A1(n_2102),
.A2(n_2103),
.B1(n_1878),
.B2(n_1862),
.Y(n_2104)
);

OAI21xp5_ASAP7_75t_L g2105 ( 
.A1(n_2102),
.A2(n_1885),
.B(n_1868),
.Y(n_2105)
);

OAI222xp33_ASAP7_75t_L g2106 ( 
.A1(n_2104),
.A2(n_1885),
.B1(n_1891),
.B2(n_1888),
.C1(n_1893),
.C2(n_1897),
.Y(n_2106)
);

OAI222xp33_ASAP7_75t_L g2107 ( 
.A1(n_2106),
.A2(n_2105),
.B1(n_1885),
.B2(n_1888),
.C1(n_1891),
.C2(n_1893),
.Y(n_2107)
);

XNOR2xp5_ASAP7_75t_L g2108 ( 
.A(n_2107),
.B(n_1754),
.Y(n_2108)
);

OAI221xp5_ASAP7_75t_L g2109 ( 
.A1(n_2108),
.A2(n_1891),
.B1(n_1893),
.B2(n_1853),
.C(n_1846),
.Y(n_2109)
);

AOI211xp5_ASAP7_75t_L g2110 ( 
.A1(n_2109),
.A2(n_1793),
.B(n_1850),
.C(n_1846),
.Y(n_2110)
);


endmodule