module fake_jpeg_18782_n_99 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_99);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_99;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx11_ASAP7_75t_SL g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_26),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

HAxp5_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_0),
.CON(n_47),
.SN(n_47)
);

OA22x2_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_39),
.B1(n_36),
.B2(n_43),
.Y(n_56)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_50),
.B(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_37),
.B(n_2),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_46),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_56),
.A2(n_58),
.B(n_60),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_42),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_40),
.C(n_44),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_61),
.B(n_63),
.C(n_65),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_41),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_64),
.A2(n_15),
.B1(n_29),
.B2(n_25),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_54),
.A2(n_17),
.B(n_32),
.Y(n_65)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_14),
.B1(n_24),
.B2(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_74),
.Y(n_77)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

AND2x6_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_10),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_13),
.B(n_22),
.C(n_20),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_72),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_75),
.A2(n_76),
.B(n_3),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_57),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_57),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_82),
.A2(n_67),
.B1(n_71),
.B2(n_76),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_86),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_87),
.A2(n_89),
.B1(n_81),
.B2(n_80),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OA21x2_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_85),
.B(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_88),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_94),
.B(n_4),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_95),
.A2(n_5),
.B(n_84),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

OAI321xp33_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_18),
.C(n_19),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_34),
.Y(n_99)
);


endmodule