module fake_jpeg_20082_n_379 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_379);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_379;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx24_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_42),
.B(n_46),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_24),
.B(n_36),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_50),
.B(n_60),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_24),
.B(n_7),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_53),
.Y(n_88)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

NAND2x1_ASAP7_75t_SL g78 ( 
.A(n_54),
.B(n_58),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_59),
.B(n_26),
.Y(n_70)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_63),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_61),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_64),
.B(n_71),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_27),
.CON(n_67),
.SN(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_52),
.B(n_37),
.C(n_39),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_63),
.A2(n_22),
.B1(n_30),
.B2(n_20),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_68),
.A2(n_76),
.B1(n_47),
.B2(n_43),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_84),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_38),
.B(n_27),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_73),
.B(n_77),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_45),
.A2(n_22),
.B1(n_30),
.B2(n_34),
.Y(n_76)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_44),
.A2(n_19),
.B(n_29),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_59),
.B(n_29),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_53),
.A2(n_22),
.B1(n_30),
.B2(n_23),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_87),
.B1(n_60),
.B2(n_89),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_34),
.B1(n_20),
.B2(n_23),
.Y(n_87)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx11_ASAP7_75t_L g131 ( 
.A(n_93),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_48),
.B(n_28),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_95),
.B(n_97),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_43),
.B(n_47),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_62),
.Y(n_119)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_57),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_35),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_49),
.A2(n_34),
.B1(n_20),
.B2(n_28),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_56),
.B1(n_55),
.B2(n_41),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

BUFx4f_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_102),
.A2(n_109),
.B1(n_83),
.B2(n_69),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_105),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_74),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_106),
.A2(n_78),
.B(n_32),
.C(n_17),
.Y(n_149)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_111),
.B(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_83),
.B1(n_69),
.B2(n_66),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_89),
.A2(n_17),
.B1(n_35),
.B2(n_32),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_79),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_115),
.Y(n_157)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_62),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_78),
.B(n_93),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_119),
.B(n_122),
.Y(n_150)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_120),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_71),
.B(n_11),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g162 ( 
.A(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_11),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_67),
.B(n_8),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_130),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_86),
.B(n_8),
.Y(n_130)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_86),
.B(n_35),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_88),
.B(n_35),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_8),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_135),
.B(n_138),
.Y(n_161)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_88),
.B(n_85),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_78),
.C(n_97),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_135),
.C(n_121),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_141),
.Y(n_192)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_133),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_147),
.A2(n_154),
.B1(n_172),
.B2(n_110),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_149),
.A2(n_165),
.B(n_173),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_101),
.Y(n_153)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_120),
.A2(n_98),
.B1(n_80),
.B2(n_72),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_0),
.B(n_1),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_119),
.A2(n_72),
.B1(n_80),
.B2(n_81),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_166),
.A2(n_167),
.B1(n_137),
.B2(n_123),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_72),
.B1(n_81),
.B2(n_32),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_108),
.B(n_12),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_169),
.B(n_108),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_136),
.A2(n_32),
.B1(n_17),
.B2(n_2),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_100),
.B(n_65),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_180),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_136),
.B(n_105),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_175),
.A2(n_179),
.B(n_183),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_182),
.B1(n_199),
.B2(n_157),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g179 ( 
.A(n_152),
.B(n_104),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_171),
.B(n_117),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_181),
.Y(n_211)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_112),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_150),
.B(n_117),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_186),
.B(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_187),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_126),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_103),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_103),
.Y(n_193)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_193),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_143),
.B(n_118),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_196),
.Y(n_213)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_195),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_143),
.B(n_134),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_173),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_203),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_162),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_130),
.B1(n_106),
.B2(n_132),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_139),
.B(n_129),
.C(n_116),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_208),
.C(n_173),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_159),
.B(n_122),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_166),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_146),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

AND2x2_ASAP7_75t_SL g208 ( 
.A(n_159),
.B(n_115),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_145),
.B(n_101),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_146),
.Y(n_210)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

AO21x1_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_149),
.B(n_161),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_234),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_218),
.B(n_196),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_198),
.B(n_190),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_220),
.B(n_240),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_192),
.A2(n_147),
.B1(n_148),
.B2(n_161),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_221),
.A2(n_225),
.B1(n_239),
.B2(n_208),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_204),
.A2(n_209),
.B(n_183),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_224),
.A2(n_226),
.B(n_210),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_192),
.A2(n_148),
.B1(n_158),
.B2(n_107),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_158),
.B(n_162),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_183),
.B(n_162),
.C(n_127),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_233),
.C(n_243),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_241),
.B1(n_197),
.B2(n_203),
.Y(n_248)
);

AO22x1_ASAP7_75t_SL g234 ( 
.A1(n_206),
.A2(n_151),
.B1(n_163),
.B2(n_142),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_131),
.B1(n_163),
.B2(n_151),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_156),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_178),
.A2(n_164),
.B1(n_131),
.B2(n_144),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_164),
.C(n_153),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_211),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_246),
.Y(n_278)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_215),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_179),
.Y(n_247)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_251),
.Y(n_287)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_219),
.Y(n_249)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_249),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_230),
.Y(n_251)
);

OA22x2_ASAP7_75t_L g252 ( 
.A1(n_238),
.A2(n_187),
.B1(n_181),
.B2(n_184),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_252),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_253),
.B(n_218),
.C(n_243),
.Y(n_277)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_255),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_232),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_185),
.Y(n_258)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_258),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_223),
.B(n_205),
.Y(n_259)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_199),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_267),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_217),
.Y(n_263)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_223),
.B(n_208),
.Y(n_265)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_216),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_266),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_234),
.Y(n_268)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_268),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_214),
.B(n_191),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_212),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_237),
.B(n_195),
.Y(n_270)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_270),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_225),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_272),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_242),
.B(n_202),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_224),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_298),
.C(n_261),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_286),
.B(n_297),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_240),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_294),
.C(n_176),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_229),
.C(n_226),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_213),
.C(n_231),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_278),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_299),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_65),
.C(n_6),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_260),
.C(n_267),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_301),
.B(n_309),
.C(n_310),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_274),
.A2(n_256),
.B1(n_271),
.B2(n_262),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_287),
.B1(n_283),
.B2(n_296),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_293),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_303),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_259),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_305),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_275),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_306),
.B(n_313),
.Y(n_330)
);

OA22x2_ASAP7_75t_L g307 ( 
.A1(n_281),
.A2(n_250),
.B1(n_273),
.B2(n_244),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_307),
.A2(n_311),
.B(n_316),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_292),
.A2(n_250),
.B(n_266),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_308),
.A2(n_279),
.B(n_286),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_253),
.C(n_269),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_294),
.B(n_265),
.C(n_252),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_292),
.A2(n_252),
.B(n_227),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_276),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_312),
.B(n_318),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_251),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_252),
.C(n_221),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_315),
.C(n_279),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_207),
.C(n_241),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_283),
.A2(n_234),
.B(n_236),
.Y(n_316)
);

OAI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_281),
.A2(n_236),
.B1(n_177),
.B2(n_176),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_317),
.A2(n_295),
.B1(n_280),
.B2(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_276),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_319),
.B(n_288),
.Y(n_322)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_321),
.B(n_324),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_328),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_297),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g331 ( 
.A(n_308),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_331),
.A2(n_15),
.B(n_14),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_333),
.B(n_335),
.C(n_5),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_314),
.A2(n_285),
.B1(n_177),
.B2(n_131),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_334),
.B(n_315),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_336),
.B(n_341),
.Y(n_355)
);

AOI21xp33_ASAP7_75t_L g337 ( 
.A1(n_325),
.A2(n_310),
.B(n_319),
.Y(n_337)
);

NAND2xp33_ASAP7_75t_L g349 ( 
.A(n_337),
.B(n_327),
.Y(n_349)
);

XNOR2x1_ASAP7_75t_L g338 ( 
.A(n_321),
.B(n_304),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_328),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_323),
.B(n_300),
.C(n_301),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_339),
.B(n_340),
.C(n_342),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_304),
.C(n_307),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_332),
.B(n_307),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_307),
.C(n_6),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_343),
.B(n_335),
.C(n_326),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_330),
.B(n_15),
.Y(n_344)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_344),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_14),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_349),
.A2(n_345),
.B(n_1),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_350),
.B(n_352),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_340),
.B(n_322),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_0),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_327),
.C(n_329),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_354),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_342),
.A2(n_324),
.B1(n_13),
.B2(n_12),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_356),
.B(n_13),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_355),
.A2(n_348),
.B1(n_338),
.B2(n_347),
.Y(n_359)
);

OAI321xp33_ASAP7_75t_L g368 ( 
.A1(n_359),
.A2(n_2),
.A3(n_3),
.B1(n_351),
.B2(n_358),
.C(n_364),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_361),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_362),
.A2(n_357),
.B(n_3),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_358),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_364),
.Y(n_370)
);

FAx1_ASAP7_75t_SL g364 ( 
.A(n_350),
.B(n_0),
.CI(n_2),
.CON(n_364),
.SN(n_364)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_365),
.B(n_3),
.Y(n_369)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_367),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_368),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g372 ( 
.A1(n_369),
.A2(n_360),
.B(n_366),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_372),
.A2(n_370),
.B(n_371),
.Y(n_375)
);

FAx1_ASAP7_75t_SL g376 ( 
.A(n_375),
.B(n_374),
.CI(n_359),
.CON(n_376),
.SN(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_376),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_377),
.B(n_376),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_378),
.A2(n_373),
.B(n_364),
.Y(n_379)
);


endmodule