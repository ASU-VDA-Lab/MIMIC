module fake_jpeg_7393_n_179 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_179);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_179;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_2),
.B(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx12f_ASAP7_75t_SL g32 ( 
.A(n_18),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_32),
.A2(n_0),
.B(n_2),
.Y(n_56)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_13),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_32),
.A2(n_23),
.B1(n_31),
.B2(n_36),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_40),
.A2(n_42),
.B1(n_47),
.B2(n_50),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_34),
.A2(n_23),
.B1(n_21),
.B2(n_26),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_23),
.B1(n_21),
.B2(n_26),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_21),
.B1(n_15),
.B2(n_26),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_53),
.A2(n_20),
.B1(n_19),
.B2(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_28),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_25),
.C(n_20),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_14),
.C(n_44),
.Y(n_60)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_57),
.B(n_58),
.Y(n_94)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_59),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_79)
);

OAI21xp33_ASAP7_75t_L g90 ( 
.A1(n_60),
.A2(n_3),
.B(n_4),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_27),
.Y(n_63)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_23),
.B1(n_28),
.B2(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_28),
.B1(n_15),
.B2(n_25),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_68),
.A2(n_19),
.B1(n_16),
.B2(n_15),
.Y(n_83)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_51),
.B(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_51),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_20),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_19),
.B1(n_16),
.B2(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_46),
.B1(n_52),
.B2(n_39),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_76),
.A2(n_77),
.B1(n_80),
.B2(n_73),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_62),
.A2(n_52),
.B1(n_51),
.B2(n_48),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_64),
.B1(n_66),
.B2(n_52),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_91),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_58),
.B1(n_57),
.B2(n_7),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_84),
.A2(n_95),
.B1(n_6),
.B2(n_7),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_92),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_67),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_88),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_67),
.B(n_49),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_93),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_3),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_72),
.B1(n_73),
.B2(n_70),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_5),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_112),
.B(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_5),
.Y(n_103)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_109),
.B(n_95),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_81),
.A2(n_61),
.B(n_11),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_76),
.Y(n_110)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_92),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_117),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_126),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_87),
.B(n_79),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_112),
.B(n_98),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_128),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_101),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_129),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_119),
.A2(n_99),
.B1(n_100),
.B2(n_111),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

FAx1_ASAP7_75t_SL g134 ( 
.A(n_118),
.B(n_113),
.CI(n_98),
.CON(n_134),
.SN(n_134)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_134),
.B(n_135),
.Y(n_147)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_121),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_136),
.A2(n_120),
.B(n_115),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_138),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_116),
.B(n_78),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_113),
.Y(n_142)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_146),
.A2(n_141),
.B(n_133),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_135),
.A2(n_127),
.B(n_129),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_107),
.C(n_128),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_82),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_125),
.C(n_124),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_153),
.A2(n_145),
.B(n_102),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_144),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_149),
.B(n_140),
.C(n_139),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_114),
.B1(n_131),
.B2(n_134),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_156),
.A2(n_152),
.B1(n_146),
.B2(n_114),
.Y(n_162)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_159),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_87),
.C(n_131),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_147),
.B(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_165),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_10),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_83),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_165),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_61),
.B1(n_11),
.B2(n_12),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_167),
.C(n_166),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_173),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_172),
.A2(n_166),
.B(n_10),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_13),
.C(n_174),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_172),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);


endmodule