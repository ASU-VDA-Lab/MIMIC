module fake_jpeg_28494_n_472 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_50),
.Y(n_128)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_53),
.Y(n_116)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_55),
.B(n_90),
.Y(n_118)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_56),
.Y(n_151)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_59),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_31),
.A2(n_16),
.B(n_2),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_60),
.B(n_29),
.C(n_28),
.Y(n_138)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_66),
.Y(n_131)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_70),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_27),
.Y(n_71)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_18),
.B(n_0),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_84),
.Y(n_100)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_32),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_76),
.Y(n_114)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_19),
.Y(n_78)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_25),
.B(n_2),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_86),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_87),
.Y(n_139)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_88),
.Y(n_149)
);

BUFx4f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_92),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_91),
.B(n_93),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_30),
.B(n_3),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_94),
.B(n_95),
.Y(n_147)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_33),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_97),
.B(n_33),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_70),
.A2(n_42),
.B1(n_48),
.B2(n_35),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_103),
.A2(n_110),
.B1(n_111),
.B2(n_117),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_50),
.A2(n_47),
.B1(n_45),
.B2(n_44),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_42),
.B1(n_48),
.B2(n_35),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_115),
.B(n_121),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_88),
.A2(n_42),
.B1(n_48),
.B2(n_35),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_45),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_74),
.A2(n_44),
.B1(n_37),
.B2(n_30),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_138),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_89),
.A2(n_42),
.B1(n_20),
.B2(n_29),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_135),
.A2(n_144),
.B1(n_146),
.B2(n_34),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_58),
.B(n_37),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_29),
.B1(n_28),
.B2(n_20),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_76),
.A2(n_20),
.B1(n_28),
.B2(n_49),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_39),
.Y(n_148)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_152),
.B(n_33),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_97),
.B1(n_94),
.B2(n_93),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_153),
.A2(n_155),
.B1(n_164),
.B2(n_170),
.Y(n_233)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_154),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_104),
.A2(n_51),
.B1(n_73),
.B2(n_90),
.Y(n_155)
);

BUFx24_ASAP7_75t_L g157 ( 
.A(n_112),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_145),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_158),
.Y(n_235)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_105),
.A2(n_34),
.B1(n_24),
.B2(n_39),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_161),
.A2(n_178),
.B1(n_182),
.B2(n_184),
.Y(n_213)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_162),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_66),
.B1(n_91),
.B2(n_87),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_101),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_165),
.B(n_176),
.Y(n_214)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_166),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_201),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_168),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_116),
.A2(n_59),
.B1(n_85),
.B2(n_81),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_120),
.Y(n_171)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_172),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_75),
.B1(n_71),
.B2(n_63),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_173),
.A2(n_130),
.B1(n_123),
.B2(n_128),
.Y(n_232)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_174),
.Y(n_205)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_175),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_101),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_108),
.Y(n_177)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_177),
.Y(n_243)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_124),
.B(n_49),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_190),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_133),
.Y(n_181)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_133),
.A2(n_46),
.B1(n_24),
.B2(n_21),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_183),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_134),
.A2(n_46),
.B1(n_21),
.B2(n_96),
.Y(n_184)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_186),
.B(n_187),
.Y(n_220)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_125),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_109),
.B(n_53),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_134),
.A2(n_22),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_191),
.A2(n_195),
.B1(n_197),
.B2(n_7),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_151),
.Y(n_192)
);

BUFx8_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_100),
.A2(n_3),
.B(n_5),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_119),
.Y(n_194)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_194),
.B(n_198),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_143),
.A2(n_22),
.B1(n_5),
.B2(n_6),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_143),
.A2(n_22),
.B1(n_7),
.B2(n_8),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_107),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_128),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_199),
.B(n_200),
.Y(n_237)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_113),
.Y(n_200)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_140),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_144),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_141),
.B(n_3),
.C(n_7),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_114),
.C(n_113),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_146),
.B(n_112),
.C(n_135),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_204),
.B(n_169),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_196),
.A2(n_142),
.B1(n_150),
.B2(n_131),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_206),
.A2(n_198),
.B1(n_192),
.B2(n_173),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_208),
.B(n_185),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_142),
.B1(n_131),
.B2(n_150),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_209),
.A2(n_232),
.B1(n_236),
.B2(n_198),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_171),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_217),
.B(n_234),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_163),
.B(n_136),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_221),
.B(n_200),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_163),
.B(n_103),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_225),
.C(n_228),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_180),
.B(n_111),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_117),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_203),
.B(n_149),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_229),
.B(n_166),
.C(n_157),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_196),
.A2(n_139),
.B(n_130),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_192),
.B(n_175),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_158),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_153),
.A2(n_123),
.B1(n_186),
.B2(n_162),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_238),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_283)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_214),
.Y(n_246)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_247),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_248),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_190),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_263),
.Y(n_289)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_250),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_251),
.Y(n_290)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_227),
.Y(n_254)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_254),
.Y(n_313)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_255),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_256),
.A2(n_271),
.B1(n_278),
.B2(n_215),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_257),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_258),
.A2(n_259),
.B(n_261),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_244),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_270),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_223),
.A2(n_183),
.B(n_201),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_177),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_226),
.B(n_189),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_264),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_216),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_265),
.Y(n_314)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_267),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_213),
.A2(n_179),
.B(n_157),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_276),
.B(n_215),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_277),
.Y(n_302)
);

FAx1_ASAP7_75t_SL g270 ( 
.A(n_221),
.B(n_194),
.CI(n_174),
.CON(n_270),
.SN(n_270)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_213),
.A2(n_172),
.B1(n_199),
.B2(n_160),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_228),
.A2(n_210),
.B1(n_233),
.B2(n_218),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_272),
.A2(n_232),
.B1(n_233),
.B2(n_238),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_159),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_154),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_208),
.B(n_168),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_281),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_204),
.A2(n_221),
.B(n_218),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_225),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_237),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_279),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_218),
.B(n_16),
.C(n_10),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_224),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_231),
.B(n_8),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_240),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_282),
.B(n_219),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_283),
.A2(n_281),
.B1(n_280),
.B2(n_268),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_242),
.C(n_207),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_284),
.B(n_315),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_285),
.B(n_297),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_244),
.B(n_207),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_288),
.A2(n_304),
.B(n_262),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_291),
.A2(n_308),
.B(n_257),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_293),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_348)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_296),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_249),
.B(n_263),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_310),
.Y(n_326)
);

OAI21xp33_ASAP7_75t_SL g304 ( 
.A1(n_259),
.A2(n_212),
.B(n_211),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_270),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_271),
.A2(n_212),
.B1(n_224),
.B2(n_230),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_211),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_269),
.C(n_277),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_272),
.A2(n_251),
.B1(n_274),
.B2(n_252),
.Y(n_310)
);

AO22x1_ASAP7_75t_L g312 ( 
.A1(n_270),
.A2(n_222),
.B1(n_230),
.B2(n_245),
.Y(n_312)
);

AO22x1_ASAP7_75t_SL g340 ( 
.A1(n_312),
.A2(n_266),
.B1(n_222),
.B2(n_219),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_246),
.B(n_235),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_320),
.B(n_307),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_289),
.B(n_278),
.CI(n_257),
.CON(n_322),
.SN(n_322)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_343),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_323),
.A2(n_330),
.B(n_336),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_296),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_324),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_275),
.C(n_261),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_325),
.B(n_328),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_327),
.B(n_292),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_253),
.C(n_279),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_301),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_331),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_290),
.A2(n_283),
.B1(n_256),
.B2(n_262),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_337),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_267),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_342),
.Y(n_368)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_300),
.Y(n_334)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_289),
.B(n_254),
.Y(n_335)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_335),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_288),
.A2(n_273),
.B(n_264),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_293),
.A2(n_260),
.B1(n_247),
.B2(n_250),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_338),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_291),
.A2(n_285),
.B1(n_308),
.B2(n_297),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_339),
.B(n_340),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_295),
.A2(n_265),
.B1(n_248),
.B2(n_282),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_341),
.B(n_347),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_310),
.B(n_235),
.C(n_255),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_286),
.A2(n_239),
.B(n_245),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_318),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_344),
.B(n_314),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_318),
.B(n_11),
.Y(n_345)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_346),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_312),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_348),
.A2(n_316),
.B1(n_306),
.B2(n_299),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_305),
.B1(n_311),
.B2(n_298),
.Y(n_350)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_350),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_321),
.A2(n_311),
.B1(n_298),
.B2(n_295),
.Y(n_353)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_354),
.B(n_322),
.C(n_287),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_331),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_375),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_347),
.A2(n_292),
.B1(n_286),
.B2(n_312),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_359),
.A2(n_339),
.B1(n_323),
.B2(n_332),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_363),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_325),
.B(n_294),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_320),
.B(n_303),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_367),
.B(n_326),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_314),
.Y(n_369)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_369),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_333),
.B(n_317),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_327),
.Y(n_378)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_372),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_319),
.A2(n_301),
.B1(n_317),
.B2(n_299),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_374),
.A2(n_345),
.B1(n_324),
.B2(n_329),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_383),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_355),
.A2(n_336),
.B(n_330),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_381),
.B(n_349),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_382),
.B(n_356),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_385),
.A2(n_390),
.B1(n_359),
.B2(n_351),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_365),
.A2(n_337),
.B1(n_329),
.B2(n_343),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_386),
.B(n_391),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_326),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_393),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_367),
.B(n_328),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_388),
.B(n_392),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_361),
.Y(n_389)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_389),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_356),
.A2(n_335),
.B1(n_342),
.B2(n_346),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g391 ( 
.A(n_360),
.B(n_322),
.CI(n_287),
.CON(n_391),
.SN(n_391)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_338),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_340),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_394),
.B(n_397),
.C(n_363),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_352),
.B(n_306),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_396),
.B(n_352),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_366),
.B(n_340),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_355),
.A2(n_370),
.B(n_364),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_398),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_364),
.Y(n_399)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_399),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_401),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_382),
.Y(n_422)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_404),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_406),
.B(n_379),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_366),
.C(n_371),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_412),
.C(n_416),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_408),
.B(n_410),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_395),
.A2(n_362),
.B1(n_373),
.B2(n_358),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_383),
.B(n_370),
.C(n_351),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_391),
.B(n_362),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_413),
.B(n_414),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_391),
.B(n_349),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_373),
.C(n_358),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_387),
.C(n_397),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_419),
.C(n_428),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_416),
.B(n_394),
.C(n_379),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_425),
.Y(n_434)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_400),
.Y(n_423)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_423),
.Y(n_433)
);

OAI221xp5_ASAP7_75t_L g427 ( 
.A1(n_411),
.A2(n_398),
.B1(n_380),
.B2(n_376),
.C(n_386),
.Y(n_427)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_427),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_392),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_412),
.B(n_377),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_430),
.B(n_420),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_415),
.B(n_378),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_431),
.B(n_425),
.C(n_428),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_399),
.Y(n_432)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_432),
.Y(n_453)
);

AOI21x1_ASAP7_75t_L g436 ( 
.A1(n_424),
.A2(n_405),
.B(n_402),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_437),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_439),
.B(n_441),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_406),
.C(n_409),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_440),
.B(n_431),
.C(n_409),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g441 ( 
.A(n_422),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_421),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_442),
.B(n_443),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_405),
.Y(n_443)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_429),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_389),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_438),
.A2(n_429),
.B1(n_419),
.B2(n_418),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_446),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_448),
.B(n_452),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_449),
.B(n_450),
.Y(n_457)
);

HAxp5_ASAP7_75t_SL g450 ( 
.A(n_436),
.B(n_441),
.CON(n_450),
.SN(n_450)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_435),
.B(n_316),
.Y(n_452)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_433),
.B(n_361),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_454),
.B(n_334),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_435),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_458),
.B(n_460),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_445),
.A2(n_440),
.B(n_437),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_461),
.C(n_447),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_453),
.B(n_300),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_457),
.A2(n_455),
.B(n_449),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_463),
.A2(n_464),
.B(n_465),
.Y(n_467)
);

OAI31xp33_ASAP7_75t_SL g464 ( 
.A1(n_455),
.A2(n_450),
.A3(n_451),
.B(n_454),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g466 ( 
.A1(n_462),
.A2(n_456),
.B(n_434),
.Y(n_466)
);

NOR3xp33_ASAP7_75t_L g468 ( 
.A(n_466),
.B(n_467),
.C(n_434),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_468),
.B(n_13),
.Y(n_469)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_16),
.B(n_14),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_15),
.B(n_344),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_15),
.Y(n_472)
);


endmodule