module real_aes_976_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_434;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_733;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_756;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_797;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g596 ( .A(n_0), .B(n_269), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_1), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g146 ( .A(n_2), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_3), .B(n_519), .Y(n_551) );
NAND2xp33_ASAP7_75t_SL g545 ( .A(n_4), .B(n_158), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_5), .B(n_165), .Y(n_261) );
INVx1_ASAP7_75t_L g538 ( .A(n_6), .Y(n_538) );
INVx1_ASAP7_75t_L g174 ( .A(n_7), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g478 ( .A(n_8), .Y(n_478) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_9), .Y(n_191) );
AND2x2_ASAP7_75t_L g549 ( .A(n_10), .B(n_218), .Y(n_549) );
INVx2_ASAP7_75t_L g135 ( .A(n_11), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_12), .Y(n_109) );
INVx1_ASAP7_75t_L g270 ( .A(n_13), .Y(n_270) );
AOI221x1_ASAP7_75t_L g541 ( .A1(n_14), .A2(n_132), .B1(n_518), .B2(n_542), .C(n_544), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_15), .B(n_519), .Y(n_527) );
INVx1_ASAP7_75t_L g113 ( .A(n_16), .Y(n_113) );
INVx1_ASAP7_75t_L g267 ( .A(n_17), .Y(n_267) );
INVx1_ASAP7_75t_SL g232 ( .A(n_18), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_19), .B(n_152), .Y(n_253) );
AOI33xp33_ASAP7_75t_L g203 ( .A1(n_20), .A2(n_51), .A3(n_141), .B1(n_150), .B2(n_204), .B3(n_205), .Y(n_203) );
AOI221xp5_ASAP7_75t_SL g517 ( .A1(n_21), .A2(n_40), .B1(n_518), .B2(n_519), .C(n_520), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_22), .A2(n_518), .B(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_23), .B(n_269), .Y(n_554) );
INVx1_ASAP7_75t_L g808 ( .A(n_24), .Y(n_808) );
INVx1_ASAP7_75t_L g183 ( .A(n_25), .Y(n_183) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_26), .A2(n_92), .B(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g166 ( .A(n_26), .B(n_92), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_27), .B(n_272), .Y(n_531) );
INVxp67_ASAP7_75t_L g540 ( .A(n_28), .Y(n_540) );
AND2x2_ASAP7_75t_L g585 ( .A(n_29), .B(n_217), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_30), .B(n_160), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_31), .A2(n_518), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_32), .B(n_272), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_33), .A2(n_43), .B1(n_798), .B2(n_799), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_33), .Y(n_798) );
INVx1_ASAP7_75t_L g140 ( .A(n_34), .Y(n_140) );
AND2x2_ASAP7_75t_L g158 ( .A(n_34), .B(n_146), .Y(n_158) );
AND2x2_ASAP7_75t_L g164 ( .A(n_34), .B(n_143), .Y(n_164) );
OR2x6_ASAP7_75t_L g111 ( .A(n_35), .B(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g186 ( .A(n_36), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_37), .B(n_160), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_38), .A2(n_133), .B1(n_165), .B2(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_39), .B(n_255), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_41), .A2(n_81), .B1(n_138), .B2(n_518), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_42), .B(n_152), .Y(n_233) );
INVx1_ASAP7_75t_L g799 ( .A(n_43), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_44), .B(n_269), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_45), .A2(n_118), .B1(n_119), .B2(n_122), .Y(n_117) );
INVx1_ASAP7_75t_L g122 ( .A(n_45), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_46), .B(n_171), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_47), .B(n_152), .Y(n_175) );
CKINVDCx5p33_ASAP7_75t_R g250 ( .A(n_48), .Y(n_250) );
AOI222xp33_ASAP7_75t_L g104 ( .A1(n_49), .A2(n_105), .B1(n_475), .B2(n_480), .C1(n_489), .C2(n_493), .Y(n_104) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_49), .A2(n_77), .B1(n_120), .B2(n_121), .Y(n_119) );
INVxp67_ASAP7_75t_L g120 ( .A(n_49), .Y(n_120) );
AND2x2_ASAP7_75t_L g599 ( .A(n_49), .B(n_217), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_50), .B(n_217), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_52), .B(n_152), .Y(n_215) );
INVx1_ASAP7_75t_L g145 ( .A(n_53), .Y(n_145) );
INVx1_ASAP7_75t_L g154 ( .A(n_53), .Y(n_154) );
AND2x2_ASAP7_75t_L g216 ( .A(n_54), .B(n_217), .Y(n_216) );
AOI221xp5_ASAP7_75t_L g172 ( .A1(n_55), .A2(n_73), .B1(n_138), .B2(n_160), .C(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_56), .B(n_160), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g584 ( .A(n_57), .B(n_519), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_58), .B(n_133), .Y(n_193) );
AOI21xp5_ASAP7_75t_SL g137 ( .A1(n_59), .A2(n_138), .B(n_147), .Y(n_137) );
AND2x2_ASAP7_75t_L g564 ( .A(n_60), .B(n_217), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_61), .B(n_272), .Y(n_597) );
INVx1_ASAP7_75t_L g264 ( .A(n_62), .Y(n_264) );
AND2x2_ASAP7_75t_SL g532 ( .A(n_63), .B(n_218), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_64), .B(n_269), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_65), .A2(n_518), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g214 ( .A(n_66), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_67), .B(n_272), .Y(n_555) );
AND2x2_ASAP7_75t_SL g570 ( .A(n_68), .B(n_171), .Y(n_570) );
OAI22xp5_ASAP7_75t_SL g468 ( .A1(n_69), .A2(n_91), .B1(n_469), .B2(n_470), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_69), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_70), .A2(n_138), .B(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g143 ( .A(n_71), .Y(n_143) );
INVx1_ASAP7_75t_L g156 ( .A(n_71), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_72), .B(n_160), .Y(n_206) );
AND2x2_ASAP7_75t_L g234 ( .A(n_74), .B(n_132), .Y(n_234) );
INVx1_ASAP7_75t_L g265 ( .A(n_75), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_76), .A2(n_138), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_78), .A2(n_138), .B(n_198), .C(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_79), .B(n_519), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g568 ( .A1(n_80), .A2(n_84), .B1(n_160), .B2(n_519), .Y(n_568) );
INVx1_ASAP7_75t_L g114 ( .A(n_82), .Y(n_114) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_83), .B(n_132), .Y(n_131) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_85), .A2(n_138), .B1(n_201), .B2(n_202), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_86), .B(n_269), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_87), .B(n_269), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_88), .B(n_473), .Y(n_472) );
XNOR2x2_ASAP7_75t_SL g795 ( .A(n_89), .B(n_796), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_90), .A2(n_518), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g470 ( .A(n_91), .Y(n_470) );
NOR2xp33_ASAP7_75t_SL g498 ( .A(n_91), .B(n_499), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_91), .A2(n_502), .B(n_503), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g504 ( .A1(n_91), .A2(n_499), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g148 ( .A(n_93), .Y(n_148) );
XNOR2xp5_ASAP7_75t_L g796 ( .A(n_94), .B(n_797), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_95), .B(n_272), .Y(n_561) );
AND2x2_ASAP7_75t_L g207 ( .A(n_96), .B(n_132), .Y(n_207) );
A2O1A1Ixp33_ASAP7_75t_L g180 ( .A1(n_97), .A2(n_181), .B(n_182), .C(n_185), .Y(n_180) );
INVxp67_ASAP7_75t_L g543 ( .A(n_98), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_99), .B(n_519), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_100), .B(n_272), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_101), .A2(n_518), .B(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g479 ( .A(n_102), .Y(n_479) );
BUFx2_ASAP7_75t_SL g486 ( .A(n_102), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_103), .B(n_152), .Y(n_151) );
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_115), .B(n_472), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
BUFx2_ASAP7_75t_L g474 ( .A(n_108), .Y(n_474) );
BUFx2_ASAP7_75t_L g488 ( .A(n_108), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x6_ASAP7_75t_SL g509 ( .A(n_109), .B(n_111), .Y(n_509) );
OR2x6_ASAP7_75t_SL g794 ( .A(n_109), .B(n_110), .Y(n_794) );
OR2x2_ASAP7_75t_L g811 ( .A(n_109), .B(n_111), .Y(n_811) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
AOI22xp33_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_117), .B1(n_123), .B2(n_471), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g471 ( .A(n_123), .Y(n_471) );
XOR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_467), .Y(n_123) );
NAND3x1_ASAP7_75t_L g124 ( .A(n_125), .B(n_357), .C(n_422), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_311), .Y(n_125) );
AOI21xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_256), .B(n_284), .Y(n_126) );
AOI21xp33_ASAP7_75t_SL g500 ( .A1(n_127), .A2(n_256), .B(n_284), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_219), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_167), .Y(n_128) );
AOI21xp33_ASAP7_75t_L g358 ( .A1(n_129), .A2(n_359), .B(n_370), .Y(n_358) );
AND2x2_ASAP7_75t_SL g393 ( .A(n_129), .B(n_300), .Y(n_393) );
AND2x2_ASAP7_75t_L g408 ( .A(n_129), .B(n_409), .Y(n_408) );
OR2x6_ASAP7_75t_L g418 ( .A(n_129), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g420 ( .A(n_129), .B(n_410), .Y(n_420) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g294 ( .A(n_130), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_130), .B(n_308), .Y(n_307) );
INVx4_ASAP7_75t_L g326 ( .A(n_130), .Y(n_326) );
AND2x2_ASAP7_75t_L g329 ( .A(n_130), .B(n_245), .Y(n_329) );
NOR2x1_ASAP7_75t_SL g332 ( .A(n_130), .B(n_260), .Y(n_332) );
AND2x4_ASAP7_75t_L g344 ( .A(n_130), .B(n_342), .Y(n_344) );
OR2x2_ASAP7_75t_L g354 ( .A(n_130), .B(n_226), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_130), .B(n_366), .Y(n_371) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_132), .A2(n_180), .B1(n_186), .B2(n_187), .Y(n_179) );
INVx3_ASAP7_75t_L g187 ( .A(n_132), .Y(n_187) );
INVx4_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_133), .B(n_190), .Y(n_189) );
AOI21x1_ASAP7_75t_L g592 ( .A1(n_133), .A2(n_593), .B(n_599), .Y(n_592) );
INVx3_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
BUFx4f_ASAP7_75t_L g171 ( .A(n_134), .Y(n_171) );
AND2x4_ASAP7_75t_L g165 ( .A(n_135), .B(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_SL g218 ( .A(n_135), .B(n_166), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_159), .B(n_165), .Y(n_136) );
INVxp67_ASAP7_75t_L g192 ( .A(n_138), .Y(n_192) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_138), .A2(n_160), .B1(n_537), .B2(n_539), .Y(n_536) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
NOR2x1p5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
INVx1_ASAP7_75t_L g205 ( .A(n_141), .Y(n_205) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
OR2x6_ASAP7_75t_L g149 ( .A(n_142), .B(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g269 ( .A(n_143), .B(n_153), .Y(n_269) );
AND2x6_ASAP7_75t_L g518 ( .A(n_144), .B(n_164), .Y(n_518) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
INVx2_ASAP7_75t_L g150 ( .A(n_145), .Y(n_150) );
AND2x4_ASAP7_75t_L g272 ( .A(n_145), .B(n_155), .Y(n_272) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_146), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_149), .B(n_151), .C(n_157), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_SL g173 ( .A1(n_149), .A2(n_157), .B(n_174), .C(n_175), .Y(n_173) );
INVxp67_ASAP7_75t_L g181 ( .A(n_149), .Y(n_181) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_149), .A2(n_157), .B(n_214), .C(n_215), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_SL g231 ( .A1(n_149), .A2(n_157), .B(n_232), .C(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g255 ( .A(n_149), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g263 ( .A1(n_149), .A2(n_184), .B1(n_264), .B2(n_265), .Y(n_263) );
AND2x2_ASAP7_75t_L g161 ( .A(n_150), .B(n_162), .Y(n_161) );
INVxp33_ASAP7_75t_L g204 ( .A(n_150), .Y(n_204) );
INVx1_ASAP7_75t_L g184 ( .A(n_152), .Y(n_184) );
AND2x4_ASAP7_75t_L g519 ( .A(n_152), .B(n_158), .Y(n_519) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_155), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g201 ( .A(n_157), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_157), .A2(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_157), .B(n_165), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_157), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_157), .A2(n_530), .B(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_157), .A2(n_554), .B(n_555), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_157), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_157), .A2(n_582), .B(n_583), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_157), .A2(n_596), .B(n_597), .Y(n_595) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_158), .Y(n_185) );
INVx1_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
INVx1_ASAP7_75t_L g248 ( .A(n_161), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_163), .Y(n_249) );
BUFx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_165), .B(n_538), .Y(n_537) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_165), .B(n_540), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_165), .B(n_543), .Y(n_542) );
NOR3xp33_ASAP7_75t_L g544 ( .A(n_165), .B(n_184), .C(n_545), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_165), .A2(n_551), .B(n_552), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_167), .A2(n_300), .B1(n_395), .B2(n_396), .Y(n_394) );
INVx1_ASAP7_75t_SL g438 ( .A(n_167), .Y(n_438) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_195), .Y(n_167) );
INVx2_ASAP7_75t_L g369 ( .A(n_168), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_168), .B(n_315), .Y(n_441) );
AND2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_177), .Y(n_168) );
BUFx3_ASAP7_75t_L g287 ( .A(n_169), .Y(n_287) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g280 ( .A(n_170), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_170), .B(n_197), .Y(n_302) );
AND2x4_ASAP7_75t_L g319 ( .A(n_170), .B(n_320), .Y(n_319) );
INVxp67_ASAP7_75t_L g335 ( .A(n_170), .Y(n_335) );
INVx2_ASAP7_75t_L g392 ( .A(n_170), .Y(n_392) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_176), .Y(n_170) );
INVx2_ASAP7_75t_SL g198 ( .A(n_171), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_171), .A2(n_527), .B(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_L g310 ( .A(n_177), .B(n_276), .Y(n_310) );
NOR2xp67_ASAP7_75t_L g356 ( .A(n_177), .B(n_279), .Y(n_356) );
AND2x2_ASAP7_75t_L g375 ( .A(n_177), .B(n_279), .Y(n_375) );
INVx2_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g237 ( .A(n_178), .Y(n_237) );
INVx1_ASAP7_75t_L g318 ( .A(n_178), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_178), .B(n_209), .Y(n_337) );
AND2x4_ASAP7_75t_L g391 ( .A(n_178), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g178 ( .A(n_179), .B(n_188), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_183), .B(n_184), .Y(n_182) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_187), .A2(n_210), .B(n_216), .Y(n_209) );
AO21x2_ASAP7_75t_L g279 ( .A1(n_187), .A2(n_210), .B(n_216), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_192), .B1(n_193), .B2(n_194), .Y(n_188) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g350 ( .A(n_195), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_195), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_208), .Y(n_195) );
AND2x2_ASAP7_75t_L g334 ( .A(n_196), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g374 ( .A(n_196), .Y(n_374) );
AND2x2_ASAP7_75t_L g379 ( .A(n_196), .B(n_279), .Y(n_379) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_197), .B(n_209), .Y(n_239) );
AO21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_207), .Y(n_197) );
AO21x2_ASAP7_75t_L g276 ( .A1(n_198), .A2(n_199), .B(n_207), .Y(n_276) );
AOI21x1_ASAP7_75t_L g566 ( .A1(n_198), .A2(n_567), .B(n_570), .Y(n_566) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_200), .B(n_206), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx3_ASAP7_75t_L g315 ( .A(n_208), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g433 ( .A(n_208), .B(n_287), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_208), .B(n_237), .Y(n_454) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_209), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_217), .Y(n_227) );
OA21x2_ASAP7_75t_L g516 ( .A1(n_217), .A2(n_517), .B(n_523), .Y(n_516) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OAI21xp33_ASAP7_75t_SL g219 ( .A1(n_220), .A2(n_235), .B(n_240), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_222), .B(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g292 ( .A(n_223), .Y(n_292) );
AND2x2_ASAP7_75t_L g306 ( .A(n_223), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g340 ( .A(n_223), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g406 ( .A(n_223), .B(n_324), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g452 ( .A(n_223), .B(n_453), .C(n_454), .Y(n_452) );
INVx3_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
HB1xp67_ASAP7_75t_L g283 ( .A(n_224), .Y(n_283) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g299 ( .A(n_226), .Y(n_299) );
AND2x2_ASAP7_75t_L g305 ( .A(n_226), .B(n_260), .Y(n_305) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_226), .Y(n_316) );
AND2x2_ASAP7_75t_L g361 ( .A(n_226), .B(n_259), .Y(n_361) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_226), .Y(n_384) );
INVx1_ASAP7_75t_L g401 ( .A(n_226), .Y(n_401) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_234), .Y(n_226) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_227), .A2(n_558), .B(n_564), .Y(n_557) );
AO21x2_ASAP7_75t_L g578 ( .A1(n_227), .A2(n_579), .B(n_585), .Y(n_578) );
AO21x2_ASAP7_75t_L g642 ( .A1(n_227), .A2(n_579), .B(n_585), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g443 ( .A(n_235), .Y(n_443) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_236), .B(n_314), .Y(n_415) );
INVx1_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g277 ( .A(n_237), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AOI211x1_ASAP7_75t_L g311 ( .A1(n_241), .A2(n_312), .B(n_321), .C(n_338), .Y(n_311) );
INVx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_SL g304 ( .A(n_242), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g364 ( .A(n_242), .B(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g300 ( .A(n_244), .B(n_259), .Y(n_300) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x4_ASAP7_75t_L g258 ( .A(n_245), .B(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_245), .Y(n_325) );
INVx1_ASAP7_75t_L g342 ( .A(n_245), .Y(n_342) );
AND2x2_ASAP7_75t_L g410 ( .A(n_245), .B(n_260), .Y(n_410) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_251), .Y(n_245) );
NOR3xp33_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .C(n_250), .Y(n_247) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_274), .B(n_281), .Y(n_256) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_257), .B(n_326), .Y(n_429) );
INVx2_ASAP7_75t_L g461 ( .A(n_257), .Y(n_461) );
INVx4_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g293 ( .A(n_258), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g366 ( .A(n_259), .Y(n_366) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
AND2x4_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_266), .B(n_273), .Y(n_262) );
OAI22xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B1(n_270), .B2(n_271), .Y(n_266) );
INVxp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
OR2x2_ASAP7_75t_L g368 ( .A(n_275), .B(n_369), .Y(n_368) );
NAND2x1_ASAP7_75t_SL g390 ( .A(n_275), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x4_ASAP7_75t_L g290 ( .A(n_276), .B(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g320 ( .A(n_276), .Y(n_320) );
INVx1_ASAP7_75t_L g444 ( .A(n_277), .Y(n_444) );
AND2x2_ASAP7_75t_L g309 ( .A(n_278), .B(n_310), .Y(n_309) );
NOR2x1_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
INVxp33_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g348 ( .A(n_283), .B(n_341), .Y(n_348) );
OAI211xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_288), .B(n_295), .C(n_303), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g372 ( .A(n_286), .B(n_373), .Y(n_372) );
NOR2xp67_ASAP7_75t_SL g377 ( .A(n_286), .B(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_287), .B(n_374), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_289), .B(n_293), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_292), .Y(n_289) );
AND2x2_ASAP7_75t_L g421 ( .A(n_290), .B(n_391), .Y(n_421) );
AOI222xp33_ASAP7_75t_L g439 ( .A1(n_293), .A2(n_440), .B1(n_442), .B2(n_445), .C1(n_446), .C2(n_449), .Y(n_439) );
INVx1_ASAP7_75t_L g403 ( .A(n_294), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_301), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
AND2x4_ASAP7_75t_SL g365 ( .A(n_299), .B(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g419 ( .A(n_300), .Y(n_419) );
AND2x2_ASAP7_75t_L g464 ( .A(n_300), .B(n_316), .Y(n_464) );
AND2x2_ASAP7_75t_L g345 ( .A(n_301), .B(n_346), .Y(n_345) );
INVx2_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g458 ( .A(n_302), .B(n_337), .Y(n_458) );
OAI21xp33_ASAP7_75t_SL g303 ( .A1(n_304), .A2(n_306), .B(n_309), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_304), .A2(n_324), .B(n_365), .Y(n_425) );
AND2x2_ASAP7_75t_L g449 ( .A(n_305), .B(n_326), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g459 ( .A(n_305), .B(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g397 ( .A(n_308), .Y(n_397) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_308), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g432 ( .A(n_310), .Y(n_432) );
INVx1_ASAP7_75t_L g499 ( .A(n_311), .Y(n_499) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_317), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AND2x2_ASAP7_75t_L g435 ( .A(n_315), .B(n_319), .Y(n_435) );
BUFx2_ASAP7_75t_L g323 ( .A(n_316), .Y(n_323) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g346 ( .A(n_318), .Y(n_346) );
INVx2_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
AND2x2_ASAP7_75t_L g388 ( .A(n_318), .B(n_379), .Y(n_388) );
AND2x4_ASAP7_75t_L g355 ( .A(n_319), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g395 ( .A(n_319), .B(n_352), .Y(n_395) );
AND2x2_ASAP7_75t_L g446 ( .A(n_319), .B(n_447), .Y(n_446) );
AOI31xp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_327), .A3(n_331), .B(n_333), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AND2x2_ASAP7_75t_L g343 ( .A(n_323), .B(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_SL g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x4_ASAP7_75t_L g341 ( .A(n_326), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g411 ( .A1(n_329), .A2(n_381), .B1(n_412), .B2(n_415), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_329), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g466 ( .A(n_329), .B(n_382), .Y(n_466) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g381 ( .A(n_332), .B(n_382), .Y(n_381) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
AND2x2_ASAP7_75t_L g404 ( .A(n_334), .B(n_375), .Y(n_404) );
INVx1_ASAP7_75t_L g414 ( .A(n_336), .Y(n_414) );
INVx2_ASAP7_75t_SL g336 ( .A(n_337), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_347), .Y(n_338) );
OAI21xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_343), .B(n_345), .Y(n_339) );
INVx1_ASAP7_75t_L g437 ( .A(n_340), .Y(n_437) );
AND2x2_ASAP7_75t_L g445 ( .A(n_341), .B(n_397), .Y(n_445) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_341), .Y(n_451) );
AND2x2_ASAP7_75t_L g396 ( .A(n_344), .B(n_397), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_349), .B1(n_353), .B2(n_355), .Y(n_347) );
NOR2xp33_ASAP7_75t_SL g349 ( .A(n_350), .B(n_351), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g462 ( .A1(n_350), .A2(n_369), .B1(n_463), .B2(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_SL g353 ( .A(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g362 ( .A(n_355), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g497 ( .A(n_357), .B(n_422), .C(n_498), .D(n_500), .Y(n_497) );
INVxp67_ASAP7_75t_L g502 ( .A(n_357), .Y(n_502) );
AND2x2_ASAP7_75t_L g357 ( .A(n_358), .B(n_385), .Y(n_357) );
OAI21xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B(n_363), .Y(n_359) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
OAI21xp33_ASAP7_75t_L g363 ( .A1(n_361), .A2(n_364), .B(n_367), .Y(n_363) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_364), .A2(n_388), .B1(n_389), .B2(n_393), .Y(n_387) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_372), .B1(n_376), .B2(n_380), .Y(n_370) );
INVx1_ASAP7_75t_L g405 ( .A(n_373), .Y(n_405) );
NAND2x1p5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NOR2xp67_ASAP7_75t_L g385 ( .A(n_386), .B(n_398), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_394), .Y(n_386) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NAND2xp33_ASAP7_75t_SL g440 ( .A(n_390), .B(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g413 ( .A(n_391), .Y(n_413) );
INVx3_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
INVxp67_ASAP7_75t_L g456 ( .A(n_396), .Y(n_456) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_399), .B(n_407), .C(n_411), .D(n_416), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_404), .B1(n_405), .B2(n_406), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
AND2x2_ASAP7_75t_L g409 ( .A(n_401), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g457 ( .A(n_405), .Y(n_457) );
NAND2xp33_ASAP7_75t_SL g412 ( .A(n_413), .B(n_414), .Y(n_412) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_420), .B(n_421), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g505 ( .A(n_422), .Y(n_505) );
AND3x2_ASAP7_75t_L g422 ( .A(n_423), .B(n_439), .C(n_450), .Y(n_422) );
AOI221x1_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_426), .B1(n_428), .B2(n_430), .C(n_436), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND2xp33_ASAP7_75t_SL g430 ( .A(n_431), .B(n_434), .Y(n_430) );
OR2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NAND2xp33_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI211xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_455), .C(n_462), .Y(n_450) );
OAI22xp5_ASAP7_75t_L g455 ( .A1(n_456), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_455) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g489 ( .A(n_474), .B(n_490), .Y(n_489) );
CKINVDCx9p33_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
OR2x2_ASAP7_75t_SL g476 ( .A(n_477), .B(n_479), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_477), .A2(n_484), .B(n_487), .Y(n_483) );
INVx2_ASAP7_75t_L g492 ( .A(n_477), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_479), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
CKINVDCx11_ASAP7_75t_R g484 ( .A(n_485), .Y(n_484) );
CKINVDCx8_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI21xp5_ASAP7_75t_SL g493 ( .A1(n_494), .A2(n_795), .B(n_800), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g495 ( .A1(n_496), .A2(n_506), .B1(n_510), .B2(n_792), .Y(n_495) );
INVx1_ASAP7_75t_L g802 ( .A(n_496), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g496 ( .A(n_497), .B(n_501), .C(n_504), .Y(n_496) );
INVx1_ASAP7_75t_L g503 ( .A(n_500), .Y(n_503) );
OAI21x1_ASAP7_75t_L g801 ( .A1(n_506), .A2(n_802), .B(n_803), .Y(n_801) );
CKINVDCx6p67_ASAP7_75t_R g506 ( .A(n_507), .Y(n_506) );
INVx3_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_509), .Y(n_508) );
NAND2x1_ASAP7_75t_SL g803 ( .A(n_510), .B(n_804), .Y(n_803) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_705), .Y(n_511) );
NAND3xp33_ASAP7_75t_SL g512 ( .A(n_513), .B(n_615), .C(n_655), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_533), .B(n_546), .C(n_571), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_514), .B(n_620), .Y(n_654) );
NOR2x1p5_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
BUFx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g590 ( .A(n_516), .Y(n_590) );
INVx2_ASAP7_75t_L g606 ( .A(n_516), .Y(n_606) );
OR2x2_ASAP7_75t_L g618 ( .A(n_516), .B(n_525), .Y(n_618) );
AND2x2_ASAP7_75t_L g632 ( .A(n_516), .B(n_591), .Y(n_632) );
INVx1_ASAP7_75t_L g660 ( .A(n_516), .Y(n_660) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_516), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_516), .B(n_525), .Y(n_766) );
OR2x2_ASAP7_75t_L g587 ( .A(n_524), .B(n_588), .Y(n_587) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_524), .Y(n_722) );
AND2x2_ASAP7_75t_L g727 ( .A(n_524), .B(n_589), .Y(n_727) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x4_ASAP7_75t_L g533 ( .A(n_525), .B(n_534), .Y(n_533) );
OR2x2_ASAP7_75t_L g586 ( .A(n_525), .B(n_535), .Y(n_586) );
OR2x2_ASAP7_75t_L g605 ( .A(n_525), .B(n_606), .Y(n_605) );
INVx2_ASAP7_75t_L g634 ( .A(n_525), .Y(n_634) );
AND2x4_ASAP7_75t_SL g673 ( .A(n_525), .B(n_535), .Y(n_673) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_525), .Y(n_677) );
OR2x2_ASAP7_75t_L g694 ( .A(n_525), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g704 ( .A(n_525), .B(n_611), .Y(n_704) );
INVx1_ASAP7_75t_L g733 ( .A(n_525), .Y(n_733) );
OR2x6_ASAP7_75t_L g525 ( .A(n_526), .B(n_532), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_533), .B(n_662), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_534), .B(n_591), .Y(n_608) );
AND2x2_ASAP7_75t_L g620 ( .A(n_534), .B(n_621), .Y(n_620) );
OR2x2_ASAP7_75t_L g638 ( .A(n_534), .B(n_605), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_534), .B(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g611 ( .A(n_535), .B(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g633 ( .A(n_535), .B(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g668 ( .A(n_535), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_535), .B(n_591), .Y(n_692) );
AND2x4_ASAP7_75t_L g535 ( .A(n_536), .B(n_541), .Y(n_535) );
AND2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_556), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_547), .B(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g641 ( .A(n_547), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_547), .B(n_557), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_547), .B(n_662), .C(n_663), .Y(n_661) );
AND2x2_ASAP7_75t_L g709 ( .A(n_547), .B(n_614), .Y(n_709) );
INVx5_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x2_ASAP7_75t_L g576 ( .A(n_548), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_SL g613 ( .A(n_548), .B(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g629 ( .A(n_548), .Y(n_629) );
OR2x2_ASAP7_75t_L g652 ( .A(n_548), .B(n_642), .Y(n_652) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_548), .Y(n_669) );
AND2x2_ASAP7_75t_SL g687 ( .A(n_548), .B(n_575), .Y(n_687) );
AND2x4_ASAP7_75t_L g702 ( .A(n_548), .B(n_578), .Y(n_702) );
AND2x2_ASAP7_75t_L g716 ( .A(n_548), .B(n_557), .Y(n_716) );
OR2x2_ASAP7_75t_L g737 ( .A(n_548), .B(n_565), .Y(n_737) );
OR2x6_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
AND2x2_ASAP7_75t_L g791 ( .A(n_556), .B(n_669), .Y(n_791) );
AND2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_565), .Y(n_556) );
AND2x4_ASAP7_75t_L g614 ( .A(n_557), .B(n_577), .Y(n_614) );
INVx2_ASAP7_75t_L g625 ( .A(n_557), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_557), .B(n_575), .Y(n_630) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_557), .Y(n_663) );
OR2x2_ASAP7_75t_L g686 ( .A(n_557), .B(n_578), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_557), .B(n_578), .Y(n_689) );
INVx1_ASAP7_75t_L g698 ( .A(n_557), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
AND2x2_ASAP7_75t_L g601 ( .A(n_565), .B(n_578), .Y(n_601) );
BUFx2_ASAP7_75t_L g650 ( .A(n_565), .Y(n_650) );
AND2x2_ASAP7_75t_L g745 ( .A(n_565), .B(n_625), .Y(n_745) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_566), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_586), .B1(n_587), .B2(n_600), .C(n_602), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_576), .Y(n_573) );
NOR2x1_ASAP7_75t_L g647 ( .A(n_574), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_574), .B(n_641), .Y(n_681) );
OR2x2_ASAP7_75t_L g693 ( .A(n_574), .B(n_689), .Y(n_693) );
OR2x2_ASAP7_75t_L g696 ( .A(n_574), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g785 ( .A(n_574), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g624 ( .A(n_575), .B(n_625), .Y(n_624) );
OA33x2_ASAP7_75t_L g657 ( .A1(n_575), .A2(n_618), .A3(n_658), .B1(n_661), .B2(n_664), .B3(n_667), .Y(n_657) );
OR2x2_ASAP7_75t_L g688 ( .A(n_575), .B(n_689), .Y(n_688) );
OR2x2_ASAP7_75t_L g712 ( .A(n_575), .B(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g720 ( .A(n_575), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g740 ( .A(n_575), .B(n_614), .Y(n_740) );
NOR2xp33_ASAP7_75t_L g778 ( .A(n_575), .B(n_629), .Y(n_778) );
INVx2_ASAP7_75t_L g648 ( .A(n_576), .Y(n_648) );
AOI322xp5_ASAP7_75t_L g718 ( .A1(n_576), .A2(n_631), .A3(n_719), .B1(n_722), .B2(n_723), .C1(n_725), .C2(n_727), .Y(n_718) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_578), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_584), .Y(n_579) );
OR2x2_ASAP7_75t_L g700 ( .A(n_586), .B(n_679), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g752 ( .A(n_586), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g773 ( .A(n_586), .Y(n_773) );
INVx1_ASAP7_75t_SL g639 ( .A(n_587), .Y(n_639) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g672 ( .A(n_589), .B(n_673), .Y(n_672) );
AND2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx2_ASAP7_75t_L g612 ( .A(n_591), .Y(n_612) );
INVx1_ASAP7_75t_L g621 ( .A(n_591), .Y(n_621) );
INVx1_ASAP7_75t_L g662 ( .A(n_591), .Y(n_662) );
OR2x2_ASAP7_75t_L g679 ( .A(n_591), .B(n_606), .Y(n_679) );
HB1xp67_ASAP7_75t_L g754 ( .A(n_591), .Y(n_754) );
INVx3_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_598), .Y(n_593) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_SL g723 ( .A(n_601), .B(n_724), .Y(n_723) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_603), .A2(n_609), .B(n_613), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_L g676 ( .A1(n_603), .A2(n_677), .B(n_678), .C(n_680), .Y(n_676) );
AND2x4_ASAP7_75t_L g603 ( .A(n_604), .B(n_607), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g741 ( .A(n_605), .B(n_742), .Y(n_741) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_606), .Y(n_610) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
OR2x2_ASAP7_75t_L g765 ( .A(n_608), .B(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
AND2x2_ASAP7_75t_SL g734 ( .A(n_611), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g742 ( .A(n_611), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_611), .B(n_733), .Y(n_750) );
INVx3_ASAP7_75t_SL g675 ( .A(n_614), .Y(n_675) );
AOI221xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_622), .B1(n_626), .B2(n_631), .C(n_635), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_621), .Y(n_666) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_624), .A2(n_651), .B(n_723), .Y(n_729) );
AND2x2_ASAP7_75t_L g755 ( .A(n_624), .B(n_702), .Y(n_755) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_625), .Y(n_643) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_629), .B(n_745), .Y(n_744) );
OR2x2_ASAP7_75t_L g764 ( .A(n_629), .B(n_686), .Y(n_764) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
INVx2_ASAP7_75t_L g713 ( .A(n_632), .Y(n_713) );
OAI21xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_640), .B(n_644), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
INVx1_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx2_ASAP7_75t_L g786 ( .A(n_641), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_642), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g715 ( .A(n_642), .B(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_643), .B(n_665), .Y(n_664) );
OAI31xp33_ASAP7_75t_SL g644 ( .A1(n_645), .A2(n_647), .A3(n_649), .B(n_653), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_648), .B(n_675), .Y(n_674) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
OR2x2_ASAP7_75t_L g726 ( .A(n_650), .B(n_652), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_650), .B(n_702), .Y(n_781) );
INVx1_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR5xp2_ASAP7_75t_L g655 ( .A(n_656), .B(n_670), .C(n_682), .D(n_691), .E(n_699), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_660), .B(n_662), .Y(n_695) );
INVx1_ASAP7_75t_L g735 ( .A(n_660), .Y(n_735) );
INVxp67_ASAP7_75t_SL g772 ( .A(n_660), .Y(n_772) );
INVx1_ASAP7_75t_L g724 ( .A(n_663), .Y(n_724) );
INVxp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND2xp33_ASAP7_75t_SL g667 ( .A(n_668), .B(n_669), .Y(n_667) );
OAI321xp33_ASAP7_75t_L g707 ( .A1(n_668), .A2(n_708), .A3(n_710), .B1(n_714), .B2(n_717), .C(n_718), .Y(n_707) );
INVx1_ASAP7_75t_L g761 ( .A(n_669), .Y(n_761) );
OAI21xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_674), .B(n_676), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_672), .A2(n_745), .B1(n_752), .B2(n_755), .Y(n_751) );
AND2x2_ASAP7_75t_L g780 ( .A(n_673), .B(n_754), .Y(n_780) );
INVx1_ASAP7_75t_L g690 ( .A(n_678), .Y(n_690) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_688), .B(n_690), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_689), .A2(n_700), .B1(n_701), .B2(n_703), .Y(n_699) );
INVx1_ASAP7_75t_L g762 ( .A(n_689), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_694), .B2(n_696), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_698), .B(n_702), .Y(n_701) );
OAI221xp5_ASAP7_75t_L g776 ( .A1(n_700), .A2(n_777), .B1(n_779), .B2(n_781), .C(n_782), .Y(n_776) );
INVx1_ASAP7_75t_L g783 ( .A(n_700), .Y(n_783) );
OAI221xp5_ASAP7_75t_L g757 ( .A1(n_701), .A2(n_758), .B1(n_765), .B2(n_767), .C(n_768), .Y(n_757) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_703), .A2(n_729), .B(n_730), .Y(n_728) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_756), .Y(n_705) );
NOR3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_728), .C(n_746), .Y(n_706) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
HB1xp67_ASAP7_75t_L g775 ( .A(n_709), .Y(n_775) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx3_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g774 ( .A(n_717), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_719), .B(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g767 ( .A(n_727), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_736), .B(n_738), .Y(n_730) );
INVxp67_ASAP7_75t_L g788 ( .A(n_731), .Y(n_788) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_SL g743 ( .A(n_734), .Y(n_743) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
OAI22xp33_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_738) );
INVx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
OAI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_748), .B(n_751), .Y(n_746) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g789 ( .A(n_752), .Y(n_789) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
NOR3xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_776), .C(n_787), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_763), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
OAI21xp5_ASAP7_75t_SL g768 ( .A1(n_769), .A2(n_774), .B(n_775), .Y(n_768) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVxp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g782 ( .A1(n_780), .A2(n_783), .B(n_784), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
AOI21xp33_ASAP7_75t_L g787 ( .A1(n_788), .A2(n_789), .B(n_790), .Y(n_787) );
INVx1_ASAP7_75t_SL g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g806 ( .A(n_793), .Y(n_806) );
CKINVDCx11_ASAP7_75t_R g793 ( .A(n_794), .Y(n_793) );
AOI21xp33_ASAP7_75t_SL g800 ( .A1(n_795), .A2(n_801), .B(n_807), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_805), .Y(n_804) );
BUFx4f_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
NOR2xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_809), .Y(n_807) );
INVx1_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
INVx2_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
endmodule