module real_jpeg_19559_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_333, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_333;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_103),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_0),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_0),
.A2(n_51),
.B1(n_52),
.B2(n_103),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_103),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_0),
.A2(n_28),
.B1(n_32),
.B2(n_103),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_1),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_1),
.B(n_22),
.Y(n_137)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_16),
.B(n_51),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_106),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_1),
.A2(n_85),
.B1(n_86),
.B2(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_62),
.Y(n_178)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_1),
.A2(n_25),
.B(n_196),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_2),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_97),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_97),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_2),
.A2(n_28),
.B1(n_32),
.B2(n_97),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_28),
.B1(n_32),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_3),
.A2(n_47),
.B1(n_48),
.B2(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_67),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_3),
.A2(n_24),
.B1(n_25),
.B2(n_67),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_4),
.A2(n_28),
.B1(n_32),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_4),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_108),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_47),
.B1(n_48),
.B2(n_108),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_4),
.A2(n_51),
.B1(n_52),
.B2(n_108),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_5),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_5),
.A2(n_28),
.B1(n_32),
.B2(n_101),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_51),
.B1(n_52),
.B2(n_101),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_101),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_28),
.B1(n_32),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_6),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_6),
.A2(n_51),
.B1(n_52),
.B2(n_70),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_70),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_70),
.Y(n_281)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_8),
.A2(n_28),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_24),
.B1(n_25),
.B2(n_36),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_8),
.A2(n_36),
.B1(n_51),
.B2(n_52),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_8),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_268)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_9),
.Y(n_86)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_10),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_31),
.B1(n_47),
.B2(n_48),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_10),
.A2(n_31),
.B1(n_51),
.B2(n_52),
.Y(n_233)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_13),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_13),
.A2(n_51),
.B1(n_52),
.B2(n_91),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_91),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_13),
.A2(n_28),
.B1(n_32),
.B2(n_91),
.Y(n_289)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_58),
.Y(n_60)
);

OAI32xp33_ASAP7_75t_L g190 ( 
.A1(n_14),
.A2(n_25),
.A3(n_48),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_16),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_16),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_37),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_30),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B(n_28),
.C(n_29),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_22),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_22),
.A2(n_27),
.B1(n_35),
.B2(n_74),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_22),
.A2(n_27),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_22),
.A2(n_27),
.B1(n_288),
.B2(n_289),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_28),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_23),
.B(n_25),
.Y(n_120)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_24),
.A2(n_58),
.B(n_59),
.C(n_60),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_58),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_24),
.A2(n_29),
.B1(n_105),
.B2(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_24),
.B(n_106),
.Y(n_192)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_28),
.B(n_106),
.CON(n_105),
.SN(n_105)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_34),
.B(n_41),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_75),
.B(n_331),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_71),
.C(n_73),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_42),
.A2(n_43),
.B1(n_327),
.B2(n_329),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_54),
.C(n_63),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_44),
.A2(n_298),
.B1(n_299),
.B2(n_301),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_44),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_44),
.A2(n_54),
.B1(n_301),
.B2(n_314),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_50),
.B(n_53),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_45),
.A2(n_50),
.B1(n_90),
.B2(n_92),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_45),
.A2(n_50),
.B1(n_90),
.B2(n_96),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_45),
.A2(n_50),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_45),
.A2(n_50),
.B1(n_161),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_45),
.A2(n_50),
.B1(n_181),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_45),
.A2(n_50),
.B1(n_96),
.B2(n_199),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_45),
.A2(n_50),
.B1(n_92),
.B2(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_45),
.A2(n_50),
.B1(n_235),
.B2(n_268),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_45),
.A2(n_50),
.B1(n_53),
.B2(n_268),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_50),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_47),
.B(n_58),
.Y(n_191)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_48),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_48),
.A2(n_49),
.B(n_106),
.C(n_157),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_50),
.B(n_106),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_51),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_52),
.B(n_169),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_54),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_61),
.B2(n_62),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_55),
.A2(n_56),
.B1(n_62),
.B2(n_300),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_56),
.A2(n_61),
.B(n_62),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_56),
.A2(n_62),
.B1(n_134),
.B2(n_136),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_56),
.A2(n_62),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_60),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_57),
.A2(n_60),
.B1(n_102),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_57),
.A2(n_60),
.B1(n_135),
.B2(n_195),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_57),
.A2(n_60),
.B1(n_116),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_57),
.A2(n_60),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_63),
.A2(n_64),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_65),
.A2(n_68),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_65),
.A2(n_68),
.B1(n_114),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_65),
.A2(n_68),
.B1(n_242),
.B2(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_69),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_328),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_73),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_324),
.B(n_330),
.Y(n_75)
);

OAI321xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_293),
.A3(n_316),
.B1(n_322),
.B2(n_323),
.C(n_333),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_272),
.B(n_292),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_79),
.A2(n_248),
.B(n_271),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_141),
.B(n_224),
.C(n_247),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_126),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_81),
.B(n_126),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_109),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_93),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_83),
.B(n_93),
.C(n_109),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_84),
.B(n_89),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_85),
.A2(n_87),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_85),
.A2(n_86),
.B1(n_122),
.B2(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_85),
.A2(n_123),
.B1(n_151),
.B2(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_85),
.A2(n_86),
.B1(n_153),
.B2(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_85),
.A2(n_86),
.B1(n_140),
.B2(n_183),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_85),
.A2(n_88),
.B1(n_125),
.B2(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_85),
.A2(n_86),
.B(n_233),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_86),
.B(n_106),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_98),
.C(n_104),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_94),
.A2(n_95),
.B1(n_98),
.B2(n_99),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g109 ( 
.A(n_110),
.B(n_118),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_117),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_111),
.B(n_117),
.C(n_118),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_115),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_121),
.Y(n_130)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_148)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.C(n_131),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_127),
.B(n_221),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_129),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.C(n_138),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_133),
.B(n_209),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_223),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_218),
.B(n_222),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_204),
.B(n_217),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_185),
.B(n_203),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_173),
.B(n_184),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_162),
.B(n_172),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_154),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_148),
.B(n_154),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_158),
.B2(n_159),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_158),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_167),
.B(n_171),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_166),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_174),
.B(n_175),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_177),
.B(n_180),
.C(n_182),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_193),
.B1(n_201),
.B2(n_202),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_188),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_190),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_192),
.Y(n_196)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_194),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_200),
.C(n_201),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_205),
.B(n_206),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_214),
.C(n_215),
.Y(n_219)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_213),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_219),
.B(n_220),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_225),
.B(n_226),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_229),
.B2(n_246),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_227),
.Y(n_246)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_236),
.B2(n_237),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_230),
.B(n_237),
.C(n_246),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_234),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_234),
.Y(n_254)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_240),
.C(n_245),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_243),
.B2(n_245),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_243),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_249),
.B(n_250),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_270),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_263),
.B2(n_264),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_264),
.C(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_256),
.C(n_260),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_259),
.B2(n_260),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_258),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_262),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_269),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_265),
.A2(n_266),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_267),
.Y(n_284)
);

AOI21xp33_ASAP7_75t_L g307 ( 
.A1(n_266),
.A2(n_284),
.B(n_287),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_267),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_273),
.B(n_274),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_290),
.B2(n_291),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_283),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_277),
.B(n_283),
.C(n_291),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B(n_282),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_281),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_282),
.B(n_295),
.C(n_306),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_282),
.A2(n_295),
.B1(n_296),
.B2(n_321),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_282),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_289),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_290),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_308),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_302),
.B1(n_304),
.B2(n_305),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_297),
.Y(n_304)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_299),
.B(n_301),
.C(n_302),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_302),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_302),
.A2(n_305),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_310),
.C(n_315),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_306),
.A2(n_307),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_315),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_318),
.Y(n_322)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_326),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_327),
.Y(n_329)
);


endmodule