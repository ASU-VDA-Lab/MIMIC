module real_jpeg_26185_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_15;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx3_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_1),
.A2(n_35),
.B1(n_40),
.B2(n_44),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_1),
.A2(n_35),
.B1(n_67),
.B2(n_69),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_1),
.A2(n_35),
.B1(n_55),
.B2(n_56),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_2),
.A2(n_40),
.B1(n_44),
.B2(n_47),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_2),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_2),
.A2(n_47),
.B1(n_55),
.B2(n_56),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_47),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_2),
.A2(n_59),
.B(n_107),
.C(n_108),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_2),
.A2(n_47),
.B1(n_62),
.B2(n_67),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_2),
.B(n_54),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_2),
.A2(n_56),
.B(n_75),
.C(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_24),
.C(n_43),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_2),
.B(n_132),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_2),
.B(n_90),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_2),
.B(n_45),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_4),
.A2(n_26),
.B1(n_40),
.B2(n_44),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_55),
.B1(n_56),
.B2(n_63),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_7),
.A2(n_40),
.B1(n_44),
.B2(n_63),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_63),
.Y(n_188)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_8),
.Y(n_76)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_11),
.Y(n_91)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_11),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_135),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_133),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_111),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_15),
.B(n_111),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_95),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_82),
.B2(n_83),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_50),
.B2(n_51),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_36),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_21),
.B(n_36),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_27),
.B(n_29),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_22),
.A2(n_94),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_23),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_24),
.B(n_200),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_27),
.B(n_34),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_27),
.B(n_93),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_27),
.A2(n_93),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_27),
.B(n_187),
.Y(n_186)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_30),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_30),
.B(n_186),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_48),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_37),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_46),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_38),
.B(n_49),
.Y(n_87)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_38),
.B(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_45),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_39)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_40),
.A2(n_44),
.B1(n_75),
.B2(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_40),
.B(n_176),
.Y(n_175)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_44),
.A2(n_47),
.B(n_77),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_45),
.B(n_156),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_46),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g107 ( 
.A1(n_47),
.A2(n_56),
.B(n_58),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_48),
.B(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_71),
.B1(n_72),
.B2(n_81),
.Y(n_51)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_64),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_53),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_68),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_58),
.B2(n_59),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_55),
.A2(n_56),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_58),
.A2(n_59),
.B1(n_62),
.B2(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_60),
.B(n_65),
.Y(n_99)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_65),
.B(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_78),
.B(n_79),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_73),
.B(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_73),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_78),
.B(n_79),
.Y(n_104)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_78),
.B(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_80),
.B(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_88),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_86),
.B(n_87),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_85),
.A2(n_125),
.B(n_126),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_85),
.B(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_87),
.B(n_173),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_94),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_89),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_94),
.B(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_100),
.C(n_105),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_97),
.B1(n_100),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_100),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_109),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_117),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_112),
.A2(n_113),
.B1(n_230),
.B2(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_116),
.Y(n_232)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_127),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_119),
.A2(n_120),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_123),
.A2(n_124),
.B1(n_127),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_214),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_233),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_227),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_167),
.B(n_226),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_157),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_139),
.B(n_157),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.C(n_152),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_140),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_145),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_142),
.B(n_143),
.C(n_145),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_144),
.B(n_202),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_147),
.B(n_152),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_148),
.A2(n_150),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_148),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_150),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

INVxp33_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_161),
.C(n_162),
.Y(n_228)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_221),
.B(n_225),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_209),
.B(n_220),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_190),
.B(n_208),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_177),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_171),
.B(n_177),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_172),
.A2(n_174),
.B1(n_175),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_184),
.B2(n_189),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_180),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_183),
.C(n_189),
.Y(n_210)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_188),
.B(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_191),
.A2(n_197),
.B(n_207),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_192),
.B(n_195),
.Y(n_207)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_193),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_203),
.B(n_206),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_210),
.B(n_211),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_217),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_216),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_216),
.C(n_217),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_222),
.B(n_223),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_229),
.Y(n_233)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);


endmodule