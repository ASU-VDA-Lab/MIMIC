module fake_jpeg_4146_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_152;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_40),
.Y(n_42)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_7),
.Y(n_38)
);

OR2x4_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_21),
.B(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_21),
.B1(n_16),
.B2(n_22),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_43),
.A2(n_52),
.B1(n_55),
.B2(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_48),
.Y(n_61)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_45),
.A2(n_35),
.B1(n_24),
.B2(n_31),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_46),
.B(n_60),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_38),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_47),
.Y(n_79)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_54),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_32),
.B1(n_22),
.B2(n_16),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_22),
.B1(n_21),
.B2(n_16),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_53),
.A2(n_23),
.B(n_18),
.Y(n_88)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_34),
.A2(n_32),
.B1(n_17),
.B2(n_27),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_39),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_24),
.B1(n_35),
.B2(n_37),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_87),
.B1(n_41),
.B2(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_65),
.Y(n_95)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_68),
.Y(n_94)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_67),
.Y(n_101)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_70),
.A2(n_85),
.B(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_34),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_25),
.Y(n_92)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_28),
.B1(n_30),
.B2(n_26),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_41),
.B1(n_20),
.B2(n_18),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_86),
.Y(n_104)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_60),
.A2(n_40),
.B(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_41),
.A2(n_40),
.B1(n_28),
.B2(n_17),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_79),
.B(n_30),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_89),
.B(n_93),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_72),
.B(n_49),
.C(n_48),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_91),
.C(n_99),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_54),
.C(n_59),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_108),
.B1(n_18),
.B2(n_29),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_61),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_71),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_25),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_86),
.Y(n_119)
);

MAJx2_ASAP7_75t_L g99 ( 
.A(n_63),
.B(n_39),
.C(n_33),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_111),
.B1(n_69),
.B2(n_76),
.Y(n_121)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_85),
.B(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_56),
.B1(n_25),
.B2(n_29),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_83),
.A2(n_20),
.B1(n_18),
.B2(n_25),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_39),
.C(n_33),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_56),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_63),
.B1(n_88),
.B2(n_64),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_115),
.B(n_116),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_117),
.B(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_122),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_84),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_130),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_137),
.B1(n_140),
.B2(n_107),
.Y(n_149)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_124),
.B(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_95),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_92),
.A2(n_80),
.B1(n_68),
.B2(n_66),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_131),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_25),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_96),
.B(n_62),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_132),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_97),
.A2(n_69),
.B1(n_25),
.B2(n_39),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_62),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

INVx13_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_100),
.A2(n_29),
.B1(n_20),
.B2(n_18),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_91),
.Y(n_138)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

OR2x4_ASAP7_75t_L g139 ( 
.A(n_99),
.B(n_109),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_141),
.B(n_126),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_110),
.A2(n_9),
.B(n_1),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_29),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_119),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_148),
.B(n_151),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_149),
.A2(n_171),
.B1(n_122),
.B2(n_131),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_100),
.Y(n_151)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_139),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_154),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_134),
.B(n_90),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_193)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_115),
.Y(n_157)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.C(n_4),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_114),
.C(n_104),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_104),
.B(n_106),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_1),
.B(n_5),
.Y(n_195)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_127),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_164),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_112),
.C(n_99),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_163),
.B(n_128),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_120),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_165),
.B(n_166),
.Y(n_188)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_133),
.B(n_108),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_167),
.A2(n_19),
.B(n_2),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_124),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_123),
.A2(n_89),
.B1(n_101),
.B2(n_19),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_175),
.C(n_177),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_117),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_117),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_178),
.A2(n_192),
.B1(n_195),
.B2(n_151),
.Y(n_210)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_180),
.B(n_181),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_161),
.B(n_125),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_144),
.A2(n_116),
.B1(n_136),
.B2(n_101),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_183),
.B1(n_191),
.B2(n_164),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_116),
.B1(n_19),
.B2(n_0),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_150),
.B(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_190),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_189),
.Y(n_214)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_145),
.A2(n_19),
.B1(n_3),
.B2(n_5),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_153),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_194),
.B(n_165),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_148),
.B(n_6),
.Y(n_196)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_196),
.Y(n_204)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_166),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_200),
.A2(n_202),
.B(n_207),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_150),
.Y(n_202)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_173),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_208),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_147),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_209),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_210),
.A2(n_212),
.B1(n_190),
.B2(n_158),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_147),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_215),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_192),
.A2(n_169),
.B1(n_162),
.B2(n_163),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_217),
.Y(n_220)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_211),
.B(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_219),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_193),
.C(n_177),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_217),
.C(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_193),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_232),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_SL g225 ( 
.A(n_203),
.B(n_160),
.C(n_154),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_167),
.B1(n_179),
.B2(n_168),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_230),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_175),
.Y(n_231)
);

FAx1_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_201),
.CI(n_200),
.CON(n_237),
.SN(n_237)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_195),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_171),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_207),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_240),
.C(n_243),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_229),
.A2(n_215),
.B1(n_208),
.B2(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_235),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_237),
.A2(n_219),
.B(n_225),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_227),
.A2(n_203),
.B1(n_198),
.B2(n_214),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_232),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_220),
.C(n_224),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_226),
.B(n_204),
.C(n_206),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_238),
.B(n_205),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_250),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_233),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_252),
.C(n_253),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_204),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_228),
.C(n_231),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_239),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_236),
.B(n_221),
.C(n_218),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_236),
.C(n_237),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_251),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_8),
.Y(n_267)
);

AO21x1_ASAP7_75t_L g257 ( 
.A1(n_248),
.A2(n_245),
.B(n_237),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_262),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_253),
.B1(n_249),
.B2(n_252),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_263),
.C(n_8),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_143),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_218),
.C(n_152),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_266),
.C(n_268),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_262),
.A2(n_156),
.B(n_143),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_269),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_260),
.A2(n_8),
.B(n_9),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_258),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);

OAI31xp33_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_9),
.A3(n_10),
.B(n_12),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_12),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_275),
.B(n_272),
.C(n_14),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_274),
.B(n_14),
.Y(n_277)
);

OAI31xp33_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_13),
.A3(n_15),
.B(n_273),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_15),
.Y(n_279)
);


endmodule