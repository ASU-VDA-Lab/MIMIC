module fake_netlist_5_2591_n_1480 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1480);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1480;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1370;
wire n_1292;
wire n_1360;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1097;
wire n_1036;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1419;
wire n_693;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

INVx1_ASAP7_75t_L g371 ( 
.A(n_326),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_135),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_168),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_343),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_272),
.B(n_98),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_121),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_110),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_366),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_303),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_367),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_201),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_287),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_163),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_105),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_196),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_347),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_190),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_306),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_162),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_64),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_161),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_159),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_19),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_14),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_93),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_362),
.Y(n_398)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_40),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_248),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_128),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_314),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_319),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_36),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_238),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_55),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_212),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_255),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g409 ( 
.A(n_80),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_209),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_262),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_88),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_97),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_296),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_222),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_121),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_361),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_270),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_L g420 ( 
.A(n_74),
.B(n_297),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_193),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_66),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_75),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_195),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_365),
.Y(n_425)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_241),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_52),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_169),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_286),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_57),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_48),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_300),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_302),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_143),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_259),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_245),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_36),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_304),
.B(n_82),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_311),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_203),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_250),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_41),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_233),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_206),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_288),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_281),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_112),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_252),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_109),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_43),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_100),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_145),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_52),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_251),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g457 ( 
.A(n_357),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_140),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_147),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_89),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_119),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_256),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_182),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_282),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_50),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_277),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_352),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_231),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_185),
.Y(n_469)
);

BUFx5_ASAP7_75t_L g470 ( 
.A(n_146),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_170),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_338),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_349),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_68),
.Y(n_474)
);

CKINVDCx14_ASAP7_75t_R g475 ( 
.A(n_214),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_254),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_74),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_3),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_200),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_27),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_118),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_229),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_63),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_165),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_340),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_348),
.Y(n_486)
);

CKINVDCx14_ASAP7_75t_R g487 ( 
.A(n_312),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_25),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_102),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_58),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_184),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_316),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_86),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g494 ( 
.A(n_305),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_166),
.B(n_197),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_230),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_44),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_310),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_204),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_125),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_315),
.B(n_358),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_235),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_198),
.B(n_242),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_336),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_178),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_127),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_268),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_39),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_226),
.Y(n_509)
);

HB1xp67_ASAP7_75t_L g510 ( 
.A(n_354),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_301),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_313),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_57),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_101),
.Y(n_514)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_202),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_249),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_23),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_137),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_299),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_171),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_351),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_95),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_45),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_263),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_264),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_298),
.B(n_56),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_329),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_149),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_324),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_67),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_70),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_188),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_174),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_65),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_156),
.Y(n_535)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_12),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_220),
.Y(n_537)
);

NOR2xp67_ASAP7_75t_L g538 ( 
.A(n_323),
.B(n_83),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_211),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_3),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_16),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_158),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_216),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_356),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_79),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_84),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_120),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_54),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_71),
.Y(n_549)
);

INVxp67_ASAP7_75t_SL g550 ( 
.A(n_225),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_164),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_317),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_232),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_322),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_76),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_258),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_399),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_409),
.B(n_0),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_409),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_406),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_406),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_138),
.B(n_136),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_520),
.B(n_0),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_406),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_473),
.B(n_1),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_536),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_SL g567 ( 
.A(n_390),
.B(n_436),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_467),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_473),
.B(n_510),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_426),
.B(n_139),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g571 ( 
.A1(n_377),
.A2(n_392),
.B1(n_404),
.B2(n_523),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_L g572 ( 
.A1(n_378),
.A2(n_5),
.B1(n_2),
.B2(n_4),
.Y(n_572)
);

OAI22x1_ASAP7_75t_SL g573 ( 
.A1(n_372),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_510),
.B(n_6),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_504),
.B(n_7),
.Y(n_575)
);

INVxp33_ASAP7_75t_SL g576 ( 
.A(n_396),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_483),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_523),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_460),
.A2(n_514),
.B1(n_376),
.B2(n_449),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_483),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_401),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_426),
.Y(n_582)
);

BUFx12f_ASAP7_75t_L g583 ( 
.A(n_399),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

INVx6_ASAP7_75t_L g585 ( 
.A(n_467),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_545),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_393),
.B(n_8),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_470),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_426),
.Y(n_589)
);

NAND2x1_ASAP7_75t_L g590 ( 
.A(n_426),
.B(n_141),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_466),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_546),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_376),
.A2(n_449),
.B1(n_378),
.B2(n_489),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_547),
.Y(n_594)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_422),
.A2(n_433),
.B1(n_452),
.B2(n_423),
.Y(n_595)
);

CKINVDCx16_ASAP7_75t_R g596 ( 
.A(n_491),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_414),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_470),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_470),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_386),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_457),
.B(n_9),
.Y(n_601)
);

BUFx8_ASAP7_75t_L g602 ( 
.A(n_526),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_466),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_395),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_397),
.Y(n_605)
);

INVx5_ASAP7_75t_L g606 ( 
.A(n_466),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_459),
.B(n_10),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_466),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_412),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_413),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_416),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_492),
.Y(n_612)
);

AOI22x1_ASAP7_75t_SL g613 ( 
.A1(n_455),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_428),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_419),
.Y(n_615)
);

OA21x2_ASAP7_75t_L g616 ( 
.A1(n_371),
.A2(n_375),
.B(n_374),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_398),
.B(n_435),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_432),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g619 ( 
.A1(n_447),
.A2(n_471),
.B(n_448),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_439),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_444),
.Y(n_622)
);

NAND2x1_ASAP7_75t_L g623 ( 
.A(n_492),
.B(n_142),
.Y(n_623)
);

BUFx6f_ASAP7_75t_L g624 ( 
.A(n_492),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_484),
.B(n_11),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_496),
.B(n_14),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_451),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_524),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_453),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_465),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_478),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_480),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_535),
.B(n_15),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_481),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_454),
.B(n_15),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_498),
.B(n_16),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_457),
.B(n_17),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_597),
.B(n_615),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_582),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_560),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_564),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_570),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_559),
.B(n_475),
.Y(n_644)
);

AOI22xp33_ASAP7_75t_L g645 ( 
.A1(n_569),
.A2(n_487),
.B1(n_475),
.B2(n_464),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_617),
.B(n_487),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_616),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_617),
.B(n_379),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_616),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_561),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_585),
.Y(n_651)
);

OR2x6_ASAP7_75t_L g652 ( 
.A(n_569),
.B(n_420),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_606),
.B(n_601),
.Y(n_653)
);

AND3x2_ASAP7_75t_L g654 ( 
.A(n_558),
.B(n_435),
.C(n_398),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_594),
.B(n_494),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_524),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_585),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_606),
.B(n_380),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_568),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_619),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_570),
.Y(n_661)
);

AND2x6_ASAP7_75t_L g662 ( 
.A(n_635),
.B(n_503),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_582),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_606),
.B(n_381),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_567),
.B(n_515),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_596),
.B(n_594),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_635),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_583),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_582),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_581),
.B(n_490),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_579),
.B(n_474),
.C(n_461),
.Y(n_671)
);

INVx2_ASAP7_75t_SL g672 ( 
.A(n_637),
.Y(n_672)
);

BUFx10_ASAP7_75t_L g673 ( 
.A(n_637),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_584),
.B(n_493),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_576),
.B(n_550),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_557),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_589),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_565),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_586),
.Y(n_679)
);

INVx5_ASAP7_75t_L g680 ( 
.A(n_570),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_589),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_575),
.B(n_517),
.C(n_477),
.Y(n_682)
);

AOI22xp5_ASAP7_75t_L g683 ( 
.A1(n_567),
.A2(n_394),
.B1(n_402),
.B2(n_388),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_593),
.B(n_440),
.Y(n_684)
);

INVx4_ASAP7_75t_L g685 ( 
.A(n_570),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_577),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_565),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_563),
.B(n_530),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_563),
.B(n_531),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_592),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_589),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_595),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_603),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_591),
.B(n_385),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_666),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_646),
.Y(n_696)
);

INVx2_ASAP7_75t_SL g697 ( 
.A(n_651),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_645),
.B(n_593),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_655),
.B(n_595),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_663),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_651),
.Y(n_701)
);

INVx2_ASAP7_75t_SL g702 ( 
.A(n_651),
.Y(n_702)
);

HB1xp67_ASAP7_75t_L g703 ( 
.A(n_655),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_675),
.B(n_579),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_672),
.B(n_591),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_672),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_653),
.B(n_580),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_678),
.B(n_495),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_678),
.B(n_603),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_687),
.B(n_501),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_687),
.B(n_603),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_662),
.B(n_608),
.Y(n_712)
);

INVx4_ASAP7_75t_L g713 ( 
.A(n_693),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_662),
.B(n_608),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_684),
.B(n_574),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_681),
.Y(n_716)
);

O2A1O1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_648),
.A2(n_607),
.B(n_587),
.C(n_625),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_669),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_644),
.B(n_634),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_640),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_659),
.Y(n_721)
);

NOR2x2_ASAP7_75t_L g722 ( 
.A(n_652),
.B(n_573),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_670),
.B(n_620),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_668),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_640),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_639),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_676),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_684),
.B(n_607),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_669),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_662),
.B(n_608),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_662),
.B(n_612),
.Y(n_731)
);

AND3x1_ASAP7_75t_L g732 ( 
.A(n_683),
.B(n_566),
.C(n_578),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_652),
.B(n_626),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_657),
.B(n_652),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_691),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_662),
.B(n_612),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_657),
.B(n_652),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_667),
.B(n_636),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_662),
.A2(n_633),
.B1(n_500),
.B2(n_506),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_667),
.B(n_604),
.Y(n_740)
);

OR2x2_ASAP7_75t_L g741 ( 
.A(n_692),
.B(n_571),
.Y(n_741)
);

NOR2xp67_ASAP7_75t_L g742 ( 
.A(n_690),
.B(n_373),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_640),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_689),
.B(n_612),
.Y(n_744)
);

OAI21xp5_ASAP7_75t_L g745 ( 
.A1(n_647),
.A2(n_562),
.B(n_550),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_677),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_647),
.A2(n_508),
.B1(n_513),
.B2(n_497),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_689),
.B(n_677),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_677),
.B(n_621),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_691),
.Y(n_750)
);

NAND2x1p5_ASAP7_75t_L g751 ( 
.A(n_680),
.B(n_590),
.Y(n_751)
);

A2O1A1Ixp33_ASAP7_75t_L g752 ( 
.A1(n_649),
.A2(n_588),
.B(n_599),
.C(n_598),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_671),
.B(n_602),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_656),
.B(n_621),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_L g755 ( 
.A(n_694),
.B(n_602),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_656),
.B(n_621),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_649),
.B(n_624),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_693),
.B(n_624),
.Y(n_758)
);

OR2x6_ASAP7_75t_L g759 ( 
.A(n_665),
.B(n_572),
.Y(n_759)
);

NOR3xp33_ASAP7_75t_L g760 ( 
.A(n_665),
.B(n_572),
.C(n_566),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_679),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_641),
.B(n_642),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_679),
.B(n_600),
.Y(n_763)
);

AOI21xp5_ASAP7_75t_L g764 ( 
.A1(n_660),
.A2(n_664),
.B(n_658),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_654),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_650),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_641),
.B(n_628),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_681),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_682),
.B(n_628),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_728),
.B(n_673),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_696),
.B(n_660),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_728),
.A2(n_688),
.B(n_503),
.C(n_538),
.Y(n_772)
);

OAI21xp5_ASAP7_75t_L g773 ( 
.A1(n_745),
.A2(n_661),
.B(n_643),
.Y(n_773)
);

OAI21xp5_ASAP7_75t_L g774 ( 
.A1(n_752),
.A2(n_661),
.B(n_643),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_696),
.B(n_673),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_715),
.B(n_673),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_715),
.B(n_685),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_739),
.B(n_685),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_716),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_739),
.B(n_685),
.Y(n_780)
);

NAND2x1p5_ASAP7_75t_L g781 ( 
.A(n_695),
.B(n_680),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_747),
.B(n_688),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_766),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_717),
.A2(n_623),
.B(n_400),
.C(n_408),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_747),
.B(n_703),
.Y(n_785)
);

BUFx2_ASAP7_75t_L g786 ( 
.A(n_727),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_704),
.A2(n_537),
.B1(n_539),
.B2(n_442),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_703),
.A2(n_543),
.B1(n_391),
.B2(n_411),
.Y(n_788)
);

NOR2xp33_ASAP7_75t_SL g789 ( 
.A(n_701),
.B(n_382),
.Y(n_789)
);

O2A1O1Ixp5_ASAP7_75t_L g790 ( 
.A1(n_757),
.A2(n_708),
.B(n_710),
.C(n_748),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_760),
.A2(n_417),
.B1(n_418),
.B2(n_415),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_730),
.A2(n_736),
.B(n_731),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_733),
.A2(n_424),
.B1(n_425),
.B2(n_421),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_706),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_706),
.B(n_690),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_719),
.B(n_670),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_726),
.B(n_709),
.Y(n_797)
);

INVx3_ASAP7_75t_L g798 ( 
.A(n_723),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_698),
.A2(n_674),
.B(n_534),
.C(n_540),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_700),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_762),
.Y(n_801)
);

OAI21xp5_ASAP7_75t_L g802 ( 
.A1(n_764),
.A2(n_429),
.B(n_427),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_711),
.B(n_740),
.Y(n_803)
);

OR2x6_ASAP7_75t_SL g804 ( 
.A(n_741),
.B(n_555),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_698),
.A2(n_431),
.B1(n_434),
.B2(n_430),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_699),
.B(n_383),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_708),
.B(n_686),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_710),
.B(n_571),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_SL g809 ( 
.A(n_721),
.B(n_384),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_723),
.Y(n_810)
);

O2A1O1Ixp33_ASAP7_75t_L g811 ( 
.A1(n_760),
.A2(n_674),
.B(n_548),
.C(n_549),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_705),
.A2(n_441),
.B1(n_445),
.B2(n_437),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_R g813 ( 
.A(n_724),
.B(n_387),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_707),
.B(n_446),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_759),
.A2(n_578),
.B(n_605),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_738),
.B(n_609),
.Y(n_816)
);

OR2x6_ASAP7_75t_SL g817 ( 
.A(n_722),
.B(n_573),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_769),
.A2(n_522),
.B(n_611),
.C(n_610),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_718),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_763),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_734),
.A2(n_403),
.B1(n_405),
.B2(n_389),
.Y(n_821)
);

NAND2x1p5_ASAP7_75t_L g822 ( 
.A(n_697),
.B(n_618),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_737),
.B(n_407),
.Y(n_823)
);

O2A1O1Ixp33_ASAP7_75t_L g824 ( 
.A1(n_744),
.A2(n_759),
.B(n_756),
.C(n_754),
.Y(n_824)
);

AND2x4_ASAP7_75t_L g825 ( 
.A(n_713),
.B(n_627),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_758),
.A2(n_458),
.B(n_456),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_720),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_759),
.A2(n_630),
.B(n_631),
.C(n_629),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_742),
.B(n_462),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_753),
.A2(n_732),
.B1(n_755),
.B2(n_765),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_729),
.B(n_463),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_749),
.A2(n_472),
.B(n_469),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_702),
.B(n_410),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_735),
.B(n_476),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_767),
.A2(n_482),
.B(n_479),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_716),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_763),
.B(n_753),
.C(n_632),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_750),
.B(n_486),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_725),
.A2(n_505),
.B(n_499),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_716),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_743),
.A2(n_511),
.B(n_509),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_746),
.A2(n_516),
.B(n_512),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_751),
.A2(n_519),
.B1(n_521),
.B2(n_518),
.Y(n_843)
);

OAI22x1_ASAP7_75t_L g844 ( 
.A1(n_768),
.A2(n_613),
.B1(n_528),
.B2(n_542),
.Y(n_844)
);

OR2x6_ASAP7_75t_L g845 ( 
.A(n_751),
.B(n_614),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_716),
.B(n_525),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_739),
.A2(n_551),
.B1(n_553),
.B2(n_544),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_728),
.A2(n_556),
.B(n_554),
.C(n_614),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_712),
.A2(n_443),
.B(n_438),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_761),
.B(n_622),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_696),
.B(n_450),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_696),
.B(n_468),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_706),
.B(n_485),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_766),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_706),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_696),
.B(n_502),
.Y(n_856)
);

OR2x6_ASAP7_75t_SL g857 ( 
.A(n_741),
.B(n_507),
.Y(n_857)
);

BUFx3_ASAP7_75t_L g858 ( 
.A(n_761),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_728),
.B(n_527),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_706),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_739),
.A2(n_532),
.B1(n_533),
.B2(n_529),
.Y(n_861)
);

OR2x6_ASAP7_75t_L g862 ( 
.A(n_721),
.B(n_17),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_728),
.A2(n_552),
.B(n_20),
.C(n_18),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_728),
.A2(n_20),
.B(n_18),
.C(n_19),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_706),
.Y(n_865)
);

OAI22xp5_ASAP7_75t_L g866 ( 
.A1(n_739),
.A2(n_148),
.B1(n_150),
.B2(n_144),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_695),
.B(n_151),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_712),
.A2(n_153),
.B(n_152),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_716),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_696),
.B(n_21),
.Y(n_870)
);

INVxp67_ASAP7_75t_SL g871 ( 
.A(n_779),
.Y(n_871)
);

A2O1A1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_772),
.A2(n_808),
.B(n_782),
.C(n_824),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_790),
.A2(n_23),
.B(n_21),
.C(n_22),
.Y(n_873)
);

AO31x2_ASAP7_75t_L g874 ( 
.A1(n_784),
.A2(n_25),
.A3(n_22),
.B(n_24),
.Y(n_874)
);

AO31x2_ASAP7_75t_L g875 ( 
.A1(n_792),
.A2(n_29),
.A3(n_26),
.B(n_28),
.Y(n_875)
);

OA21x2_ASAP7_75t_L g876 ( 
.A1(n_773),
.A2(n_155),
.B(n_154),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_777),
.A2(n_774),
.B(n_778),
.Y(n_877)
);

BUFx10_ASAP7_75t_L g878 ( 
.A(n_852),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_801),
.B(n_28),
.Y(n_879)
);

OAI21xp5_ASAP7_75t_L g880 ( 
.A1(n_780),
.A2(n_160),
.B(n_157),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_803),
.B(n_820),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_786),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_783),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_785),
.A2(n_31),
.B(n_29),
.C(n_30),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_797),
.B(n_30),
.Y(n_885)
);

AOI22xp5_ASAP7_75t_L g886 ( 
.A1(n_830),
.A2(n_172),
.B1(n_173),
.B2(n_167),
.Y(n_886)
);

INVx5_ASAP7_75t_L g887 ( 
.A(n_779),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_811),
.A2(n_33),
.B(n_31),
.C(n_32),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_787),
.A2(n_176),
.B1(n_177),
.B2(n_175),
.Y(n_889)
);

OAI21x1_ASAP7_75t_SL g890 ( 
.A1(n_802),
.A2(n_180),
.B(n_179),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_865),
.Y(n_891)
);

AOI21xp33_ASAP7_75t_L g892 ( 
.A1(n_859),
.A2(n_32),
.B(n_33),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_810),
.B(n_181),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_813),
.Y(n_894)
);

INVx3_ASAP7_75t_SL g895 ( 
.A(n_862),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_794),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_858),
.B(n_183),
.Y(n_897)
);

BUFx12f_ASAP7_75t_L g898 ( 
.A(n_862),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_850),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_771),
.B(n_34),
.Y(n_900)
);

AOI31xp67_ASAP7_75t_L g901 ( 
.A1(n_800),
.A2(n_187),
.A3(n_189),
.B(n_186),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_854),
.Y(n_902)
);

AOI221x1_ASAP7_75t_L g903 ( 
.A1(n_805),
.A2(n_194),
.B1(n_199),
.B2(n_192),
.C(n_191),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_799),
.A2(n_37),
.B(n_34),
.C(n_35),
.Y(n_904)
);

AO31x2_ASAP7_75t_L g905 ( 
.A1(n_793),
.A2(n_38),
.A3(n_35),
.B(n_37),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_798),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_850),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_SL g908 ( 
.A1(n_863),
.A2(n_40),
.B(n_38),
.C(n_39),
.Y(n_908)
);

AOI221x1_ASAP7_75t_L g909 ( 
.A1(n_848),
.A2(n_208),
.B1(n_210),
.B2(n_207),
.C(n_205),
.Y(n_909)
);

AO31x2_ASAP7_75t_L g910 ( 
.A1(n_866),
.A2(n_43),
.A3(n_41),
.B(n_42),
.Y(n_910)
);

AO32x2_ASAP7_75t_L g911 ( 
.A1(n_788),
.A2(n_42),
.A3(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_796),
.B(n_46),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_770),
.A2(n_837),
.B(n_847),
.Y(n_913)
);

INVxp67_ASAP7_75t_L g914 ( 
.A(n_870),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_795),
.Y(n_915)
);

CKINVDCx20_ASAP7_75t_R g916 ( 
.A(n_806),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_816),
.B(n_47),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_855),
.Y(n_918)
);

OAI22xp33_ASAP7_75t_L g919 ( 
.A1(n_775),
.A2(n_809),
.B1(n_856),
.B2(n_851),
.Y(n_919)
);

O2A1O1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_864),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_860),
.Y(n_921)
);

A2O1A1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_828),
.A2(n_54),
.B(n_51),
.C(n_53),
.Y(n_922)
);

A2O1A1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_815),
.A2(n_56),
.B(n_53),
.C(n_55),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_822),
.Y(n_924)
);

OAI21xp5_ASAP7_75t_SL g925 ( 
.A1(n_791),
.A2(n_58),
.B(n_59),
.Y(n_925)
);

AO31x2_ASAP7_75t_L g926 ( 
.A1(n_846),
.A2(n_62),
.A3(n_60),
.B(n_61),
.Y(n_926)
);

INVx3_ASAP7_75t_SL g927 ( 
.A(n_833),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_819),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_L g929 ( 
.A(n_853),
.B(n_65),
.C(n_66),
.Y(n_929)
);

AO21x2_ASAP7_75t_L g930 ( 
.A1(n_823),
.A2(n_215),
.B(n_213),
.Y(n_930)
);

AO21x1_ASAP7_75t_L g931 ( 
.A1(n_861),
.A2(n_67),
.B(n_68),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_821),
.B(n_69),
.C(n_70),
.Y(n_932)
);

O2A1O1Ixp5_ASAP7_75t_L g933 ( 
.A1(n_814),
.A2(n_218),
.B(n_219),
.C(n_217),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_825),
.B(n_221),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_807),
.A2(n_224),
.B(n_223),
.Y(n_935)
);

AO31x2_ASAP7_75t_L g936 ( 
.A1(n_812),
.A2(n_72),
.A3(n_69),
.B(n_71),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_789),
.B(n_72),
.C(n_73),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_825),
.A2(n_76),
.B(n_73),
.C(n_75),
.Y(n_938)
);

CKINVDCx11_ASAP7_75t_R g939 ( 
.A(n_817),
.Y(n_939)
);

INVx5_ASAP7_75t_L g940 ( 
.A(n_836),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_818),
.A2(n_829),
.B(n_826),
.C(n_831),
.Y(n_941)
);

AND2x4_ASAP7_75t_L g942 ( 
.A(n_827),
.B(n_227),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_840),
.B(n_228),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_857),
.B(n_77),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_834),
.A2(n_79),
.B(n_77),
.C(n_78),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_804),
.B(n_78),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_840),
.A2(n_236),
.B(n_234),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_840),
.A2(n_239),
.B(n_237),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_869),
.B(n_240),
.Y(n_949)
);

OAI22xp5_ASAP7_75t_L g950 ( 
.A1(n_845),
.A2(n_285),
.B1(n_369),
.B2(n_368),
.Y(n_950)
);

AO32x2_ASAP7_75t_L g951 ( 
.A1(n_843),
.A2(n_81),
.A3(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_951)
);

AO32x2_ASAP7_75t_L g952 ( 
.A1(n_844),
.A2(n_81),
.A3(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_952)
);

OAI22x1_ASAP7_75t_L g953 ( 
.A1(n_867),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_953)
);

OAI21xp5_ASAP7_75t_L g954 ( 
.A1(n_849),
.A2(n_244),
.B(n_243),
.Y(n_954)
);

INVx1_ASAP7_75t_SL g955 ( 
.A(n_838),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_832),
.A2(n_89),
.B(n_90),
.C(n_91),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_845),
.Y(n_957)
);

OA21x2_ASAP7_75t_L g958 ( 
.A1(n_835),
.A2(n_247),
.B(n_246),
.Y(n_958)
);

AND2x4_ASAP7_75t_L g959 ( 
.A(n_868),
.B(n_253),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_781),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_839),
.B(n_90),
.Y(n_961)
);

BUFx10_ASAP7_75t_L g962 ( 
.A(n_841),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_842),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_810),
.B(n_257),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_786),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_790),
.A2(n_261),
.B(n_260),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_796),
.B(n_92),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_786),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_792),
.A2(n_266),
.B(n_265),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_783),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_783),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_787),
.B(n_94),
.Y(n_972)
);

CKINVDCx16_ASAP7_75t_R g973 ( 
.A(n_813),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_801),
.B(n_94),
.Y(n_974)
);

INVx8_ASAP7_75t_L g975 ( 
.A(n_825),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_790),
.A2(n_269),
.B(n_267),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_801),
.B(n_95),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_790),
.A2(n_273),
.B(n_271),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_865),
.Y(n_979)
);

AO21x2_ASAP7_75t_L g980 ( 
.A1(n_773),
.A2(n_275),
.B(n_274),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_801),
.B(n_96),
.Y(n_981)
);

AO31x2_ASAP7_75t_L g982 ( 
.A1(n_784),
.A2(n_99),
.A3(n_100),
.B(n_101),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_810),
.B(n_276),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_813),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_792),
.A2(n_279),
.B(n_278),
.Y(n_985)
);

NOR4xp25_ASAP7_75t_L g986 ( 
.A(n_772),
.B(n_99),
.C(n_102),
.D(n_103),
.Y(n_986)
);

A2O1A1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_772),
.A2(n_103),
.B(n_104),
.C(n_105),
.Y(n_987)
);

AO31x2_ASAP7_75t_L g988 ( 
.A1(n_784),
.A2(n_104),
.A3(n_106),
.B(n_107),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_786),
.Y(n_989)
);

INVx3_ASAP7_75t_L g990 ( 
.A(n_810),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_SL g991 ( 
.A(n_786),
.B(n_280),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_801),
.B(n_106),
.Y(n_992)
);

INVx6_ASAP7_75t_L g993 ( 
.A(n_862),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_786),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_776),
.B(n_283),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_783),
.Y(n_996)
);

AO21x2_ASAP7_75t_L g997 ( 
.A1(n_773),
.A2(n_309),
.B(n_364),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_801),
.B(n_107),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_801),
.B(n_108),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_810),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_786),
.Y(n_1001)
);

OA21x2_ASAP7_75t_L g1002 ( 
.A1(n_773),
.A2(n_308),
.B(n_363),
.Y(n_1002)
);

BUFx6f_ASAP7_75t_L g1003 ( 
.A(n_810),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_810),
.Y(n_1004)
);

AO31x2_ASAP7_75t_L g1005 ( 
.A1(n_784),
.A2(n_108),
.A3(n_109),
.B(n_110),
.Y(n_1005)
);

AOI221xp5_ASAP7_75t_L g1006 ( 
.A1(n_815),
.A2(n_111),
.B1(n_112),
.B2(n_113),
.C(n_114),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_790),
.A2(n_318),
.B(n_360),
.Y(n_1007)
);

NOR2x1_ASAP7_75t_L g1008 ( 
.A(n_776),
.B(n_284),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_786),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_783),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_790),
.A2(n_307),
.B(n_359),
.Y(n_1011)
);

NOR2x1_ASAP7_75t_R g1012 ( 
.A(n_894),
.B(n_111),
.Y(n_1012)
);

AOI22xp33_ASAP7_75t_L g1013 ( 
.A1(n_972),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_881),
.B(n_115),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_883),
.Y(n_1015)
);

INVx2_ASAP7_75t_L g1016 ( 
.A(n_902),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_914),
.B(n_116),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_955),
.B(n_116),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_919),
.B(n_117),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_970),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_879),
.B(n_117),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_973),
.Y(n_1022)
);

NAND3xp33_ASAP7_75t_SL g1023 ( 
.A(n_1006),
.B(n_118),
.C(n_119),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_971),
.Y(n_1024)
);

HB1xp67_ASAP7_75t_L g1025 ( 
.A(n_965),
.Y(n_1025)
);

BUFx8_ASAP7_75t_L g1026 ( 
.A(n_989),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_899),
.B(n_893),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_887),
.Y(n_1028)
);

NAND3xp33_ASAP7_75t_L g1029 ( 
.A(n_892),
.B(n_120),
.C(n_122),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_878),
.B(n_122),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_915),
.B(n_123),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_996),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_1010),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_913),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_1034)
);

AO21x2_ASAP7_75t_L g1035 ( 
.A1(n_978),
.A2(n_1011),
.B(n_1007),
.Y(n_1035)
);

OA21x2_ASAP7_75t_L g1036 ( 
.A1(n_880),
.A2(n_320),
.B(n_353),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_974),
.B(n_124),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_977),
.B(n_126),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_994),
.Y(n_1039)
);

NAND2x1p5_ASAP7_75t_L g1040 ( 
.A(n_940),
.B(n_295),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_928),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_1009),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_981),
.B(n_992),
.Y(n_1043)
);

AO31x2_ASAP7_75t_L g1044 ( 
.A1(n_873),
.A2(n_126),
.A3(n_127),
.B(n_128),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_964),
.B(n_325),
.Y(n_1045)
);

NAND2x1p5_ASAP7_75t_L g1046 ( 
.A(n_940),
.B(n_328),
.Y(n_1046)
);

AOI22xp33_ASAP7_75t_L g1047 ( 
.A1(n_932),
.A2(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_906),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_975),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_998),
.B(n_129),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_1001),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_900),
.A2(n_321),
.B(n_350),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_921),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_SL g1054 ( 
.A(n_898),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_SL g1055 ( 
.A(n_984),
.B(n_130),
.C(n_131),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_999),
.B(n_885),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_882),
.B(n_132),
.Y(n_1057)
);

AO21x2_ASAP7_75t_L g1058 ( 
.A1(n_890),
.A2(n_935),
.B(n_980),
.Y(n_1058)
);

NAND2x1p5_ASAP7_75t_L g1059 ( 
.A(n_1003),
.B(n_330),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_975),
.Y(n_1060)
);

AO31x2_ASAP7_75t_L g1061 ( 
.A1(n_909),
.A2(n_133),
.A3(n_134),
.B(n_135),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_891),
.B(n_979),
.Y(n_1062)
);

HB1xp67_ASAP7_75t_L g1063 ( 
.A(n_968),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_916),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_912),
.A2(n_289),
.B(n_290),
.C(n_291),
.Y(n_1065)
);

CKINVDCx20_ASAP7_75t_R g1066 ( 
.A(n_939),
.Y(n_1066)
);

INVx2_ASAP7_75t_SL g1067 ( 
.A(n_896),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_967),
.B(n_292),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_942),
.Y(n_1069)
);

OAI21xp33_ASAP7_75t_SL g1070 ( 
.A1(n_917),
.A2(n_293),
.B(n_294),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_918),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_941),
.A2(n_331),
.B(n_332),
.Y(n_1072)
);

INVx2_ASAP7_75t_SL g1073 ( 
.A(n_993),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_871),
.A2(n_333),
.B(n_334),
.Y(n_1074)
);

NOR2x1_ASAP7_75t_SL g1075 ( 
.A(n_997),
.B(n_335),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_SL g1076 ( 
.A1(n_991),
.A2(n_337),
.B1(n_341),
.B2(n_344),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_934),
.B(n_370),
.Y(n_1077)
);

AND2x4_ASAP7_75t_L g1078 ( 
.A(n_983),
.B(n_345),
.Y(n_1078)
);

CKINVDCx11_ASAP7_75t_R g1079 ( 
.A(n_895),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_963),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_990),
.B(n_1000),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_897),
.B(n_923),
.Y(n_1082)
);

AO31x2_ASAP7_75t_L g1083 ( 
.A1(n_903),
.A2(n_931),
.A3(n_987),
.B(n_904),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_995),
.A2(n_933),
.B(n_1008),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_876),
.A2(n_1002),
.B(n_954),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_1003),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_907),
.Y(n_1087)
);

AND2x6_ASAP7_75t_L g1088 ( 
.A(n_886),
.B(n_959),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_962),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_960),
.B(n_925),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_924),
.B(n_1004),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_874),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_927),
.B(n_1004),
.Y(n_1093)
);

OAI21xp33_ASAP7_75t_SL g1094 ( 
.A1(n_889),
.A2(n_961),
.B(n_943),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_993),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_949),
.A2(n_958),
.B(n_950),
.Y(n_1096)
);

AND2x4_ASAP7_75t_L g1097 ( 
.A(n_957),
.B(n_929),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_938),
.B(n_945),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_944),
.B(n_946),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_920),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_930),
.B(n_937),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_908),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_874),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_952),
.B(n_953),
.Y(n_1104)
);

INVx4_ASAP7_75t_SL g1105 ( 
.A(n_905),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_922),
.B(n_1005),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_982),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_986),
.B(n_888),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_910),
.B(n_956),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_901),
.A2(n_947),
.B(n_948),
.Y(n_1110)
);

AO21x2_ASAP7_75t_L g1111 ( 
.A1(n_884),
.A2(n_875),
.B(n_1005),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_875),
.A2(n_988),
.A3(n_982),
.B(n_910),
.Y(n_1112)
);

INVx1_ASAP7_75t_SL g1113 ( 
.A(n_952),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_905),
.Y(n_1114)
);

NAND2x1p5_ASAP7_75t_L g1115 ( 
.A(n_911),
.B(n_951),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_936),
.Y(n_1116)
);

OR2x2_ASAP7_75t_L g1117 ( 
.A(n_936),
.B(n_926),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_911),
.B(n_951),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_926),
.B(n_899),
.Y(n_1119)
);

BUFx12f_ASAP7_75t_L g1120 ( 
.A(n_965),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_915),
.B(n_796),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_881),
.B(n_728),
.Y(n_1122)
);

INVxp67_ASAP7_75t_L g1123 ( 
.A(n_891),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_SL g1124 ( 
.A1(n_916),
.A2(n_808),
.B1(n_787),
.B2(n_830),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_883),
.Y(n_1125)
);

INVx4_ASAP7_75t_SL g1126 ( 
.A(n_927),
.Y(n_1126)
);

A2O1A1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_872),
.A2(n_728),
.B(n_715),
.C(n_808),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_915),
.B(n_796),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_877),
.A2(n_773),
.B(n_714),
.Y(n_1129)
);

AOI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_919),
.A2(n_715),
.B1(n_830),
.B2(n_728),
.Y(n_1130)
);

NAND2x1p5_ASAP7_75t_L g1131 ( 
.A(n_887),
.B(n_940),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_877),
.A2(n_773),
.B(n_714),
.Y(n_1132)
);

OAI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_872),
.A2(n_877),
.B(n_777),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_883),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_969),
.A2(n_792),
.B(n_985),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_881),
.B(n_728),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_965),
.Y(n_1137)
);

AND2x4_ASAP7_75t_L g1138 ( 
.A(n_899),
.B(n_893),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_881),
.B(n_728),
.Y(n_1139)
);

AO21x2_ASAP7_75t_L g1140 ( 
.A1(n_877),
.A2(n_976),
.B(n_966),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_881),
.B(n_728),
.Y(n_1141)
);

AO21x2_ASAP7_75t_L g1142 ( 
.A1(n_877),
.A2(n_976),
.B(n_966),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_899),
.B(n_893),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_916),
.A2(n_808),
.B1(n_787),
.B2(n_830),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_883),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_883),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_881),
.B(n_728),
.Y(n_1147)
);

OAI21xp33_ASAP7_75t_L g1148 ( 
.A1(n_881),
.A2(n_715),
.B(n_728),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_881),
.B(n_728),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_877),
.A2(n_976),
.B(n_966),
.Y(n_1150)
);

AO21x2_ASAP7_75t_L g1151 ( 
.A1(n_1085),
.A2(n_1133),
.B(n_1132),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1137),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_1121),
.B(n_1128),
.Y(n_1153)
);

AO21x2_ASAP7_75t_L g1154 ( 
.A1(n_1129),
.A2(n_1110),
.B(n_1096),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1025),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1015),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1020),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1024),
.Y(n_1158)
);

OR2x6_ASAP7_75t_L g1159 ( 
.A(n_1045),
.B(n_1078),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1032),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1033),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1122),
.B(n_1136),
.Y(n_1162)
);

AND2x2_ASAP7_75t_L g1163 ( 
.A(n_1124),
.B(n_1144),
.Y(n_1163)
);

HB1xp67_ASAP7_75t_L g1164 ( 
.A(n_1039),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1041),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_1139),
.B(n_1141),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1125),
.Y(n_1167)
);

AOI221xp5_ASAP7_75t_L g1168 ( 
.A1(n_1099),
.A2(n_1127),
.B1(n_1023),
.B2(n_1148),
.C(n_1013),
.Y(n_1168)
);

INVx2_ASAP7_75t_SL g1169 ( 
.A(n_1063),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1031),
.B(n_1147),
.Y(n_1170)
);

OAI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1130),
.A2(n_1149),
.B1(n_1082),
.B2(n_1090),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1051),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_1062),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1071),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_1067),
.Y(n_1175)
);

AO21x2_ASAP7_75t_L g1176 ( 
.A1(n_1140),
.A2(n_1142),
.B(n_1084),
.Y(n_1176)
);

OA21x2_ASAP7_75t_L g1177 ( 
.A1(n_1116),
.A2(n_1103),
.B(n_1092),
.Y(n_1177)
);

AO21x2_ASAP7_75t_L g1178 ( 
.A1(n_1035),
.A2(n_1058),
.B(n_1135),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1097),
.B(n_1091),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1104),
.B(n_1056),
.Y(n_1180)
);

INVx2_ASAP7_75t_SL g1181 ( 
.A(n_1042),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1134),
.Y(n_1182)
);

OA21x2_ASAP7_75t_L g1183 ( 
.A1(n_1109),
.A2(n_1072),
.B(n_1117),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_1028),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1086),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1123),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1145),
.Y(n_1187)
);

AND2x4_ASAP7_75t_L g1188 ( 
.A(n_1027),
.B(n_1138),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1131),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1146),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1043),
.B(n_1014),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1026),
.Y(n_1192)
);

AND2x2_ASAP7_75t_L g1193 ( 
.A(n_1138),
.B(n_1143),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1143),
.B(n_1045),
.Y(n_1194)
);

OR2x2_ASAP7_75t_L g1195 ( 
.A(n_1064),
.B(n_1053),
.Y(n_1195)
);

INVx2_ASAP7_75t_SL g1196 ( 
.A(n_1120),
.Y(n_1196)
);

OR2x6_ASAP7_75t_L g1197 ( 
.A(n_1078),
.B(n_1060),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1026),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1100),
.B(n_1098),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_1126),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1102),
.B(n_1016),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1126),
.Y(n_1202)
);

OA21x2_ASAP7_75t_L g1203 ( 
.A1(n_1108),
.A2(n_1107),
.B(n_1114),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_1028),
.Y(n_1204)
);

NOR2xp33_ASAP7_75t_SL g1205 ( 
.A(n_1022),
.B(n_1093),
.Y(n_1205)
);

OR2x6_ASAP7_75t_L g1206 ( 
.A(n_1060),
.B(n_1089),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1048),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1081),
.B(n_1017),
.Y(n_1208)
);

AND2x4_ASAP7_75t_L g1209 ( 
.A(n_1069),
.B(n_1049),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1018),
.B(n_1057),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1119),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1019),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1112),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1112),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1049),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1087),
.B(n_1038),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1030),
.B(n_1037),
.Y(n_1217)
);

AO21x2_ASAP7_75t_L g1218 ( 
.A1(n_1075),
.A2(n_1111),
.B(n_1052),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1021),
.Y(n_1219)
);

BUFx12f_ASAP7_75t_L g1220 ( 
.A(n_1079),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1050),
.B(n_1047),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1106),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1073),
.B(n_1095),
.Y(n_1223)
);

AND2x2_ASAP7_75t_L g1224 ( 
.A(n_1106),
.B(n_1083),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1094),
.A2(n_1068),
.B(n_1101),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1049),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1088),
.A2(n_1070),
.B(n_1150),
.Y(n_1227)
);

INVx4_ASAP7_75t_L g1228 ( 
.A(n_1088),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1044),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1105),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1065),
.A2(n_1074),
.B(n_1118),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1113),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1088),
.B(n_1034),
.Y(n_1233)
);

OR2x6_ASAP7_75t_L g1234 ( 
.A(n_1040),
.B(n_1046),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_1054),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1059),
.B(n_1077),
.Y(n_1236)
);

OR2x6_ASAP7_75t_L g1237 ( 
.A(n_1029),
.B(n_1115),
.Y(n_1237)
);

INVx4_ASAP7_75t_L g1238 ( 
.A(n_1088),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1076),
.B(n_1083),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1012),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1083),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1061),
.B(n_1036),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1061),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1055),
.B(n_1061),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1066),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1015),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1025),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_1080),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1015),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1080),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1121),
.B(n_1128),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1121),
.B(n_1128),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1121),
.B(n_1128),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1180),
.B(n_1163),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1156),
.Y(n_1255)
);

AND2x2_ASAP7_75t_L g1256 ( 
.A(n_1180),
.B(n_1199),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1199),
.B(n_1224),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1224),
.B(n_1221),
.Y(n_1258)
);

AND2x4_ASAP7_75t_L g1259 ( 
.A(n_1228),
.B(n_1238),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1157),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1158),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1155),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1162),
.B(n_1191),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1160),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1152),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1201),
.B(n_1170),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1161),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1165),
.Y(n_1268)
);

AND2x2_ASAP7_75t_L g1269 ( 
.A(n_1201),
.B(n_1222),
.Y(n_1269)
);

AND2x4_ASAP7_75t_L g1270 ( 
.A(n_1228),
.B(n_1238),
.Y(n_1270)
);

INVxp67_ASAP7_75t_SL g1271 ( 
.A(n_1248),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1222),
.B(n_1219),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1167),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1212),
.B(n_1171),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1182),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1187),
.Y(n_1276)
);

INVxp67_ASAP7_75t_L g1277 ( 
.A(n_1155),
.Y(n_1277)
);

OR2x2_ASAP7_75t_L g1278 ( 
.A(n_1232),
.B(n_1241),
.Y(n_1278)
);

HB1xp67_ASAP7_75t_L g1279 ( 
.A(n_1164),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1250),
.B(n_1166),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_L g1281 ( 
.A1(n_1168),
.A2(n_1233),
.B1(n_1217),
.B2(n_1225),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_L g1282 ( 
.A(n_1195),
.B(n_1153),
.Y(n_1282)
);

HB1xp67_ASAP7_75t_L g1283 ( 
.A(n_1164),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1190),
.Y(n_1284)
);

BUFx8_ASAP7_75t_SL g1285 ( 
.A(n_1220),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1246),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1177),
.Y(n_1287)
);

HB1xp67_ASAP7_75t_L g1288 ( 
.A(n_1172),
.Y(n_1288)
);

HB1xp67_ASAP7_75t_L g1289 ( 
.A(n_1172),
.Y(n_1289)
);

HB1xp67_ASAP7_75t_L g1290 ( 
.A(n_1247),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1251),
.B(n_1252),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1237),
.A2(n_1210),
.B1(n_1239),
.B2(n_1179),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1253),
.B(n_1173),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1241),
.B(n_1203),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1159),
.B(n_1211),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1247),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1237),
.B(n_1249),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1237),
.B(n_1236),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1203),
.B(n_1244),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1173),
.B(n_1208),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1205),
.B(n_1186),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1207),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1227),
.A2(n_1231),
.B1(n_1151),
.B2(n_1186),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1215),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_1215),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1174),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1174),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1229),
.B(n_1242),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1216),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1204),
.Y(n_1310)
);

INVx5_ASAP7_75t_L g1311 ( 
.A(n_1234),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1204),
.Y(n_1312)
);

HB1xp67_ASAP7_75t_L g1313 ( 
.A(n_1175),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1175),
.Y(n_1314)
);

CKINVDCx8_ASAP7_75t_R g1315 ( 
.A(n_1200),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1203),
.B(n_1183),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1184),
.B(n_1213),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1214),
.B(n_1243),
.Y(n_1318)
);

AND2x2_ASAP7_75t_L g1319 ( 
.A(n_1230),
.B(n_1183),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1183),
.B(n_1194),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1257),
.B(n_1151),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1257),
.B(n_1258),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1263),
.B(n_1169),
.Y(n_1323)
);

AOI33xp33_ASAP7_75t_L g1324 ( 
.A1(n_1281),
.A2(n_1169),
.A3(n_1185),
.B1(n_1181),
.B2(n_1196),
.B3(n_1245),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1306),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1258),
.B(n_1176),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1279),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1256),
.B(n_1176),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1287),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1307),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1311),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1271),
.Y(n_1332)
);

BUFx2_ASAP7_75t_SL g1333 ( 
.A(n_1315),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1255),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1260),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1261),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_L g1337 ( 
.A(n_1280),
.B(n_1188),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1264),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1283),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1320),
.B(n_1254),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1299),
.B(n_1154),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1280),
.B(n_1188),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1294),
.B(n_1154),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1267),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1259),
.B(n_1270),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1291),
.B(n_1245),
.Y(n_1346)
);

INVx3_ASAP7_75t_L g1347 ( 
.A(n_1259),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1297),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1300),
.B(n_1188),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1268),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1273),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1288),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1297),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1275),
.Y(n_1354)
);

HB1xp67_ASAP7_75t_L g1355 ( 
.A(n_1289),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1308),
.B(n_1231),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1276),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1269),
.B(n_1178),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1284),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1290),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1286),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1266),
.B(n_1193),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1310),
.Y(n_1363)
);

BUFx2_ASAP7_75t_L g1364 ( 
.A(n_1319),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1312),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1313),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1269),
.B(n_1218),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1314),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1278),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1340),
.B(n_1319),
.Y(n_1370)
);

OR2x2_ASAP7_75t_L g1371 ( 
.A(n_1364),
.B(n_1316),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1325),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1340),
.B(n_1318),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1330),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1321),
.B(n_1318),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1329),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1334),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1327),
.B(n_1274),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1321),
.B(n_1303),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1335),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1336),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1328),
.B(n_1298),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1338),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1328),
.B(n_1298),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1344),
.Y(n_1385)
);

NOR3xp33_ASAP7_75t_L g1386 ( 
.A(n_1324),
.B(n_1274),
.C(n_1301),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1350),
.Y(n_1387)
);

HB1xp67_ASAP7_75t_L g1388 ( 
.A(n_1366),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1339),
.B(n_1309),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1351),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1326),
.B(n_1317),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1354),
.Y(n_1392)
);

INVx2_ASAP7_75t_SL g1393 ( 
.A(n_1368),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1352),
.B(n_1355),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1357),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1360),
.B(n_1266),
.Y(n_1396)
);

NAND2x1p5_ASAP7_75t_L g1397 ( 
.A(n_1331),
.B(n_1311),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1358),
.B(n_1316),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1322),
.B(n_1272),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1322),
.B(n_1323),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1359),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1361),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1348),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1348),
.B(n_1270),
.Y(n_1404)
);

OR2x2_ASAP7_75t_L g1405 ( 
.A(n_1398),
.B(n_1343),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1393),
.B(n_1388),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1371),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1398),
.B(n_1343),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1394),
.B(n_1332),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1377),
.Y(n_1410)
);

INVxp67_ASAP7_75t_SL g1411 ( 
.A(n_1371),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1378),
.B(n_1353),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1400),
.B(n_1346),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1393),
.B(n_1353),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1380),
.Y(n_1415)
);

AND2x2_ASAP7_75t_SL g1416 ( 
.A(n_1386),
.B(n_1324),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1389),
.B(n_1367),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1379),
.B(n_1292),
.C(n_1282),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1382),
.B(n_1367),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_SL g1420 ( 
.A1(n_1396),
.A2(n_1315),
.B1(n_1349),
.B2(n_1365),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1384),
.B(n_1341),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1384),
.B(n_1341),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1370),
.B(n_1356),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1376),
.Y(n_1424)
);

INVx1_ASAP7_75t_SL g1425 ( 
.A(n_1404),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1373),
.B(n_1369),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1370),
.B(n_1356),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1403),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1381),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1410),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1415),
.Y(n_1431)
);

INVxp67_ASAP7_75t_L g1432 ( 
.A(n_1414),
.Y(n_1432)
);

AOI22xp5_ASAP7_75t_L g1433 ( 
.A1(n_1416),
.A2(n_1270),
.B1(n_1379),
.B2(n_1345),
.Y(n_1433)
);

AOI221xp5_ASAP7_75t_L g1434 ( 
.A1(n_1418),
.A2(n_1262),
.B1(n_1277),
.B2(n_1296),
.C(n_1401),
.Y(n_1434)
);

INVxp33_ASAP7_75t_L g1435 ( 
.A(n_1413),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_SL g1436 ( 
.A(n_1416),
.B(n_1345),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1417),
.B(n_1373),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1406),
.A2(n_1333),
.B(n_1198),
.C(n_1403),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1429),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1423),
.B(n_1375),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1420),
.A2(n_1293),
.B(n_1304),
.C(n_1363),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1426),
.A2(n_1342),
.B1(n_1337),
.B2(n_1399),
.Y(n_1442)
);

AOI21xp33_ASAP7_75t_L g1443 ( 
.A1(n_1409),
.A2(n_1385),
.B(n_1383),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1412),
.B(n_1375),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1425),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1424),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1427),
.B(n_1391),
.Y(n_1447)
);

OAI21xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1433),
.A2(n_1192),
.B(n_1397),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1430),
.Y(n_1449)
);

AOI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1436),
.A2(n_1345),
.B1(n_1404),
.B2(n_1347),
.Y(n_1450)
);

OAI221xp5_ASAP7_75t_L g1451 ( 
.A1(n_1434),
.A2(n_1438),
.B1(n_1441),
.B2(n_1432),
.C(n_1443),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1431),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1447),
.B(n_1421),
.Y(n_1453)
);

NAND3xp33_ASAP7_75t_L g1454 ( 
.A(n_1442),
.B(n_1428),
.C(n_1374),
.Y(n_1454)
);

OAI322xp33_ASAP7_75t_L g1455 ( 
.A1(n_1451),
.A2(n_1442),
.A3(n_1439),
.B1(n_1446),
.B2(n_1411),
.C1(n_1407),
.C2(n_1428),
.Y(n_1455)
);

AOI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1448),
.A2(n_1435),
.B(n_1372),
.C(n_1411),
.Y(n_1456)
);

AOI211xp5_ASAP7_75t_L g1457 ( 
.A1(n_1454),
.A2(n_1407),
.B(n_1390),
.C(n_1402),
.Y(n_1457)
);

OAI221xp5_ASAP7_75t_L g1458 ( 
.A1(n_1450),
.A2(n_1452),
.B1(n_1449),
.B2(n_1196),
.C(n_1453),
.Y(n_1458)
);

AOI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1451),
.A2(n_1437),
.B1(n_1444),
.B2(n_1387),
.C(n_1392),
.Y(n_1459)
);

NAND4xp25_ASAP7_75t_L g1460 ( 
.A(n_1459),
.B(n_1240),
.C(n_1362),
.D(n_1265),
.Y(n_1460)
);

AOI211xp5_ASAP7_75t_L g1461 ( 
.A1(n_1455),
.A2(n_1198),
.B(n_1202),
.C(n_1395),
.Y(n_1461)
);

AOI221xp5_ASAP7_75t_L g1462 ( 
.A1(n_1456),
.A2(n_1445),
.B1(n_1265),
.B2(n_1419),
.C(n_1424),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1457),
.B(n_1440),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1458),
.A2(n_1445),
.B1(n_1408),
.B2(n_1405),
.Y(n_1464)
);

OAI211xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1459),
.A2(n_1223),
.B(n_1181),
.C(n_1185),
.Y(n_1465)
);

NAND4xp25_ASAP7_75t_L g1466 ( 
.A(n_1461),
.B(n_1235),
.C(n_1295),
.D(n_1302),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1463),
.B(n_1422),
.Y(n_1467)
);

OAI221xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1462),
.A2(n_1197),
.B1(n_1234),
.B2(n_1206),
.C(n_1235),
.Y(n_1468)
);

NOR3xp33_ASAP7_75t_SL g1469 ( 
.A(n_1468),
.B(n_1460),
.C(n_1465),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1467),
.Y(n_1470)
);

XNOR2xp5_ASAP7_75t_L g1471 ( 
.A(n_1469),
.B(n_1466),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1471),
.B(n_1470),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1472),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1472),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_SL g1475 ( 
.A(n_1473),
.B(n_1220),
.Y(n_1475)
);

AOI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1474),
.A2(n_1464),
.B1(n_1304),
.B2(n_1305),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1475),
.A2(n_1285),
.B(n_1226),
.Y(n_1477)
);

OAI22xp5_ASAP7_75t_L g1478 ( 
.A1(n_1476),
.A2(n_1285),
.B1(n_1305),
.B2(n_1226),
.Y(n_1478)
);

OR2x6_ASAP7_75t_L g1479 ( 
.A(n_1477),
.B(n_1197),
.Y(n_1479)
);

AOI211xp5_ASAP7_75t_L g1480 ( 
.A1(n_1479),
.A2(n_1478),
.B(n_1209),
.C(n_1189),
.Y(n_1480)
);


endmodule