module fake_jpeg_11090_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_38),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_46),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_54),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_1),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_38),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_42),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_52),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_3),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_51),
.B(n_2),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_20),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_41),
.C(n_39),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_47),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_66),
.B(n_67),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_64),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_65),
.A2(n_39),
.B1(n_37),
.B2(n_48),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_7),
.Y(n_80)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_26),
.Y(n_87)
);

AO22x1_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_43),
.B1(n_35),
.B2(n_37),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_75),
.A2(n_7),
.B(n_8),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_62),
.A2(n_43),
.B1(n_4),
.B2(n_5),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_23),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_6),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_80),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_81),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_83),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_66),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_87),
.B(n_89),
.Y(n_93)
);

OA22x2_ASAP7_75t_SL g86 ( 
.A1(n_75),
.A2(n_74),
.B1(n_76),
.B2(n_69),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_86),
.Y(n_95)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_68),
.B(n_8),
.C(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_10),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_33),
.B1(n_19),
.B2(n_21),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_92),
.A2(n_87),
.B(n_85),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_92),
.C(n_90),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_97),
.A2(n_99),
.B(n_85),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_93),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_101),
.C(n_96),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_94),
.B(n_91),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_103),
.Y(n_104)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_86),
.A3(n_88),
.B1(n_28),
.B2(n_30),
.C1(n_18),
.C2(n_31),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_27),
.Y(n_106)
);


endmodule