module fake_aes_1238_n_1431 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_39, n_279, n_303, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_137, n_277, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_241, n_95, n_238, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_210, n_184, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1431);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_39;
input n_279;
input n_303;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_241;
input n_95;
input n_238;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_210;
input n_184;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1431;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_311;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_312;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_314;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_319;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_315;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_327;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_487;
wire n_451;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_310;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_329;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_317;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_323;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_316;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_321;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_313;
wire n_322;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_328;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_326;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1132;
wire n_1389;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_318;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_935;
wire n_910;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_320;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1411;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_325;
wire n_349;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
HB1xp67_ASAP7_75t_L g310 ( .A(n_236), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_66), .Y(n_311) );
CKINVDCx5p33_ASAP7_75t_R g312 ( .A(n_64), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_225), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_294), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_254), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_9), .Y(n_316) );
BUFx3_ASAP7_75t_L g317 ( .A(n_162), .Y(n_317) );
INVxp67_ASAP7_75t_SL g318 ( .A(n_194), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_131), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_88), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_15), .Y(n_321) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_47), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_63), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_189), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_21), .Y(n_325) );
INVxp67_ASAP7_75t_SL g326 ( .A(n_179), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_231), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_98), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_27), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_173), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_214), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_100), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_15), .Y(n_333) );
BUFx10_ASAP7_75t_L g334 ( .A(n_227), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_185), .Y(n_335) );
CKINVDCx16_ASAP7_75t_R g336 ( .A(n_164), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_114), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_70), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_84), .Y(n_339) );
CKINVDCx16_ASAP7_75t_R g340 ( .A(n_14), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_222), .Y(n_341) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_94), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_291), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_58), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_83), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_72), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_43), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_304), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_237), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_252), .Y(n_350) );
BUFx3_ASAP7_75t_L g351 ( .A(n_187), .Y(n_351) );
INVxp33_ASAP7_75t_L g352 ( .A(n_309), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_188), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_279), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_150), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_119), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_308), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_263), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_107), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_75), .Y(n_360) );
INVx2_ASAP7_75t_L g361 ( .A(n_307), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_149), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_82), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_92), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_42), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_77), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_33), .Y(n_367) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_57), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_172), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_264), .Y(n_370) );
HB1xp67_ASAP7_75t_L g371 ( .A(n_277), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_103), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_191), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_155), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_67), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_253), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_306), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_106), .Y(n_378) );
CKINVDCx20_ASAP7_75t_R g379 ( .A(n_176), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_18), .Y(n_380) );
BUFx6f_ASAP7_75t_L g381 ( .A(n_47), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_111), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_40), .Y(n_383) );
INVx2_ASAP7_75t_SL g384 ( .A(n_52), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_302), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_271), .Y(n_386) );
CKINVDCx14_ASAP7_75t_R g387 ( .A(n_174), .Y(n_387) );
CKINVDCx20_ASAP7_75t_R g388 ( .A(n_127), .Y(n_388) );
INVxp67_ASAP7_75t_L g389 ( .A(n_69), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_295), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_257), .Y(n_391) );
INVxp67_ASAP7_75t_L g392 ( .A(n_239), .Y(n_392) );
CKINVDCx11_ASAP7_75t_R g393 ( .A(n_68), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_18), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_1), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_13), .B(n_160), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_126), .Y(n_397) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_283), .Y(n_398) );
BUFx3_ASAP7_75t_L g399 ( .A(n_167), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_68), .Y(n_400) );
CKINVDCx5p33_ASAP7_75t_R g401 ( .A(n_12), .Y(n_401) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_81), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_211), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_73), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_288), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_207), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_224), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_130), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_31), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g410 ( .A(n_244), .Y(n_410) );
CKINVDCx14_ASAP7_75t_R g411 ( .A(n_180), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_274), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_124), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_23), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_161), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_2), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_243), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_204), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_76), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_101), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_200), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_238), .Y(n_422) );
INVxp33_ASAP7_75t_SL g423 ( .A(n_206), .Y(n_423) );
CKINVDCx5p33_ASAP7_75t_R g424 ( .A(n_136), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_190), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_258), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_2), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_299), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_286), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_289), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g431 ( .A(n_297), .Y(n_431) );
INVxp33_ASAP7_75t_SL g432 ( .A(n_245), .Y(n_432) );
BUFx3_ASAP7_75t_L g433 ( .A(n_70), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_249), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_44), .Y(n_435) );
INVxp67_ASAP7_75t_SL g436 ( .A(n_27), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_74), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_133), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_58), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_13), .Y(n_440) );
INVxp33_ASAP7_75t_SL g441 ( .A(n_212), .Y(n_441) );
INVxp67_ASAP7_75t_L g442 ( .A(n_265), .Y(n_442) );
BUFx3_ASAP7_75t_L g443 ( .A(n_113), .Y(n_443) );
CKINVDCx14_ASAP7_75t_R g444 ( .A(n_290), .Y(n_444) );
CKINVDCx16_ASAP7_75t_R g445 ( .A(n_40), .Y(n_445) );
INVxp67_ASAP7_75t_L g446 ( .A(n_115), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_270), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_165), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_141), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_230), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_273), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_73), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_300), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_122), .Y(n_454) );
BUFx6f_ASAP7_75t_L g455 ( .A(n_32), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_117), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_217), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_42), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_137), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_30), .Y(n_460) );
BUFx2_ASAP7_75t_SL g461 ( .A(n_298), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g462 ( .A(n_145), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_281), .Y(n_463) );
CKINVDCx5p33_ASAP7_75t_R g464 ( .A(n_213), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_334), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_338), .B(n_365), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_398), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_398), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_334), .Y(n_469) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_340), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_338), .B(n_0), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_398), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_384), .B(n_3), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_365), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_398), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_402), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_402), .Y(n_477) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_384), .B(n_4), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_395), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_395), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_433), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g483 ( .A(n_336), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_310), .B(n_4), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_433), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_402), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_342), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_319), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_342), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_352), .B(n_5), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_320), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_324), .Y(n_492) );
OAI21x1_ASAP7_75t_L g493 ( .A1(n_313), .A2(n_79), .B(n_78), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_327), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_313), .Y(n_495) );
BUFx6f_ASAP7_75t_L g496 ( .A(n_317), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_328), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_330), .Y(n_498) );
OA21x2_ASAP7_75t_L g499 ( .A1(n_332), .A2(n_85), .B(n_80), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_379), .Y(n_500) );
INVx4_ASAP7_75t_L g501 ( .A(n_471), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_469), .B(n_352), .Y(n_502) );
INVx4_ASAP7_75t_L g503 ( .A(n_471), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_495), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_496), .Y(n_505) );
OR2x2_ASAP7_75t_SL g506 ( .A(n_484), .B(n_445), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_496), .Y(n_507) );
INVx1_ASAP7_75t_SL g508 ( .A(n_483), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_469), .B(n_314), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_496), .Y(n_510) );
INVx3_ASAP7_75t_L g511 ( .A(n_471), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_484), .B(n_311), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_495), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_469), .B(n_315), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_465), .B(n_371), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_495), .Y(n_516) );
INVx3_ASAP7_75t_L g517 ( .A(n_471), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_471), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_467), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_467), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_467), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_490), .A2(n_316), .B1(n_323), .B2(n_321), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_468), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_469), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_468), .Y(n_526) );
INVx3_ASAP7_75t_L g527 ( .A(n_466), .Y(n_527) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_465), .B(n_419), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_465), .B(n_355), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_469), .B(n_312), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_465), .B(n_312), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_496), .Y(n_532) );
OAI21xp5_ASAP7_75t_L g533 ( .A1(n_493), .A2(n_350), .B(n_332), .Y(n_533) );
XNOR2xp5_ASAP7_75t_L g534 ( .A(n_487), .B(n_435), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_468), .Y(n_535) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_489), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_472), .Y(n_537) );
AND2x6_ASAP7_75t_L g538 ( .A(n_490), .B(n_317), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_472), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_488), .B(n_392), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_472), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_475), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_500), .Y(n_543) );
BUFx3_ASAP7_75t_L g544 ( .A(n_496), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_475), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_488), .B(n_383), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_491), .B(n_442), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_502), .B(n_491), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_508), .B(n_466), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_509), .B(n_335), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_509), .B(n_492), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g552 ( .A(n_534), .Y(n_552) );
NAND3xp33_ASAP7_75t_SL g553 ( .A(n_543), .B(n_470), .C(n_386), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_531), .B(n_492), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_527), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_527), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_527), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_509), .B(n_335), .Y(n_558) );
CKINVDCx6p67_ASAP7_75t_R g559 ( .A(n_509), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_514), .B(n_494), .Y(n_560) );
AO22x2_ASAP7_75t_L g561 ( .A1(n_512), .A2(n_470), .B1(n_479), .B2(n_473), .Y(n_561) );
INVx3_ASAP7_75t_L g562 ( .A(n_501), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_518), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_518), .Y(n_564) );
OAI21xp5_ASAP7_75t_L g565 ( .A1(n_533), .A2(n_493), .B(n_499), .Y(n_565) );
AND2x4_ASAP7_75t_L g566 ( .A(n_501), .B(n_466), .Y(n_566) );
NAND3xp33_ASAP7_75t_SL g567 ( .A(n_536), .B(n_386), .C(n_379), .Y(n_567) );
AND2x4_ASAP7_75t_L g568 ( .A(n_501), .B(n_466), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_501), .Y(n_569) );
NOR3xp33_ASAP7_75t_SL g570 ( .A(n_536), .B(n_394), .C(n_383), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_512), .B(n_322), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_530), .B(n_494), .Y(n_572) );
AO22x1_ASAP7_75t_L g573 ( .A1(n_538), .A2(n_432), .B1(n_441), .B2(n_423), .Y(n_573) );
OR2x6_ASAP7_75t_L g574 ( .A(n_546), .B(n_473), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_515), .B(n_497), .Y(n_575) );
NOR2x1p5_ASAP7_75t_L g576 ( .A(n_534), .B(n_394), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_528), .B(n_497), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_525), .B(n_498), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_529), .B(n_498), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_540), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_503), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_547), .B(n_479), .Y(n_582) );
INVx6_ASAP7_75t_L g583 ( .A(n_503), .Y(n_583) );
NAND2xp33_ASAP7_75t_SL g584 ( .A(n_503), .B(n_388), .Y(n_584) );
AND2x4_ASAP7_75t_L g585 ( .A(n_503), .B(n_466), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_511), .B(n_482), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_544), .Y(n_587) );
A2O1A1Ixp33_ASAP7_75t_L g588 ( .A1(n_511), .A2(n_485), .B(n_482), .C(n_493), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_522), .B(n_354), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g590 ( .A1(n_511), .A2(n_435), .B1(n_388), .B2(n_405), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_504), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_504), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_517), .B(n_485), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_513), .Y(n_594) );
OR2x6_ASAP7_75t_L g595 ( .A(n_517), .B(n_375), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_517), .B(n_354), .Y(n_596) );
NAND2x1p5_ASAP7_75t_L g597 ( .A(n_513), .B(n_325), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_516), .Y(n_598) );
BUFx3_ASAP7_75t_L g599 ( .A(n_516), .Y(n_599) );
HB1xp67_ASAP7_75t_SL g600 ( .A(n_538), .Y(n_600) );
INVx4_ASAP7_75t_L g601 ( .A(n_538), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_544), .B(n_329), .Y(n_602) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_506), .B(n_378), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_538), .B(n_405), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_506), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_538), .B(n_378), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_538), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_519), .Y(n_608) );
BUFx3_ASAP7_75t_L g609 ( .A(n_538), .Y(n_609) );
NOR3xp33_ASAP7_75t_SL g610 ( .A(n_519), .B(n_416), .C(n_401), .Y(n_610) );
BUFx8_ASAP7_75t_L g611 ( .A(n_520), .Y(n_611) );
INVx5_ASAP7_75t_L g612 ( .A(n_524), .Y(n_612) );
OR2x6_ASAP7_75t_L g613 ( .A(n_505), .B(n_461), .Y(n_613) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_505), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g615 ( .A1(n_520), .A2(n_389), .B(n_480), .C(n_474), .Y(n_615) );
NAND2xp33_ASAP7_75t_SL g616 ( .A(n_507), .B(n_410), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g617 ( .A1(n_507), .A2(n_499), .B(n_358), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_521), .Y(n_618) );
BUFx6f_ASAP7_75t_L g619 ( .A(n_510), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_510), .B(n_410), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_545), .A2(n_416), .B1(n_401), .B2(n_368), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g622 ( .A1(n_521), .A2(n_367), .B1(n_432), .B2(n_423), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g623 ( .A1(n_532), .A2(n_441), .B1(n_436), .B2(n_411), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_523), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_523), .Y(n_625) );
OR2x2_ASAP7_75t_L g626 ( .A(n_545), .B(n_474), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_526), .A2(n_344), .B1(n_346), .B2(n_333), .Y(n_627) );
NAND3xp33_ASAP7_75t_SL g628 ( .A(n_526), .B(n_413), .C(n_412), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_535), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_535), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g631 ( .A(n_532), .Y(n_631) );
NAND2xp33_ASAP7_75t_R g632 ( .A(n_537), .B(n_499), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_537), .B(n_412), .Y(n_633) );
NOR2xp33_ASAP7_75t_L g634 ( .A(n_539), .B(n_446), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_539), .B(n_413), .Y(n_635) );
AO22x1_ASAP7_75t_L g636 ( .A1(n_542), .A2(n_424), .B1(n_431), .B2(n_421), .Y(n_636) );
BUFx4f_ASAP7_75t_L g637 ( .A(n_559), .Y(n_637) );
INVx3_ASAP7_75t_L g638 ( .A(n_599), .Y(n_638) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_601), .Y(n_639) );
INVx3_ASAP7_75t_L g640 ( .A(n_583), .Y(n_640) );
BUFx2_ASAP7_75t_L g641 ( .A(n_611), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_566), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_583), .Y(n_643) );
OR2x6_ASAP7_75t_L g644 ( .A(n_595), .B(n_347), .Y(n_644) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_595), .Y(n_645) );
INVx2_ASAP7_75t_SL g646 ( .A(n_611), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_580), .B(n_393), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_600), .A2(n_400), .B1(n_404), .B2(n_380), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g649 ( .A(n_605), .B(n_393), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_561), .A2(n_387), .B1(n_444), .B2(n_411), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_575), .B(n_409), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_566), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_574), .B(n_414), .Y(n_653) );
INVx5_ASAP7_75t_L g654 ( .A(n_601), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_574), .B(n_427), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_562), .Y(n_656) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_587), .Y(n_657) );
AOI21xp5_ASAP7_75t_L g658 ( .A1(n_565), .A2(n_499), .B(n_541), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_568), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_571), .B(n_437), .Y(n_660) );
NAND3xp33_ASAP7_75t_L g661 ( .A(n_588), .B(n_496), .C(n_499), .Y(n_661) );
BUFx2_ASAP7_75t_L g662 ( .A(n_549), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_561), .B(n_480), .Y(n_663) );
O2A1O1Ixp5_ASAP7_75t_L g664 ( .A1(n_617), .A2(n_326), .B(n_318), .C(n_396), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_548), .B(n_439), .Y(n_665) );
BUFx2_ASAP7_75t_L g666 ( .A(n_584), .Y(n_666) );
AND2x4_ASAP7_75t_L g667 ( .A(n_568), .B(n_440), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_569), .Y(n_668) );
BUFx4f_ASAP7_75t_L g669 ( .A(n_597), .Y(n_669) );
AND2x4_ASAP7_75t_L g670 ( .A(n_585), .B(n_452), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_585), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_591), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_554), .B(n_458), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_569), .Y(n_674) );
INVx6_ASAP7_75t_L g675 ( .A(n_576), .Y(n_675) );
BUFx3_ASAP7_75t_L g676 ( .A(n_614), .Y(n_676) );
NOR2xp33_ASAP7_75t_SL g677 ( .A(n_609), .B(n_421), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_581), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_572), .A2(n_542), .B(n_541), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_592), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_592), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_560), .B(n_481), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_604), .A2(n_444), .B1(n_387), .B2(n_431), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_594), .Y(n_684) );
INVx2_ASAP7_75t_L g685 ( .A(n_626), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_552), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_604), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_550), .A2(n_457), .B1(n_462), .B2(n_424), .Y(n_688) );
O2A1O1Ixp33_ASAP7_75t_L g689 ( .A1(n_577), .A2(n_481), .B(n_460), .C(n_337), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_555), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_556), .Y(n_691) );
INVx3_ASAP7_75t_L g692 ( .A(n_602), .Y(n_692) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_587), .Y(n_693) );
INVx2_ASAP7_75t_L g694 ( .A(n_625), .Y(n_694) );
AOI21xp5_ASAP7_75t_L g695 ( .A1(n_579), .A2(n_339), .B(n_331), .Y(n_695) );
OAI22xp5_ASAP7_75t_SL g696 ( .A1(n_553), .A2(n_462), .B1(n_464), .B2(n_457), .Y(n_696) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_567), .Y(n_697) );
INVx3_ASAP7_75t_L g698 ( .A(n_598), .Y(n_698) );
BUFx8_ASAP7_75t_L g699 ( .A(n_590), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_557), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_586), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_582), .A2(n_343), .B(n_341), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_563), .A2(n_345), .B1(n_349), .B2(n_348), .Y(n_703) );
O2A1O1Ixp5_ASAP7_75t_L g704 ( .A1(n_573), .A2(n_350), .B(n_361), .C(n_358), .Y(n_704) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_636), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_551), .B(n_464), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_593), .Y(n_707) );
CKINVDCx5p33_ASAP7_75t_R g708 ( .A(n_570), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_564), .A2(n_356), .B(n_353), .Y(n_709) );
OR2x6_ASAP7_75t_L g710 ( .A(n_558), .B(n_381), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_625), .Y(n_711) );
BUFx2_ASAP7_75t_L g712 ( .A(n_613), .Y(n_712) );
O2A1O1Ixp5_ASAP7_75t_L g713 ( .A1(n_603), .A2(n_616), .B(n_620), .C(n_606), .Y(n_713) );
BUFx8_ASAP7_75t_SL g714 ( .A(n_613), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_630), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_589), .B(n_334), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g717 ( .A(n_622), .B(n_373), .Y(n_717) );
BUFx6f_ASAP7_75t_L g718 ( .A(n_587), .Y(n_718) );
OR2x6_ASAP7_75t_L g719 ( .A(n_615), .B(n_381), .Y(n_719) );
AO21x1_ASAP7_75t_L g720 ( .A1(n_632), .A2(n_359), .B(n_357), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_578), .A2(n_360), .B1(n_363), .B2(n_362), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_630), .B(n_364), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_629), .Y(n_723) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_612), .Y(n_724) );
INVx2_ASAP7_75t_SL g725 ( .A(n_621), .Y(n_725) );
BUFx8_ASAP7_75t_SL g726 ( .A(n_633), .Y(n_726) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_623), .B(n_382), .Y(n_727) );
O2A1O1Ixp33_ASAP7_75t_L g728 ( .A1(n_596), .A2(n_369), .B(n_370), .C(n_366), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_608), .Y(n_729) );
BUFx3_ASAP7_75t_L g730 ( .A(n_624), .Y(n_730) );
BUFx3_ASAP7_75t_L g731 ( .A(n_618), .Y(n_731) );
BUFx3_ASAP7_75t_L g732 ( .A(n_631), .Y(n_732) );
INVxp67_ASAP7_75t_SL g733 ( .A(n_635), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g734 ( .A1(n_607), .A2(n_374), .B(n_372), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_610), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_627), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_634), .Y(n_737) );
BUFx3_ASAP7_75t_L g738 ( .A(n_612), .Y(n_738) );
INVx3_ASAP7_75t_L g739 ( .A(n_612), .Y(n_739) );
AND2x4_ASAP7_75t_L g740 ( .A(n_619), .B(n_376), .Y(n_740) );
INVx1_ASAP7_75t_SL g741 ( .A(n_619), .Y(n_741) );
BUFx6f_ASAP7_75t_L g742 ( .A(n_619), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_628), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_566), .Y(n_744) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_611), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_599), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_599), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_559), .A2(n_455), .B1(n_381), .B2(n_385), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_571), .B(n_381), .Y(n_749) );
OAI221xp5_ASAP7_75t_L g750 ( .A1(n_551), .A2(n_430), .B1(n_453), .B2(n_377), .C(n_390), .Y(n_750) );
INVxp67_ASAP7_75t_L g751 ( .A(n_595), .Y(n_751) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_595), .Y(n_752) );
NOR2x1_ASAP7_75t_L g753 ( .A(n_628), .B(n_391), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_559), .A2(n_403), .B1(n_406), .B2(n_397), .Y(n_754) );
AND2x4_ASAP7_75t_L g755 ( .A(n_595), .B(n_407), .Y(n_755) );
INVx4_ASAP7_75t_L g756 ( .A(n_559), .Y(n_756) );
OR2x6_ASAP7_75t_L g757 ( .A(n_595), .B(n_455), .Y(n_757) );
OAI21xp33_ASAP7_75t_L g758 ( .A1(n_575), .A2(n_417), .B(n_415), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_566), .Y(n_759) );
BUFx2_ASAP7_75t_L g760 ( .A(n_559), .Y(n_760) );
O2A1O1Ixp33_ASAP7_75t_L g761 ( .A1(n_577), .A2(n_420), .B(n_422), .C(n_418), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g762 ( .A1(n_561), .A2(n_455), .B1(n_496), .B2(n_428), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g763 ( .A(n_559), .B(n_426), .Y(n_763) );
INVx1_ASAP7_75t_SL g764 ( .A(n_559), .Y(n_764) );
INVx1_ASAP7_75t_SL g765 ( .A(n_559), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_685), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_714), .Y(n_767) );
OAI21x1_ASAP7_75t_L g768 ( .A1(n_658), .A2(n_408), .B(n_361), .Y(n_768) );
OAI21x1_ASAP7_75t_SL g769 ( .A1(n_681), .A2(n_425), .B(n_408), .Y(n_769) );
INVx2_ASAP7_75t_SL g770 ( .A(n_637), .Y(n_770) );
INVx6_ASAP7_75t_L g771 ( .A(n_756), .Y(n_771) );
AO21x2_ASAP7_75t_L g772 ( .A1(n_661), .A2(n_434), .B(n_429), .Y(n_772) );
INVx6_ASAP7_75t_L g773 ( .A(n_756), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_667), .Y(n_774) );
AND2x4_ASAP7_75t_L g775 ( .A(n_757), .B(n_438), .Y(n_775) );
INVx2_ASAP7_75t_SL g776 ( .A(n_637), .Y(n_776) );
OAI21x1_ASAP7_75t_L g777 ( .A1(n_658), .A2(n_448), .B(n_425), .Y(n_777) );
OAI21x1_ASAP7_75t_L g778 ( .A1(n_661), .A2(n_454), .B(n_448), .Y(n_778) );
OAI21x1_ASAP7_75t_L g779 ( .A1(n_664), .A2(n_454), .B(n_449), .Y(n_779) );
OAI21x1_ASAP7_75t_L g780 ( .A1(n_720), .A2(n_450), .B(n_447), .Y(n_780) );
OAI21x1_ASAP7_75t_SL g781 ( .A1(n_694), .A2(n_456), .B(n_451), .Y(n_781) );
OAI21x1_ASAP7_75t_L g782 ( .A1(n_762), .A2(n_463), .B(n_459), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_711), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_644), .B(n_455), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_715), .Y(n_785) );
BUFx10_ASAP7_75t_L g786 ( .A(n_757), .Y(n_786) );
INVx1_ASAP7_75t_SL g787 ( .A(n_644), .Y(n_787) );
BUFx2_ASAP7_75t_L g788 ( .A(n_757), .Y(n_788) );
AO21x2_ASAP7_75t_L g789 ( .A1(n_734), .A2(n_476), .B(n_475), .Y(n_789) );
OAI21x1_ASAP7_75t_L g790 ( .A1(n_734), .A2(n_477), .B(n_476), .Y(n_790) );
BUFx2_ASAP7_75t_L g791 ( .A(n_644), .Y(n_791) );
NAND2x1p5_ASAP7_75t_L g792 ( .A(n_669), .B(n_351), .Y(n_792) );
BUFx2_ASAP7_75t_L g793 ( .A(n_676), .Y(n_793) );
AND2x4_ASAP7_75t_L g794 ( .A(n_723), .B(n_351), .Y(n_794) );
OAI21x1_ASAP7_75t_L g795 ( .A1(n_704), .A2(n_722), .B(n_713), .Y(n_795) );
OAI222xp33_ASAP7_75t_L g796 ( .A1(n_650), .A2(n_399), .B1(n_443), .B2(n_476), .C1(n_477), .C2(n_486), .Y(n_796) );
AOI21xp5_ASAP7_75t_SL g797 ( .A1(n_648), .A2(n_443), .B(n_399), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_736), .A2(n_486), .B1(n_477), .B2(n_478), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_667), .Y(n_799) );
NAND2xp33_ASAP7_75t_SL g800 ( .A(n_705), .B(n_478), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_680), .Y(n_801) );
OA21x2_ASAP7_75t_L g802 ( .A1(n_722), .A2(n_486), .B(n_478), .Y(n_802) );
NAND2x1p5_ASAP7_75t_L g803 ( .A(n_669), .B(n_478), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_670), .Y(n_804) );
OAI21x1_ASAP7_75t_SL g805 ( .A1(n_648), .A2(n_5), .B(n_6), .Y(n_805) );
INVx1_ASAP7_75t_L g806 ( .A(n_670), .Y(n_806) );
AND2x2_ASAP7_75t_L g807 ( .A(n_653), .B(n_6), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_682), .Y(n_808) );
OA21x2_ASAP7_75t_L g809 ( .A1(n_695), .A2(n_478), .B(n_524), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g810 ( .A(n_725), .B(n_7), .Y(n_810) );
O2A1O1Ixp33_ASAP7_75t_L g811 ( .A1(n_761), .A2(n_7), .B(n_8), .C(n_9), .Y(n_811) );
OAI21x1_ASAP7_75t_L g812 ( .A1(n_709), .A2(n_478), .B(n_524), .Y(n_812) );
AO21x2_ASAP7_75t_L g813 ( .A1(n_709), .A2(n_524), .B(n_87), .Y(n_813) );
AO21x2_ASAP7_75t_L g814 ( .A1(n_695), .A2(n_524), .B(n_89), .Y(n_814) );
AOI21xp33_ASAP7_75t_L g815 ( .A1(n_647), .A2(n_8), .B(n_10), .Y(n_815) );
NOR2xp67_ASAP7_75t_L g816 ( .A(n_646), .B(n_10), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_663), .A2(n_11), .B1(n_12), .B2(n_14), .Y(n_817) );
AO21x2_ASAP7_75t_L g818 ( .A1(n_702), .A2(n_90), .B(n_86), .Y(n_818) );
INVx2_ASAP7_75t_SL g819 ( .A(n_641), .Y(n_819) );
CKINVDCx11_ASAP7_75t_R g820 ( .A(n_764), .Y(n_820) );
O2A1O1Ixp33_ASAP7_75t_L g821 ( .A1(n_761), .A2(n_11), .B(n_16), .C(n_17), .Y(n_821) );
OAI21x1_ASAP7_75t_L g822 ( .A1(n_679), .A2(n_93), .B(n_91), .Y(n_822) );
AO21x2_ASAP7_75t_L g823 ( .A1(n_702), .A2(n_96), .B(n_95), .Y(n_823) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_645), .Y(n_824) );
AOI21xp5_ASAP7_75t_L g825 ( .A1(n_733), .A2(n_99), .B(n_97), .Y(n_825) );
BUFx2_ASAP7_75t_L g826 ( .A(n_752), .Y(n_826) );
OAI21x1_ASAP7_75t_L g827 ( .A1(n_679), .A2(n_104), .B(n_102), .Y(n_827) );
BUFx3_ASAP7_75t_L g828 ( .A(n_724), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_737), .B(n_16), .Y(n_829) );
NOR2xp33_ASAP7_75t_SL g830 ( .A(n_745), .B(n_17), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_698), .A2(n_108), .B(n_105), .Y(n_831) );
OAI21x1_ASAP7_75t_L g832 ( .A1(n_698), .A2(n_110), .B(n_109), .Y(n_832) );
OAI21x1_ASAP7_75t_L g833 ( .A1(n_689), .A2(n_116), .B(n_112), .Y(n_833) );
A2O1A1Ixp33_ASAP7_75t_L g834 ( .A1(n_689), .A2(n_19), .B(n_20), .C(n_21), .Y(n_834) );
INVx8_ASAP7_75t_L g835 ( .A(n_724), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_668), .Y(n_836) );
OAI21x1_ASAP7_75t_L g837 ( .A1(n_672), .A2(n_120), .B(n_118), .Y(n_837) );
INVx2_ASAP7_75t_SL g838 ( .A(n_760), .Y(n_838) );
OAI21x1_ASAP7_75t_L g839 ( .A1(n_672), .A2(n_123), .B(n_121), .Y(n_839) );
OAI21xp5_ASAP7_75t_L g840 ( .A1(n_701), .A2(n_128), .B(n_125), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_674), .Y(n_841) );
INVx2_ASAP7_75t_L g842 ( .A(n_684), .Y(n_842) );
NAND2x1p5_ASAP7_75t_L g843 ( .A(n_638), .B(n_692), .Y(n_843) );
INVx1_ASAP7_75t_L g844 ( .A(n_749), .Y(n_844) );
INVx1_ASAP7_75t_L g845 ( .A(n_678), .Y(n_845) );
OR2x2_ASAP7_75t_L g846 ( .A(n_751), .B(n_19), .Y(n_846) );
CKINVDCx20_ASAP7_75t_R g847 ( .A(n_699), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_690), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_653), .B(n_20), .Y(n_849) );
OAI21x1_ASAP7_75t_L g850 ( .A1(n_753), .A2(n_132), .B(n_129), .Y(n_850) );
AND2x2_ASAP7_75t_L g851 ( .A(n_655), .B(n_22), .Y(n_851) );
NOR2xp33_ASAP7_75t_L g852 ( .A(n_687), .B(n_22), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_642), .B(n_23), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g854 ( .A1(n_707), .A2(n_24), .B1(n_25), .B2(n_26), .Y(n_854) );
INVx2_ASAP7_75t_L g855 ( .A(n_729), .Y(n_855) );
OAI21x1_ASAP7_75t_L g856 ( .A1(n_728), .A2(n_135), .B(n_134), .Y(n_856) );
INVx3_ASAP7_75t_L g857 ( .A(n_724), .Y(n_857) );
BUFx2_ASAP7_75t_L g858 ( .A(n_699), .Y(n_858) );
INVx2_ASAP7_75t_L g859 ( .A(n_742), .Y(n_859) );
AND2x4_ASAP7_75t_L g860 ( .A(n_652), .B(n_24), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g861 ( .A(n_659), .B(n_25), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_719), .A2(n_26), .B1(n_28), .B2(n_29), .Y(n_862) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_671), .B(n_28), .Y(n_863) );
INVx1_ASAP7_75t_L g864 ( .A(n_691), .Y(n_864) );
OAI21x1_ASAP7_75t_L g865 ( .A1(n_703), .A2(n_739), .B(n_700), .Y(n_865) );
AO22x2_ASAP7_75t_L g866 ( .A1(n_754), .A2(n_743), .B1(n_755), .B2(n_655), .Y(n_866) );
OAI21x1_ASAP7_75t_SL g867 ( .A1(n_754), .A2(n_29), .B(n_30), .Y(n_867) );
INVx1_ASAP7_75t_L g868 ( .A(n_744), .Y(n_868) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_730), .A2(n_31), .B1(n_32), .B2(n_33), .Y(n_869) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_750), .A2(n_34), .B1(n_35), .B2(n_36), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_759), .Y(n_871) );
OR2x6_ASAP7_75t_L g872 ( .A(n_675), .B(n_34), .Y(n_872) );
OAI21x1_ASAP7_75t_SL g873 ( .A1(n_683), .A2(n_35), .B(n_36), .Y(n_873) );
INVx3_ASAP7_75t_SL g874 ( .A(n_764), .Y(n_874) );
INVx3_ASAP7_75t_L g875 ( .A(n_638), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_731), .Y(n_876) );
INVx3_ASAP7_75t_L g877 ( .A(n_738), .Y(n_877) );
OA21x2_ASAP7_75t_L g878 ( .A1(n_758), .A2(n_192), .B(n_303), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_703), .A2(n_186), .B(n_301), .Y(n_879) );
AND2x4_ASAP7_75t_L g880 ( .A(n_692), .B(n_37), .Y(n_880) );
OAI21xp5_ASAP7_75t_L g881 ( .A1(n_706), .A2(n_184), .B(n_296), .Y(n_881) );
OAI21x1_ASAP7_75t_L g882 ( .A1(n_739), .A2(n_183), .B(n_293), .Y(n_882) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_673), .A2(n_182), .B(n_292), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_765), .Y(n_884) );
OAI21x1_ASAP7_75t_L g885 ( .A1(n_665), .A2(n_181), .B(n_287), .Y(n_885) );
BUFx3_ASAP7_75t_L g886 ( .A(n_657), .Y(n_886) );
OAI21x1_ASAP7_75t_L g887 ( .A1(n_665), .A2(n_178), .B(n_285), .Y(n_887) );
OAI211xp5_ASAP7_75t_SL g888 ( .A1(n_649), .A2(n_37), .B(n_38), .C(n_39), .Y(n_888) );
AO21x2_ASAP7_75t_L g889 ( .A1(n_651), .A2(n_193), .B(n_284), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_706), .B(n_38), .Y(n_890) );
AOI22xp33_ASAP7_75t_SL g891 ( .A1(n_696), .A2(n_39), .B1(n_41), .B2(n_43), .Y(n_891) );
OAI21x1_ASAP7_75t_L g892 ( .A1(n_673), .A2(n_195), .B(n_282), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_717), .B(n_41), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_742), .Y(n_894) );
OAI21x1_ASAP7_75t_SL g895 ( .A1(n_746), .A2(n_44), .B(n_45), .Y(n_895) );
OAI21x1_ASAP7_75t_L g896 ( .A1(n_651), .A2(n_177), .B(n_280), .Y(n_896) );
INVxp67_ASAP7_75t_L g897 ( .A(n_662), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_660), .B(n_45), .Y(n_898) );
OA21x2_ASAP7_75t_L g899 ( .A1(n_740), .A2(n_196), .B(n_278), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_742), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_712), .Y(n_901) );
AO31x2_ASAP7_75t_L g902 ( .A1(n_666), .A2(n_46), .A3(n_48), .B(n_49), .Y(n_902) );
AO21x2_ASAP7_75t_L g903 ( .A1(n_750), .A2(n_175), .B(n_276), .Y(n_903) );
OAI21x1_ASAP7_75t_L g904 ( .A1(n_656), .A2(n_171), .B(n_275), .Y(n_904) );
OAI21x1_ASAP7_75t_L g905 ( .A1(n_747), .A2(n_170), .B(n_272), .Y(n_905) );
NAND2xp5_ASAP7_75t_SL g906 ( .A(n_639), .B(n_138), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g907 ( .A1(n_719), .A2(n_46), .B1(n_48), .B2(n_49), .Y(n_907) );
INVx3_ASAP7_75t_L g908 ( .A(n_639), .Y(n_908) );
OAI222xp33_ASAP7_75t_L g909 ( .A1(n_872), .A2(n_719), .B1(n_710), .B2(n_697), .C1(n_735), .C2(n_765), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g910 ( .A1(n_777), .A2(n_741), .B(n_677), .Y(n_910) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_866), .A2(n_893), .B1(n_755), .B2(n_860), .Y(n_911) );
INVx2_ASAP7_75t_L g912 ( .A(n_801), .Y(n_912) );
BUFx2_ASAP7_75t_L g913 ( .A(n_791), .Y(n_913) );
AOI22xp33_ASAP7_75t_SL g914 ( .A1(n_866), .A2(n_732), .B1(n_675), .B2(n_710), .Y(n_914) );
NAND2xp5_ASAP7_75t_L g915 ( .A(n_808), .B(n_721), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_866), .A2(n_710), .B1(n_763), .B2(n_727), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_801), .Y(n_917) );
OA21x2_ASAP7_75t_L g918 ( .A1(n_778), .A2(n_740), .B(n_741), .Y(n_918) );
AOI21xp5_ASAP7_75t_L g919 ( .A1(n_777), .A2(n_677), .B(n_718), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_766), .B(n_708), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_893), .A2(n_686), .B1(n_716), .B2(n_688), .Y(n_921) );
INVx2_ASAP7_75t_L g922 ( .A(n_783), .Y(n_922) );
OAI221xp5_ASAP7_75t_L g923 ( .A1(n_898), .A2(n_640), .B1(n_643), .B2(n_726), .C(n_654), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_810), .A2(n_748), .B1(n_640), .B2(n_643), .Y(n_924) );
BUFx3_ASAP7_75t_L g925 ( .A(n_874), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g926 ( .A1(n_810), .A2(n_639), .B1(n_654), .B2(n_657), .Y(n_926) );
INVx2_ASAP7_75t_SL g927 ( .A(n_771), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_848), .Y(n_928) );
AO21x2_ASAP7_75t_L g929 ( .A1(n_778), .A2(n_718), .B(n_693), .Y(n_929) );
NAND2xp5_ASAP7_75t_L g930 ( .A(n_774), .B(n_657), .Y(n_930) );
AO22x1_ASAP7_75t_L g931 ( .A1(n_858), .A2(n_654), .B1(n_718), .B2(n_693), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_783), .Y(n_932) );
BUFx2_ASAP7_75t_L g933 ( .A(n_874), .Y(n_933) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_830), .A2(n_654), .B1(n_693), .B2(n_52), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_872), .A2(n_50), .B1(n_51), .B2(n_53), .Y(n_935) );
OAI21xp33_ASAP7_75t_L g936 ( .A1(n_862), .A2(n_50), .B(n_51), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g937 ( .A1(n_860), .A2(n_907), .B1(n_862), .B2(n_788), .Y(n_937) );
NOR2xp33_ASAP7_75t_L g938 ( .A(n_787), .B(n_53), .Y(n_938) );
A2O1A1Ixp33_ASAP7_75t_L g939 ( .A1(n_811), .A2(n_54), .B(n_55), .C(n_56), .Y(n_939) );
OAI21x1_ASAP7_75t_L g940 ( .A1(n_768), .A2(n_201), .B(n_269), .Y(n_940) );
OA21x2_ASAP7_75t_L g941 ( .A1(n_812), .A2(n_199), .B(n_268), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g942 ( .A1(n_860), .A2(n_54), .B1(n_55), .B2(n_56), .Y(n_942) );
AO21x2_ASAP7_75t_L g943 ( .A1(n_772), .A2(n_769), .B(n_780), .Y(n_943) );
OAI21xp5_ASAP7_75t_L g944 ( .A1(n_780), .A2(n_57), .B(n_59), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_775), .A2(n_59), .B1(n_60), .B2(n_61), .Y(n_945) );
INVx2_ASAP7_75t_L g946 ( .A(n_785), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_775), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_947) );
AO21x2_ASAP7_75t_L g948 ( .A1(n_772), .A2(n_205), .B(n_267), .Y(n_948) );
OAI221xp5_ASAP7_75t_L g949 ( .A1(n_815), .A2(n_62), .B1(n_63), .B2(n_64), .C(n_65), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g950 ( .A1(n_870), .A2(n_65), .B1(n_66), .B2(n_67), .C(n_69), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_807), .B(n_71), .Y(n_951) );
OAI21xp33_ASAP7_75t_L g952 ( .A1(n_907), .A2(n_71), .B(n_72), .Y(n_952) );
BUFx4f_ASAP7_75t_SL g953 ( .A(n_767), .Y(n_953) );
OA21x2_ASAP7_75t_L g954 ( .A1(n_812), .A2(n_216), .B(n_139), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_864), .Y(n_955) );
AND2x2_ASAP7_75t_L g956 ( .A(n_849), .B(n_74), .Y(n_956) );
BUFx3_ASAP7_75t_L g957 ( .A(n_820), .Y(n_957) );
NAND3xp33_ASAP7_75t_L g958 ( .A(n_888), .B(n_140), .C(n_142), .Y(n_958) );
AOI22xp33_ASAP7_75t_L g959 ( .A1(n_775), .A2(n_143), .B1(n_144), .B2(n_146), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g960 ( .A1(n_852), .A2(n_147), .B1(n_148), .B2(n_151), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_890), .A2(n_152), .B(n_153), .Y(n_961) );
INVx1_ASAP7_75t_L g962 ( .A(n_845), .Y(n_962) );
INVx2_ASAP7_75t_L g963 ( .A(n_785), .Y(n_963) );
INVx1_ASAP7_75t_SL g964 ( .A(n_820), .Y(n_964) );
AOI21xp5_ASAP7_75t_L g965 ( .A1(n_809), .A2(n_154), .B(n_156), .Y(n_965) );
INVx1_ASAP7_75t_L g966 ( .A(n_868), .Y(n_966) );
A2O1A1Ixp33_ASAP7_75t_L g967 ( .A1(n_821), .A2(n_865), .B(n_834), .C(n_852), .Y(n_967) );
INVx1_ASAP7_75t_L g968 ( .A(n_871), .Y(n_968) );
AOI222xp33_ASAP7_75t_L g969 ( .A1(n_847), .A2(n_157), .B1(n_158), .B2(n_159), .C1(n_163), .C2(n_166), .Y(n_969) );
AOI22xp5_ASAP7_75t_L g970 ( .A1(n_880), .A2(n_168), .B1(n_169), .B2(n_197), .Y(n_970) );
OAI211xp5_ASAP7_75t_SL g971 ( .A1(n_891), .A2(n_305), .B(n_202), .C(n_203), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_799), .B(n_198), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_804), .B(n_266), .Y(n_973) );
INVx1_ASAP7_75t_L g974 ( .A(n_880), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_829), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_975) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_806), .B(n_262), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_880), .Y(n_977) );
NAND2xp5_ASAP7_75t_SL g978 ( .A(n_786), .B(n_215), .Y(n_978) );
AND2x2_ASAP7_75t_L g979 ( .A(n_851), .B(n_218), .Y(n_979) );
A2O1A1Ixp33_ASAP7_75t_L g980 ( .A1(n_865), .A2(n_219), .B(n_220), .C(n_221), .Y(n_980) );
NOR2xp33_ASAP7_75t_L g981 ( .A(n_826), .B(n_223), .Y(n_981) );
NOR2x1p5_ASAP7_75t_L g982 ( .A(n_767), .B(n_226), .Y(n_982) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_844), .A2(n_228), .B1(n_229), .B2(n_232), .Y(n_983) );
OAI211xp5_ASAP7_75t_SL g984 ( .A1(n_846), .A2(n_233), .B(n_234), .C(n_235), .Y(n_984) );
AND2x2_ASAP7_75t_L g985 ( .A(n_884), .B(n_240), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_853), .Y(n_986) );
INVx1_ASAP7_75t_L g987 ( .A(n_861), .Y(n_987) );
OAI21xp5_ASAP7_75t_L g988 ( .A1(n_795), .A2(n_241), .B(n_242), .Y(n_988) );
OAI22xp5_ASAP7_75t_L g989 ( .A1(n_817), .A2(n_246), .B1(n_247), .B2(n_248), .Y(n_989) );
OAI22xp33_ASAP7_75t_L g990 ( .A1(n_872), .A2(n_250), .B1(n_251), .B2(n_255), .Y(n_990) );
O2A1O1Ixp33_ASAP7_75t_SL g991 ( .A1(n_906), .A2(n_256), .B(n_259), .C(n_260), .Y(n_991) );
INVx2_ASAP7_75t_L g992 ( .A(n_836), .Y(n_992) );
OR2x2_ASAP7_75t_L g993 ( .A(n_897), .B(n_261), .Y(n_993) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_784), .A2(n_794), .B1(n_793), .B2(n_819), .Y(n_994) );
OA21x2_ASAP7_75t_L g995 ( .A1(n_892), .A2(n_887), .B(n_885), .Y(n_995) );
INVx3_ASAP7_75t_L g996 ( .A(n_835), .Y(n_996) );
INVx2_ASAP7_75t_SL g997 ( .A(n_771), .Y(n_997) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_867), .A2(n_805), .B1(n_817), .B2(n_873), .Y(n_998) );
A2O1A1Ixp33_ASAP7_75t_L g999 ( .A1(n_834), .A2(n_782), .B(n_833), .C(n_881), .Y(n_999) );
INVx3_ASAP7_75t_L g1000 ( .A(n_835), .Y(n_1000) );
AND2x2_ASAP7_75t_L g1001 ( .A(n_884), .B(n_897), .Y(n_1001) );
NAND2xp5_ASAP7_75t_L g1002 ( .A(n_876), .B(n_824), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1003 ( .A1(n_847), .A2(n_838), .B1(n_824), .B2(n_901), .Y(n_1003) );
NOR2x1_ASAP7_75t_SL g1004 ( .A(n_828), .B(n_886), .Y(n_1004) );
OA21x2_ASAP7_75t_L g1005 ( .A1(n_892), .A2(n_887), .B(n_885), .Y(n_1005) );
A2O1A1Ixp33_ASAP7_75t_L g1006 ( .A1(n_782), .A2(n_833), .B(n_795), .C(n_856), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1007 ( .A1(n_836), .A2(n_841), .B1(n_797), .B2(n_855), .Y(n_1007) );
OAI21xp5_ASAP7_75t_L g1008 ( .A1(n_779), .A2(n_863), .B(n_796), .Y(n_1008) );
INVx3_ASAP7_75t_L g1009 ( .A(n_835), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1010 ( .A(n_794), .B(n_841), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_792), .B(n_794), .Y(n_1011) );
AOI21xp5_ASAP7_75t_L g1012 ( .A1(n_809), .A2(n_779), .B(n_800), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_854), .Y(n_1013) );
A2O1A1Ixp33_ASAP7_75t_L g1014 ( .A1(n_856), .A2(n_879), .B(n_825), .C(n_800), .Y(n_1014) );
AO31x2_ASAP7_75t_L g1015 ( .A1(n_883), .A2(n_900), .A3(n_894), .B(n_859), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1016 ( .A1(n_869), .A2(n_781), .B1(n_895), .B2(n_770), .C(n_776), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_842), .Y(n_1017) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_842), .A2(n_855), .B1(n_803), .B2(n_792), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_843), .B(n_771), .Y(n_1019) );
INVx3_ASAP7_75t_L g1020 ( .A(n_828), .Y(n_1020) );
BUFx3_ASAP7_75t_L g1021 ( .A(n_773), .Y(n_1021) );
AOI22xp33_ASAP7_75t_SL g1022 ( .A1(n_786), .A2(n_903), .B1(n_879), .B2(n_773), .Y(n_1022) );
AOI21xp5_ASAP7_75t_L g1023 ( .A1(n_809), .A2(n_802), .B(n_790), .Y(n_1023) );
OAI22xp33_ASAP7_75t_L g1024 ( .A1(n_816), .A2(n_803), .B1(n_840), .B2(n_899), .Y(n_1024) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_773), .A2(n_843), .B1(n_798), .B2(n_875), .C(n_877), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_877), .B(n_875), .Y(n_1026) );
AND2x2_ASAP7_75t_L g1027 ( .A(n_786), .B(n_857), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_903), .A2(n_823), .B1(n_818), .B2(n_789), .Y(n_1028) );
AND2x4_ASAP7_75t_L g1029 ( .A(n_857), .B(n_908), .Y(n_1029) );
AOI21xp33_ASAP7_75t_L g1030 ( .A1(n_908), .A2(n_789), .B(n_823), .Y(n_1030) );
INVx2_ASAP7_75t_L g1031 ( .A(n_886), .Y(n_1031) );
BUFx10_ASAP7_75t_L g1032 ( .A(n_902), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_902), .B(n_798), .Y(n_1033) );
AND2x4_ASAP7_75t_L g1034 ( .A(n_859), .B(n_900), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1035 ( .A(n_902), .B(n_818), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1036 ( .A(n_902), .B(n_894), .Y(n_1036) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_814), .B(n_790), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1038 ( .A(n_832), .Y(n_1038) );
INVx2_ASAP7_75t_SL g1039 ( .A(n_925), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_928), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_955), .Y(n_1041) );
INVxp67_ASAP7_75t_L g1042 ( .A(n_933), .Y(n_1042) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_1013), .A2(n_899), .B1(n_889), .B2(n_850), .Y(n_1043) );
BUFx3_ASAP7_75t_L g1044 ( .A(n_996), .Y(n_1044) );
INVxp67_ASAP7_75t_L g1045 ( .A(n_1001), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_912), .B(n_850), .Y(n_1046) );
INVx1_ASAP7_75t_L g1047 ( .A(n_962), .Y(n_1047) );
INVx1_ASAP7_75t_L g1048 ( .A(n_966), .Y(n_1048) );
OR2x2_ASAP7_75t_L g1049 ( .A(n_1002), .B(n_889), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_913), .B(n_899), .Y(n_1050) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_917), .B(n_896), .Y(n_1051) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_996), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_968), .Y(n_1053) );
OR2x2_ASAP7_75t_L g1054 ( .A(n_1010), .B(n_896), .Y(n_1054) );
INVxp67_ASAP7_75t_SL g1055 ( .A(n_922), .Y(n_1055) );
OR2x2_ASAP7_75t_L g1056 ( .A(n_951), .B(n_832), .Y(n_1056) );
INVxp67_ASAP7_75t_L g1057 ( .A(n_920), .Y(n_1057) );
AOI22xp33_ASAP7_75t_SL g1058 ( .A1(n_937), .A2(n_878), .B1(n_882), .B2(n_813), .Y(n_1058) );
INVxp67_ASAP7_75t_SL g1059 ( .A(n_932), .Y(n_1059) );
INVx2_ASAP7_75t_L g1060 ( .A(n_946), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_1017), .B(n_882), .Y(n_1061) );
INVx1_ASAP7_75t_L g1062 ( .A(n_963), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_992), .Y(n_1063) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_986), .B(n_822), .Y(n_1064) );
INVx1_ASAP7_75t_L g1065 ( .A(n_956), .Y(n_1065) );
INVx3_ASAP7_75t_L g1066 ( .A(n_1000), .Y(n_1066) );
BUFx6f_ASAP7_75t_L g1067 ( .A(n_1029), .Y(n_1067) );
INVx1_ASAP7_75t_L g1068 ( .A(n_993), .Y(n_1068) );
BUFx3_ASAP7_75t_L g1069 ( .A(n_1000), .Y(n_1069) );
AND2x4_ASAP7_75t_L g1070 ( .A(n_974), .B(n_831), .Y(n_1070) );
INVx1_ASAP7_75t_L g1071 ( .A(n_977), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_915), .B(n_827), .Y(n_1072) );
BUFx6f_ASAP7_75t_L g1073 ( .A(n_1029), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_935), .Y(n_1074) );
BUFx3_ASAP7_75t_L g1075 ( .A(n_1009), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1076 ( .A(n_987), .B(n_878), .Y(n_1076) );
OR2x6_ASAP7_75t_L g1077 ( .A(n_982), .B(n_837), .Y(n_1077) );
INVx1_ASAP7_75t_L g1078 ( .A(n_935), .Y(n_1078) );
OR2x2_ASAP7_75t_L g1079 ( .A(n_1011), .B(n_839), .Y(n_1079) );
OR2x6_ASAP7_75t_L g1080 ( .A(n_931), .B(n_905), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1026), .Y(n_1081) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_911), .B(n_878), .Y(n_1082) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_1009), .Y(n_1083) );
INVx2_ASAP7_75t_L g1084 ( .A(n_941), .Y(n_1084) );
INVx1_ASAP7_75t_L g1085 ( .A(n_930), .Y(n_1085) );
AND2x4_ASAP7_75t_L g1086 ( .A(n_1034), .B(n_904), .Y(n_1086) );
OAI33xp33_ASAP7_75t_L g1087 ( .A1(n_990), .A2(n_952), .A3(n_936), .B1(n_1018), .B2(n_1024), .B3(n_1036), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_944), .Y(n_1088) );
INVx2_ASAP7_75t_L g1089 ( .A(n_941), .Y(n_1089) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1007), .Y(n_1090) );
INVx2_ASAP7_75t_L g1091 ( .A(n_954), .Y(n_1091) );
AND2x2_ASAP7_75t_L g1092 ( .A(n_994), .B(n_1019), .Y(n_1092) );
AND2x2_ASAP7_75t_L g1093 ( .A(n_938), .B(n_1021), .Y(n_1093) );
INVx2_ASAP7_75t_L g1094 ( .A(n_954), .Y(n_1094) );
NAND2xp5_ASAP7_75t_L g1095 ( .A(n_921), .B(n_1003), .Y(n_1095) );
OAI22xp33_ASAP7_75t_L g1096 ( .A1(n_990), .A2(n_950), .B1(n_949), .B2(n_1025), .Y(n_1096) );
OR2x2_ASAP7_75t_L g1097 ( .A(n_927), .B(n_997), .Y(n_1097) );
BUFx2_ASAP7_75t_L g1098 ( .A(n_957), .Y(n_1098) );
AND2x2_ASAP7_75t_L g1099 ( .A(n_1035), .B(n_985), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_914), .B(n_1020), .Y(n_1100) );
INVx5_ASAP7_75t_L g1101 ( .A(n_1020), .Y(n_1101) );
INVx2_ASAP7_75t_L g1102 ( .A(n_929), .Y(n_1102) );
AND2x4_ASAP7_75t_SL g1103 ( .A(n_1027), .B(n_979), .Y(n_1103) );
INVx1_ASAP7_75t_L g1104 ( .A(n_1032), .Y(n_1104) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_914), .B(n_916), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1106 ( .A(n_981), .B(n_964), .Y(n_1106) );
OR2x2_ASAP7_75t_L g1107 ( .A(n_916), .B(n_923), .Y(n_1107) );
BUFx2_ASAP7_75t_L g1108 ( .A(n_953), .Y(n_1108) );
AND2x4_ASAP7_75t_L g1109 ( .A(n_1034), .B(n_1031), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1032), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_950), .Y(n_1111) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_998), .B(n_942), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_972), .Y(n_1113) );
HB1xp67_ASAP7_75t_L g1114 ( .A(n_1038), .Y(n_1114) );
OR2x2_ASAP7_75t_L g1115 ( .A(n_945), .B(n_947), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_973), .Y(n_1116) );
INVx1_ASAP7_75t_L g1117 ( .A(n_976), .Y(n_1117) );
AND2x2_ASAP7_75t_L g1118 ( .A(n_998), .B(n_967), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_969), .B(n_934), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_939), .B(n_1016), .Y(n_1120) );
BUFx6f_ASAP7_75t_L g1121 ( .A(n_918), .Y(n_1121) );
AND2x4_ASAP7_75t_L g1122 ( .A(n_1004), .B(n_1015), .Y(n_1122) );
INVx2_ASAP7_75t_L g1123 ( .A(n_929), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_934), .B(n_1033), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_943), .B(n_1022), .Y(n_1125) );
INVx4_ASAP7_75t_L g1126 ( .A(n_953), .Y(n_1126) );
INVx1_ASAP7_75t_L g1127 ( .A(n_970), .Y(n_1127) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1016), .B(n_924), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1129 ( .A(n_943), .B(n_1022), .Y(n_1129) );
INVx2_ASAP7_75t_L g1130 ( .A(n_1015), .Y(n_1130) );
NAND4xp25_ASAP7_75t_L g1131 ( .A(n_1028), .B(n_924), .C(n_960), .D(n_999), .Y(n_1131) );
AOI22xp33_ASAP7_75t_SL g1132 ( .A1(n_989), .A2(n_909), .B1(n_958), .B2(n_1038), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1133 ( .A(n_926), .B(n_960), .Y(n_1133) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_926), .B(n_1028), .Y(n_1134) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1008), .B(n_978), .Y(n_1135) );
INVx3_ASAP7_75t_L g1136 ( .A(n_1015), .Y(n_1136) );
AND2x4_ASAP7_75t_L g1137 ( .A(n_1015), .B(n_980), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_948), .B(n_983), .Y(n_1138) );
NAND2xp5_ASAP7_75t_L g1139 ( .A(n_961), .B(n_975), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_1023), .Y(n_1140) );
BUFx2_ASAP7_75t_L g1141 ( .A(n_940), .Y(n_1141) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_971), .A2(n_984), .B1(n_1030), .B2(n_983), .Y(n_1142) );
OR2x2_ASAP7_75t_L g1143 ( .A(n_1023), .B(n_909), .Y(n_1143) );
HB1xp67_ASAP7_75t_L g1144 ( .A(n_1045), .Y(n_1144) );
BUFx2_ASAP7_75t_SL g1145 ( .A(n_1101), .Y(n_1145) );
INVx2_ASAP7_75t_SL g1146 ( .A(n_1101), .Y(n_1146) );
BUFx2_ASAP7_75t_L g1147 ( .A(n_1122), .Y(n_1147) );
OAI221xp5_ASAP7_75t_L g1148 ( .A1(n_1095), .A2(n_971), .B1(n_984), .B2(n_975), .C(n_1014), .Y(n_1148) );
AND2x2_ASAP7_75t_L g1149 ( .A(n_1118), .B(n_995), .Y(n_1149) );
AOI33xp33_ASAP7_75t_L g1150 ( .A1(n_1065), .A2(n_959), .A3(n_991), .B1(n_948), .B2(n_1005), .B3(n_995), .Y(n_1150) );
OAI22xp5_ASAP7_75t_L g1151 ( .A1(n_1119), .A2(n_965), .B1(n_1006), .B2(n_1012), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1152 ( .A(n_1118), .B(n_1005), .Y(n_1152) );
INVxp67_ASAP7_75t_SL g1153 ( .A(n_1055), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1099), .B(n_918), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1155 ( .A(n_1122), .Y(n_1155) );
INVx2_ASAP7_75t_SL g1156 ( .A(n_1101), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1099), .B(n_988), .Y(n_1157) );
HB1xp67_ASAP7_75t_L g1158 ( .A(n_1059), .Y(n_1158) );
NAND2xp5_ASAP7_75t_L g1159 ( .A(n_1040), .B(n_961), .Y(n_1159) );
BUFx2_ASAP7_75t_L g1160 ( .A(n_1122), .Y(n_1160) );
INVx2_ASAP7_75t_SL g1161 ( .A(n_1101), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1162 ( .A(n_1057), .B(n_965), .Y(n_1162) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1041), .B(n_910), .Y(n_1163) );
AOI33xp33_ASAP7_75t_L g1164 ( .A1(n_1119), .A2(n_919), .A3(n_1037), .B1(n_1053), .B2(n_1048), .B3(n_1081), .Y(n_1164) );
BUFx2_ASAP7_75t_L g1165 ( .A(n_1114), .Y(n_1165) );
OR2x6_ASAP7_75t_L g1166 ( .A(n_1077), .B(n_1100), .Y(n_1166) );
OAI221xp5_ASAP7_75t_L g1167 ( .A1(n_1111), .A2(n_1107), .B1(n_1042), .B2(n_1120), .C(n_1128), .Y(n_1167) );
BUFx3_ASAP7_75t_L g1168 ( .A(n_1044), .Y(n_1168) );
INVx5_ASAP7_75t_L g1169 ( .A(n_1077), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1170 ( .A(n_1124), .B(n_1060), .Y(n_1170) );
OAI21xp33_ASAP7_75t_L g1171 ( .A1(n_1105), .A2(n_1143), .B(n_1131), .Y(n_1171) );
INVx2_ASAP7_75t_L g1172 ( .A(n_1130), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1124), .B(n_1060), .Y(n_1173) );
OAI31xp33_ASAP7_75t_L g1174 ( .A1(n_1096), .A2(n_1112), .A3(n_1074), .B(n_1078), .Y(n_1174) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1140), .Y(n_1175) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1092), .B(n_1100), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1140), .Y(n_1177) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1063), .B(n_1134), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1063), .B(n_1134), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1114), .Y(n_1180) );
NOR2xp33_ASAP7_75t_L g1181 ( .A(n_1098), .B(n_1126), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1125), .B(n_1129), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1183 ( .A(n_1104), .B(n_1110), .Y(n_1183) );
BUFx3_ASAP7_75t_L g1184 ( .A(n_1044), .Y(n_1184) );
INVxp67_ASAP7_75t_R g1185 ( .A(n_1093), .Y(n_1185) );
NAND2x1_ASAP7_75t_L g1186 ( .A(n_1077), .B(n_1080), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1049), .B(n_1112), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1061), .Y(n_1188) );
INVx2_ASAP7_75t_L g1189 ( .A(n_1136), .Y(n_1189) );
INVx4_ASAP7_75t_L g1190 ( .A(n_1103), .Y(n_1190) );
INVx5_ASAP7_75t_L g1191 ( .A(n_1080), .Y(n_1191) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1061), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1125), .B(n_1129), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1062), .B(n_1047), .Y(n_1194) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1136), .Y(n_1195) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_1127), .A2(n_1115), .B1(n_1096), .B2(n_1087), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1076), .Y(n_1197) );
OAI31xp33_ASAP7_75t_L g1198 ( .A1(n_1103), .A2(n_1068), .A3(n_1133), .B(n_1113), .Y(n_1198) );
HB1xp67_ASAP7_75t_L g1199 ( .A(n_1039), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1200 ( .A(n_1082), .B(n_1076), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1082), .B(n_1071), .Y(n_1201) );
OAI33xp33_ASAP7_75t_L g1202 ( .A1(n_1097), .A2(n_1050), .A3(n_1088), .B1(n_1056), .B2(n_1085), .B3(n_1117), .Y(n_1202) );
HB1xp67_ASAP7_75t_L g1203 ( .A(n_1039), .Y(n_1203) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1072), .B(n_1054), .Y(n_1204) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1136), .Y(n_1205) );
INVxp67_ASAP7_75t_SL g1206 ( .A(n_1051), .Y(n_1206) );
AOI22xp5_ASAP7_75t_L g1207 ( .A1(n_1106), .A2(n_1116), .B1(n_1126), .B2(n_1139), .Y(n_1207) );
INVxp67_ASAP7_75t_SL g1208 ( .A(n_1051), .Y(n_1208) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1064), .B(n_1046), .Y(n_1209) );
OR2x2_ASAP7_75t_L g1210 ( .A(n_1109), .B(n_1079), .Y(n_1210) );
INVxp67_ASAP7_75t_SL g1211 ( .A(n_1046), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1064), .B(n_1109), .Y(n_1212) );
NAND2xp5_ASAP7_75t_SL g1213 ( .A(n_1052), .B(n_1083), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1214 ( .A(n_1109), .B(n_1138), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1138), .B(n_1070), .Y(n_1215) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1102), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1069), .B(n_1075), .Y(n_1217) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1069), .B(n_1075), .Y(n_1218) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1090), .B(n_1123), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1070), .B(n_1137), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1123), .Y(n_1221) );
HB1xp67_ASAP7_75t_L g1222 ( .A(n_1158), .Y(n_1222) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1187), .B(n_1090), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1174), .B(n_1067), .Y(n_1224) );
INVx2_ASAP7_75t_SL g1225 ( .A(n_1147), .Y(n_1225) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1187), .B(n_1121), .Y(n_1226) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1194), .Y(n_1227) );
AND2x4_ASAP7_75t_SL g1228 ( .A(n_1190), .B(n_1126), .Y(n_1228) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1194), .Y(n_1229) );
AOI21xp5_ASAP7_75t_L g1230 ( .A1(n_1153), .A2(n_1142), .B(n_1080), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1182), .B(n_1137), .Y(n_1231) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1144), .B(n_1067), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1196), .B(n_1067), .Y(n_1233) );
INVx2_ASAP7_75t_L g1234 ( .A(n_1172), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_1182), .B(n_1137), .Y(n_1235) );
NOR2x1_ASAP7_75t_L g1236 ( .A(n_1190), .B(n_1108), .Y(n_1236) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1199), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1238 ( .A(n_1181), .B(n_1066), .Y(n_1238) );
NOR3xp33_ASAP7_75t_SL g1239 ( .A(n_1167), .B(n_1135), .C(n_1132), .Y(n_1239) );
INVxp67_ASAP7_75t_L g1240 ( .A(n_1203), .Y(n_1240) );
NOR3xp33_ASAP7_75t_SL g1241 ( .A(n_1171), .B(n_1067), .C(n_1073), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1193), .B(n_1121), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1193), .B(n_1121), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1244 ( .A(n_1209), .B(n_1121), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1209), .B(n_1070), .Y(n_1245) );
INVx1_ASAP7_75t_L g1246 ( .A(n_1180), .Y(n_1246) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1214), .B(n_1086), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1248 ( .A(n_1214), .B(n_1086), .Y(n_1248) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_1162), .A2(n_1073), .B1(n_1086), .B2(n_1066), .Y(n_1249) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1176), .B(n_1089), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1201), .B(n_1084), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1212), .B(n_1091), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1170), .B(n_1073), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1212), .B(n_1094), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1200), .B(n_1043), .Y(n_1255) );
NAND2xp5_ASAP7_75t_SL g1256 ( .A(n_1190), .B(n_1073), .Y(n_1256) );
NOR3xp33_ASAP7_75t_SL g1257 ( .A(n_1198), .B(n_1148), .C(n_1202), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1200), .B(n_1043), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1215), .B(n_1058), .Y(n_1259) );
INVx1_ASAP7_75t_L g1260 ( .A(n_1180), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1215), .B(n_1141), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1149), .B(n_1142), .Y(n_1262) );
INVx2_ASAP7_75t_SL g1263 ( .A(n_1147), .Y(n_1263) );
HB1xp67_ASAP7_75t_L g1264 ( .A(n_1165), .Y(n_1264) );
BUFx2_ASAP7_75t_L g1265 ( .A(n_1155), .Y(n_1265) );
NOR2x1_ASAP7_75t_L g1266 ( .A(n_1145), .B(n_1066), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1183), .Y(n_1267) );
BUFx2_ASAP7_75t_L g1268 ( .A(n_1155), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1269 ( .A(n_1170), .B(n_1173), .Y(n_1269) );
OR2x2_ASAP7_75t_L g1270 ( .A(n_1176), .B(n_1173), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1183), .Y(n_1271) );
OR2x2_ASAP7_75t_L g1272 ( .A(n_1178), .B(n_1179), .Y(n_1272) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_1169), .B(n_1160), .Y(n_1273) );
OR2x2_ASAP7_75t_L g1274 ( .A(n_1178), .B(n_1179), .Y(n_1274) );
OR2x2_ASAP7_75t_L g1275 ( .A(n_1160), .B(n_1192), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1276 ( .A(n_1188), .B(n_1192), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1277 ( .A(n_1188), .B(n_1204), .Y(n_1277) );
AOI22xp33_ASAP7_75t_SL g1278 ( .A1(n_1145), .A2(n_1169), .B1(n_1166), .B2(n_1168), .Y(n_1278) );
NOR2xp33_ASAP7_75t_L g1279 ( .A(n_1207), .B(n_1217), .Y(n_1279) );
NOR2x1_ASAP7_75t_L g1280 ( .A(n_1168), .B(n_1184), .Y(n_1280) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1204), .B(n_1165), .Y(n_1281) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1149), .B(n_1152), .Y(n_1282) );
AOI21xp33_ASAP7_75t_L g1283 ( .A1(n_1159), .A2(n_1146), .B(n_1156), .Y(n_1283) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1210), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1152), .B(n_1154), .Y(n_1285) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1222), .Y(n_1286) );
INVx1_ASAP7_75t_SL g1287 ( .A(n_1228), .Y(n_1287) );
AND2x4_ASAP7_75t_SL g1288 ( .A(n_1241), .B(n_1166), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1285), .B(n_1154), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1285), .B(n_1220), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1282), .B(n_1220), .Y(n_1291) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1276), .Y(n_1292) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1270), .B(n_1177), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1267), .B(n_1164), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1282), .B(n_1166), .Y(n_1295) );
NAND2xp5_ASAP7_75t_SL g1296 ( .A(n_1280), .B(n_1169), .Y(n_1296) );
NOR2xp33_ASAP7_75t_L g1297 ( .A(n_1240), .B(n_1184), .Y(n_1297) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1277), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1242), .B(n_1166), .Y(n_1299) );
INVx2_ASAP7_75t_L g1300 ( .A(n_1234), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1242), .B(n_1197), .Y(n_1301) );
OR2x2_ASAP7_75t_L g1302 ( .A(n_1270), .B(n_1175), .Y(n_1302) );
OAI21xp5_ASAP7_75t_L g1303 ( .A1(n_1257), .A2(n_1146), .B(n_1161), .Y(n_1303) );
AND2x4_ASAP7_75t_L g1304 ( .A(n_1273), .B(n_1169), .Y(n_1304) );
OR2x2_ASAP7_75t_L g1305 ( .A(n_1272), .B(n_1175), .Y(n_1305) );
INVx1_ASAP7_75t_SL g1306 ( .A(n_1228), .Y(n_1306) );
NOR2xp33_ASAP7_75t_L g1307 ( .A(n_1227), .B(n_1218), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1271), .B(n_1197), .Y(n_1308) );
HB1xp67_ASAP7_75t_L g1309 ( .A(n_1264), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1277), .Y(n_1310) );
OR2x2_ASAP7_75t_L g1311 ( .A(n_1272), .B(n_1177), .Y(n_1311) );
INVx1_ASAP7_75t_L g1312 ( .A(n_1281), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1281), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1314 ( .A1(n_1279), .A2(n_1157), .B1(n_1151), .B2(n_1210), .Y(n_1314) );
OR2x2_ASAP7_75t_L g1315 ( .A(n_1274), .B(n_1163), .Y(n_1315) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1229), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1246), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1243), .B(n_1211), .Y(n_1318) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1260), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1237), .Y(n_1320) );
INVx2_ASAP7_75t_L g1321 ( .A(n_1234), .Y(n_1321) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1284), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1323 ( .A(n_1274), .B(n_1223), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1324 ( .A(n_1243), .B(n_1208), .Y(n_1324) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1275), .Y(n_1325) );
NAND2xp5_ASAP7_75t_L g1326 ( .A(n_1269), .B(n_1157), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1275), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1223), .B(n_1219), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1262), .B(n_1206), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1231), .B(n_1205), .Y(n_1330) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1250), .Y(n_1331) );
AOI21xp5_ASAP7_75t_L g1332 ( .A1(n_1296), .A2(n_1186), .B(n_1266), .Y(n_1332) );
INVx2_ASAP7_75t_SL g1333 ( .A(n_1287), .Y(n_1333) );
OA21x2_ASAP7_75t_L g1334 ( .A1(n_1294), .A2(n_1230), .B(n_1283), .Y(n_1334) );
INVx1_ASAP7_75t_SL g1335 ( .A(n_1306), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1312), .B(n_1262), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1337 ( .A(n_1290), .B(n_1245), .Y(n_1337) );
AOI22xp5_ASAP7_75t_L g1338 ( .A1(n_1314), .A2(n_1239), .B1(n_1224), .B2(n_1259), .Y(n_1338) );
AOI21xp5_ASAP7_75t_L g1339 ( .A1(n_1296), .A2(n_1186), .B(n_1256), .Y(n_1339) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1323), .Y(n_1340) );
OAI31xp33_ASAP7_75t_L g1341 ( .A1(n_1288), .A2(n_1268), .A3(n_1265), .B(n_1238), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1323), .Y(n_1342) );
INVx1_ASAP7_75t_L g1343 ( .A(n_1305), .Y(n_1343) );
INVx2_ASAP7_75t_SL g1344 ( .A(n_1304), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1313), .B(n_1255), .Y(n_1345) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1289), .B(n_1244), .Y(n_1346) );
INVxp67_ASAP7_75t_SL g1347 ( .A(n_1309), .Y(n_1347) );
INVxp67_ASAP7_75t_L g1348 ( .A(n_1297), .Y(n_1348) );
OAI22xp5_ASAP7_75t_L g1349 ( .A1(n_1303), .A2(n_1236), .B1(n_1185), .B2(n_1278), .Y(n_1349) );
INVxp67_ASAP7_75t_L g1350 ( .A(n_1286), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1305), .Y(n_1351) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1311), .Y(n_1352) );
OAI322xp33_ASAP7_75t_L g1353 ( .A1(n_1315), .A2(n_1250), .A3(n_1226), .B1(n_1232), .B2(n_1233), .C1(n_1263), .C2(n_1225), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1289), .B(n_1244), .Y(n_1354) );
XOR2xp5_ASAP7_75t_L g1355 ( .A(n_1315), .B(n_1253), .Y(n_1355) );
AOI22xp5_ASAP7_75t_L g1356 ( .A1(n_1307), .A2(n_1259), .B1(n_1258), .B2(n_1255), .Y(n_1356) );
NAND2xp5_ASAP7_75t_SL g1357 ( .A(n_1288), .B(n_1169), .Y(n_1357) );
NOR2xp33_ASAP7_75t_L g1358 ( .A(n_1320), .B(n_1213), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1292), .B(n_1258), .Y(n_1359) );
OAI21xp5_ASAP7_75t_L g1360 ( .A1(n_1311), .A2(n_1161), .B(n_1156), .Y(n_1360) );
NOR2xp33_ASAP7_75t_L g1361 ( .A(n_1316), .B(n_1231), .Y(n_1361) );
INVx2_ASAP7_75t_L g1362 ( .A(n_1300), .Y(n_1362) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1340), .B(n_1328), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1356), .B(n_1292), .Y(n_1364) );
INVx1_ASAP7_75t_L g1365 ( .A(n_1362), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1346), .B(n_1290), .Y(n_1366) );
A2O1A1Ixp33_ASAP7_75t_L g1367 ( .A1(n_1341), .A2(n_1295), .B(n_1265), .C(n_1268), .Y(n_1367) );
NOR2xp33_ASAP7_75t_L g1368 ( .A(n_1348), .B(n_1310), .Y(n_1368) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1342), .Y(n_1369) );
HB1xp67_ASAP7_75t_L g1370 ( .A(n_1347), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_1343), .B(n_1301), .Y(n_1371) );
AOI22xp5_ASAP7_75t_L g1372 ( .A1(n_1338), .A2(n_1295), .B1(n_1298), .B2(n_1329), .Y(n_1372) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1362), .Y(n_1373) );
INVxp67_ASAP7_75t_L g1374 ( .A(n_1333), .Y(n_1374) );
INVx2_ASAP7_75t_L g1375 ( .A(n_1351), .Y(n_1375) );
NAND2xp5_ASAP7_75t_SL g1376 ( .A(n_1349), .B(n_1304), .Y(n_1376) );
O2A1O1Ixp33_ASAP7_75t_L g1377 ( .A1(n_1350), .A2(n_1333), .B(n_1335), .C(n_1334), .Y(n_1377) );
OAI21xp33_ASAP7_75t_L g1378 ( .A1(n_1359), .A2(n_1291), .B(n_1326), .Y(n_1378) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1352), .Y(n_1379) );
INVxp33_ASAP7_75t_L g1380 ( .A(n_1357), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1336), .Y(n_1381) );
INVxp67_ASAP7_75t_L g1382 ( .A(n_1358), .Y(n_1382) );
INVx2_ASAP7_75t_L g1383 ( .A(n_1346), .Y(n_1383) );
OAI311xp33_ASAP7_75t_L g1384 ( .A1(n_1377), .A2(n_1360), .A3(n_1249), .B1(n_1328), .C1(n_1302), .Y(n_1384) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1370), .Y(n_1385) );
AOI322xp5_ASAP7_75t_L g1386 ( .A1(n_1376), .A2(n_1361), .A3(n_1345), .B1(n_1354), .B2(n_1337), .C1(n_1291), .C2(n_1344), .Y(n_1386) );
A2O1A1Ixp33_ASAP7_75t_SL g1387 ( .A1(n_1374), .A2(n_1358), .B(n_1332), .C(n_1339), .Y(n_1387) );
INVx3_ASAP7_75t_SL g1388 ( .A(n_1363), .Y(n_1388) );
AOI21xp5_ASAP7_75t_L g1389 ( .A1(n_1367), .A2(n_1357), .B(n_1353), .Y(n_1389) );
AOI22xp5_ASAP7_75t_L g1390 ( .A1(n_1372), .A2(n_1334), .B1(n_1361), .B2(n_1344), .Y(n_1390) );
AOI211xp5_ASAP7_75t_L g1391 ( .A1(n_1380), .A2(n_1185), .B(n_1293), .C(n_1302), .Y(n_1391) );
OAI32xp33_ASAP7_75t_L g1392 ( .A1(n_1380), .A2(n_1355), .A3(n_1293), .B1(n_1354), .B2(n_1325), .Y(n_1392) );
O2A1O1Ixp33_ASAP7_75t_L g1393 ( .A1(n_1382), .A2(n_1334), .B(n_1322), .C(n_1319), .Y(n_1393) );
AOI221xp5_ASAP7_75t_L g1394 ( .A1(n_1368), .A2(n_1327), .B1(n_1331), .B2(n_1308), .C(n_1317), .Y(n_1394) );
AOI21xp33_ASAP7_75t_SL g1395 ( .A1(n_1364), .A2(n_1225), .B(n_1263), .Y(n_1395) );
AOI22xp5_ASAP7_75t_L g1396 ( .A1(n_1381), .A2(n_1331), .B1(n_1301), .B2(n_1330), .Y(n_1396) );
AOI221xp5_ASAP7_75t_L g1397 ( .A1(n_1378), .A2(n_1235), .B1(n_1330), .B2(n_1324), .C(n_1318), .Y(n_1397) );
AOI221xp5_ASAP7_75t_L g1398 ( .A1(n_1384), .A2(n_1369), .B1(n_1379), .B2(n_1375), .C(n_1383), .Y(n_1398) );
NOR3xp33_ASAP7_75t_SL g1399 ( .A(n_1389), .B(n_1371), .C(n_1373), .Y(n_1399) );
AOI21xp33_ASAP7_75t_L g1400 ( .A1(n_1387), .A2(n_1379), .B(n_1375), .Y(n_1400) );
OAI211xp5_ASAP7_75t_SL g1401 ( .A1(n_1386), .A2(n_1363), .B(n_1383), .C(n_1365), .Y(n_1401) );
NAND5xp2_ASAP7_75t_SL g1402 ( .A(n_1390), .B(n_1366), .C(n_1299), .D(n_1324), .E(n_1318), .Y(n_1402) );
XOR2xp5_ASAP7_75t_L g1403 ( .A(n_1385), .B(n_1226), .Y(n_1403) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1388), .Y(n_1404) );
AOI211xp5_ASAP7_75t_L g1405 ( .A1(n_1392), .A2(n_1366), .B(n_1304), .C(n_1299), .Y(n_1405) );
AOI221xp5_ASAP7_75t_L g1406 ( .A1(n_1393), .A2(n_1373), .B1(n_1365), .B2(n_1235), .C(n_1245), .Y(n_1406) );
NOR2x1p5_ASAP7_75t_L g1407 ( .A(n_1404), .B(n_1395), .Y(n_1407) );
INVx2_ASAP7_75t_L g1408 ( .A(n_1403), .Y(n_1408) );
BUFx3_ASAP7_75t_L g1409 ( .A(n_1402), .Y(n_1409) );
INVx2_ASAP7_75t_L g1410 ( .A(n_1400), .Y(n_1410) );
INVx2_ASAP7_75t_L g1411 ( .A(n_1398), .Y(n_1411) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1399), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1401), .Y(n_1413) );
OR3x1_ASAP7_75t_L g1414 ( .A(n_1412), .B(n_1405), .C(n_1391), .Y(n_1414) );
NOR5xp2_ASAP7_75t_L g1415 ( .A(n_1413), .B(n_1406), .C(n_1394), .D(n_1397), .E(n_1396), .Y(n_1415) );
NOR5xp2_ASAP7_75t_L g1416 ( .A(n_1410), .B(n_1205), .C(n_1221), .D(n_1216), .E(n_1150), .Y(n_1416) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1407), .Y(n_1417) );
NOR3xp33_ASAP7_75t_L g1418 ( .A(n_1410), .B(n_1273), .C(n_1195), .Y(n_1418) );
NOR2x1_ASAP7_75t_L g1419 ( .A(n_1417), .B(n_1409), .Y(n_1419) );
OAI31xp33_ASAP7_75t_L g1420 ( .A1(n_1415), .A2(n_1411), .A3(n_1409), .B(n_1408), .Y(n_1420) );
INVxp67_ASAP7_75t_L g1421 ( .A(n_1418), .Y(n_1421) );
INVx1_ASAP7_75t_L g1422 ( .A(n_1414), .Y(n_1422) );
OAI22xp5_ASAP7_75t_SL g1423 ( .A1(n_1422), .A2(n_1408), .B1(n_1416), .B2(n_1191), .Y(n_1423) );
XOR2x2_ASAP7_75t_L g1424 ( .A(n_1419), .B(n_1273), .Y(n_1424) );
OAI22xp5_ASAP7_75t_SL g1425 ( .A1(n_1420), .A2(n_1191), .B1(n_1300), .B2(n_1321), .Y(n_1425) );
OAI21xp5_ASAP7_75t_L g1426 ( .A1(n_1424), .A2(n_1421), .B(n_1191), .Y(n_1426) );
XNOR2xp5_ASAP7_75t_L g1427 ( .A(n_1425), .B(n_1261), .Y(n_1427) );
OAI22xp5_ASAP7_75t_L g1428 ( .A1(n_1423), .A2(n_1191), .B1(n_1321), .B2(n_1219), .Y(n_1428) );
AOI222xp33_ASAP7_75t_L g1429 ( .A1(n_1426), .A2(n_1427), .B1(n_1428), .B2(n_1191), .C1(n_1221), .C2(n_1216), .Y(n_1429) );
AOI22x1_ASAP7_75t_L g1430 ( .A1(n_1429), .A2(n_1189), .B1(n_1261), .B2(n_1248), .Y(n_1430) );
AOI221xp5_ASAP7_75t_L g1431 ( .A1(n_1430), .A2(n_1247), .B1(n_1252), .B2(n_1254), .C(n_1251), .Y(n_1431) );
endmodule