module real_aes_2524_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_564;
wire n_638;
wire n_519;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_817;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_146;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_762;
wire n_325;
wire n_575;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_0), .B(n_137), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_1), .A2(n_119), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_2), .B(n_792), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_3), .A2(n_11), .B1(n_807), .B2(n_808), .Y(n_806) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_3), .Y(n_808) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_4), .B(n_127), .Y(n_183) );
INVx1_ASAP7_75t_L g124 ( .A(n_5), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_6), .B(n_127), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_7), .B(n_114), .Y(n_464) );
INVx1_ASAP7_75t_L g492 ( .A(n_8), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g792 ( .A(n_9), .Y(n_792) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_10), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_11), .Y(n_807) );
NAND2xp33_ASAP7_75t_L g164 ( .A(n_12), .B(n_131), .Y(n_164) );
INVx2_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
AOI221x1_ASAP7_75t_L g206 ( .A1(n_14), .A2(n_27), .B1(n_119), .B2(n_137), .C(n_207), .Y(n_206) );
CKINVDCx16_ASAP7_75t_R g427 ( .A(n_15), .Y(n_427) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_16), .B(n_137), .Y(n_160) );
AO21x2_ASAP7_75t_L g157 ( .A1(n_17), .A2(n_158), .B(n_159), .Y(n_157) );
INVx1_ASAP7_75t_L g473 ( .A(n_18), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g814 ( .A(n_19), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_20), .B(n_150), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_21), .B(n_127), .Y(n_126) );
AO21x1_ASAP7_75t_L g178 ( .A1(n_22), .A2(n_137), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_L g430 ( .A(n_23), .Y(n_430) );
INVx1_ASAP7_75t_L g471 ( .A(n_24), .Y(n_471) );
INVx1_ASAP7_75t_SL g457 ( .A(n_25), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_26), .B(n_138), .Y(n_551) );
NAND2x1_ASAP7_75t_L g192 ( .A(n_28), .B(n_127), .Y(n_192) );
AOI33xp33_ASAP7_75t_L g519 ( .A1(n_29), .A2(n_55), .A3(n_447), .B1(n_454), .B2(n_520), .B3(n_521), .Y(n_519) );
NAND2x1_ASAP7_75t_L g146 ( .A(n_30), .B(n_131), .Y(n_146) );
INVx1_ASAP7_75t_L g501 ( .A(n_31), .Y(n_501) );
OR2x2_ASAP7_75t_L g115 ( .A(n_32), .B(n_88), .Y(n_115) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_32), .A2(n_88), .B(n_116), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_33), .B(n_445), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_34), .B(n_131), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_35), .B(n_127), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_36), .B(n_131), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_37), .A2(n_119), .B(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g120 ( .A(n_38), .B(n_121), .Y(n_120) );
AND2x2_ASAP7_75t_L g135 ( .A(n_38), .B(n_124), .Y(n_135) );
INVx1_ASAP7_75t_L g453 ( .A(n_38), .Y(n_453) );
OR2x6_ASAP7_75t_L g428 ( .A(n_39), .B(n_429), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_40), .Y(n_503) );
XNOR2xp5_ASAP7_75t_L g773 ( .A(n_41), .B(n_774), .Y(n_773) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_42), .B(n_137), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_43), .B(n_445), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_44), .A2(n_114), .B1(n_154), .B2(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_45), .B(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_46), .A2(n_773), .B1(n_778), .B2(n_782), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_47), .B(n_138), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g140 ( .A(n_48), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_49), .B(n_131), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_50), .B(n_158), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_51), .B(n_138), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_52), .A2(n_119), .B(n_145), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g548 ( .A(n_53), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_54), .B(n_131), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_56), .B(n_138), .Y(n_531) );
INVx1_ASAP7_75t_L g123 ( .A(n_57), .Y(n_123) );
INVx1_ASAP7_75t_L g133 ( .A(n_57), .Y(n_133) );
AND2x2_ASAP7_75t_L g532 ( .A(n_58), .B(n_150), .Y(n_532) );
AOI221xp5_ASAP7_75t_L g490 ( .A1(n_59), .A2(n_76), .B1(n_445), .B2(n_451), .C(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_60), .B(n_445), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_61), .B(n_127), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_62), .B(n_154), .Y(n_509) );
AOI21xp5_ASAP7_75t_SL g481 ( .A1(n_63), .A2(n_451), .B(n_482), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_64), .A2(n_119), .B(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g467 ( .A(n_65), .Y(n_467) );
AO21x1_ASAP7_75t_L g180 ( .A1(n_66), .A2(n_119), .B(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_67), .B(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g530 ( .A(n_68), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_69), .B(n_137), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_70), .A2(n_451), .B(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g229 ( .A(n_71), .B(n_151), .Y(n_229) );
INVx1_ASAP7_75t_L g121 ( .A(n_72), .Y(n_121) );
INVx1_ASAP7_75t_L g129 ( .A(n_72), .Y(n_129) );
AOI22xp5_ASAP7_75t_L g774 ( .A1(n_73), .A2(n_98), .B1(n_775), .B2(n_776), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g775 ( .A(n_73), .Y(n_775) );
AND2x2_ASAP7_75t_L g152 ( .A(n_74), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_75), .B(n_445), .Y(n_522) );
AND2x2_ASAP7_75t_L g460 ( .A(n_77), .B(n_153), .Y(n_460) );
INVx1_ASAP7_75t_L g468 ( .A(n_78), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_79), .A2(n_451), .B(n_456), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g549 ( .A1(n_80), .A2(n_451), .B(n_514), .C(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g431 ( .A(n_81), .Y(n_431) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_82), .B(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g166 ( .A(n_83), .B(n_153), .Y(n_166) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_84), .B(n_153), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_85), .A2(n_451), .B1(n_517), .B2(n_518), .Y(n_516) );
AOI222xp33_ASAP7_75t_L g102 ( .A1(n_86), .A2(n_103), .B1(n_785), .B2(n_796), .C1(n_815), .C2(n_817), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g803 ( .A1(n_86), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
CKINVDCx20_ASAP7_75t_R g804 ( .A(n_86), .Y(n_804) );
AND2x2_ASAP7_75t_L g179 ( .A(n_87), .B(n_114), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_89), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g196 ( .A(n_90), .B(n_153), .Y(n_196) );
INVx1_ASAP7_75t_L g483 ( .A(n_91), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_92), .B(n_127), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_93), .A2(n_119), .B(n_125), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_94), .B(n_131), .Y(n_208) );
AND2x2_ASAP7_75t_L g523 ( .A(n_95), .B(n_153), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_96), .B(n_127), .Y(n_171) );
A2O1A1Ixp33_ASAP7_75t_L g498 ( .A1(n_97), .A2(n_499), .B(n_500), .C(n_502), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g776 ( .A(n_98), .Y(n_776) );
BUFx2_ASAP7_75t_L g793 ( .A(n_99), .Y(n_793) );
BUFx2_ASAP7_75t_SL g821 ( .A(n_99), .Y(n_821) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_100), .A2(n_119), .B(n_162), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_101), .B(n_138), .Y(n_484) );
OAI21xp5_ASAP7_75t_SL g103 ( .A1(n_104), .A2(n_773), .B(n_777), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
OAI22xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_423), .B1(n_432), .B2(n_436), .Y(n_105) );
INVx2_ASAP7_75t_L g779 ( .A(n_106), .Y(n_779) );
XNOR2x1_ASAP7_75t_L g802 ( .A(n_106), .B(n_803), .Y(n_802) );
OR2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_321), .Y(n_106) );
NAND3xp33_ASAP7_75t_SL g107 ( .A(n_108), .B(n_233), .C(n_288), .Y(n_107) );
AOI221xp5_ASAP7_75t_L g108 ( .A1(n_109), .A2(n_173), .B1(n_197), .B2(n_201), .C(n_211), .Y(n_108) );
AND2x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_156), .Y(n_109) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_110), .B(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g232 ( .A(n_110), .Y(n_232) );
AND2x2_ASAP7_75t_L g277 ( .A(n_110), .B(n_214), .Y(n_277) );
AND2x4_ASAP7_75t_L g110 ( .A(n_111), .B(n_141), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_L g265 ( .A(n_112), .Y(n_265) );
INVx1_ASAP7_75t_L g275 ( .A(n_112), .Y(n_275) );
AO21x2_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_139), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_113), .B(n_140), .Y(n_139) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_113), .A2(n_117), .B(n_139), .Y(n_239) );
INVx1_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_114), .A2(n_160), .B(n_161), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_114), .B(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_114), .B(n_134), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_114), .A2(n_481), .B(n_485), .Y(n_480) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_115), .B(n_116), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_118), .B(n_136), .Y(n_117) );
AND2x6_ASAP7_75t_L g119 ( .A(n_120), .B(n_122), .Y(n_119) );
BUFx3_ASAP7_75t_L g449 ( .A(n_120), .Y(n_449) );
AND2x6_ASAP7_75t_L g131 ( .A(n_121), .B(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g455 ( .A(n_121), .Y(n_455) );
AND2x4_ASAP7_75t_L g451 ( .A(n_122), .B(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
AND2x4_ASAP7_75t_L g127 ( .A(n_123), .B(n_128), .Y(n_127) );
INVx2_ASAP7_75t_L g447 ( .A(n_123), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_124), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_130), .B(n_134), .Y(n_125) );
INVxp67_ASAP7_75t_L g474 ( .A(n_127), .Y(n_474) );
AND2x4_ASAP7_75t_L g138 ( .A(n_128), .B(n_132), .Y(n_138) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVxp67_ASAP7_75t_L g472 ( .A(n_131), .Y(n_472) );
INVx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_134), .A2(n_146), .B(n_147), .Y(n_145) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_134), .A2(n_163), .B(n_164), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_134), .A2(n_171), .B(n_172), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_134), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_134), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_134), .A2(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_134), .A2(n_226), .B(n_227), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_SL g456 ( .A1(n_134), .A2(n_457), .B(n_458), .C(n_459), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_134), .A2(n_458), .B(n_483), .C(n_484), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_134), .A2(n_458), .B(n_492), .C(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g517 ( .A(n_134), .Y(n_517) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_134), .A2(n_458), .B(n_530), .C(n_531), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_134), .A2(n_551), .B(n_552), .Y(n_550) );
INVx5_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g137 ( .A(n_135), .B(n_138), .Y(n_137) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_135), .Y(n_502) );
INVx1_ASAP7_75t_L g469 ( .A(n_138), .Y(n_469) );
OR2x2_ASAP7_75t_L g254 ( .A(n_141), .B(n_157), .Y(n_254) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_141), .B(n_200), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_141), .B(n_165), .Y(n_298) );
INVx2_ASAP7_75t_L g307 ( .A(n_141), .Y(n_307) );
AND2x2_ASAP7_75t_L g328 ( .A(n_141), .B(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g412 ( .A(n_141), .B(n_231), .Y(n_412) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g240 ( .A(n_142), .B(n_165), .Y(n_240) );
AND2x2_ASAP7_75t_L g373 ( .A(n_142), .B(n_200), .Y(n_373) );
HB1xp67_ASAP7_75t_L g399 ( .A(n_142), .Y(n_399) );
AO21x2_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_149), .B(n_152), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_144), .B(n_148), .Y(n_143) );
AO21x2_ASAP7_75t_L g442 ( .A1(n_149), .A2(n_443), .B(n_460), .Y(n_442) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_150), .Y(n_149) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_150), .A2(n_168), .B(n_169), .Y(n_167) );
OA21x2_ASAP7_75t_L g205 ( .A1(n_150), .A2(n_206), .B(n_210), .Y(n_205) );
OA21x2_ASAP7_75t_L g217 ( .A1(n_150), .A2(n_206), .B(n_210), .Y(n_217) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx3_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_153), .A2(n_195), .B1(n_498), .B2(n_503), .Y(n_497) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_154), .B(n_506), .Y(n_505) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx4f_ASAP7_75t_L g158 ( .A(n_155), .Y(n_158) );
AND2x4_ASAP7_75t_L g327 ( .A(n_156), .B(n_328), .Y(n_327) );
AOI321xp33_ASAP7_75t_L g341 ( .A1(n_156), .A2(n_270), .A3(n_271), .B1(n_303), .B2(n_342), .C(n_345), .Y(n_341) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_165), .Y(n_156) );
BUFx3_ASAP7_75t_L g198 ( .A(n_157), .Y(n_198) );
INVx2_ASAP7_75t_L g231 ( .A(n_157), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_157), .B(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g264 ( .A(n_157), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g297 ( .A(n_157), .Y(n_297) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_158), .A2(n_490), .B(n_494), .Y(n_489) );
INVx2_ASAP7_75t_SL g514 ( .A(n_158), .Y(n_514) );
INVx5_ASAP7_75t_L g200 ( .A(n_165), .Y(n_200) );
NOR2x1_ASAP7_75t_SL g249 ( .A(n_165), .B(n_239), .Y(n_249) );
BUFx2_ASAP7_75t_L g344 ( .A(n_165), .Y(n_344) );
OR2x6_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVxp67_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_186), .Y(n_174) );
NOR2xp33_ASAP7_75t_SL g242 ( .A(n_175), .B(n_243), .Y(n_242) );
NOR4xp25_ASAP7_75t_L g345 ( .A(n_175), .B(n_339), .C(n_343), .D(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g383 ( .A(n_175), .Y(n_383) );
AND2x2_ASAP7_75t_L g417 ( .A(n_175), .B(n_357), .Y(n_417) );
BUFx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g218 ( .A(n_176), .Y(n_218) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g272 ( .A(n_177), .Y(n_272) );
OAI21x1_ASAP7_75t_SL g177 ( .A1(n_178), .A2(n_180), .B(n_184), .Y(n_177) );
INVx1_ASAP7_75t_L g185 ( .A(n_179), .Y(n_185) );
AOI33xp33_ASAP7_75t_L g413 ( .A1(n_186), .A2(n_215), .A3(n_246), .B1(n_262), .B2(n_368), .B3(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
AND2x2_ASAP7_75t_L g203 ( .A(n_187), .B(n_204), .Y(n_203) );
AND2x4_ASAP7_75t_L g213 ( .A(n_187), .B(n_214), .Y(n_213) );
BUFx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx2_ASAP7_75t_L g220 ( .A(n_188), .Y(n_220) );
INVxp67_ASAP7_75t_L g301 ( .A(n_188), .Y(n_301) );
AND2x2_ASAP7_75t_L g357 ( .A(n_188), .B(n_222), .Y(n_357) );
AO21x2_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_188) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_189), .A2(n_195), .B(n_196), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_190), .B(n_194), .Y(n_189) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_195), .A2(n_223), .B(n_229), .Y(n_222) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_195), .A2(n_223), .B(n_229), .Y(n_258) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_195), .A2(n_526), .B(n_532), .Y(n_525) );
AO21x2_ASAP7_75t_L g563 ( .A1(n_195), .A2(n_526), .B(n_532), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_197), .A2(n_379), .B(n_380), .Y(n_378) );
AND2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
AND2x2_ASAP7_75t_L g366 ( .A(n_198), .B(n_240), .Y(n_366) );
AND3x2_ASAP7_75t_L g368 ( .A(n_198), .B(n_252), .C(n_307), .Y(n_368) );
INVx3_ASAP7_75t_SL g320 ( .A(n_199), .Y(n_320) );
INVx4_ASAP7_75t_L g214 ( .A(n_200), .Y(n_214) );
AND2x2_ASAP7_75t_L g252 ( .A(n_200), .B(n_239), .Y(n_252) );
INVxp67_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
BUFx2_ASAP7_75t_L g246 ( .A(n_204), .Y(n_246) );
AND2x4_ASAP7_75t_L g271 ( .A(n_204), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g334 ( .A(n_204), .B(n_222), .Y(n_334) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g304 ( .A(n_205), .Y(n_304) );
HB1xp67_ASAP7_75t_L g326 ( .A(n_205), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_R g211 ( .A1(n_212), .A2(n_215), .B(n_219), .C(n_230), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g212 ( .A(n_213), .Y(n_212) );
AND2x2_ASAP7_75t_L g263 ( .A(n_214), .B(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_214), .B(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_214), .B(n_231), .Y(n_392) );
INVx1_ASAP7_75t_SL g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g374 ( .A(n_216), .B(n_364), .Y(n_374) );
AND2x2_ASAP7_75t_SL g216 ( .A(n_217), .B(n_218), .Y(n_216) );
AND2x2_ASAP7_75t_L g221 ( .A(n_217), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g243 ( .A(n_217), .B(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g259 ( .A(n_217), .B(n_260), .Y(n_259) );
AND2x4_ASAP7_75t_L g292 ( .A(n_217), .B(n_272), .Y(n_292) );
AND2x4_ASAP7_75t_L g257 ( .A(n_218), .B(n_258), .Y(n_257) );
OR2x2_ASAP7_75t_L g281 ( .A(n_218), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g319 ( .A(n_218), .B(n_244), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
AND2x2_ASAP7_75t_L g247 ( .A(n_220), .B(n_244), .Y(n_247) );
AND2x2_ASAP7_75t_L g262 ( .A(n_220), .B(n_222), .Y(n_262) );
BUFx2_ASAP7_75t_L g318 ( .A(n_220), .Y(n_318) );
AND2x2_ASAP7_75t_L g332 ( .A(n_220), .B(n_243), .Y(n_332) );
INVx2_ASAP7_75t_L g244 ( .A(n_222), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_224), .B(n_228), .Y(n_223) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_230), .A2(n_281), .B1(n_283), .B2(n_287), .Y(n_280) );
INVx2_ASAP7_75t_SL g311 ( .A(n_230), .Y(n_311) );
OR2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
AND2x2_ASAP7_75t_L g286 ( .A(n_231), .B(n_239), .Y(n_286) );
INVx1_ASAP7_75t_L g393 ( .A(n_232), .Y(n_393) );
NOR3xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_266), .C(n_280), .Y(n_233) );
OAI221xp5_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_241), .B1(n_245), .B2(n_248), .C(n_250), .Y(n_234) );
INVx1_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_240), .Y(n_236) );
INVxp67_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g294 ( .A(n_238), .Y(n_294) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_238), .Y(n_422) );
INVx1_ASAP7_75t_L g385 ( .A(n_240), .Y(n_385) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_240), .B(n_264), .Y(n_395) );
INVxp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_244), .B(n_272), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_246), .B(n_247), .Y(n_245) );
OR2x2_ASAP7_75t_L g278 ( .A(n_246), .B(n_279), .Y(n_278) );
INVx1_ASAP7_75t_L g356 ( .A(n_246), .Y(n_356) );
AND2x2_ASAP7_75t_L g291 ( .A(n_247), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g337 ( .A(n_249), .B(n_297), .Y(n_337) );
AND2x2_ASAP7_75t_L g414 ( .A(n_249), .B(n_412), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_255), .B1(n_262), .B2(n_263), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g273 ( .A(n_254), .B(n_274), .Y(n_273) );
INVx1_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_259), .Y(n_256) );
INVx2_ASAP7_75t_L g279 ( .A(n_257), .Y(n_279) );
AND2x4_ASAP7_75t_L g303 ( .A(n_257), .B(n_304), .Y(n_303) );
OAI21xp33_ASAP7_75t_SL g333 ( .A1(n_257), .A2(n_334), .B(n_335), .Y(n_333) );
AND2x2_ASAP7_75t_L g360 ( .A(n_257), .B(n_318), .Y(n_360) );
INVx2_ASAP7_75t_L g282 ( .A(n_258), .Y(n_282) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_258), .Y(n_315) );
INVx1_ASAP7_75t_SL g339 ( .A(n_259), .Y(n_339) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
BUFx2_ASAP7_75t_L g270 ( .A(n_261), .Y(n_270) );
AND2x4_ASAP7_75t_SL g364 ( .A(n_261), .B(n_282), .Y(n_364) );
AND2x2_ASAP7_75t_L g361 ( .A(n_264), .B(n_307), .Y(n_361) );
AND2x2_ASAP7_75t_L g387 ( .A(n_264), .B(n_373), .Y(n_387) );
HB1xp67_ASAP7_75t_L g309 ( .A(n_265), .Y(n_309) );
INVx1_ASAP7_75t_L g329 ( .A(n_265), .Y(n_329) );
OAI22xp33_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_273), .B1(n_276), .B2(n_278), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_269), .B(n_271), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_271), .B(n_282), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_271), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g410 ( .A(n_271), .Y(n_410) );
INVx2_ASAP7_75t_SL g335 ( .A(n_273), .Y(n_335) );
AND2x2_ASAP7_75t_L g347 ( .A(n_275), .B(n_307), .Y(n_347) );
INVx2_ASAP7_75t_L g353 ( .A(n_275), .Y(n_353) );
INVxp33_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g312 ( .A(n_278), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_281), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_L g403 ( .A(n_281), .Y(n_403) );
INVx1_ASAP7_75t_L g331 ( .A(n_283), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_284), .B(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g342 ( .A(n_286), .B(n_343), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_286), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_415) );
NOR3xp33_ASAP7_75t_L g288 ( .A(n_289), .B(n_310), .C(n_313), .Y(n_288) );
OAI221xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_293), .B1(n_295), .B2(n_299), .C(n_302), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_SL g408 ( .A(n_293), .Y(n_408) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g377 ( .A(n_294), .B(n_343), .Y(n_377) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g308 ( .A(n_297), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g379 ( .A(n_299), .Y(n_379) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g376 ( .A(n_300), .Y(n_376) );
INVx1_ASAP7_75t_L g382 ( .A(n_301), .Y(n_382) );
OR2x2_ASAP7_75t_L g405 ( .A(n_301), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
INVx1_ASAP7_75t_SL g314 ( .A(n_304), .Y(n_314) );
AND2x2_ASAP7_75t_L g384 ( .A(n_304), .B(n_364), .Y(n_384) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_304), .B(n_317), .Y(n_416) );
INVx1_ASAP7_75t_SL g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g421 ( .A(n_307), .Y(n_421) );
INVx1_ASAP7_75t_L g371 ( .A(n_309), .Y(n_371) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
O2A1O1Ixp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B(n_316), .C(n_320), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_314), .B(n_364), .Y(n_388) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_317), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x2_ASAP7_75t_L g325 ( .A(n_319), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g406 ( .A(n_319), .Y(n_406) );
NAND4xp75_ASAP7_75t_L g321 ( .A(n_322), .B(n_378), .C(n_394), .D(n_415), .Y(n_321) );
NOR3x1_ASAP7_75t_L g322 ( .A(n_323), .B(n_340), .C(n_362), .Y(n_322) );
NAND4xp75_ASAP7_75t_L g323 ( .A(n_324), .B(n_330), .C(n_333), .D(n_336), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_325), .B(n_327), .Y(n_324) );
AND2x2_ASAP7_75t_L g375 ( .A(n_326), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g400 ( .A(n_327), .Y(n_400) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_SL g389 ( .A(n_332), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_341), .B(n_348), .Y(n_340) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_344), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_354), .B(n_358), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OAI322xp33_ASAP7_75t_L g380 ( .A1(n_352), .A2(n_381), .A3(n_385), .B1(n_386), .B2(n_388), .C1(n_389), .C2(n_390), .Y(n_380) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_353), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_356), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_357), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
OAI211xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_365), .B(n_367), .C(n_369), .Y(n_362) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_374), .B1(n_375), .B2(n_377), .Y(n_369) );
NOR2xp33_ASAP7_75t_SL g370 ( .A(n_371), .B(n_372), .Y(n_370) );
INVx2_ASAP7_75t_SL g372 ( .A(n_373), .Y(n_372) );
AOI21xp5_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_383), .B(n_384), .Y(n_381) );
INVxp67_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g419 ( .A(n_387), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_SL g390 ( .A(n_391), .B(n_393), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g397 ( .A(n_392), .B(n_398), .Y(n_397) );
O2A1O1Ixp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_396), .B(n_401), .C(n_404), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g396 ( .A(n_397), .B(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI221xp5_ASAP7_75t_SL g404 ( .A1(n_405), .A2(n_407), .B1(n_409), .B2(n_411), .C(n_413), .Y(n_404) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
CKINVDCx6p67_ASAP7_75t_R g423 ( .A(n_424), .Y(n_423) );
INVx4_ASAP7_75t_SL g780 ( .A(n_424), .Y(n_780) );
INVx3_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_426), .Y(n_425) );
AND2x6_ASAP7_75t_SL g426 ( .A(n_427), .B(n_428), .Y(n_426) );
OR2x6_ASAP7_75t_SL g434 ( .A(n_427), .B(n_435), .Y(n_434) );
OR2x2_ASAP7_75t_L g784 ( .A(n_427), .B(n_428), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_427), .B(n_435), .Y(n_795) );
CKINVDCx5p33_ASAP7_75t_R g435 ( .A(n_428), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
CKINVDCx11_ASAP7_75t_R g433 ( .A(n_434), .Y(n_433) );
OAI22x1_ASAP7_75t_L g778 ( .A1(n_434), .A2(n_779), .B1(n_780), .B2(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_436), .Y(n_781) );
OR3x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_638), .C(n_709), .Y(n_436) );
NAND3x1_ASAP7_75t_SL g437 ( .A(n_438), .B(n_565), .C(n_587), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_555), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_486), .B1(n_533), .B2(n_537), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_440), .A2(n_741), .B1(n_742), .B2(n_744), .Y(n_740) );
AND2x2_ASAP7_75t_L g440 ( .A(n_441), .B(n_461), .Y(n_440) );
AND2x2_ASAP7_75t_L g556 ( .A(n_441), .B(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_441), .B(n_603), .Y(n_622) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g540 ( .A(n_442), .Y(n_540) );
AND2x2_ASAP7_75t_L g590 ( .A(n_442), .B(n_463), .Y(n_590) );
INVx1_ASAP7_75t_L g629 ( .A(n_442), .Y(n_629) );
OR2x2_ASAP7_75t_L g666 ( .A(n_442), .B(n_478), .Y(n_666) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_442), .Y(n_678) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_442), .Y(n_702) );
AND2x2_ASAP7_75t_L g759 ( .A(n_442), .B(n_586), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_444), .B(n_450), .Y(n_443) );
INVx1_ASAP7_75t_L g510 ( .A(n_445), .Y(n_510) );
AND2x4_ASAP7_75t_L g445 ( .A(n_446), .B(n_449), .Y(n_445) );
INVx1_ASAP7_75t_L g546 ( .A(n_446), .Y(n_546) );
AND2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_448), .Y(n_446) );
OR2x6_ASAP7_75t_L g458 ( .A(n_447), .B(n_455), .Y(n_458) );
INVxp33_ASAP7_75t_L g520 ( .A(n_447), .Y(n_520) );
INVx1_ASAP7_75t_L g547 ( .A(n_449), .Y(n_547) );
INVxp67_ASAP7_75t_L g508 ( .A(n_451), .Y(n_508) );
NOR2x1p5_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx1_ASAP7_75t_L g521 ( .A(n_454), .Y(n_521) );
INVx3_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_458), .A2(n_467), .B1(n_468), .B2(n_469), .Y(n_466) );
INVxp67_ASAP7_75t_L g499 ( .A(n_458), .Y(n_499) );
INVx2_ASAP7_75t_L g553 ( .A(n_458), .Y(n_553) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_476), .Y(n_461) );
INVx1_ASAP7_75t_L g634 ( .A(n_462), .Y(n_634) );
AND2x2_ASAP7_75t_L g660 ( .A(n_462), .B(n_478), .Y(n_660) );
NAND2x1_ASAP7_75t_L g676 ( .A(n_462), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g557 ( .A(n_463), .B(n_543), .Y(n_557) );
INVx3_ASAP7_75t_L g586 ( .A(n_463), .Y(n_586) );
NOR2x1_ASAP7_75t_SL g705 ( .A(n_463), .B(n_478), .Y(n_705) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_470), .B(n_475), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_469), .B(n_501), .Y(n_500) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_472), .B1(n_473), .B2(n_474), .Y(n_470) );
NOR2x1_ASAP7_75t_L g613 ( .A(n_476), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g584 ( .A(n_477), .B(n_585), .Y(n_584) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx4_ASAP7_75t_L g554 ( .A(n_478), .Y(n_554) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_478), .Y(n_599) );
AND2x2_ASAP7_75t_L g671 ( .A(n_478), .B(n_543), .Y(n_671) );
AND2x4_ASAP7_75t_L g688 ( .A(n_478), .B(n_632), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g735 ( .A(n_478), .B(n_630), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_478), .B(n_539), .Y(n_764) );
OR2x6_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_486), .A2(n_581), .B1(n_652), .B2(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_511), .Y(n_486) );
INVx2_ASAP7_75t_L g654 ( .A(n_487), .Y(n_654) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_495), .Y(n_487) );
BUFx3_ASAP7_75t_L g644 ( .A(n_488), .Y(n_644) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_489), .B(n_513), .Y(n_536) );
INVx2_ASAP7_75t_L g560 ( .A(n_489), .Y(n_560) );
INVx1_ASAP7_75t_L g572 ( .A(n_489), .Y(n_572) );
AND2x4_ASAP7_75t_L g579 ( .A(n_489), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g596 ( .A(n_489), .B(n_496), .Y(n_596) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_489), .Y(n_610) );
INVxp67_ASAP7_75t_L g618 ( .A(n_489), .Y(n_618) );
AND2x2_ASAP7_75t_L g647 ( .A(n_495), .B(n_563), .Y(n_647) );
AND2x2_ASAP7_75t_L g663 ( .A(n_495), .B(n_564), .Y(n_663) );
NOR2xp67_ASAP7_75t_L g750 ( .A(n_495), .B(n_563), .Y(n_750) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x4_ASAP7_75t_L g559 ( .A(n_496), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g570 ( .A(n_496), .Y(n_570) );
INVx1_ASAP7_75t_L g583 ( .A(n_496), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_496), .B(n_525), .Y(n_620) );
OR2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_504), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_508), .B1(n_509), .B2(n_510), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g743 ( .A(n_511), .Y(n_743) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_524), .Y(n_511) );
AND2x2_ASAP7_75t_L g617 ( .A(n_512), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g646 ( .A(n_512), .Y(n_646) );
AND2x2_ASAP7_75t_L g748 ( .A(n_512), .B(n_563), .Y(n_748) );
INVx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_513), .B(n_525), .Y(n_608) );
AO21x2_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B(n_523), .Y(n_513) );
AO21x2_ASAP7_75t_L g564 ( .A1(n_514), .A2(n_515), .B(n_523), .Y(n_564) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g534 ( .A(n_524), .Y(n_534) );
NAND2x1p5_ASAP7_75t_L g723 ( .A(n_524), .B(n_644), .Y(n_723) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_525), .Y(n_637) );
AND2x2_ASAP7_75t_L g664 ( .A(n_525), .B(n_610), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_528), .Y(n_526) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g578 ( .A(n_534), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g594 ( .A(n_534), .Y(n_594) );
AND2x2_ASAP7_75t_L g682 ( .A(n_534), .B(n_559), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_534), .B(n_702), .Y(n_707) );
AND2x2_ASAP7_75t_L g717 ( .A(n_534), .B(n_596), .Y(n_717) );
OR2x2_ASAP7_75t_L g754 ( .A(n_534), .B(n_654), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_535), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g714 ( .A(n_535), .B(n_570), .Y(n_714) );
AND2x2_ASAP7_75t_L g730 ( .A(n_535), .B(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g724 ( .A(n_536), .B(n_620), .Y(n_724) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_541), .Y(n_537) );
INVx1_ASAP7_75t_L g606 ( .A(n_538), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_538), .B(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g704 ( .A(n_538), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_538), .B(n_585), .Y(n_729) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_539), .Y(n_576) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_540), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_541), .A2(n_574), .B1(n_592), .B2(n_595), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_541), .B(n_676), .Y(n_675) );
INVx2_ASAP7_75t_SL g708 ( .A(n_541), .Y(n_708) );
AND2x4_ASAP7_75t_SL g541 ( .A(n_542), .B(n_554), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g585 ( .A(n_543), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g605 ( .A(n_543), .Y(n_605) );
INVx1_ASAP7_75t_L g632 ( .A(n_543), .Y(n_632) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_549), .Y(n_543) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .C(n_548), .Y(n_545) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_554), .Y(n_574) );
AND2x4_ASAP7_75t_L g631 ( .A(n_554), .B(n_632), .Y(n_631) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_554), .B(n_661), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
AND2x2_ASAP7_75t_L g656 ( .A(n_556), .B(n_599), .Y(n_656) );
OAI21xp5_ASAP7_75t_L g736 ( .A1(n_556), .A2(n_737), .B(n_738), .Y(n_736) );
INVx2_ASAP7_75t_L g614 ( .A(n_557), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_558), .A2(n_668), .B1(n_672), .B2(n_675), .Y(n_667) );
AND2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_561), .Y(n_558) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_559), .Y(n_625) );
AND2x2_ASAP7_75t_L g635 ( .A(n_559), .B(n_636), .Y(n_635) );
INVx3_ASAP7_75t_L g674 ( .A(n_559), .Y(n_674) );
NAND2x1_ASAP7_75t_SL g699 ( .A(n_559), .B(n_568), .Y(n_699) );
AND2x2_ASAP7_75t_L g595 ( .A(n_561), .B(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_563), .B(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g568 ( .A(n_564), .Y(n_568) );
INVx2_ASAP7_75t_L g580 ( .A(n_564), .Y(n_580) );
AOI21xp5_ASAP7_75t_SL g565 ( .A1(n_566), .A2(n_573), .B(n_577), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_568), .B(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_569), .A2(n_658), .B1(n_662), .B2(n_665), .Y(n_657) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
BUFx2_ASAP7_75t_L g762 ( .A(n_570), .Y(n_762) );
INVx1_ASAP7_75t_SL g769 ( .A(n_570), .Y(n_769) );
HB1xp67_ASAP7_75t_L g732 ( .A(n_571), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_581), .B(n_584), .Y(n_577) );
AND2x2_ASAP7_75t_L g581 ( .A(n_579), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g623 ( .A(n_579), .B(n_619), .Y(n_623) );
AND2x2_ASAP7_75t_L g738 ( .A(n_579), .B(n_636), .Y(n_738) );
AND2x2_ASAP7_75t_L g741 ( .A(n_579), .B(n_647), .Y(n_741) );
AND2x4_ASAP7_75t_L g749 ( .A(n_579), .B(n_750), .Y(n_749) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_581), .A2(n_704), .B(n_706), .Y(n_703) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g731 ( .A(n_583), .Y(n_731) );
AND2x2_ASAP7_75t_L g747 ( .A(n_583), .B(n_748), .Y(n_747) );
INVx4_ASAP7_75t_L g661 ( .A(n_585), .Y(n_661) );
INVx1_ASAP7_75t_L g630 ( .A(n_586), .Y(n_630) );
AND2x2_ASAP7_75t_L g652 ( .A(n_586), .B(n_605), .Y(n_652) );
NOR2x1_ASAP7_75t_L g587 ( .A(n_588), .B(n_611), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_591), .B(n_597), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g598 ( .A(n_590), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_SL g751 ( .A(n_590), .B(n_603), .Y(n_751) );
AND2x2_ASAP7_75t_L g772 ( .A(n_590), .B(n_688), .Y(n_772) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g698 ( .A(n_595), .Y(n_698) );
OAI21xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_600), .B(n_607), .Y(n_597) );
OR2x6_ASAP7_75t_L g650 ( .A(n_599), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_602), .B(n_606), .Y(n_601) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
OR2x2_ASAP7_75t_L g673 ( .A(n_608), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g770 ( .A(n_608), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_609), .B(n_743), .Y(n_742) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_624), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B1(n_621), .B2(n_623), .Y(n_612) );
OR2x2_ASAP7_75t_L g684 ( .A(n_614), .B(n_685), .Y(n_684) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
HB1xp67_ASAP7_75t_L g641 ( .A(n_616), .Y(n_641) );
NAND2x1p5_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .Y(n_616) );
INVx1_ASAP7_75t_L g690 ( .A(n_619), .Y(n_690) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
INVxp67_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_633), .B2(n_635), .Y(n_624) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_631), .Y(n_627) );
AND2x4_ASAP7_75t_SL g628 ( .A(n_629), .B(n_630), .Y(n_628) );
AND2x2_ASAP7_75t_L g633 ( .A(n_631), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g694 ( .A(n_634), .B(n_688), .Y(n_694) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_639), .B(n_679), .Y(n_638) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_640), .B(n_653), .Y(n_639) );
AOI21xp33_ASAP7_75t_SL g640 ( .A1(n_641), .A2(n_642), .B(n_648), .Y(n_640) );
OR2x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
INVx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2x1p5_ASAP7_75t_L g645 ( .A(n_646), .B(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
OAI22xp33_ASAP7_75t_SL g718 ( .A1(n_650), .A2(n_719), .B1(n_721), .B2(n_724), .Y(n_718) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_651), .B(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g701 ( .A(n_652), .B(n_702), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_655), .B(n_657), .C(n_667), .Y(n_653) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp33_ASAP7_75t_SL g658 ( .A(n_659), .B(n_661), .Y(n_658) );
INVxp33_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g670 ( .A(n_661), .Y(n_670) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_662), .A2(n_682), .B1(n_683), .B2(n_686), .C(n_689), .Y(n_681) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx1_ASAP7_75t_L g722 ( .A(n_663), .Y(n_722) );
INVx2_ASAP7_75t_SL g720 ( .A(n_666), .Y(n_720) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
NAND2x1_ASAP7_75t_L g719 ( .A(n_670), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g716 ( .A(n_676), .Y(n_716) );
INVx1_ASAP7_75t_L g745 ( .A(n_677), .Y(n_745) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
NOR2x1_ASAP7_75t_L g679 ( .A(n_680), .B(n_695), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_693), .Y(n_680) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g734 ( .A(n_685), .Y(n_734) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g755 ( .A(n_688), .B(n_756), .Y(n_755) );
INVx2_ASAP7_75t_L g760 ( .A(n_688), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
INVxp33_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx2_ASAP7_75t_L g713 ( .A(n_692), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g695 ( .A1(n_696), .A2(n_700), .B(n_703), .Y(n_695) );
INVxp67_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g756 ( .A(n_702), .Y(n_756) );
AND2x2_ASAP7_75t_L g744 ( .A(n_705), .B(n_745), .Y(n_744) );
NOR2xp33_ASAP7_75t_R g706 ( .A(n_707), .B(n_708), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_725), .C(n_752), .Y(n_709) );
NOR2xp33_ASAP7_75t_L g710 ( .A(n_711), .B(n_718), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_712), .B(n_715), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
OR2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_723), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_726), .B(n_739), .Y(n_725) );
NAND2xp5_ASAP7_75t_SL g726 ( .A(n_727), .B(n_736), .Y(n_726) );
AOI22xp33_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_730), .B1(n_732), .B2(n_733), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVxp67_ASAP7_75t_SL g737 ( .A(n_735), .Y(n_737) );
NAND2xp5_ASAP7_75t_SL g739 ( .A(n_740), .B(n_746), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B(n_751), .Y(n_746) );
INVx1_ASAP7_75t_L g765 ( .A(n_749), .Y(n_765) );
AOI211xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_755), .B(n_757), .C(n_766), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g757 ( .A1(n_758), .A2(n_761), .B1(n_763), .B2(n_765), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
HB1xp67_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_767), .B(n_771), .Y(n_766) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
INVxp67_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
BUFx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g787 ( .A(n_788), .B(n_794), .Y(n_787) );
INVxp67_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_790), .B(n_793), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
OR2x2_ASAP7_75t_SL g816 ( .A(n_791), .B(n_793), .Y(n_816) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_791), .A2(n_819), .B(n_822), .Y(n_818) );
BUFx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx2_ASAP7_75t_R g800 ( .A(n_795), .Y(n_800) );
BUFx3_ASAP7_75t_L g813 ( .A(n_795), .Y(n_813) );
BUFx2_ASAP7_75t_L g823 ( .A(n_795), .Y(n_823) );
INVxp33_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_801), .B(n_809), .Y(n_797) );
INVx1_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
CKINVDCx20_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
NOR2xp33_ASAP7_75t_SL g809 ( .A(n_810), .B(n_814), .Y(n_809) );
INVx1_ASAP7_75t_SL g810 ( .A(n_811), .Y(n_810) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
INVx1_ASAP7_75t_SL g817 ( .A(n_818), .Y(n_817) );
CKINVDCx11_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
CKINVDCx8_ASAP7_75t_R g820 ( .A(n_821), .Y(n_820) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
endmodule